module basic_2500_25000_3000_20_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
nand U0 (N_0,In_2243,In_2177);
xnor U1 (N_1,In_677,In_2217);
nand U2 (N_2,In_1782,In_423);
xor U3 (N_3,In_892,In_1000);
nand U4 (N_4,In_1309,In_2061);
nor U5 (N_5,In_1852,In_866);
nand U6 (N_6,In_1461,In_2241);
or U7 (N_7,In_991,In_2419);
nor U8 (N_8,In_1666,In_535);
nand U9 (N_9,In_1975,In_2411);
nand U10 (N_10,In_561,In_327);
nand U11 (N_11,In_941,In_753);
nand U12 (N_12,In_859,In_1277);
nor U13 (N_13,In_161,In_40);
nand U14 (N_14,In_108,In_17);
or U15 (N_15,In_2308,In_1516);
or U16 (N_16,In_545,In_1158);
nand U17 (N_17,In_2418,In_2227);
or U18 (N_18,In_780,In_169);
and U19 (N_19,In_1134,In_1676);
and U20 (N_20,In_1818,In_1577);
xor U21 (N_21,In_2303,In_2468);
or U22 (N_22,In_1179,In_2181);
xor U23 (N_23,In_928,In_2461);
nand U24 (N_24,In_1026,In_1282);
nor U25 (N_25,In_246,In_673);
nor U26 (N_26,In_860,In_874);
nor U27 (N_27,In_1702,In_661);
and U28 (N_28,In_412,In_1426);
or U29 (N_29,In_1028,In_1694);
nor U30 (N_30,In_585,In_1456);
or U31 (N_31,In_1332,In_482);
nor U32 (N_32,In_1752,In_1020);
or U33 (N_33,In_1249,In_1418);
or U34 (N_34,In_121,In_362);
nand U35 (N_35,In_1692,In_1596);
xnor U36 (N_36,In_95,In_1485);
or U37 (N_37,In_1019,In_1403);
and U38 (N_38,In_2380,In_2148);
or U39 (N_39,In_675,In_1711);
or U40 (N_40,In_557,In_2037);
xnor U41 (N_41,In_1725,In_1305);
nand U42 (N_42,In_1992,In_666);
or U43 (N_43,In_767,In_578);
or U44 (N_44,In_1447,In_2162);
or U45 (N_45,In_1776,In_1270);
nor U46 (N_46,In_2230,In_2004);
nand U47 (N_47,In_1371,In_225);
xnor U48 (N_48,In_875,In_354);
and U49 (N_49,In_91,In_1482);
and U50 (N_50,In_2363,In_1192);
nand U51 (N_51,In_850,In_1664);
or U52 (N_52,In_1651,In_182);
nor U53 (N_53,In_1040,In_1677);
nand U54 (N_54,In_2280,In_278);
nand U55 (N_55,In_1204,In_387);
xnor U56 (N_56,In_747,In_708);
nor U57 (N_57,In_956,In_1458);
and U58 (N_58,In_397,In_490);
nor U59 (N_59,In_1759,In_1015);
or U60 (N_60,In_1377,In_349);
and U61 (N_61,In_867,In_712);
nand U62 (N_62,In_119,In_1048);
and U63 (N_63,In_2034,In_757);
or U64 (N_64,In_717,In_1);
nor U65 (N_65,In_21,In_101);
nor U66 (N_66,In_605,In_378);
nor U67 (N_67,In_1671,In_2111);
nor U68 (N_68,In_319,In_1727);
or U69 (N_69,In_313,In_250);
xnor U70 (N_70,In_614,In_2385);
nand U71 (N_71,In_32,In_220);
and U72 (N_72,In_152,In_1295);
nor U73 (N_73,In_1720,In_1369);
nand U74 (N_74,In_1036,In_18);
and U75 (N_75,In_1043,In_1423);
nand U76 (N_76,In_832,In_2134);
nor U77 (N_77,In_120,In_587);
nand U78 (N_78,In_1566,In_2142);
nor U79 (N_79,In_2095,In_2193);
or U80 (N_80,In_758,In_751);
nor U81 (N_81,In_1092,In_694);
nor U82 (N_82,In_157,In_2174);
nor U83 (N_83,In_524,In_2469);
nand U84 (N_84,In_1935,In_573);
xor U85 (N_85,In_1500,In_174);
or U86 (N_86,In_392,In_2222);
and U87 (N_87,In_744,In_986);
nand U88 (N_88,In_1216,In_2291);
nor U89 (N_89,In_1652,In_176);
xnor U90 (N_90,In_809,In_2027);
nand U91 (N_91,In_238,In_1874);
nor U92 (N_92,In_2208,In_2321);
and U93 (N_93,In_623,In_1308);
nor U94 (N_94,In_1261,In_1795);
xnor U95 (N_95,In_510,In_1140);
and U96 (N_96,In_248,In_632);
xnor U97 (N_97,In_1153,In_416);
xor U98 (N_98,In_1001,In_418);
nand U99 (N_99,In_1582,In_1044);
or U100 (N_100,In_94,In_1053);
and U101 (N_101,In_555,In_78);
nand U102 (N_102,In_224,In_2078);
or U103 (N_103,In_1990,In_330);
nand U104 (N_104,In_797,In_343);
nand U105 (N_105,In_664,In_1619);
or U106 (N_106,In_500,In_1122);
and U107 (N_107,In_1487,In_1733);
nand U108 (N_108,In_1494,In_864);
and U109 (N_109,In_1382,In_1824);
and U110 (N_110,In_1235,In_1521);
xnor U111 (N_111,In_749,In_1346);
xor U112 (N_112,In_1835,In_1062);
xor U113 (N_113,In_1114,In_2190);
nor U114 (N_114,In_1334,In_1252);
and U115 (N_115,In_612,In_1735);
and U116 (N_116,In_2338,In_1680);
nor U117 (N_117,In_1004,In_1430);
or U118 (N_118,In_16,In_1258);
xnor U119 (N_119,In_1579,In_1643);
or U120 (N_120,In_1221,In_52);
xnor U121 (N_121,In_1862,In_2480);
nor U122 (N_122,In_630,In_400);
and U123 (N_123,In_854,In_266);
nor U124 (N_124,In_1368,In_2156);
or U125 (N_125,In_1289,In_787);
nor U126 (N_126,In_714,In_2220);
or U127 (N_127,In_1663,In_985);
nor U128 (N_128,In_1945,In_1478);
nand U129 (N_129,In_2441,In_1182);
xor U130 (N_130,In_214,In_1265);
nand U131 (N_131,In_1683,In_1262);
and U132 (N_132,In_764,In_1201);
xnor U133 (N_133,In_1223,In_1675);
or U134 (N_134,In_1095,In_1699);
xnor U135 (N_135,In_276,In_2015);
nand U136 (N_136,In_610,In_1564);
nor U137 (N_137,In_1187,In_1799);
nor U138 (N_138,In_2276,In_2149);
or U139 (N_139,In_2250,In_316);
nor U140 (N_140,In_2214,In_29);
nor U141 (N_141,In_1546,In_2347);
nand U142 (N_142,In_2056,In_766);
and U143 (N_143,In_1867,In_1137);
xor U144 (N_144,In_1833,In_2185);
nor U145 (N_145,In_1748,In_1061);
nand U146 (N_146,In_215,In_2284);
xnor U147 (N_147,In_1803,In_2368);
xor U148 (N_148,In_1805,In_639);
and U149 (N_149,In_1836,In_885);
nand U150 (N_150,In_1218,In_1467);
and U151 (N_151,In_2483,In_813);
xor U152 (N_152,In_1452,In_348);
xor U153 (N_153,In_2274,In_2235);
and U154 (N_154,In_922,In_242);
and U155 (N_155,In_56,In_329);
or U156 (N_156,In_73,In_116);
and U157 (N_157,In_1072,In_721);
nor U158 (N_158,In_1294,In_964);
nand U159 (N_159,In_1373,In_2163);
and U160 (N_160,In_1356,In_2332);
nor U161 (N_161,In_1076,In_754);
nand U162 (N_162,In_1339,In_2075);
and U163 (N_163,In_1283,In_381);
nor U164 (N_164,In_979,In_296);
nand U165 (N_165,In_665,In_48);
nor U166 (N_166,In_1413,In_1679);
nand U167 (N_167,In_822,In_204);
xor U168 (N_168,In_2081,In_304);
nor U169 (N_169,In_1248,In_1366);
xnor U170 (N_170,In_226,In_2172);
xor U171 (N_171,In_2089,In_734);
and U172 (N_172,In_39,In_435);
and U173 (N_173,In_597,In_2209);
xnor U174 (N_174,In_1816,In_1585);
xnor U175 (N_175,In_1385,In_30);
nor U176 (N_176,In_2216,In_2012);
nand U177 (N_177,In_2481,In_801);
nor U178 (N_178,In_1657,In_1125);
or U179 (N_179,In_363,In_974);
nand U180 (N_180,In_485,In_852);
xor U181 (N_181,In_299,In_2110);
xnor U182 (N_182,In_772,In_1693);
xor U183 (N_183,In_1817,In_1988);
nand U184 (N_184,In_2117,In_911);
and U185 (N_185,In_1139,In_2240);
nor U186 (N_186,In_2329,In_1572);
or U187 (N_187,In_1230,In_393);
nand U188 (N_188,In_2159,In_2327);
nand U189 (N_189,In_36,In_2470);
nor U190 (N_190,In_893,In_1082);
xnor U191 (N_191,In_105,In_306);
nand U192 (N_192,In_1200,In_762);
xor U193 (N_193,In_653,In_443);
nand U194 (N_194,In_1132,In_1673);
xor U195 (N_195,In_984,In_2266);
nor U196 (N_196,In_310,In_978);
nand U197 (N_197,In_1491,In_2350);
and U198 (N_198,In_1633,In_687);
nor U199 (N_199,In_2140,In_962);
and U200 (N_200,In_2377,In_567);
and U201 (N_201,In_1639,In_1448);
and U202 (N_202,In_541,In_2073);
xnor U203 (N_203,In_129,In_1916);
or U204 (N_204,In_2492,In_1731);
xor U205 (N_205,In_1864,In_1970);
nand U206 (N_206,In_1454,In_1925);
or U207 (N_207,In_829,In_335);
and U208 (N_208,In_2334,In_814);
xnor U209 (N_209,In_1505,In_2277);
and U210 (N_210,In_1296,In_1831);
nor U211 (N_211,In_2031,In_1495);
nor U212 (N_212,In_2044,In_1592);
and U213 (N_213,In_1987,In_124);
or U214 (N_214,In_185,In_658);
xor U215 (N_215,In_1220,In_1163);
nand U216 (N_216,In_223,In_2085);
nand U217 (N_217,In_1588,In_1736);
nor U218 (N_218,In_1996,In_861);
nand U219 (N_219,In_1597,In_2491);
xnor U220 (N_220,In_1462,In_1393);
and U221 (N_221,In_1492,In_640);
xnor U222 (N_222,In_562,In_2030);
or U223 (N_223,In_1553,In_2378);
nor U224 (N_224,In_1190,In_1707);
or U225 (N_225,In_543,In_2158);
nor U226 (N_226,In_1861,In_61);
and U227 (N_227,In_1209,In_1035);
xor U228 (N_228,In_291,In_533);
nor U229 (N_229,In_759,In_2108);
nand U230 (N_230,In_656,In_2320);
xnor U231 (N_231,In_1922,In_868);
and U232 (N_232,In_1840,In_1421);
nor U233 (N_233,In_1108,In_1018);
or U234 (N_234,In_913,In_389);
and U235 (N_235,In_1606,In_1321);
xor U236 (N_236,In_1510,In_2397);
xor U237 (N_237,In_1921,In_1515);
nand U238 (N_238,In_835,In_1376);
nand U239 (N_239,In_2169,In_147);
nor U240 (N_240,In_494,In_2290);
or U241 (N_241,In_360,In_512);
or U242 (N_242,In_1595,In_1007);
xnor U243 (N_243,In_2183,In_2428);
or U244 (N_244,In_507,In_253);
and U245 (N_245,In_473,In_1146);
or U246 (N_246,In_607,In_1744);
nor U247 (N_247,In_775,In_463);
xor U248 (N_248,In_257,In_680);
nor U249 (N_249,In_1049,In_1884);
or U250 (N_250,In_209,In_1207);
nor U251 (N_251,In_931,In_1243);
nor U252 (N_252,In_331,In_615);
nand U253 (N_253,In_583,In_1297);
xor U254 (N_254,In_647,In_830);
or U255 (N_255,In_28,In_1714);
xnor U256 (N_256,In_989,In_655);
or U257 (N_257,In_145,In_38);
xor U258 (N_258,In_1106,In_1721);
or U259 (N_259,In_1875,In_1877);
or U260 (N_260,In_12,In_47);
and U261 (N_261,In_445,In_602);
or U262 (N_262,In_1016,In_1766);
or U263 (N_263,In_2001,In_2165);
or U264 (N_264,In_1837,In_1775);
xnor U265 (N_265,In_2288,In_1934);
xor U266 (N_266,In_1199,In_2410);
nor U267 (N_267,In_1417,In_774);
nor U268 (N_268,In_2057,In_2067);
and U269 (N_269,In_847,In_200);
nand U270 (N_270,In_1710,In_409);
or U271 (N_271,In_2353,In_14);
nand U272 (N_272,In_1168,In_1617);
and U273 (N_273,In_840,In_540);
and U274 (N_274,In_1509,In_1800);
nor U275 (N_275,In_641,In_2325);
xnor U276 (N_276,In_2248,In_2166);
nor U277 (N_277,In_2053,In_2340);
nand U278 (N_278,In_342,In_2115);
nor U279 (N_279,In_83,In_1902);
and U280 (N_280,In_1056,In_340);
and U281 (N_281,In_790,In_2475);
nand U282 (N_282,In_888,In_670);
xor U283 (N_283,In_395,In_1629);
and U284 (N_284,In_1611,In_1365);
or U285 (N_285,In_2489,In_1580);
nand U286 (N_286,In_1599,In_2379);
and U287 (N_287,In_1010,In_1976);
nand U288 (N_288,In_2436,In_2023);
nor U289 (N_289,In_1656,In_2179);
nand U290 (N_290,In_1450,In_1333);
xor U291 (N_291,In_87,In_1326);
nand U292 (N_292,In_2007,In_1713);
nor U293 (N_293,In_1121,In_803);
xnor U294 (N_294,In_333,In_1507);
nor U295 (N_295,In_2074,In_1567);
xnor U296 (N_296,In_1627,In_460);
and U297 (N_297,In_77,In_290);
and U298 (N_298,In_150,In_599);
and U299 (N_299,In_195,In_122);
nand U300 (N_300,In_1436,In_943);
nand U301 (N_301,In_791,In_312);
or U302 (N_302,In_1930,In_2005);
xor U303 (N_303,In_206,In_383);
nor U304 (N_304,In_1378,In_1244);
nor U305 (N_305,In_1821,In_2096);
xnor U306 (N_306,In_2414,In_547);
nand U307 (N_307,In_1695,In_264);
nor U308 (N_308,In_2102,In_2333);
xnor U309 (N_309,In_1498,In_722);
nor U310 (N_310,In_1267,In_1463);
xor U311 (N_311,In_846,In_1685);
nand U312 (N_312,In_551,In_626);
and U313 (N_313,In_1012,In_203);
nand U314 (N_314,In_1778,In_351);
xor U315 (N_315,In_904,In_2315);
or U316 (N_316,In_593,In_1499);
and U317 (N_317,In_1425,In_74);
or U318 (N_318,In_2261,In_2259);
nor U319 (N_319,In_2197,In_422);
xnor U320 (N_320,In_272,In_1757);
nor U321 (N_321,In_1688,In_1075);
nand U322 (N_322,In_1375,In_542);
xor U323 (N_323,In_45,In_1081);
xor U324 (N_324,In_2429,In_1832);
nor U325 (N_325,In_2060,In_2354);
nand U326 (N_326,In_144,In_1374);
nor U327 (N_327,In_148,In_2297);
and U328 (N_328,In_287,In_2021);
nand U329 (N_329,In_1610,In_1900);
nand U330 (N_330,In_539,In_1931);
nor U331 (N_331,In_2038,In_1440);
nand U332 (N_332,In_824,In_235);
and U333 (N_333,In_322,In_1324);
nand U334 (N_334,In_821,In_2415);
nor U335 (N_335,In_990,In_944);
nor U336 (N_336,In_1917,In_727);
and U337 (N_337,In_2192,In_2420);
nor U338 (N_338,In_576,In_2059);
and U339 (N_339,In_2239,In_725);
nand U340 (N_340,In_111,In_62);
nand U341 (N_341,In_82,In_2402);
xnor U342 (N_342,In_1362,In_1932);
and U343 (N_343,In_1780,In_281);
nand U344 (N_344,In_743,In_2364);
xor U345 (N_345,In_1013,In_796);
and U346 (N_346,In_1660,In_1392);
or U347 (N_347,In_31,In_1647);
nand U348 (N_348,In_1136,In_477);
or U349 (N_349,In_723,In_1008);
nand U350 (N_350,In_1957,In_1213);
nand U351 (N_351,In_437,In_158);
nand U352 (N_352,In_2445,In_384);
xor U353 (N_353,In_983,In_2225);
xor U354 (N_354,In_1287,In_1330);
or U355 (N_355,In_243,In_285);
and U356 (N_356,In_433,In_871);
xor U357 (N_357,In_891,In_921);
nor U358 (N_358,In_609,In_1549);
xor U359 (N_359,In_1941,In_2395);
nor U360 (N_360,In_190,In_800);
xnor U361 (N_361,In_1341,In_498);
and U362 (N_362,In_789,In_1233);
or U363 (N_363,In_2400,In_1202);
xor U364 (N_364,In_1238,In_1111);
and U365 (N_365,In_2346,In_1077);
or U366 (N_366,In_1396,In_2446);
and U367 (N_367,In_2330,In_2127);
xor U368 (N_368,In_2485,In_509);
and U369 (N_369,In_2292,In_1506);
xnor U370 (N_370,In_259,In_2466);
nand U371 (N_371,In_2154,In_950);
nand U372 (N_372,In_1969,In_96);
nor U373 (N_373,In_1032,In_2271);
nor U374 (N_374,In_845,In_2202);
or U375 (N_375,In_1208,In_421);
and U376 (N_376,In_1118,In_2294);
nand U377 (N_377,In_2186,In_692);
xnor U378 (N_378,In_2157,In_321);
nand U379 (N_379,In_447,In_1355);
nor U380 (N_380,In_716,In_1227);
or U381 (N_381,In_2211,In_1255);
xnor U382 (N_382,In_1593,In_154);
or U383 (N_383,In_411,In_760);
nand U384 (N_384,In_429,In_2467);
nor U385 (N_385,In_1046,In_1944);
or U386 (N_386,In_1621,In_1428);
and U387 (N_387,In_1089,In_1850);
and U388 (N_388,In_1166,In_2135);
and U389 (N_389,In_579,In_2464);
or U390 (N_390,In_993,In_2370);
xnor U391 (N_391,In_1389,In_307);
xor U392 (N_392,In_439,In_188);
xor U393 (N_393,In_894,In_2025);
nand U394 (N_394,In_586,In_1409);
or U395 (N_395,In_427,In_1628);
or U396 (N_396,In_1232,In_756);
nor U397 (N_397,In_478,In_436);
nor U398 (N_398,In_1573,In_733);
and U399 (N_399,In_1550,In_1873);
nand U400 (N_400,In_731,In_1740);
nand U401 (N_401,In_2433,In_1278);
nor U402 (N_402,In_497,In_1942);
nor U403 (N_403,In_668,In_1340);
xor U404 (N_404,In_1432,In_1537);
and U405 (N_405,In_1380,In_23);
and U406 (N_406,In_650,In_2170);
nor U407 (N_407,In_838,In_532);
or U408 (N_408,In_1828,In_1039);
xor U409 (N_409,In_1556,In_1762);
xor U410 (N_410,In_657,In_2077);
xnor U411 (N_411,In_194,In_770);
nand U412 (N_412,In_213,In_1753);
xnor U413 (N_413,In_1872,In_1751);
or U414 (N_414,In_1317,In_1768);
nand U415 (N_415,In_598,In_918);
xor U416 (N_416,In_853,In_2455);
and U417 (N_417,In_633,In_1059);
xnor U418 (N_418,In_1603,In_234);
and U419 (N_419,In_2016,In_424);
xor U420 (N_420,In_2094,In_905);
or U421 (N_421,In_2002,In_451);
nor U422 (N_422,In_2396,In_1555);
or U423 (N_423,In_201,In_572);
nor U424 (N_424,In_651,In_1730);
and U425 (N_425,In_139,In_1160);
nor U426 (N_426,In_1788,In_2173);
and U427 (N_427,In_1329,In_2109);
or U428 (N_428,In_1353,In_324);
nor U429 (N_429,In_1594,In_1608);
xor U430 (N_430,In_104,In_1191);
or U431 (N_431,In_2107,In_1116);
nor U432 (N_432,In_1822,In_2484);
and U433 (N_433,In_1587,In_517);
and U434 (N_434,In_233,In_2459);
xor U435 (N_435,In_1130,In_355);
nand U436 (N_436,In_1973,In_426);
nand U437 (N_437,In_491,In_2228);
nor U438 (N_438,In_1704,In_528);
xor U439 (N_439,In_2215,In_2326);
xnor U440 (N_440,In_2176,In_64);
xor U441 (N_441,In_740,In_742);
nor U442 (N_442,In_2145,In_711);
nor U443 (N_443,In_1316,In_2201);
or U444 (N_444,In_553,In_1980);
nor U445 (N_445,In_2137,In_1384);
or U446 (N_446,In_1538,In_1503);
xnor U447 (N_447,In_1148,In_699);
xnor U448 (N_448,In_1034,In_773);
nand U449 (N_449,In_2155,In_1451);
or U450 (N_450,In_359,In_2206);
or U451 (N_451,In_1022,In_455);
nor U452 (N_452,In_1616,In_1814);
nor U453 (N_453,In_954,In_1064);
and U454 (N_454,In_1181,In_619);
and U455 (N_455,In_924,In_2118);
or U456 (N_456,In_560,In_1387);
xor U457 (N_457,In_2122,In_2255);
or U458 (N_458,In_2050,In_140);
nand U459 (N_459,In_2448,In_967);
nor U460 (N_460,In_2398,In_1437);
nor U461 (N_461,In_1149,In_876);
nor U462 (N_462,In_2458,In_1203);
and U463 (N_463,In_556,In_925);
nor U464 (N_464,In_1127,In_1484);
nor U465 (N_465,In_779,In_782);
xor U466 (N_466,In_153,In_191);
and U467 (N_467,In_1526,In_2187);
and U468 (N_468,In_237,In_710);
or U469 (N_469,In_1300,In_2082);
and U470 (N_470,In_570,In_1601);
nand U471 (N_471,In_369,In_2306);
nand U472 (N_472,In_682,In_210);
xor U473 (N_473,In_882,In_1804);
nor U474 (N_474,In_2473,In_1343);
xnor U475 (N_475,In_6,In_2126);
xnor U476 (N_476,In_608,In_2178);
xor U477 (N_477,In_1607,In_936);
and U478 (N_478,In_1263,In_2275);
or U479 (N_479,In_2006,In_75);
xnor U480 (N_480,In_1632,In_1899);
nand U481 (N_481,In_2093,In_537);
nor U482 (N_482,In_256,In_2252);
and U483 (N_483,In_1483,In_1194);
xor U484 (N_484,In_130,In_2342);
nand U485 (N_485,In_686,In_637);
xor U486 (N_486,In_170,In_901);
and U487 (N_487,In_648,In_1756);
nor U488 (N_488,In_577,In_474);
or U489 (N_489,In_2374,In_79);
nor U490 (N_490,In_1813,In_471);
and U491 (N_491,In_314,In_574);
nand U492 (N_492,In_464,In_1047);
xnor U493 (N_493,In_1274,In_450);
nand U494 (N_494,In_2101,In_2434);
and U495 (N_495,In_143,In_2472);
nand U496 (N_496,In_1551,In_350);
or U497 (N_497,In_1951,In_138);
or U498 (N_498,In_1096,In_484);
nor U499 (N_499,In_289,In_2003);
nor U500 (N_500,In_2447,In_1101);
nor U501 (N_501,In_186,In_1962);
and U502 (N_502,In_645,In_19);
nor U503 (N_503,In_536,In_164);
nor U504 (N_504,In_646,In_946);
nand U505 (N_505,In_1457,In_1854);
and U506 (N_506,In_613,In_917);
or U507 (N_507,In_1404,In_1631);
xnor U508 (N_508,In_1953,In_1678);
or U509 (N_509,In_1797,In_909);
or U510 (N_510,In_1781,In_1038);
xor U511 (N_511,In_1979,In_468);
nor U512 (N_512,In_1764,In_1767);
and U513 (N_513,In_603,In_521);
and U514 (N_514,In_807,In_1272);
xnor U515 (N_515,In_1476,In_2113);
nor U516 (N_516,In_1777,In_2008);
nor U517 (N_517,In_2451,In_914);
nand U518 (N_518,In_69,In_2175);
xor U519 (N_519,In_627,In_1578);
or U520 (N_520,In_1460,In_883);
and U521 (N_521,In_595,In_862);
xor U522 (N_522,In_2440,In_1513);
and U523 (N_523,In_523,In_2246);
and U524 (N_524,In_1911,In_624);
or U525 (N_525,In_11,In_382);
nor U526 (N_526,In_2488,In_320);
xor U527 (N_527,In_912,In_2358);
and U528 (N_528,In_1051,In_163);
nand U529 (N_529,In_1613,In_1650);
xnor U530 (N_530,In_1937,In_405);
xor U531 (N_531,In_398,In_106);
nor U532 (N_532,In_1855,In_538);
xor U533 (N_533,In_1734,In_667);
nand U534 (N_534,In_584,In_1943);
nor U535 (N_535,In_818,In_1605);
nor U536 (N_536,In_1115,In_1159);
nand U537 (N_537,In_895,In_1105);
nor U538 (N_538,In_1963,In_2355);
xnor U539 (N_539,In_1829,In_1809);
or U540 (N_540,In_1644,In_1719);
nand U541 (N_541,In_1068,In_1273);
nand U542 (N_542,In_741,In_980);
nand U543 (N_543,In_2344,In_236);
xnor U544 (N_544,In_89,In_1893);
nor U545 (N_545,In_2383,In_465);
or U546 (N_546,In_240,In_1926);
nand U547 (N_547,In_1961,In_1475);
nor U548 (N_548,In_441,In_103);
xor U549 (N_549,In_2360,In_1435);
and U550 (N_550,In_1626,In_732);
or U551 (N_551,In_318,In_877);
xor U552 (N_552,In_2221,In_2260);
and U553 (N_553,In_1966,In_1796);
nand U554 (N_554,In_366,In_881);
xnor U555 (N_555,In_344,In_1042);
or U556 (N_556,In_126,In_2043);
or U557 (N_557,In_2452,In_110);
xnor U558 (N_558,In_356,In_1489);
and U559 (N_559,In_697,In_128);
xnor U560 (N_560,In_833,In_295);
or U561 (N_561,In_408,In_125);
and U562 (N_562,In_806,In_470);
or U563 (N_563,In_1938,In_1760);
xnor U564 (N_564,In_1361,In_2055);
nor U565 (N_565,In_472,In_1882);
xnor U566 (N_566,In_596,In_440);
nand U567 (N_567,In_1469,In_662);
nor U568 (N_568,In_1946,In_1480);
nor U569 (N_569,In_693,In_502);
or U570 (N_570,In_2453,In_707);
or U571 (N_571,In_251,In_1870);
nor U572 (N_572,In_81,In_377);
nand U573 (N_573,In_1798,In_1898);
nand U574 (N_574,In_2128,In_886);
nor U575 (N_575,In_1609,In_2387);
nand U576 (N_576,In_457,In_2361);
and U577 (N_577,In_2088,In_1761);
and U578 (N_578,In_2403,In_781);
nor U579 (N_579,In_788,In_1486);
and U580 (N_580,In_1895,In_2498);
or U581 (N_581,In_2066,In_2296);
or U582 (N_582,In_505,In_1399);
nor U583 (N_583,In_1391,In_794);
nor U584 (N_584,In_1618,In_820);
nor U585 (N_585,In_2164,In_2244);
xor U586 (N_586,In_2345,In_66);
and U587 (N_587,In_37,In_1844);
nand U588 (N_588,In_1548,In_2412);
nor U589 (N_589,In_1310,In_1280);
or U590 (N_590,In_20,In_2307);
and U591 (N_591,In_1738,In_317);
and U592 (N_592,In_456,In_364);
xor U593 (N_593,In_2309,In_218);
or U594 (N_594,In_420,In_414);
or U595 (N_595,In_1971,In_932);
nor U596 (N_596,In_1841,In_1978);
xor U597 (N_597,In_2150,In_589);
nand U598 (N_598,In_865,In_1928);
nor U599 (N_599,In_496,In_431);
and U600 (N_600,In_2316,In_419);
or U601 (N_601,In_2367,In_2040);
or U602 (N_602,In_2049,In_2062);
nand U603 (N_603,In_1408,In_1856);
nor U604 (N_604,In_1453,In_1769);
nor U605 (N_605,In_910,In_1774);
nand U606 (N_606,In_1622,In_826);
nor U607 (N_607,In_2018,In_903);
xnor U608 (N_608,In_1024,In_611);
nand U609 (N_609,In_1682,In_1348);
xor U610 (N_610,In_1124,In_1242);
nor U611 (N_611,In_1859,In_1886);
nor U612 (N_612,In_1785,In_713);
or U613 (N_613,In_628,In_141);
nor U614 (N_614,In_1914,In_1156);
nor U615 (N_615,In_508,In_262);
nand U616 (N_616,In_2024,In_1497);
nor U617 (N_617,In_268,In_2389);
and U618 (N_618,In_134,In_836);
or U619 (N_619,In_2450,In_292);
and U620 (N_620,In_1755,In_488);
or U621 (N_621,In_798,In_2168);
xnor U622 (N_622,In_606,In_1128);
and U623 (N_623,In_1003,In_737);
and U624 (N_624,In_2443,In_1885);
nand U625 (N_625,In_1266,In_1269);
nor U626 (N_626,In_1465,In_113);
xor U627 (N_627,In_2408,In_2487);
and U628 (N_628,In_391,In_1226);
xor U629 (N_629,In_217,In_1887);
or U630 (N_630,In_1143,In_1225);
nand U631 (N_631,In_828,In_489);
and U632 (N_632,In_2478,In_2253);
and U633 (N_633,In_1027,In_1099);
or U634 (N_634,In_1858,In_1772);
nor U635 (N_635,In_180,In_987);
or U636 (N_636,In_162,In_1655);
xor U637 (N_637,In_2039,In_481);
nand U638 (N_638,In_575,In_793);
xor U639 (N_639,In_642,In_2184);
nand U640 (N_640,In_2314,In_1894);
nor U641 (N_641,In_629,In_558);
and U642 (N_642,In_856,In_1985);
or U643 (N_643,In_2298,In_1665);
nand U644 (N_644,In_1164,In_506);
nand U645 (N_645,In_2143,In_1364);
nor U646 (N_646,In_1901,In_211);
nand U647 (N_647,In_1256,In_1700);
nand U648 (N_648,In_57,In_55);
nand U649 (N_649,In_269,In_1552);
nand U650 (N_650,In_678,In_44);
xnor U651 (N_651,In_232,In_375);
xnor U652 (N_652,In_2017,In_1701);
and U653 (N_653,In_1011,In_288);
and U654 (N_654,In_475,In_690);
nand U655 (N_655,In_622,In_42);
and U656 (N_656,In_1995,In_1431);
xor U657 (N_657,In_1066,In_1984);
or U658 (N_658,In_2014,In_1097);
or U659 (N_659,In_1544,In_2268);
nor U660 (N_660,In_1288,In_1154);
and U661 (N_661,In_283,In_1920);
or U662 (N_662,In_953,In_2449);
xor U663 (N_663,In_1222,In_2199);
nand U664 (N_664,In_1323,In_117);
or U665 (N_665,In_2278,In_907);
and U666 (N_666,In_1747,In_1625);
nand U667 (N_667,In_1493,In_976);
xnor U668 (N_668,In_1983,In_301);
and U669 (N_669,In_142,In_156);
xnor U670 (N_670,In_1703,In_2390);
and U671 (N_671,In_2310,In_2249);
nand U672 (N_672,In_938,In_386);
or U673 (N_673,In_2097,In_305);
nor U674 (N_674,In_966,In_1879);
nor U675 (N_675,In_581,In_1801);
nand U676 (N_676,In_2041,In_1063);
and U677 (N_677,In_2213,In_1940);
nor U678 (N_678,In_1420,In_2000);
or U679 (N_679,In_2405,In_159);
xnor U680 (N_680,In_1745,In_927);
or U681 (N_681,In_263,In_2442);
nand U682 (N_682,In_270,In_1224);
or U683 (N_683,In_388,In_438);
nor U684 (N_684,In_49,In_1715);
xor U685 (N_685,In_1890,In_80);
and U686 (N_686,In_929,In_2245);
nor U687 (N_687,In_1758,In_2106);
and U688 (N_688,In_2083,In_872);
and U689 (N_689,In_1073,In_1583);
and U690 (N_690,In_963,In_1569);
nand U691 (N_691,In_1668,In_1260);
nand U692 (N_692,In_1843,In_1820);
and U693 (N_693,In_1331,In_1060);
xor U694 (N_694,In_1574,In_1180);
or U695 (N_695,In_718,In_1519);
nor U696 (N_696,In_804,In_394);
xnor U697 (N_697,In_197,In_1806);
and U698 (N_698,In_1085,In_916);
nand U699 (N_699,In_1406,In_448);
xnor U700 (N_700,In_1002,In_1427);
nor U701 (N_701,In_939,In_92);
nand U702 (N_702,In_1615,In_1271);
nand U703 (N_703,In_1057,In_808);
xnor U704 (N_704,In_683,In_831);
xnor U705 (N_705,In_1104,In_1754);
and U706 (N_706,In_1231,In_1903);
or U707 (N_707,In_50,In_68);
and U708 (N_708,In_1729,In_13);
or U709 (N_709,In_1352,In_1554);
nand U710 (N_710,In_2323,In_1598);
or U711 (N_711,In_9,In_127);
nor U712 (N_712,In_265,In_1991);
nor U713 (N_713,In_2267,In_566);
xor U714 (N_714,In_617,In_1311);
or U715 (N_715,In_1030,In_1910);
nand U716 (N_716,In_179,In_1264);
or U717 (N_717,In_1074,In_2092);
or U718 (N_718,In_298,In_495);
nand U719 (N_719,In_1994,In_1313);
xnor U720 (N_720,In_1649,In_341);
or U721 (N_721,In_1684,In_1525);
nor U722 (N_722,In_739,In_688);
or U723 (N_723,In_216,In_2099);
nor U724 (N_724,In_880,In_1520);
nand U725 (N_725,In_1189,In_2349);
nor U726 (N_726,In_1658,In_410);
xor U727 (N_727,In_1742,In_2229);
nor U728 (N_728,In_196,In_444);
xnor U729 (N_729,In_59,In_1591);
nor U730 (N_730,In_136,In_1697);
nand U731 (N_731,In_1790,In_2242);
and U732 (N_732,In_189,In_2265);
xor U733 (N_733,In_1414,In_2424);
nand U734 (N_734,In_1173,In_900);
and U735 (N_735,In_65,In_2357);
nor U736 (N_736,In_2191,In_534);
or U737 (N_737,In_1183,In_459);
and U738 (N_738,In_1069,In_825);
nor U739 (N_739,In_100,In_527);
nand U740 (N_740,In_1712,In_2339);
nor U741 (N_741,In_1982,In_616);
nor U742 (N_742,In_2404,In_1576);
or U743 (N_743,In_1383,In_1986);
or U744 (N_744,In_275,In_332);
and U745 (N_745,In_2421,In_2372);
nor U746 (N_746,In_1690,In_869);
nor U747 (N_747,In_385,In_663);
xnor U748 (N_748,In_1743,In_2139);
or U749 (N_749,In_1279,In_2430);
nor U750 (N_750,In_15,In_1948);
or U751 (N_751,In_2153,In_1284);
and U752 (N_752,In_2289,In_620);
xor U753 (N_753,In_591,In_1119);
and U754 (N_754,In_1722,In_249);
xor U755 (N_755,In_1006,In_1045);
and U756 (N_756,In_2371,In_1342);
or U757 (N_757,In_1562,In_1094);
or U758 (N_758,In_2300,In_300);
nor U759 (N_759,In_476,In_960);
nand U760 (N_760,In_2324,In_2151);
or U761 (N_761,In_1411,In_2028);
nand U762 (N_762,In_652,In_2223);
nand U763 (N_763,In_168,In_2063);
or U764 (N_764,In_1291,In_1842);
nand U765 (N_765,In_112,In_1892);
and U766 (N_766,In_1783,In_1749);
and U767 (N_767,In_2132,In_2281);
nor U768 (N_768,In_1681,In_1254);
nor U769 (N_769,In_1344,In_601);
nor U770 (N_770,In_1653,In_2036);
or U771 (N_771,In_2254,In_1819);
xnor U772 (N_772,In_4,In_1691);
xnor U773 (N_773,In_2079,In_568);
or U774 (N_774,In_1998,In_768);
nand U775 (N_775,In_571,In_544);
nand U776 (N_776,In_1318,In_115);
and U777 (N_777,In_415,In_2218);
and U778 (N_778,In_2328,In_1696);
nor U779 (N_779,In_192,In_923);
or U780 (N_780,In_2282,In_520);
xnor U781 (N_781,In_1741,In_254);
xor U782 (N_782,In_1614,In_368);
nor U783 (N_783,In_8,In_467);
or U784 (N_784,In_1918,In_1337);
or U785 (N_785,In_2116,In_1210);
nand U786 (N_786,In_1087,In_1023);
nand U787 (N_787,In_279,In_41);
and U788 (N_788,In_526,In_644);
xnor U789 (N_789,In_771,In_2460);
nand U790 (N_790,In_952,In_1386);
or U791 (N_791,In_487,In_1839);
nor U792 (N_792,In_2373,In_1135);
nand U793 (N_793,In_2381,In_636);
or U794 (N_794,In_46,In_347);
and U795 (N_795,In_1102,In_1939);
nor U796 (N_796,In_786,In_2069);
and U797 (N_797,In_3,In_1602);
xor U798 (N_798,In_634,In_729);
xor U799 (N_799,In_2204,In_2131);
or U800 (N_800,In_2463,In_255);
nand U801 (N_801,In_1299,In_973);
or U802 (N_802,In_2322,In_1502);
and U803 (N_803,In_769,In_302);
or U804 (N_804,In_1871,In_580);
and U805 (N_805,In_1123,In_1670);
nor U806 (N_806,In_784,In_1960);
nor U807 (N_807,In_403,In_1737);
nor U808 (N_808,In_1709,In_2080);
nor U809 (N_809,In_1641,In_1952);
and U810 (N_810,In_2384,In_2032);
nand U811 (N_811,In_2188,In_2465);
and U812 (N_812,In_221,In_706);
and U813 (N_813,In_1113,In_1239);
and U814 (N_814,In_107,In_999);
and U815 (N_815,In_1320,In_1445);
and U816 (N_816,In_548,In_1357);
and U817 (N_817,In_778,In_172);
or U818 (N_818,In_933,In_2212);
or U819 (N_819,In_2343,In_1360);
nor U820 (N_820,In_0,In_1950);
and U821 (N_821,In_1247,In_1205);
xor U822 (N_822,In_816,In_1534);
or U823 (N_823,In_1142,In_594);
or U824 (N_824,In_2119,In_434);
xor U825 (N_825,In_1470,In_63);
and U826 (N_826,In_915,In_2301);
nor U827 (N_827,In_748,In_1792);
nand U828 (N_828,In_930,In_1147);
and U829 (N_829,In_54,In_1512);
nand U830 (N_830,In_2352,In_2125);
and U831 (N_831,In_454,In_2194);
or U832 (N_832,In_805,In_1708);
nand U833 (N_833,In_1455,In_149);
and U834 (N_834,In_212,In_2295);
nand U835 (N_835,In_1446,In_515);
or U836 (N_836,In_373,In_1328);
xor U837 (N_837,In_22,In_2417);
xnor U838 (N_838,In_2141,In_315);
xnor U839 (N_839,In_531,In_483);
nor U840 (N_840,In_1312,In_241);
nand U841 (N_841,In_1786,In_1474);
or U842 (N_842,In_1236,In_2076);
nor U843 (N_843,In_2196,In_948);
nor U844 (N_844,In_1541,In_2112);
or U845 (N_845,In_2046,In_1955);
nor U846 (N_846,In_2129,In_404);
xnor U847 (N_847,In_1802,In_671);
xnor U848 (N_848,In_2136,In_1586);
nor U849 (N_849,In_2086,In_701);
or U850 (N_850,In_942,In_546);
nor U851 (N_851,In_406,In_1449);
and U852 (N_852,In_2318,In_1964);
nand U853 (N_853,In_88,In_795);
nand U854 (N_854,In_2285,In_1634);
xnor U855 (N_855,In_2237,In_1091);
or U856 (N_856,In_1186,In_649);
nor U857 (N_857,In_660,In_267);
xor U858 (N_858,In_1390,In_1876);
nor U859 (N_859,In_529,In_2203);
xor U860 (N_860,In_2477,In_1155);
xor U861 (N_861,In_207,In_361);
xnor U862 (N_862,In_2123,In_2256);
nand U863 (N_863,In_323,In_689);
and U864 (N_864,In_1109,In_681);
or U865 (N_865,In_1419,In_93);
and U866 (N_866,In_2161,In_1172);
xor U867 (N_867,In_1989,In_2105);
nand U868 (N_868,In_1698,In_1501);
and U869 (N_869,In_2091,In_1464);
xor U870 (N_870,In_674,In_2022);
nor U871 (N_871,In_1812,In_1904);
nand U872 (N_872,In_1705,In_1635);
xor U873 (N_873,In_1176,In_2146);
xor U874 (N_874,In_1370,In_1345);
or U875 (N_875,In_244,In_1372);
xnor U876 (N_876,In_1529,In_1098);
or U877 (N_877,In_638,In_1228);
xor U878 (N_878,In_1084,In_1286);
nand U879 (N_879,In_2432,In_1834);
and U880 (N_880,In_691,In_271);
nand U881 (N_881,In_1746,In_1958);
nand U882 (N_882,In_184,In_2013);
xnor U883 (N_883,In_2495,In_992);
nand U884 (N_884,In_1093,In_994);
and U885 (N_885,In_97,In_995);
or U886 (N_886,In_949,In_98);
nor U887 (N_887,In_1794,In_413);
and U888 (N_888,In_247,In_2388);
nand U889 (N_889,In_1468,In_1351);
and U890 (N_890,In_849,In_728);
nor U891 (N_891,In_2494,In_1070);
nand U892 (N_892,In_982,In_1150);
and U893 (N_893,In_1825,In_750);
and U894 (N_894,In_1424,In_920);
nand U895 (N_895,In_1661,In_337);
xnor U896 (N_896,In_1897,In_1161);
nor U897 (N_897,In_1528,In_1954);
and U898 (N_898,In_1581,In_446);
nand U899 (N_899,In_761,In_1739);
nand U900 (N_900,In_1849,In_2456);
xnor U901 (N_901,In_839,In_530);
nor U902 (N_902,In_1993,In_1545);
nand U903 (N_903,In_565,In_696);
xnor U904 (N_904,In_1770,In_792);
and U905 (N_905,In_1211,In_1477);
nand U906 (N_906,In_187,In_1866);
nand U907 (N_907,In_1686,In_492);
xnor U908 (N_908,In_2407,In_114);
nand U909 (N_909,In_765,In_1584);
nand U910 (N_910,In_1648,In_1138);
xnor U911 (N_911,In_60,In_72);
nand U912 (N_912,In_2231,In_1251);
xor U913 (N_913,In_1315,In_1335);
nor U914 (N_914,In_996,In_1245);
and U915 (N_915,In_906,In_1915);
nand U916 (N_916,In_1530,In_2413);
nor U917 (N_917,In_2219,In_1646);
or U918 (N_918,In_2051,In_294);
and U919 (N_919,In_947,In_2011);
nand U920 (N_920,In_131,In_934);
nand U921 (N_921,In_1214,In_592);
nand U922 (N_922,In_53,In_898);
nand U923 (N_923,In_1765,In_2476);
and U924 (N_924,In_2386,In_273);
xor U925 (N_925,In_1518,In_199);
nand U926 (N_926,In_308,In_1559);
xnor U927 (N_927,In_1913,In_625);
or U928 (N_928,In_518,In_2331);
nor U929 (N_929,In_2279,In_752);
nor U930 (N_930,In_1354,In_1246);
xor U931 (N_931,In_1784,In_325);
xor U932 (N_932,In_286,In_1100);
nor U933 (N_933,In_2009,In_2335);
or U934 (N_934,In_1416,In_676);
xnor U935 (N_935,In_1878,In_1394);
nor U936 (N_936,In_2189,In_2029);
nand U937 (N_937,In_926,In_2121);
nor U938 (N_938,In_27,In_1133);
nor U939 (N_939,In_709,In_1367);
xor U940 (N_940,In_2336,In_503);
nand U941 (N_941,In_802,In_1379);
nor U942 (N_942,In_1869,In_940);
xor U943 (N_943,In_1575,In_1883);
and U944 (N_944,In_2457,In_1444);
nand U945 (N_945,In_873,In_1977);
xnor U946 (N_946,In_812,In_2205);
nand U947 (N_947,In_695,In_133);
and U948 (N_948,In_2232,In_1275);
xnor U949 (N_949,In_280,In_1479);
xnor U950 (N_950,In_2054,In_1732);
xor U951 (N_951,In_2391,In_245);
or U952 (N_952,In_86,In_1086);
nand U953 (N_953,In_2369,In_1302);
and U954 (N_954,In_1604,In_1145);
xor U955 (N_955,In_2133,In_1750);
and U956 (N_956,In_2234,In_1217);
and U957 (N_957,In_2269,In_2399);
or U958 (N_958,In_151,In_1144);
nor U959 (N_959,In_230,In_1923);
nor U960 (N_960,In_1481,In_2160);
xor U961 (N_961,In_937,In_1589);
and U962 (N_962,In_1845,In_1846);
nand U963 (N_963,In_357,In_205);
nand U964 (N_964,In_1195,In_972);
xnor U965 (N_965,In_1117,In_198);
and U966 (N_966,In_1031,In_1071);
or U967 (N_967,In_2182,In_1687);
xor U968 (N_968,In_1823,In_1388);
nor U969 (N_969,In_1723,In_1257);
nor U970 (N_970,In_178,In_1490);
and U971 (N_971,In_897,In_258);
and U972 (N_972,In_71,In_1909);
or U973 (N_973,In_1322,In_2098);
and U974 (N_974,In_1496,In_1600);
nand U975 (N_975,In_1088,In_1908);
nor U976 (N_976,In_2409,In_559);
nand U977 (N_977,In_2090,In_1624);
nor U978 (N_978,In_2238,In_1531);
nor U979 (N_979,In_1522,In_2270);
and U980 (N_980,In_1523,In_461);
or U981 (N_981,In_685,In_458);
nand U982 (N_982,In_1126,In_1929);
and U983 (N_983,In_2283,In_1141);
or U984 (N_984,In_499,In_1407);
nor U985 (N_985,In_2337,In_1415);
nand U986 (N_986,In_1547,In_26);
or U987 (N_987,In_827,In_1674);
or U988 (N_988,In_2401,In_297);
nand U989 (N_989,In_1290,In_1307);
and U990 (N_990,In_1151,In_1363);
nand U991 (N_991,In_2406,In_2195);
xnor U992 (N_992,In_219,In_2431);
xor U993 (N_993,In_858,In_2226);
or U994 (N_994,In_1868,In_600);
nand U995 (N_995,In_1234,In_2486);
and U996 (N_996,In_58,In_1268);
xnor U997 (N_997,In_1129,In_746);
nor U998 (N_998,In_2048,In_1466);
xnor U999 (N_999,In_1571,In_334);
or U1000 (N_1000,In_698,In_511);
or U1001 (N_1001,In_1488,In_2497);
or U1002 (N_1002,In_842,In_425);
or U1003 (N_1003,In_1459,In_2287);
xnor U1004 (N_1004,In_70,In_851);
or U1005 (N_1005,In_1927,In_834);
nand U1006 (N_1006,In_102,In_2152);
or U1007 (N_1007,In_783,In_1293);
and U1008 (N_1008,In_726,In_284);
xor U1009 (N_1009,In_1933,In_1471);
xnor U1010 (N_1010,In_2264,In_2376);
nand U1011 (N_1011,In_1527,In_2180);
and U1012 (N_1012,In_303,In_1949);
nand U1013 (N_1013,In_810,In_177);
or U1014 (N_1014,In_1669,In_1429);
nor U1015 (N_1015,In_705,In_228);
nor U1016 (N_1016,In_1347,In_1301);
xor U1017 (N_1017,In_2479,In_1285);
and U1018 (N_1018,In_1511,In_1157);
xnor U1019 (N_1019,In_452,In_1405);
nor U1020 (N_1020,In_7,In_1078);
and U1021 (N_1021,In_669,In_1936);
xor U1022 (N_1022,In_965,In_550);
nor U1023 (N_1023,In_1240,In_1029);
nand U1024 (N_1024,In_1924,In_2263);
or U1025 (N_1025,In_181,In_2305);
or U1026 (N_1026,In_1659,In_971);
nand U1027 (N_1027,In_339,In_1956);
nor U1028 (N_1028,In_1401,In_2068);
nor U1029 (N_1029,In_277,In_1981);
and U1030 (N_1030,In_2438,In_777);
xnor U1031 (N_1031,In_988,In_776);
and U1032 (N_1032,In_193,In_1612);
or U1033 (N_1033,In_785,In_1350);
nor U1034 (N_1034,In_1410,In_261);
and U1035 (N_1035,In_2299,In_1033);
nand U1036 (N_1036,In_2064,In_2319);
or U1037 (N_1037,In_90,In_202);
nor U1038 (N_1038,In_260,In_1080);
xnor U1039 (N_1039,In_2262,In_2351);
nand U1040 (N_1040,In_165,In_430);
and U1041 (N_1041,In_525,In_2382);
and U1042 (N_1042,In_1237,In_968);
nor U1043 (N_1043,In_552,In_1906);
and U1044 (N_1044,In_961,In_2035);
nand U1045 (N_1045,In_1808,In_1472);
nor U1046 (N_1046,In_724,In_1206);
and U1047 (N_1047,In_311,In_1717);
xnor U1048 (N_1048,In_1662,In_2224);
nand U1049 (N_1049,In_479,In_879);
xnor U1050 (N_1050,In_1397,In_428);
and U1051 (N_1051,In_715,In_604);
or U1052 (N_1052,In_958,In_1863);
or U1053 (N_1053,In_1787,In_183);
xnor U1054 (N_1054,In_2313,In_2144);
xor U1055 (N_1055,In_998,In_99);
xor U1056 (N_1056,In_1560,In_2065);
xnor U1057 (N_1057,In_755,In_407);
or U1058 (N_1058,In_336,In_1381);
or U1059 (N_1059,In_1997,In_1815);
or U1060 (N_1060,In_173,In_745);
and U1061 (N_1061,In_1620,In_884);
or U1062 (N_1062,In_1167,In_1184);
or U1063 (N_1063,In_2499,In_1131);
nor U1064 (N_1064,In_338,In_2071);
or U1065 (N_1065,In_1789,In_519);
or U1066 (N_1066,In_631,In_730);
nor U1067 (N_1067,In_442,In_969);
and U1068 (N_1068,In_399,In_345);
nand U1069 (N_1069,In_1319,In_815);
nand U1070 (N_1070,In_1967,In_1017);
xnor U1071 (N_1071,In_229,In_955);
xor U1072 (N_1072,In_841,In_2072);
nor U1073 (N_1073,In_380,In_1165);
or U1074 (N_1074,In_1303,In_1630);
nand U1075 (N_1075,In_919,In_621);
or U1076 (N_1076,In_2104,In_1504);
xor U1077 (N_1077,In_1219,In_1968);
and U1078 (N_1078,In_1590,In_2444);
xnor U1079 (N_1079,In_1400,In_1853);
or U1080 (N_1080,In_702,In_811);
nor U1081 (N_1081,In_1972,In_1198);
nor U1082 (N_1082,In_684,In_2496);
and U1083 (N_1083,In_1919,In_1830);
nand U1084 (N_1084,In_1827,In_2207);
or U1085 (N_1085,In_1439,In_1771);
nor U1086 (N_1086,In_374,In_1107);
nor U1087 (N_1087,In_1079,In_1014);
nand U1088 (N_1088,In_167,In_643);
nor U1089 (N_1089,In_863,In_2058);
and U1090 (N_1090,In_1152,In_2042);
or U1091 (N_1091,In_1889,In_155);
nor U1092 (N_1092,In_1838,In_449);
nor U1093 (N_1093,In_309,In_1514);
and U1094 (N_1094,In_2084,In_2247);
xor U1095 (N_1095,In_1112,In_1174);
xor U1096 (N_1096,In_1947,In_1298);
and U1097 (N_1097,In_2273,In_1178);
nor U1098 (N_1098,In_1557,In_2233);
nand U1099 (N_1099,In_2251,In_635);
xnor U1100 (N_1100,In_1259,In_1169);
nor U1101 (N_1101,In_549,In_935);
or U1102 (N_1102,In_2020,In_1532);
xnor U1103 (N_1103,In_2348,In_24);
xor U1104 (N_1104,In_1103,In_1395);
nand U1105 (N_1105,In_1175,In_977);
and U1106 (N_1106,In_889,In_945);
nand U1107 (N_1107,In_1865,In_899);
or U1108 (N_1108,In_1791,In_2356);
or U1109 (N_1109,In_2393,In_1054);
nand U1110 (N_1110,In_1542,In_2258);
nor U1111 (N_1111,In_1640,In_569);
or U1112 (N_1112,In_504,In_2416);
or U1113 (N_1113,In_1565,In_1642);
or U1114 (N_1114,In_1197,In_2359);
nor U1115 (N_1115,In_1473,In_590);
nor U1116 (N_1116,In_1229,In_878);
xor U1117 (N_1117,In_10,In_35);
and U1118 (N_1118,In_1067,In_1338);
or U1119 (N_1119,In_2435,In_1726);
or U1120 (N_1120,In_2426,In_1851);
xor U1121 (N_1121,In_2033,In_2302);
nand U1122 (N_1122,In_1773,In_2312);
xnor U1123 (N_1123,In_2394,In_1276);
xnor U1124 (N_1124,In_1905,In_1826);
and U1125 (N_1125,In_252,In_2427);
nand U1126 (N_1126,In_896,In_76);
nand U1127 (N_1127,In_2293,In_1314);
or U1128 (N_1128,In_1570,In_1718);
xor U1129 (N_1129,In_2147,In_390);
xor U1130 (N_1130,In_981,In_736);
xor U1131 (N_1131,In_466,In_371);
xnor U1132 (N_1132,In_2026,In_2304);
nand U1133 (N_1133,In_2375,In_137);
nand U1134 (N_1134,In_346,In_1422);
xnor U1135 (N_1135,In_2493,In_2462);
xnor U1136 (N_1136,In_2341,In_328);
nand U1137 (N_1137,In_2070,In_2052);
nor U1138 (N_1138,In_208,In_2200);
or U1139 (N_1139,In_659,In_1517);
or U1140 (N_1140,In_951,In_2019);
xnor U1141 (N_1141,In_1083,In_1636);
nand U1142 (N_1142,In_2423,In_365);
and U1143 (N_1143,In_2138,In_1442);
nor U1144 (N_1144,In_231,In_2130);
nand U1145 (N_1145,In_704,In_43);
nor U1146 (N_1146,In_1021,In_1847);
xor U1147 (N_1147,In_2120,In_1349);
nand U1148 (N_1148,In_1037,In_887);
nor U1149 (N_1149,In_401,In_1543);
xor U1150 (N_1150,In_282,In_417);
nor U1151 (N_1151,In_123,In_379);
nand U1152 (N_1152,In_1689,In_1336);
or U1153 (N_1153,In_1058,In_2437);
nor U1154 (N_1154,In_1563,In_1009);
xor U1155 (N_1155,In_493,In_1793);
or U1156 (N_1156,In_1912,In_2087);
or U1157 (N_1157,In_51,In_1974);
nand U1158 (N_1158,In_1999,In_353);
and U1159 (N_1159,In_1568,In_2482);
nor U1160 (N_1160,In_857,In_462);
or U1161 (N_1161,In_2454,In_997);
nor U1162 (N_1162,In_1763,In_396);
or U1163 (N_1163,In_1533,In_84);
or U1164 (N_1164,In_855,In_132);
xor U1165 (N_1165,In_1443,In_1881);
nor U1166 (N_1166,In_222,In_823);
xnor U1167 (N_1167,In_2490,In_1807);
xnor U1168 (N_1168,In_514,In_367);
xnor U1169 (N_1169,In_67,In_1724);
nor U1170 (N_1170,In_2366,In_1327);
nand U1171 (N_1171,In_554,In_1965);
and U1172 (N_1172,In_2471,In_1860);
nor U1173 (N_1173,In_171,In_959);
xor U1174 (N_1174,In_1212,In_2439);
and U1175 (N_1175,In_1359,In_2114);
or U1176 (N_1176,In_1623,In_175);
and U1177 (N_1177,In_1438,In_735);
xnor U1178 (N_1178,In_166,In_618);
nand U1179 (N_1179,In_817,In_1848);
xor U1180 (N_1180,In_352,In_25);
nand U1181 (N_1181,In_1215,In_2045);
nor U1182 (N_1182,In_376,In_1716);
xor U1183 (N_1183,In_85,In_1637);
xor U1184 (N_1184,In_848,In_358);
or U1185 (N_1185,In_469,In_1050);
xnor U1186 (N_1186,In_672,In_1398);
nor U1187 (N_1187,In_522,In_719);
and U1188 (N_1188,In_2425,In_1654);
nor U1189 (N_1189,In_2124,In_679);
nand U1190 (N_1190,In_2198,In_1358);
or U1191 (N_1191,In_564,In_763);
xor U1192 (N_1192,In_1524,In_326);
and U1193 (N_1193,In_2365,In_2474);
nand U1194 (N_1194,In_908,In_453);
and U1195 (N_1195,In_1433,In_582);
nor U1196 (N_1196,In_870,In_160);
nand U1197 (N_1197,In_1706,In_513);
nor U1198 (N_1198,In_1811,In_1402);
nor U1199 (N_1199,In_1090,In_1250);
nor U1200 (N_1200,In_720,In_2);
nand U1201 (N_1201,In_2171,In_2236);
nand U1202 (N_1202,In_1120,In_1880);
nor U1203 (N_1203,In_5,In_1540);
nand U1204 (N_1204,In_1728,In_837);
and U1205 (N_1205,In_372,In_370);
nand U1206 (N_1206,In_1025,In_700);
or U1207 (N_1207,In_799,In_2317);
or U1208 (N_1208,In_1857,In_738);
nor U1209 (N_1209,In_1535,In_588);
nand U1210 (N_1210,In_1041,In_1005);
and U1211 (N_1211,In_501,In_1959);
nor U1212 (N_1212,In_1539,In_2103);
nor U1213 (N_1213,In_2422,In_2272);
xnor U1214 (N_1214,In_1325,In_1667);
xnor U1215 (N_1215,In_135,In_902);
xnor U1216 (N_1216,In_1561,In_109);
xnor U1217 (N_1217,In_1185,In_890);
xor U1218 (N_1218,In_1907,In_1891);
nand U1219 (N_1219,In_819,In_563);
nand U1220 (N_1220,In_843,In_1177);
nand U1221 (N_1221,In_274,In_1536);
xnor U1222 (N_1222,In_654,In_1162);
or U1223 (N_1223,In_1281,In_2392);
and U1224 (N_1224,In_970,In_239);
nor U1225 (N_1225,In_1441,In_1188);
or U1226 (N_1226,In_1779,In_1896);
and U1227 (N_1227,In_1672,In_1888);
nand U1228 (N_1228,In_1434,In_2047);
xor U1229 (N_1229,In_2167,In_227);
and U1230 (N_1230,In_402,In_1171);
or U1231 (N_1231,In_2362,In_1508);
xnor U1232 (N_1232,In_118,In_1110);
nand U1233 (N_1233,In_432,In_480);
xor U1234 (N_1234,In_2210,In_2010);
nand U1235 (N_1235,In_146,In_1638);
nor U1236 (N_1236,In_1052,In_1292);
and U1237 (N_1237,In_1241,In_1304);
or U1238 (N_1238,In_1253,In_975);
nand U1239 (N_1239,In_2100,In_486);
xor U1240 (N_1240,In_1193,In_2257);
xnor U1241 (N_1241,In_34,In_1196);
xor U1242 (N_1242,In_1065,In_1645);
nor U1243 (N_1243,In_1558,In_2311);
xnor U1244 (N_1244,In_1170,In_1810);
nor U1245 (N_1245,In_844,In_293);
and U1246 (N_1246,In_703,In_516);
xor U1247 (N_1247,In_957,In_2286);
xnor U1248 (N_1248,In_1412,In_33);
xor U1249 (N_1249,In_1306,In_1055);
nor U1250 (N_1250,N_281,N_1026);
or U1251 (N_1251,N_352,N_1178);
nor U1252 (N_1252,N_99,N_930);
xor U1253 (N_1253,N_378,N_934);
nor U1254 (N_1254,N_231,N_827);
nand U1255 (N_1255,N_936,N_731);
nand U1256 (N_1256,N_479,N_1069);
nand U1257 (N_1257,N_496,N_311);
nand U1258 (N_1258,N_996,N_928);
nand U1259 (N_1259,N_22,N_236);
and U1260 (N_1260,N_1226,N_192);
nand U1261 (N_1261,N_332,N_675);
nand U1262 (N_1262,N_611,N_112);
nand U1263 (N_1263,N_1154,N_1074);
nand U1264 (N_1264,N_620,N_596);
xor U1265 (N_1265,N_1221,N_128);
or U1266 (N_1266,N_599,N_14);
nor U1267 (N_1267,N_328,N_1138);
or U1268 (N_1268,N_960,N_243);
or U1269 (N_1269,N_628,N_641);
or U1270 (N_1270,N_768,N_673);
and U1271 (N_1271,N_935,N_1222);
or U1272 (N_1272,N_652,N_105);
nor U1273 (N_1273,N_143,N_882);
xnor U1274 (N_1274,N_849,N_10);
nand U1275 (N_1275,N_726,N_1088);
and U1276 (N_1276,N_371,N_1077);
and U1277 (N_1277,N_485,N_300);
nand U1278 (N_1278,N_1140,N_737);
xor U1279 (N_1279,N_877,N_924);
or U1280 (N_1280,N_216,N_981);
or U1281 (N_1281,N_843,N_563);
xor U1282 (N_1282,N_211,N_1212);
or U1283 (N_1283,N_1202,N_585);
nand U1284 (N_1284,N_627,N_537);
xor U1285 (N_1285,N_402,N_1240);
and U1286 (N_1286,N_473,N_672);
nand U1287 (N_1287,N_983,N_1177);
or U1288 (N_1288,N_535,N_248);
and U1289 (N_1289,N_1115,N_478);
nor U1290 (N_1290,N_511,N_490);
or U1291 (N_1291,N_1169,N_1080);
and U1292 (N_1292,N_1249,N_270);
xnor U1293 (N_1293,N_529,N_578);
or U1294 (N_1294,N_1033,N_839);
and U1295 (N_1295,N_125,N_891);
nand U1296 (N_1296,N_422,N_580);
xor U1297 (N_1297,N_342,N_476);
or U1298 (N_1298,N_742,N_439);
xor U1299 (N_1299,N_669,N_845);
or U1300 (N_1300,N_517,N_622);
xor U1301 (N_1301,N_897,N_165);
xnor U1302 (N_1302,N_259,N_213);
or U1303 (N_1303,N_1204,N_1158);
nand U1304 (N_1304,N_944,N_539);
or U1305 (N_1305,N_296,N_867);
xor U1306 (N_1306,N_114,N_179);
xnor U1307 (N_1307,N_483,N_974);
and U1308 (N_1308,N_133,N_127);
or U1309 (N_1309,N_832,N_102);
nor U1310 (N_1310,N_288,N_607);
xnor U1311 (N_1311,N_925,N_844);
and U1312 (N_1312,N_985,N_526);
xor U1313 (N_1313,N_634,N_180);
xor U1314 (N_1314,N_1165,N_235);
nor U1315 (N_1315,N_234,N_427);
or U1316 (N_1316,N_1164,N_1246);
xnor U1317 (N_1317,N_25,N_84);
and U1318 (N_1318,N_804,N_467);
xnor U1319 (N_1319,N_140,N_168);
or U1320 (N_1320,N_501,N_584);
nand U1321 (N_1321,N_681,N_724);
and U1322 (N_1322,N_376,N_282);
nand U1323 (N_1323,N_818,N_347);
nand U1324 (N_1324,N_5,N_258);
and U1325 (N_1325,N_540,N_75);
nand U1326 (N_1326,N_838,N_462);
or U1327 (N_1327,N_1139,N_315);
nor U1328 (N_1328,N_70,N_1061);
xnor U1329 (N_1329,N_209,N_290);
and U1330 (N_1330,N_624,N_561);
and U1331 (N_1331,N_1027,N_1228);
xnor U1332 (N_1332,N_448,N_821);
or U1333 (N_1333,N_664,N_772);
or U1334 (N_1334,N_1189,N_423);
nor U1335 (N_1335,N_1067,N_257);
and U1336 (N_1336,N_39,N_692);
nor U1337 (N_1337,N_629,N_1034);
nand U1338 (N_1338,N_174,N_824);
xor U1339 (N_1339,N_1052,N_156);
nor U1340 (N_1340,N_227,N_811);
nand U1341 (N_1341,N_878,N_1076);
xnor U1342 (N_1342,N_906,N_791);
nor U1343 (N_1343,N_1110,N_119);
and U1344 (N_1344,N_876,N_788);
and U1345 (N_1345,N_339,N_565);
and U1346 (N_1346,N_558,N_157);
or U1347 (N_1347,N_765,N_287);
xnor U1348 (N_1348,N_326,N_1116);
and U1349 (N_1349,N_727,N_244);
nor U1350 (N_1350,N_68,N_569);
nor U1351 (N_1351,N_1196,N_103);
or U1352 (N_1352,N_90,N_458);
xor U1353 (N_1353,N_106,N_266);
nor U1354 (N_1354,N_1145,N_1043);
xnor U1355 (N_1355,N_813,N_1144);
and U1356 (N_1356,N_530,N_677);
nor U1357 (N_1357,N_1185,N_1100);
nor U1358 (N_1358,N_639,N_405);
and U1359 (N_1359,N_815,N_1120);
or U1360 (N_1360,N_0,N_587);
nor U1361 (N_1361,N_253,N_1133);
nor U1362 (N_1362,N_836,N_1223);
xor U1363 (N_1363,N_592,N_626);
and U1364 (N_1364,N_531,N_278);
and U1365 (N_1365,N_226,N_637);
and U1366 (N_1366,N_1233,N_250);
xnor U1367 (N_1367,N_916,N_754);
nor U1368 (N_1368,N_481,N_447);
nand U1369 (N_1369,N_1095,N_1159);
or U1370 (N_1370,N_294,N_1029);
or U1371 (N_1371,N_256,N_993);
or U1372 (N_1372,N_881,N_1130);
nor U1373 (N_1373,N_873,N_575);
or U1374 (N_1374,N_514,N_407);
nand U1375 (N_1375,N_397,N_745);
and U1376 (N_1376,N_358,N_1168);
and U1377 (N_1377,N_861,N_953);
or U1378 (N_1378,N_733,N_1079);
and U1379 (N_1379,N_619,N_577);
xor U1380 (N_1380,N_1219,N_702);
nand U1381 (N_1381,N_606,N_360);
and U1382 (N_1382,N_1224,N_848);
xnor U1383 (N_1383,N_500,N_96);
nand U1384 (N_1384,N_45,N_1241);
nand U1385 (N_1385,N_908,N_145);
nand U1386 (N_1386,N_572,N_970);
and U1387 (N_1387,N_412,N_30);
or U1388 (N_1388,N_203,N_1227);
xnor U1389 (N_1389,N_710,N_375);
and U1390 (N_1390,N_803,N_703);
nand U1391 (N_1391,N_4,N_670);
xnor U1392 (N_1392,N_783,N_55);
and U1393 (N_1393,N_954,N_76);
nand U1394 (N_1394,N_206,N_609);
and U1395 (N_1395,N_828,N_428);
nand U1396 (N_1396,N_313,N_1111);
nand U1397 (N_1397,N_1010,N_1048);
or U1398 (N_1398,N_732,N_15);
and U1399 (N_1399,N_905,N_225);
nor U1400 (N_1400,N_1191,N_969);
nor U1401 (N_1401,N_217,N_420);
xor U1402 (N_1402,N_108,N_190);
xor U1403 (N_1403,N_210,N_303);
nor U1404 (N_1404,N_777,N_1109);
nor U1405 (N_1405,N_1096,N_495);
xnor U1406 (N_1406,N_755,N_921);
and U1407 (N_1407,N_666,N_453);
nand U1408 (N_1408,N_207,N_1137);
xor U1409 (N_1409,N_1086,N_834);
and U1410 (N_1410,N_1049,N_349);
xor U1411 (N_1411,N_1143,N_605);
nor U1412 (N_1412,N_1024,N_498);
xor U1413 (N_1413,N_194,N_1036);
xor U1414 (N_1414,N_997,N_991);
and U1415 (N_1415,N_130,N_459);
xor U1416 (N_1416,N_7,N_736);
nand U1417 (N_1417,N_568,N_382);
nand U1418 (N_1418,N_551,N_268);
nand U1419 (N_1419,N_220,N_1215);
and U1420 (N_1420,N_1,N_868);
nand U1421 (N_1421,N_1066,N_571);
nand U1422 (N_1422,N_950,N_1012);
nand U1423 (N_1423,N_1247,N_1009);
and U1424 (N_1424,N_150,N_390);
and U1425 (N_1425,N_379,N_766);
nand U1426 (N_1426,N_1211,N_446);
nor U1427 (N_1427,N_917,N_385);
nor U1428 (N_1428,N_651,N_532);
or U1429 (N_1429,N_264,N_931);
nand U1430 (N_1430,N_17,N_716);
or U1431 (N_1431,N_602,N_434);
and U1432 (N_1432,N_583,N_761);
and U1433 (N_1433,N_926,N_154);
and U1434 (N_1434,N_380,N_682);
nand U1435 (N_1435,N_262,N_136);
and U1436 (N_1436,N_645,N_680);
xnor U1437 (N_1437,N_1016,N_1184);
nor U1438 (N_1438,N_764,N_322);
nand U1439 (N_1439,N_416,N_355);
nor U1440 (N_1440,N_335,N_919);
or U1441 (N_1441,N_904,N_798);
or U1442 (N_1442,N_576,N_690);
or U1443 (N_1443,N_151,N_171);
xnor U1444 (N_1444,N_1148,N_888);
or U1445 (N_1445,N_107,N_920);
nand U1446 (N_1446,N_437,N_31);
or U1447 (N_1447,N_756,N_77);
nor U1448 (N_1448,N_384,N_212);
nand U1449 (N_1449,N_292,N_1243);
or U1450 (N_1450,N_1070,N_787);
and U1451 (N_1451,N_635,N_1023);
nor U1452 (N_1452,N_1045,N_1060);
xnor U1453 (N_1453,N_493,N_973);
nand U1454 (N_1454,N_693,N_586);
nand U1455 (N_1455,N_562,N_509);
nand U1456 (N_1456,N_833,N_477);
nor U1457 (N_1457,N_441,N_1207);
nor U1458 (N_1458,N_173,N_169);
and U1459 (N_1459,N_1238,N_721);
nand U1460 (N_1460,N_749,N_126);
nand U1461 (N_1461,N_1030,N_612);
xor U1462 (N_1462,N_567,N_631);
and U1463 (N_1463,N_116,N_224);
nor U1464 (N_1464,N_242,N_792);
and U1465 (N_1465,N_489,N_187);
nor U1466 (N_1466,N_510,N_715);
or U1467 (N_1467,N_475,N_527);
xor U1468 (N_1468,N_915,N_524);
and U1469 (N_1469,N_884,N_35);
xor U1470 (N_1470,N_336,N_1237);
nand U1471 (N_1471,N_310,N_740);
and U1472 (N_1472,N_488,N_318);
xnor U1473 (N_1473,N_719,N_1098);
nor U1474 (N_1474,N_41,N_840);
and U1475 (N_1475,N_223,N_1141);
and U1476 (N_1476,N_1190,N_701);
nand U1477 (N_1477,N_158,N_879);
nand U1478 (N_1478,N_1213,N_545);
and U1479 (N_1479,N_780,N_676);
nand U1480 (N_1480,N_1150,N_520);
and U1481 (N_1481,N_1073,N_43);
nand U1482 (N_1482,N_1163,N_301);
or U1483 (N_1483,N_990,N_404);
xor U1484 (N_1484,N_121,N_809);
or U1485 (N_1485,N_131,N_53);
xnor U1486 (N_1486,N_377,N_135);
or U1487 (N_1487,N_1239,N_946);
xor U1488 (N_1488,N_753,N_272);
nor U1489 (N_1489,N_1149,N_72);
nor U1490 (N_1490,N_1008,N_314);
nand U1491 (N_1491,N_419,N_598);
xnor U1492 (N_1492,N_1142,N_482);
nand U1493 (N_1493,N_542,N_880);
nand U1494 (N_1494,N_938,N_78);
or U1495 (N_1495,N_132,N_771);
nand U1496 (N_1496,N_1087,N_730);
xnor U1497 (N_1497,N_718,N_361);
and U1498 (N_1498,N_1063,N_329);
xor U1499 (N_1499,N_874,N_999);
nand U1500 (N_1500,N_1231,N_699);
xor U1501 (N_1501,N_741,N_308);
nor U1502 (N_1502,N_47,N_850);
nor U1503 (N_1503,N_679,N_646);
nand U1504 (N_1504,N_474,N_353);
nand U1505 (N_1505,N_1245,N_383);
nor U1506 (N_1506,N_432,N_1195);
xor U1507 (N_1507,N_502,N_784);
nor U1508 (N_1508,N_431,N_623);
and U1509 (N_1509,N_994,N_170);
or U1510 (N_1510,N_164,N_890);
or U1511 (N_1511,N_1183,N_239);
xor U1512 (N_1512,N_260,N_221);
xor U1513 (N_1513,N_232,N_518);
xnor U1514 (N_1514,N_464,N_189);
and U1515 (N_1515,N_331,N_320);
or U1516 (N_1516,N_302,N_704);
and U1517 (N_1517,N_512,N_1071);
nand U1518 (N_1518,N_175,N_1121);
and U1519 (N_1519,N_966,N_396);
and U1520 (N_1520,N_33,N_471);
xnor U1521 (N_1521,N_1055,N_1153);
or U1522 (N_1522,N_276,N_1106);
nand U1523 (N_1523,N_621,N_1068);
xor U1524 (N_1524,N_417,N_748);
nor U1525 (N_1525,N_34,N_548);
and U1526 (N_1526,N_705,N_110);
nand U1527 (N_1527,N_129,N_823);
xnor U1528 (N_1528,N_57,N_297);
and U1529 (N_1529,N_451,N_65);
nand U1530 (N_1530,N_365,N_883);
nor U1531 (N_1531,N_83,N_337);
and U1532 (N_1532,N_13,N_642);
xor U1533 (N_1533,N_37,N_348);
and U1534 (N_1534,N_1059,N_654);
or U1535 (N_1535,N_148,N_708);
xnor U1536 (N_1536,N_418,N_141);
or U1537 (N_1537,N_713,N_1216);
xor U1538 (N_1538,N_866,N_245);
or U1539 (N_1539,N_433,N_685);
nor U1540 (N_1540,N_781,N_847);
and U1541 (N_1541,N_435,N_1051);
and U1542 (N_1542,N_237,N_111);
nand U1543 (N_1543,N_364,N_1218);
xor U1544 (N_1544,N_374,N_746);
and U1545 (N_1545,N_1242,N_947);
nand U1546 (N_1546,N_751,N_1235);
xnor U1547 (N_1547,N_875,N_1021);
xor U1548 (N_1548,N_660,N_1032);
nand U1549 (N_1549,N_610,N_429);
or U1550 (N_1550,N_1125,N_182);
and U1551 (N_1551,N_980,N_604);
nand U1552 (N_1552,N_694,N_265);
or U1553 (N_1553,N_1001,N_89);
nand U1554 (N_1554,N_1200,N_120);
and U1555 (N_1555,N_608,N_647);
and U1556 (N_1556,N_796,N_1044);
nor U1557 (N_1557,N_929,N_1161);
nand U1558 (N_1558,N_40,N_507);
nand U1559 (N_1559,N_238,N_909);
and U1560 (N_1560,N_900,N_965);
xor U1561 (N_1561,N_214,N_413);
nand U1562 (N_1562,N_269,N_504);
xor U1563 (N_1563,N_176,N_1025);
or U1564 (N_1564,N_505,N_319);
or U1565 (N_1565,N_113,N_9);
nand U1566 (N_1566,N_862,N_340);
nand U1567 (N_1567,N_949,N_864);
xor U1568 (N_1568,N_962,N_1146);
or U1569 (N_1569,N_549,N_138);
xor U1570 (N_1570,N_344,N_797);
or U1571 (N_1571,N_678,N_1135);
nand U1572 (N_1572,N_50,N_415);
xnor U1573 (N_1573,N_85,N_293);
nor U1574 (N_1574,N_802,N_142);
nand U1575 (N_1575,N_444,N_689);
or U1576 (N_1576,N_492,N_286);
xor U1577 (N_1577,N_1017,N_829);
xor U1578 (N_1578,N_445,N_555);
and U1579 (N_1579,N_1078,N_92);
xnor U1580 (N_1580,N_263,N_1038);
nand U1581 (N_1581,N_393,N_202);
or U1582 (N_1582,N_414,N_109);
xor U1583 (N_1583,N_316,N_559);
nand U1584 (N_1584,N_893,N_240);
or U1585 (N_1585,N_289,N_937);
and U1586 (N_1586,N_747,N_152);
nand U1587 (N_1587,N_468,N_852);
or U1588 (N_1588,N_146,N_387);
or U1589 (N_1589,N_149,N_769);
and U1590 (N_1590,N_714,N_1208);
or U1591 (N_1591,N_570,N_650);
nor U1592 (N_1592,N_686,N_1217);
and U1593 (N_1593,N_986,N_167);
nor U1594 (N_1594,N_709,N_369);
nand U1595 (N_1595,N_1103,N_421);
nor U1596 (N_1596,N_1187,N_1056);
nand U1597 (N_1597,N_889,N_858);
xor U1598 (N_1598,N_457,N_406);
or U1599 (N_1599,N_362,N_1047);
and U1600 (N_1600,N_74,N_892);
nand U1601 (N_1601,N_307,N_1209);
or U1602 (N_1602,N_794,N_60);
xnor U1603 (N_1603,N_1229,N_759);
and U1604 (N_1604,N_279,N_191);
xnor U1605 (N_1605,N_341,N_3);
nor U1606 (N_1606,N_630,N_494);
or U1607 (N_1607,N_616,N_1151);
xnor U1608 (N_1608,N_988,N_744);
xnor U1609 (N_1609,N_399,N_480);
nand U1610 (N_1610,N_400,N_82);
or U1611 (N_1611,N_497,N_48);
and U1612 (N_1612,N_770,N_800);
nand U1613 (N_1613,N_1020,N_1129);
or U1614 (N_1614,N_367,N_1205);
nor U1615 (N_1615,N_951,N_321);
nor U1616 (N_1616,N_854,N_1089);
xor U1617 (N_1617,N_773,N_1085);
nand U1618 (N_1618,N_215,N_816);
or U1619 (N_1619,N_443,N_295);
and U1620 (N_1620,N_918,N_247);
or U1621 (N_1621,N_774,N_273);
nand U1622 (N_1622,N_304,N_546);
and U1623 (N_1623,N_1022,N_323);
and U1624 (N_1624,N_430,N_684);
xor U1625 (N_1625,N_1210,N_697);
or U1626 (N_1626,N_1006,N_452);
xnor U1627 (N_1627,N_557,N_591);
xnor U1628 (N_1628,N_820,N_1197);
and U1629 (N_1629,N_73,N_28);
nand U1630 (N_1630,N_998,N_312);
and U1631 (N_1631,N_1248,N_27);
nor U1632 (N_1632,N_21,N_1124);
nor U1633 (N_1633,N_653,N_1157);
and U1634 (N_1634,N_723,N_776);
xnor U1635 (N_1635,N_508,N_544);
nor U1636 (N_1636,N_808,N_760);
or U1637 (N_1637,N_1105,N_1155);
and U1638 (N_1638,N_671,N_1199);
xor U1639 (N_1639,N_59,N_52);
or U1640 (N_1640,N_1014,N_343);
nor U1641 (N_1641,N_667,N_327);
xnor U1642 (N_1642,N_846,N_1181);
nand U1643 (N_1643,N_208,N_24);
xnor U1644 (N_1644,N_178,N_1175);
nor U1645 (N_1645,N_16,N_855);
nand U1646 (N_1646,N_372,N_71);
or U1647 (N_1647,N_722,N_160);
nor U1648 (N_1648,N_933,N_466);
and U1649 (N_1649,N_246,N_144);
nor U1650 (N_1650,N_359,N_573);
nand U1651 (N_1651,N_1113,N_426);
or U1652 (N_1652,N_594,N_181);
or U1653 (N_1653,N_298,N_856);
or U1654 (N_1654,N_657,N_1003);
nand U1655 (N_1655,N_706,N_199);
xor U1656 (N_1656,N_391,N_841);
and U1657 (N_1657,N_687,N_819);
and U1658 (N_1658,N_1174,N_19);
nor U1659 (N_1659,N_470,N_674);
and U1660 (N_1660,N_939,N_648);
xor U1661 (N_1661,N_1039,N_1194);
nor U1662 (N_1662,N_600,N_56);
nor U1663 (N_1663,N_381,N_885);
nand U1664 (N_1664,N_1091,N_560);
nor U1665 (N_1665,N_860,N_218);
xnor U1666 (N_1666,N_987,N_979);
nand U1667 (N_1667,N_1013,N_638);
nand U1668 (N_1668,N_325,N_1002);
or U1669 (N_1669,N_219,N_961);
and U1670 (N_1670,N_806,N_636);
xnor U1671 (N_1671,N_588,N_762);
nor U1672 (N_1672,N_801,N_943);
and U1673 (N_1673,N_1094,N_166);
and U1674 (N_1674,N_277,N_799);
nand U1675 (N_1675,N_197,N_728);
nand U1676 (N_1676,N_449,N_603);
and U1677 (N_1677,N_363,N_1090);
nor U1678 (N_1678,N_1000,N_830);
or U1679 (N_1679,N_456,N_734);
xnor U1680 (N_1680,N_865,N_691);
nand U1681 (N_1681,N_1031,N_521);
and U1682 (N_1682,N_354,N_392);
nand U1683 (N_1683,N_1011,N_61);
nor U1684 (N_1684,N_100,N_280);
xnor U1685 (N_1685,N_333,N_556);
or U1686 (N_1686,N_411,N_1037);
xnor U1687 (N_1687,N_1107,N_32);
xor U1688 (N_1688,N_1128,N_1123);
or U1689 (N_1689,N_291,N_177);
and U1690 (N_1690,N_945,N_117);
or U1691 (N_1691,N_401,N_1118);
xnor U1692 (N_1692,N_155,N_886);
nand U1693 (N_1693,N_717,N_533);
and U1694 (N_1694,N_79,N_285);
and U1695 (N_1695,N_38,N_484);
or U1696 (N_1696,N_859,N_118);
nor U1697 (N_1697,N_1131,N_1112);
or U1698 (N_1698,N_205,N_968);
nand U1699 (N_1699,N_894,N_94);
nand U1700 (N_1700,N_463,N_63);
nor U1701 (N_1701,N_992,N_1188);
nor U1702 (N_1702,N_870,N_632);
and U1703 (N_1703,N_29,N_1005);
or U1704 (N_1704,N_752,N_857);
nor U1705 (N_1705,N_1234,N_552);
or U1706 (N_1706,N_388,N_1004);
nor U1707 (N_1707,N_750,N_1166);
nor U1708 (N_1708,N_519,N_538);
and U1709 (N_1709,N_186,N_1046);
and U1710 (N_1710,N_698,N_370);
xor U1711 (N_1711,N_454,N_513);
nor U1712 (N_1712,N_324,N_617);
nor U1713 (N_1713,N_895,N_779);
or U1714 (N_1714,N_255,N_440);
nor U1715 (N_1715,N_1173,N_967);
nand U1716 (N_1716,N_1041,N_460);
nand U1717 (N_1717,N_436,N_1040);
nand U1718 (N_1718,N_499,N_515);
xor U1719 (N_1719,N_438,N_1081);
and U1720 (N_1720,N_1176,N_64);
and U1721 (N_1721,N_487,N_707);
nor U1722 (N_1722,N_534,N_408);
nor U1723 (N_1723,N_368,N_46);
nand U1724 (N_1724,N_2,N_516);
nand U1725 (N_1725,N_907,N_712);
xnor U1726 (N_1726,N_455,N_283);
or U1727 (N_1727,N_902,N_851);
nand U1728 (N_1728,N_1180,N_625);
nor U1729 (N_1729,N_1083,N_995);
or U1730 (N_1730,N_147,N_782);
nand U1731 (N_1731,N_124,N_1122);
and U1732 (N_1732,N_1136,N_134);
nand U1733 (N_1733,N_1082,N_241);
xor U1734 (N_1734,N_595,N_835);
xor U1735 (N_1735,N_249,N_1230);
xnor U1736 (N_1736,N_486,N_553);
nand U1737 (N_1737,N_566,N_88);
nor U1738 (N_1738,N_299,N_658);
nor U1739 (N_1739,N_597,N_601);
or U1740 (N_1740,N_640,N_159);
or U1741 (N_1741,N_941,N_795);
nor U1742 (N_1742,N_506,N_825);
xnor U1743 (N_1743,N_153,N_1053);
and U1744 (N_1744,N_948,N_1057);
xor U1745 (N_1745,N_842,N_1084);
xnor U1746 (N_1746,N_1192,N_1042);
xor U1747 (N_1747,N_899,N_725);
nand U1748 (N_1748,N_1225,N_1232);
nand U1749 (N_1749,N_785,N_989);
and U1750 (N_1750,N_54,N_743);
and U1751 (N_1751,N_1170,N_81);
and U1752 (N_1752,N_688,N_758);
nand U1753 (N_1753,N_20,N_188);
and U1754 (N_1754,N_1127,N_659);
xnor U1755 (N_1755,N_351,N_86);
nand U1756 (N_1756,N_163,N_1186);
xor U1757 (N_1757,N_1075,N_1152);
nand U1758 (N_1758,N_959,N_872);
and U1759 (N_1759,N_1171,N_115);
nand U1760 (N_1760,N_1062,N_810);
and U1761 (N_1761,N_922,N_978);
nor U1762 (N_1762,N_122,N_1117);
and U1763 (N_1763,N_12,N_757);
nand U1764 (N_1764,N_683,N_1201);
and U1765 (N_1765,N_228,N_200);
or U1766 (N_1766,N_261,N_403);
nor U1767 (N_1767,N_1064,N_729);
and U1768 (N_1768,N_101,N_80);
nand U1769 (N_1769,N_957,N_976);
nor U1770 (N_1770,N_196,N_317);
or U1771 (N_1771,N_1119,N_695);
xor U1772 (N_1772,N_137,N_655);
or U1773 (N_1773,N_442,N_618);
or U1774 (N_1774,N_267,N_582);
nor U1775 (N_1775,N_1160,N_284);
xnor U1776 (N_1776,N_58,N_665);
and U1777 (N_1777,N_614,N_62);
nand U1778 (N_1778,N_386,N_984);
and U1779 (N_1779,N_49,N_11);
nand U1780 (N_1780,N_1092,N_184);
or U1781 (N_1781,N_1054,N_338);
or U1782 (N_1782,N_104,N_643);
xor U1783 (N_1783,N_161,N_927);
xnor U1784 (N_1784,N_409,N_23);
and U1785 (N_1785,N_1015,N_523);
or U1786 (N_1786,N_554,N_1236);
nor U1787 (N_1787,N_778,N_656);
or U1788 (N_1788,N_345,N_233);
xnor U1789 (N_1789,N_91,N_633);
or U1790 (N_1790,N_528,N_1007);
nand U1791 (N_1791,N_826,N_185);
xor U1792 (N_1792,N_398,N_1167);
and U1793 (N_1793,N_550,N_1182);
or U1794 (N_1794,N_275,N_956);
or U1795 (N_1795,N_1134,N_547);
and U1796 (N_1796,N_649,N_910);
and U1797 (N_1797,N_581,N_720);
and U1798 (N_1798,N_977,N_543);
nand U1799 (N_1799,N_230,N_36);
or U1800 (N_1800,N_346,N_1220);
and U1801 (N_1801,N_469,N_51);
xnor U1802 (N_1802,N_42,N_503);
nand U1803 (N_1803,N_942,N_395);
or U1804 (N_1804,N_952,N_923);
xor U1805 (N_1805,N_139,N_696);
xor U1806 (N_1806,N_350,N_1179);
or U1807 (N_1807,N_87,N_869);
xnor U1808 (N_1808,N_913,N_198);
and U1809 (N_1809,N_807,N_932);
xor U1810 (N_1810,N_1019,N_564);
nor U1811 (N_1811,N_373,N_98);
and U1812 (N_1812,N_700,N_309);
nor U1813 (N_1813,N_95,N_424);
nor U1814 (N_1814,N_982,N_274);
and U1815 (N_1815,N_898,N_1099);
xor U1816 (N_1816,N_44,N_805);
and U1817 (N_1817,N_1126,N_366);
and U1818 (N_1818,N_790,N_222);
or U1819 (N_1819,N_1206,N_775);
xor U1820 (N_1820,N_1172,N_1214);
or U1821 (N_1821,N_887,N_1104);
and U1822 (N_1822,N_593,N_123);
and U1823 (N_1823,N_67,N_901);
nand U1824 (N_1824,N_465,N_525);
nor U1825 (N_1825,N_786,N_472);
or U1826 (N_1826,N_183,N_863);
or U1827 (N_1827,N_793,N_955);
nand U1828 (N_1828,N_739,N_1072);
xnor U1829 (N_1829,N_450,N_1198);
nor U1830 (N_1830,N_1065,N_661);
xor U1831 (N_1831,N_972,N_69);
and U1832 (N_1832,N_1132,N_8);
and U1833 (N_1833,N_26,N_896);
or U1834 (N_1834,N_662,N_254);
and U1835 (N_1835,N_1108,N_93);
and U1836 (N_1836,N_964,N_903);
or U1837 (N_1837,N_963,N_271);
or U1838 (N_1838,N_252,N_410);
xnor U1839 (N_1839,N_1244,N_812);
or U1840 (N_1840,N_306,N_914);
or U1841 (N_1841,N_663,N_912);
and U1842 (N_1842,N_357,N_536);
and U1843 (N_1843,N_644,N_822);
nor U1844 (N_1844,N_330,N_389);
or U1845 (N_1845,N_1058,N_97);
and U1846 (N_1846,N_172,N_574);
or U1847 (N_1847,N_356,N_579);
and U1848 (N_1848,N_1028,N_195);
nor U1849 (N_1849,N_305,N_613);
nor U1850 (N_1850,N_1203,N_767);
nand U1851 (N_1851,N_668,N_491);
xnor U1852 (N_1852,N_425,N_971);
nor U1853 (N_1853,N_837,N_958);
or U1854 (N_1854,N_1035,N_831);
nand U1855 (N_1855,N_334,N_1101);
xor U1856 (N_1856,N_735,N_193);
and U1857 (N_1857,N_1193,N_394);
xnor U1858 (N_1858,N_1097,N_1050);
or U1859 (N_1859,N_590,N_1162);
xor U1860 (N_1860,N_541,N_522);
or U1861 (N_1861,N_1114,N_1018);
or U1862 (N_1862,N_162,N_763);
and U1863 (N_1863,N_814,N_738);
nor U1864 (N_1864,N_201,N_1156);
or U1865 (N_1865,N_853,N_229);
xnor U1866 (N_1866,N_204,N_1102);
and U1867 (N_1867,N_817,N_1093);
nand U1868 (N_1868,N_615,N_66);
xor U1869 (N_1869,N_940,N_789);
nand U1870 (N_1870,N_1147,N_461);
and U1871 (N_1871,N_711,N_911);
or U1872 (N_1872,N_871,N_589);
and U1873 (N_1873,N_975,N_6);
xnor U1874 (N_1874,N_251,N_18);
xor U1875 (N_1875,N_314,N_551);
nor U1876 (N_1876,N_543,N_1137);
nor U1877 (N_1877,N_117,N_1192);
or U1878 (N_1878,N_855,N_129);
xnor U1879 (N_1879,N_235,N_290);
nor U1880 (N_1880,N_1099,N_477);
and U1881 (N_1881,N_101,N_1110);
nand U1882 (N_1882,N_485,N_706);
nand U1883 (N_1883,N_837,N_146);
nand U1884 (N_1884,N_443,N_310);
xnor U1885 (N_1885,N_1152,N_312);
or U1886 (N_1886,N_1224,N_92);
or U1887 (N_1887,N_295,N_738);
nand U1888 (N_1888,N_968,N_423);
nand U1889 (N_1889,N_987,N_1034);
and U1890 (N_1890,N_1019,N_876);
nor U1891 (N_1891,N_1172,N_75);
and U1892 (N_1892,N_415,N_1066);
and U1893 (N_1893,N_952,N_882);
or U1894 (N_1894,N_20,N_562);
xnor U1895 (N_1895,N_576,N_26);
nand U1896 (N_1896,N_1073,N_73);
or U1897 (N_1897,N_534,N_571);
xnor U1898 (N_1898,N_210,N_1208);
and U1899 (N_1899,N_307,N_374);
nor U1900 (N_1900,N_630,N_182);
or U1901 (N_1901,N_264,N_317);
xnor U1902 (N_1902,N_733,N_1226);
nand U1903 (N_1903,N_1111,N_758);
and U1904 (N_1904,N_381,N_1032);
nand U1905 (N_1905,N_320,N_563);
nand U1906 (N_1906,N_128,N_211);
nor U1907 (N_1907,N_259,N_515);
or U1908 (N_1908,N_165,N_524);
nor U1909 (N_1909,N_1085,N_772);
nor U1910 (N_1910,N_555,N_131);
nand U1911 (N_1911,N_756,N_148);
nor U1912 (N_1912,N_13,N_748);
or U1913 (N_1913,N_800,N_1074);
xor U1914 (N_1914,N_804,N_802);
or U1915 (N_1915,N_271,N_703);
and U1916 (N_1916,N_1198,N_1194);
nor U1917 (N_1917,N_551,N_8);
nor U1918 (N_1918,N_541,N_1228);
and U1919 (N_1919,N_214,N_641);
nor U1920 (N_1920,N_766,N_1054);
and U1921 (N_1921,N_272,N_706);
and U1922 (N_1922,N_7,N_1238);
nand U1923 (N_1923,N_124,N_820);
or U1924 (N_1924,N_718,N_918);
nor U1925 (N_1925,N_726,N_292);
nor U1926 (N_1926,N_475,N_561);
nor U1927 (N_1927,N_979,N_604);
xnor U1928 (N_1928,N_883,N_493);
and U1929 (N_1929,N_1182,N_146);
and U1930 (N_1930,N_267,N_744);
nor U1931 (N_1931,N_154,N_611);
nand U1932 (N_1932,N_1167,N_79);
xnor U1933 (N_1933,N_243,N_55);
nor U1934 (N_1934,N_214,N_494);
or U1935 (N_1935,N_577,N_873);
xnor U1936 (N_1936,N_825,N_923);
xnor U1937 (N_1937,N_721,N_433);
nand U1938 (N_1938,N_442,N_1219);
nor U1939 (N_1939,N_648,N_476);
xor U1940 (N_1940,N_705,N_37);
and U1941 (N_1941,N_232,N_105);
or U1942 (N_1942,N_375,N_664);
xnor U1943 (N_1943,N_848,N_260);
nand U1944 (N_1944,N_23,N_151);
nand U1945 (N_1945,N_824,N_641);
and U1946 (N_1946,N_311,N_34);
nand U1947 (N_1947,N_182,N_544);
nand U1948 (N_1948,N_709,N_330);
nand U1949 (N_1949,N_1172,N_106);
or U1950 (N_1950,N_250,N_118);
nor U1951 (N_1951,N_166,N_992);
nand U1952 (N_1952,N_925,N_891);
nand U1953 (N_1953,N_1114,N_465);
nor U1954 (N_1954,N_459,N_666);
xnor U1955 (N_1955,N_46,N_1115);
and U1956 (N_1956,N_30,N_1161);
and U1957 (N_1957,N_44,N_186);
nor U1958 (N_1958,N_250,N_557);
xnor U1959 (N_1959,N_452,N_48);
xor U1960 (N_1960,N_35,N_949);
xnor U1961 (N_1961,N_184,N_225);
nand U1962 (N_1962,N_1172,N_293);
and U1963 (N_1963,N_812,N_263);
nor U1964 (N_1964,N_662,N_723);
xnor U1965 (N_1965,N_445,N_476);
nand U1966 (N_1966,N_796,N_40);
xor U1967 (N_1967,N_273,N_609);
nand U1968 (N_1968,N_269,N_291);
or U1969 (N_1969,N_798,N_27);
or U1970 (N_1970,N_666,N_674);
and U1971 (N_1971,N_924,N_568);
nor U1972 (N_1972,N_205,N_1108);
nand U1973 (N_1973,N_544,N_826);
and U1974 (N_1974,N_1122,N_383);
xnor U1975 (N_1975,N_886,N_1001);
and U1976 (N_1976,N_834,N_371);
xnor U1977 (N_1977,N_1062,N_1218);
nor U1978 (N_1978,N_186,N_1063);
nand U1979 (N_1979,N_1174,N_436);
and U1980 (N_1980,N_631,N_487);
nand U1981 (N_1981,N_1126,N_533);
and U1982 (N_1982,N_503,N_1109);
nand U1983 (N_1983,N_1208,N_153);
or U1984 (N_1984,N_169,N_188);
or U1985 (N_1985,N_12,N_979);
and U1986 (N_1986,N_92,N_589);
and U1987 (N_1987,N_305,N_999);
xnor U1988 (N_1988,N_408,N_563);
or U1989 (N_1989,N_366,N_749);
nand U1990 (N_1990,N_173,N_1078);
and U1991 (N_1991,N_1220,N_34);
xor U1992 (N_1992,N_808,N_1139);
nand U1993 (N_1993,N_363,N_921);
nand U1994 (N_1994,N_949,N_836);
xnor U1995 (N_1995,N_342,N_708);
xnor U1996 (N_1996,N_844,N_300);
and U1997 (N_1997,N_1021,N_488);
nor U1998 (N_1998,N_1066,N_522);
nand U1999 (N_1999,N_164,N_999);
nand U2000 (N_2000,N_113,N_860);
or U2001 (N_2001,N_790,N_502);
nor U2002 (N_2002,N_62,N_696);
nand U2003 (N_2003,N_958,N_933);
or U2004 (N_2004,N_570,N_972);
or U2005 (N_2005,N_509,N_280);
or U2006 (N_2006,N_209,N_446);
or U2007 (N_2007,N_449,N_770);
or U2008 (N_2008,N_1169,N_611);
and U2009 (N_2009,N_1135,N_1173);
and U2010 (N_2010,N_1148,N_395);
xnor U2011 (N_2011,N_105,N_524);
nor U2012 (N_2012,N_941,N_391);
or U2013 (N_2013,N_764,N_954);
nor U2014 (N_2014,N_454,N_1108);
nor U2015 (N_2015,N_249,N_976);
xor U2016 (N_2016,N_381,N_783);
xnor U2017 (N_2017,N_1113,N_815);
nor U2018 (N_2018,N_392,N_522);
and U2019 (N_2019,N_1210,N_37);
nand U2020 (N_2020,N_1094,N_127);
and U2021 (N_2021,N_25,N_866);
nor U2022 (N_2022,N_773,N_184);
nor U2023 (N_2023,N_1063,N_274);
nand U2024 (N_2024,N_943,N_221);
or U2025 (N_2025,N_32,N_545);
nor U2026 (N_2026,N_145,N_119);
or U2027 (N_2027,N_1247,N_436);
nor U2028 (N_2028,N_1009,N_676);
nor U2029 (N_2029,N_238,N_313);
xor U2030 (N_2030,N_1032,N_174);
or U2031 (N_2031,N_883,N_741);
nand U2032 (N_2032,N_1191,N_1179);
nor U2033 (N_2033,N_934,N_98);
xor U2034 (N_2034,N_470,N_258);
nor U2035 (N_2035,N_197,N_856);
nand U2036 (N_2036,N_663,N_736);
nand U2037 (N_2037,N_377,N_963);
or U2038 (N_2038,N_387,N_460);
xor U2039 (N_2039,N_653,N_85);
and U2040 (N_2040,N_791,N_830);
nand U2041 (N_2041,N_733,N_1019);
nand U2042 (N_2042,N_1114,N_581);
or U2043 (N_2043,N_74,N_520);
or U2044 (N_2044,N_484,N_979);
xor U2045 (N_2045,N_160,N_56);
or U2046 (N_2046,N_249,N_844);
xor U2047 (N_2047,N_1200,N_351);
nor U2048 (N_2048,N_69,N_530);
xnor U2049 (N_2049,N_309,N_974);
or U2050 (N_2050,N_812,N_492);
xor U2051 (N_2051,N_254,N_50);
nor U2052 (N_2052,N_638,N_724);
nor U2053 (N_2053,N_1057,N_438);
nand U2054 (N_2054,N_1010,N_404);
nand U2055 (N_2055,N_13,N_1167);
nor U2056 (N_2056,N_20,N_553);
and U2057 (N_2057,N_969,N_414);
nand U2058 (N_2058,N_790,N_181);
or U2059 (N_2059,N_996,N_1248);
xnor U2060 (N_2060,N_778,N_501);
nand U2061 (N_2061,N_960,N_677);
or U2062 (N_2062,N_119,N_173);
nor U2063 (N_2063,N_1075,N_330);
nand U2064 (N_2064,N_379,N_1119);
nor U2065 (N_2065,N_849,N_468);
nand U2066 (N_2066,N_234,N_688);
and U2067 (N_2067,N_862,N_77);
and U2068 (N_2068,N_681,N_1083);
xnor U2069 (N_2069,N_689,N_838);
nand U2070 (N_2070,N_837,N_1157);
xor U2071 (N_2071,N_242,N_210);
nor U2072 (N_2072,N_76,N_210);
nand U2073 (N_2073,N_254,N_221);
or U2074 (N_2074,N_691,N_1125);
xor U2075 (N_2075,N_1192,N_688);
and U2076 (N_2076,N_744,N_1233);
and U2077 (N_2077,N_35,N_701);
nand U2078 (N_2078,N_884,N_1051);
or U2079 (N_2079,N_159,N_690);
or U2080 (N_2080,N_278,N_304);
and U2081 (N_2081,N_715,N_500);
or U2082 (N_2082,N_614,N_4);
nand U2083 (N_2083,N_239,N_1094);
or U2084 (N_2084,N_982,N_1222);
nor U2085 (N_2085,N_794,N_96);
and U2086 (N_2086,N_874,N_162);
nor U2087 (N_2087,N_278,N_452);
nor U2088 (N_2088,N_795,N_246);
and U2089 (N_2089,N_700,N_243);
and U2090 (N_2090,N_293,N_69);
nand U2091 (N_2091,N_1041,N_404);
and U2092 (N_2092,N_837,N_338);
nor U2093 (N_2093,N_150,N_303);
or U2094 (N_2094,N_465,N_399);
or U2095 (N_2095,N_418,N_95);
xnor U2096 (N_2096,N_107,N_498);
nor U2097 (N_2097,N_721,N_1248);
nand U2098 (N_2098,N_391,N_305);
nand U2099 (N_2099,N_532,N_72);
xnor U2100 (N_2100,N_1145,N_530);
nand U2101 (N_2101,N_309,N_872);
and U2102 (N_2102,N_1140,N_804);
nor U2103 (N_2103,N_618,N_418);
and U2104 (N_2104,N_728,N_225);
xnor U2105 (N_2105,N_46,N_150);
xnor U2106 (N_2106,N_531,N_187);
or U2107 (N_2107,N_1212,N_978);
xnor U2108 (N_2108,N_835,N_857);
or U2109 (N_2109,N_1126,N_25);
nor U2110 (N_2110,N_440,N_798);
nand U2111 (N_2111,N_242,N_1202);
or U2112 (N_2112,N_972,N_1125);
and U2113 (N_2113,N_615,N_790);
nand U2114 (N_2114,N_954,N_1189);
and U2115 (N_2115,N_1162,N_230);
and U2116 (N_2116,N_667,N_357);
nand U2117 (N_2117,N_170,N_930);
xor U2118 (N_2118,N_768,N_1087);
and U2119 (N_2119,N_379,N_357);
nor U2120 (N_2120,N_620,N_289);
nand U2121 (N_2121,N_1008,N_44);
nor U2122 (N_2122,N_346,N_676);
or U2123 (N_2123,N_660,N_473);
xor U2124 (N_2124,N_618,N_655);
nand U2125 (N_2125,N_435,N_482);
nor U2126 (N_2126,N_413,N_647);
and U2127 (N_2127,N_88,N_160);
and U2128 (N_2128,N_1171,N_595);
xnor U2129 (N_2129,N_146,N_90);
nor U2130 (N_2130,N_468,N_712);
xnor U2131 (N_2131,N_269,N_769);
nand U2132 (N_2132,N_275,N_391);
xnor U2133 (N_2133,N_1030,N_348);
nor U2134 (N_2134,N_807,N_420);
nand U2135 (N_2135,N_206,N_683);
nor U2136 (N_2136,N_234,N_352);
or U2137 (N_2137,N_892,N_552);
nand U2138 (N_2138,N_281,N_212);
nand U2139 (N_2139,N_719,N_85);
or U2140 (N_2140,N_41,N_160);
or U2141 (N_2141,N_474,N_72);
nor U2142 (N_2142,N_1170,N_413);
nor U2143 (N_2143,N_332,N_645);
xor U2144 (N_2144,N_574,N_1154);
nand U2145 (N_2145,N_1150,N_779);
and U2146 (N_2146,N_233,N_303);
nand U2147 (N_2147,N_704,N_528);
nor U2148 (N_2148,N_1104,N_1084);
and U2149 (N_2149,N_1209,N_571);
xor U2150 (N_2150,N_168,N_1);
xnor U2151 (N_2151,N_1153,N_132);
and U2152 (N_2152,N_144,N_153);
nor U2153 (N_2153,N_220,N_190);
nor U2154 (N_2154,N_120,N_847);
or U2155 (N_2155,N_788,N_1072);
nand U2156 (N_2156,N_523,N_1007);
nand U2157 (N_2157,N_904,N_777);
nor U2158 (N_2158,N_804,N_545);
xnor U2159 (N_2159,N_1078,N_669);
nor U2160 (N_2160,N_614,N_187);
and U2161 (N_2161,N_62,N_69);
nand U2162 (N_2162,N_599,N_521);
nand U2163 (N_2163,N_70,N_528);
or U2164 (N_2164,N_177,N_839);
xor U2165 (N_2165,N_878,N_135);
and U2166 (N_2166,N_657,N_1077);
xnor U2167 (N_2167,N_217,N_28);
nor U2168 (N_2168,N_999,N_77);
nor U2169 (N_2169,N_5,N_1221);
and U2170 (N_2170,N_67,N_1062);
xnor U2171 (N_2171,N_325,N_235);
nand U2172 (N_2172,N_639,N_1178);
xnor U2173 (N_2173,N_251,N_3);
xor U2174 (N_2174,N_604,N_264);
nor U2175 (N_2175,N_240,N_1136);
xor U2176 (N_2176,N_1151,N_706);
nand U2177 (N_2177,N_1007,N_867);
nor U2178 (N_2178,N_687,N_360);
and U2179 (N_2179,N_879,N_992);
nor U2180 (N_2180,N_389,N_995);
xor U2181 (N_2181,N_875,N_293);
xnor U2182 (N_2182,N_317,N_675);
and U2183 (N_2183,N_892,N_763);
xor U2184 (N_2184,N_345,N_837);
nand U2185 (N_2185,N_663,N_1178);
and U2186 (N_2186,N_473,N_857);
nor U2187 (N_2187,N_119,N_303);
nor U2188 (N_2188,N_1235,N_753);
and U2189 (N_2189,N_1083,N_945);
and U2190 (N_2190,N_1027,N_823);
and U2191 (N_2191,N_626,N_312);
xor U2192 (N_2192,N_923,N_647);
nor U2193 (N_2193,N_673,N_885);
and U2194 (N_2194,N_1096,N_562);
and U2195 (N_2195,N_960,N_419);
and U2196 (N_2196,N_512,N_534);
or U2197 (N_2197,N_32,N_194);
xnor U2198 (N_2198,N_720,N_1118);
xnor U2199 (N_2199,N_178,N_223);
and U2200 (N_2200,N_1017,N_713);
nand U2201 (N_2201,N_321,N_1119);
nand U2202 (N_2202,N_12,N_626);
and U2203 (N_2203,N_129,N_199);
or U2204 (N_2204,N_933,N_586);
nor U2205 (N_2205,N_531,N_916);
and U2206 (N_2206,N_816,N_788);
and U2207 (N_2207,N_134,N_847);
xnor U2208 (N_2208,N_1011,N_1226);
xor U2209 (N_2209,N_254,N_287);
and U2210 (N_2210,N_295,N_322);
nand U2211 (N_2211,N_314,N_769);
nand U2212 (N_2212,N_296,N_64);
xor U2213 (N_2213,N_1109,N_199);
nand U2214 (N_2214,N_402,N_910);
xnor U2215 (N_2215,N_692,N_812);
or U2216 (N_2216,N_168,N_1072);
xnor U2217 (N_2217,N_78,N_1038);
or U2218 (N_2218,N_545,N_910);
nor U2219 (N_2219,N_737,N_211);
or U2220 (N_2220,N_1115,N_121);
or U2221 (N_2221,N_854,N_592);
nor U2222 (N_2222,N_536,N_614);
and U2223 (N_2223,N_282,N_1107);
nor U2224 (N_2224,N_983,N_393);
or U2225 (N_2225,N_108,N_1051);
xor U2226 (N_2226,N_174,N_460);
nor U2227 (N_2227,N_30,N_225);
nand U2228 (N_2228,N_742,N_207);
nor U2229 (N_2229,N_40,N_454);
and U2230 (N_2230,N_1147,N_210);
and U2231 (N_2231,N_271,N_569);
nor U2232 (N_2232,N_1059,N_536);
nand U2233 (N_2233,N_85,N_1134);
and U2234 (N_2234,N_441,N_33);
xor U2235 (N_2235,N_558,N_863);
nor U2236 (N_2236,N_704,N_721);
nor U2237 (N_2237,N_644,N_545);
and U2238 (N_2238,N_812,N_808);
and U2239 (N_2239,N_906,N_746);
xnor U2240 (N_2240,N_346,N_471);
and U2241 (N_2241,N_72,N_373);
and U2242 (N_2242,N_184,N_190);
nor U2243 (N_2243,N_242,N_354);
or U2244 (N_2244,N_1205,N_771);
nor U2245 (N_2245,N_798,N_178);
xnor U2246 (N_2246,N_1057,N_625);
nand U2247 (N_2247,N_811,N_891);
and U2248 (N_2248,N_540,N_476);
nor U2249 (N_2249,N_819,N_716);
nand U2250 (N_2250,N_215,N_726);
and U2251 (N_2251,N_1195,N_687);
xor U2252 (N_2252,N_747,N_18);
nor U2253 (N_2253,N_89,N_398);
nand U2254 (N_2254,N_669,N_41);
or U2255 (N_2255,N_1063,N_905);
and U2256 (N_2256,N_1051,N_768);
nor U2257 (N_2257,N_788,N_197);
nand U2258 (N_2258,N_498,N_442);
or U2259 (N_2259,N_1128,N_806);
nor U2260 (N_2260,N_266,N_1087);
nor U2261 (N_2261,N_636,N_362);
and U2262 (N_2262,N_822,N_444);
xnor U2263 (N_2263,N_221,N_1126);
or U2264 (N_2264,N_1116,N_891);
nand U2265 (N_2265,N_953,N_272);
nor U2266 (N_2266,N_508,N_162);
and U2267 (N_2267,N_454,N_1136);
and U2268 (N_2268,N_1218,N_1079);
and U2269 (N_2269,N_252,N_325);
xnor U2270 (N_2270,N_532,N_597);
nor U2271 (N_2271,N_754,N_389);
or U2272 (N_2272,N_554,N_1183);
nand U2273 (N_2273,N_516,N_29);
and U2274 (N_2274,N_989,N_132);
or U2275 (N_2275,N_535,N_686);
or U2276 (N_2276,N_221,N_1116);
nor U2277 (N_2277,N_349,N_289);
nor U2278 (N_2278,N_568,N_946);
nand U2279 (N_2279,N_144,N_1099);
or U2280 (N_2280,N_627,N_8);
or U2281 (N_2281,N_358,N_790);
nor U2282 (N_2282,N_82,N_698);
or U2283 (N_2283,N_488,N_812);
xnor U2284 (N_2284,N_337,N_1175);
and U2285 (N_2285,N_200,N_1106);
nor U2286 (N_2286,N_101,N_848);
nor U2287 (N_2287,N_0,N_871);
or U2288 (N_2288,N_303,N_432);
xor U2289 (N_2289,N_835,N_273);
nor U2290 (N_2290,N_635,N_185);
and U2291 (N_2291,N_256,N_67);
nand U2292 (N_2292,N_317,N_908);
and U2293 (N_2293,N_550,N_433);
nand U2294 (N_2294,N_456,N_733);
xnor U2295 (N_2295,N_353,N_1063);
and U2296 (N_2296,N_8,N_1243);
or U2297 (N_2297,N_1079,N_1110);
and U2298 (N_2298,N_349,N_420);
or U2299 (N_2299,N_623,N_673);
nor U2300 (N_2300,N_735,N_829);
or U2301 (N_2301,N_603,N_837);
and U2302 (N_2302,N_1042,N_1242);
or U2303 (N_2303,N_1077,N_945);
nor U2304 (N_2304,N_1170,N_1245);
or U2305 (N_2305,N_559,N_1065);
and U2306 (N_2306,N_923,N_780);
xor U2307 (N_2307,N_375,N_629);
xor U2308 (N_2308,N_389,N_186);
nor U2309 (N_2309,N_750,N_1117);
nor U2310 (N_2310,N_502,N_709);
and U2311 (N_2311,N_369,N_1143);
and U2312 (N_2312,N_1042,N_394);
nand U2313 (N_2313,N_1131,N_520);
nor U2314 (N_2314,N_659,N_845);
nand U2315 (N_2315,N_453,N_248);
nand U2316 (N_2316,N_1172,N_302);
nor U2317 (N_2317,N_197,N_1043);
and U2318 (N_2318,N_781,N_759);
and U2319 (N_2319,N_492,N_185);
nand U2320 (N_2320,N_1057,N_161);
nand U2321 (N_2321,N_513,N_869);
nor U2322 (N_2322,N_70,N_1);
or U2323 (N_2323,N_624,N_838);
nand U2324 (N_2324,N_45,N_63);
and U2325 (N_2325,N_1190,N_963);
xor U2326 (N_2326,N_934,N_760);
or U2327 (N_2327,N_1106,N_407);
or U2328 (N_2328,N_1178,N_1121);
and U2329 (N_2329,N_1097,N_749);
nand U2330 (N_2330,N_1147,N_44);
or U2331 (N_2331,N_1158,N_1110);
xor U2332 (N_2332,N_683,N_543);
xnor U2333 (N_2333,N_921,N_189);
xor U2334 (N_2334,N_498,N_911);
and U2335 (N_2335,N_317,N_100);
nand U2336 (N_2336,N_460,N_1204);
or U2337 (N_2337,N_300,N_942);
xor U2338 (N_2338,N_71,N_1202);
or U2339 (N_2339,N_527,N_136);
nand U2340 (N_2340,N_245,N_941);
and U2341 (N_2341,N_744,N_287);
nand U2342 (N_2342,N_1219,N_234);
and U2343 (N_2343,N_192,N_1138);
xnor U2344 (N_2344,N_206,N_379);
or U2345 (N_2345,N_538,N_86);
nor U2346 (N_2346,N_679,N_674);
or U2347 (N_2347,N_732,N_774);
and U2348 (N_2348,N_924,N_222);
or U2349 (N_2349,N_410,N_1019);
or U2350 (N_2350,N_294,N_427);
nor U2351 (N_2351,N_1220,N_620);
or U2352 (N_2352,N_716,N_537);
or U2353 (N_2353,N_886,N_78);
nand U2354 (N_2354,N_55,N_252);
xor U2355 (N_2355,N_246,N_1094);
nor U2356 (N_2356,N_959,N_31);
nand U2357 (N_2357,N_162,N_663);
nand U2358 (N_2358,N_690,N_1032);
xnor U2359 (N_2359,N_1008,N_676);
xor U2360 (N_2360,N_878,N_531);
xor U2361 (N_2361,N_300,N_480);
nor U2362 (N_2362,N_229,N_614);
nand U2363 (N_2363,N_270,N_336);
nor U2364 (N_2364,N_979,N_761);
xnor U2365 (N_2365,N_818,N_962);
or U2366 (N_2366,N_336,N_445);
xnor U2367 (N_2367,N_211,N_801);
nand U2368 (N_2368,N_16,N_1153);
xnor U2369 (N_2369,N_134,N_882);
nor U2370 (N_2370,N_84,N_225);
nand U2371 (N_2371,N_1146,N_322);
xor U2372 (N_2372,N_3,N_1124);
nor U2373 (N_2373,N_163,N_1003);
xor U2374 (N_2374,N_1030,N_422);
or U2375 (N_2375,N_890,N_1014);
nand U2376 (N_2376,N_90,N_305);
nand U2377 (N_2377,N_576,N_293);
xor U2378 (N_2378,N_453,N_75);
or U2379 (N_2379,N_133,N_771);
nand U2380 (N_2380,N_345,N_40);
nand U2381 (N_2381,N_287,N_441);
and U2382 (N_2382,N_1139,N_161);
nor U2383 (N_2383,N_845,N_303);
xnor U2384 (N_2384,N_831,N_97);
nand U2385 (N_2385,N_606,N_166);
or U2386 (N_2386,N_678,N_1183);
xor U2387 (N_2387,N_1078,N_846);
and U2388 (N_2388,N_884,N_970);
xor U2389 (N_2389,N_517,N_947);
and U2390 (N_2390,N_1186,N_816);
or U2391 (N_2391,N_739,N_831);
nor U2392 (N_2392,N_1120,N_1181);
or U2393 (N_2393,N_666,N_500);
xnor U2394 (N_2394,N_819,N_441);
nor U2395 (N_2395,N_182,N_169);
nor U2396 (N_2396,N_441,N_891);
and U2397 (N_2397,N_365,N_898);
and U2398 (N_2398,N_72,N_625);
nand U2399 (N_2399,N_879,N_794);
or U2400 (N_2400,N_676,N_87);
or U2401 (N_2401,N_838,N_439);
and U2402 (N_2402,N_586,N_375);
or U2403 (N_2403,N_0,N_70);
nand U2404 (N_2404,N_848,N_718);
nand U2405 (N_2405,N_484,N_1002);
or U2406 (N_2406,N_145,N_756);
nor U2407 (N_2407,N_991,N_1194);
xor U2408 (N_2408,N_423,N_396);
and U2409 (N_2409,N_835,N_220);
nor U2410 (N_2410,N_272,N_944);
nand U2411 (N_2411,N_281,N_418);
xnor U2412 (N_2412,N_669,N_79);
and U2413 (N_2413,N_515,N_1132);
nand U2414 (N_2414,N_510,N_851);
nor U2415 (N_2415,N_881,N_756);
xnor U2416 (N_2416,N_317,N_553);
or U2417 (N_2417,N_316,N_911);
and U2418 (N_2418,N_846,N_555);
or U2419 (N_2419,N_834,N_521);
and U2420 (N_2420,N_455,N_910);
nor U2421 (N_2421,N_623,N_667);
nor U2422 (N_2422,N_960,N_734);
or U2423 (N_2423,N_776,N_732);
nand U2424 (N_2424,N_260,N_36);
or U2425 (N_2425,N_1203,N_305);
or U2426 (N_2426,N_697,N_1124);
and U2427 (N_2427,N_238,N_884);
nand U2428 (N_2428,N_205,N_1157);
nand U2429 (N_2429,N_1131,N_807);
xor U2430 (N_2430,N_392,N_2);
xnor U2431 (N_2431,N_347,N_1090);
nand U2432 (N_2432,N_1120,N_655);
or U2433 (N_2433,N_1163,N_534);
nand U2434 (N_2434,N_596,N_933);
and U2435 (N_2435,N_932,N_834);
or U2436 (N_2436,N_142,N_106);
xnor U2437 (N_2437,N_838,N_48);
or U2438 (N_2438,N_417,N_790);
and U2439 (N_2439,N_631,N_934);
nor U2440 (N_2440,N_710,N_71);
or U2441 (N_2441,N_129,N_1065);
nor U2442 (N_2442,N_988,N_1062);
nand U2443 (N_2443,N_883,N_61);
or U2444 (N_2444,N_940,N_1044);
and U2445 (N_2445,N_915,N_916);
or U2446 (N_2446,N_534,N_1160);
nand U2447 (N_2447,N_258,N_639);
xor U2448 (N_2448,N_929,N_158);
or U2449 (N_2449,N_399,N_878);
nor U2450 (N_2450,N_876,N_458);
xor U2451 (N_2451,N_973,N_23);
nand U2452 (N_2452,N_25,N_546);
nor U2453 (N_2453,N_947,N_600);
nand U2454 (N_2454,N_498,N_300);
and U2455 (N_2455,N_497,N_693);
and U2456 (N_2456,N_917,N_978);
nor U2457 (N_2457,N_1210,N_256);
xor U2458 (N_2458,N_755,N_1128);
nand U2459 (N_2459,N_388,N_1154);
xor U2460 (N_2460,N_1144,N_1069);
nand U2461 (N_2461,N_665,N_1128);
or U2462 (N_2462,N_700,N_863);
nand U2463 (N_2463,N_78,N_914);
nand U2464 (N_2464,N_811,N_728);
and U2465 (N_2465,N_490,N_479);
nand U2466 (N_2466,N_741,N_1243);
or U2467 (N_2467,N_298,N_62);
or U2468 (N_2468,N_1181,N_1035);
or U2469 (N_2469,N_151,N_502);
and U2470 (N_2470,N_1221,N_509);
nor U2471 (N_2471,N_513,N_524);
xor U2472 (N_2472,N_565,N_595);
or U2473 (N_2473,N_1007,N_539);
or U2474 (N_2474,N_198,N_545);
nand U2475 (N_2475,N_1136,N_691);
or U2476 (N_2476,N_870,N_772);
and U2477 (N_2477,N_1112,N_229);
nand U2478 (N_2478,N_857,N_733);
or U2479 (N_2479,N_133,N_477);
and U2480 (N_2480,N_89,N_466);
nor U2481 (N_2481,N_832,N_995);
or U2482 (N_2482,N_158,N_744);
or U2483 (N_2483,N_1218,N_955);
nand U2484 (N_2484,N_149,N_1006);
and U2485 (N_2485,N_369,N_660);
nor U2486 (N_2486,N_893,N_360);
nand U2487 (N_2487,N_630,N_464);
nand U2488 (N_2488,N_544,N_1155);
and U2489 (N_2489,N_12,N_396);
xnor U2490 (N_2490,N_217,N_618);
nand U2491 (N_2491,N_1237,N_77);
and U2492 (N_2492,N_973,N_128);
or U2493 (N_2493,N_605,N_62);
or U2494 (N_2494,N_809,N_1209);
nor U2495 (N_2495,N_636,N_651);
nor U2496 (N_2496,N_37,N_1099);
nand U2497 (N_2497,N_140,N_969);
nand U2498 (N_2498,N_855,N_888);
or U2499 (N_2499,N_132,N_205);
nor U2500 (N_2500,N_2271,N_2492);
nor U2501 (N_2501,N_1493,N_1339);
or U2502 (N_2502,N_1927,N_1417);
or U2503 (N_2503,N_1982,N_1586);
nand U2504 (N_2504,N_2222,N_1364);
xor U2505 (N_2505,N_2396,N_1450);
xor U2506 (N_2506,N_1981,N_2067);
and U2507 (N_2507,N_1592,N_2055);
and U2508 (N_2508,N_1899,N_2105);
nand U2509 (N_2509,N_1837,N_2256);
xnor U2510 (N_2510,N_2143,N_1610);
or U2511 (N_2511,N_1410,N_2434);
nor U2512 (N_2512,N_2302,N_2035);
or U2513 (N_2513,N_1535,N_1994);
nand U2514 (N_2514,N_1663,N_2157);
and U2515 (N_2515,N_1840,N_1463);
and U2516 (N_2516,N_2275,N_1928);
xnor U2517 (N_2517,N_1569,N_1383);
xor U2518 (N_2518,N_1424,N_1738);
xnor U2519 (N_2519,N_1361,N_1448);
nor U2520 (N_2520,N_1748,N_2364);
and U2521 (N_2521,N_2102,N_1851);
nand U2522 (N_2522,N_2483,N_1482);
nand U2523 (N_2523,N_1646,N_1348);
or U2524 (N_2524,N_2459,N_1501);
xor U2525 (N_2525,N_1872,N_2486);
or U2526 (N_2526,N_1370,N_1519);
or U2527 (N_2527,N_1485,N_1719);
nor U2528 (N_2528,N_1309,N_2276);
nor U2529 (N_2529,N_1280,N_2120);
and U2530 (N_2530,N_1733,N_1722);
nand U2531 (N_2531,N_2285,N_2006);
nor U2532 (N_2532,N_1439,N_1785);
nor U2533 (N_2533,N_1651,N_1895);
or U2534 (N_2534,N_1746,N_1911);
nor U2535 (N_2535,N_2262,N_1403);
or U2536 (N_2536,N_1843,N_1784);
xor U2537 (N_2537,N_2401,N_1910);
xnor U2538 (N_2538,N_2233,N_2382);
xor U2539 (N_2539,N_2479,N_1452);
nor U2540 (N_2540,N_2404,N_2321);
or U2541 (N_2541,N_1625,N_1422);
nor U2542 (N_2542,N_1588,N_1270);
and U2543 (N_2543,N_1741,N_1734);
xor U2544 (N_2544,N_2489,N_1347);
nor U2545 (N_2545,N_2188,N_2448);
or U2546 (N_2546,N_2130,N_2100);
and U2547 (N_2547,N_1654,N_2094);
nor U2548 (N_2548,N_1430,N_2183);
or U2549 (N_2549,N_2449,N_2037);
nor U2550 (N_2550,N_1930,N_2219);
and U2551 (N_2551,N_1838,N_2047);
nand U2552 (N_2552,N_1626,N_2447);
xor U2553 (N_2553,N_2238,N_1753);
nand U2554 (N_2554,N_2474,N_1555);
xnor U2555 (N_2555,N_1299,N_1560);
nand U2556 (N_2556,N_1466,N_2078);
xnor U2557 (N_2557,N_1562,N_1769);
xor U2558 (N_2558,N_1997,N_1526);
nor U2559 (N_2559,N_1708,N_1804);
nand U2560 (N_2560,N_1267,N_2169);
xnor U2561 (N_2561,N_1629,N_1864);
nand U2562 (N_2562,N_1916,N_2433);
nand U2563 (N_2563,N_2394,N_2427);
nor U2564 (N_2564,N_1867,N_1824);
nor U2565 (N_2565,N_1389,N_1894);
or U2566 (N_2566,N_2191,N_2012);
xnor U2567 (N_2567,N_2263,N_1632);
nand U2568 (N_2568,N_1844,N_2186);
nand U2569 (N_2569,N_2024,N_1496);
xnor U2570 (N_2570,N_1488,N_2494);
nand U2571 (N_2571,N_2088,N_2354);
nor U2572 (N_2572,N_2310,N_2019);
and U2573 (N_2573,N_1814,N_2407);
nor U2574 (N_2574,N_2206,N_2337);
and U2575 (N_2575,N_1454,N_1457);
and U2576 (N_2576,N_2054,N_2172);
and U2577 (N_2577,N_1468,N_1856);
xor U2578 (N_2578,N_1316,N_2368);
xnor U2579 (N_2579,N_1464,N_2171);
nor U2580 (N_2580,N_1480,N_1405);
and U2581 (N_2581,N_1805,N_1566);
or U2582 (N_2582,N_1882,N_1504);
xor U2583 (N_2583,N_1444,N_1685);
nor U2584 (N_2584,N_2229,N_1888);
or U2585 (N_2585,N_1436,N_2356);
or U2586 (N_2586,N_1344,N_1826);
and U2587 (N_2587,N_1371,N_1794);
or U2588 (N_2588,N_1724,N_2376);
and U2589 (N_2589,N_1530,N_1789);
xnor U2590 (N_2590,N_1877,N_1338);
nand U2591 (N_2591,N_1540,N_2180);
or U2592 (N_2592,N_1681,N_1590);
nor U2593 (N_2593,N_2274,N_1413);
or U2594 (N_2594,N_2334,N_1622);
and U2595 (N_2595,N_2412,N_2464);
and U2596 (N_2596,N_2190,N_2252);
and U2597 (N_2597,N_1357,N_1977);
and U2598 (N_2598,N_1326,N_1500);
or U2599 (N_2599,N_1711,N_1884);
and U2600 (N_2600,N_1492,N_2142);
and U2601 (N_2601,N_2264,N_1743);
nand U2602 (N_2602,N_2410,N_1905);
xor U2603 (N_2603,N_1949,N_1935);
xor U2604 (N_2604,N_1760,N_1752);
nand U2605 (N_2605,N_1284,N_1435);
xor U2606 (N_2606,N_2445,N_2214);
or U2607 (N_2607,N_1505,N_2371);
xnor U2608 (N_2608,N_2456,N_2198);
or U2609 (N_2609,N_1281,N_1489);
xnor U2610 (N_2610,N_2195,N_2383);
and U2611 (N_2611,N_1858,N_1516);
nor U2612 (N_2612,N_1276,N_2452);
and U2613 (N_2613,N_1465,N_2044);
nor U2614 (N_2614,N_1534,N_1809);
and U2615 (N_2615,N_2081,N_1922);
xnor U2616 (N_2616,N_1635,N_2090);
xor U2617 (N_2617,N_2493,N_1472);
and U2618 (N_2618,N_2418,N_2341);
or U2619 (N_2619,N_2103,N_1958);
and U2620 (N_2620,N_1307,N_1513);
nor U2621 (N_2621,N_1664,N_1407);
nor U2622 (N_2622,N_2478,N_1522);
nor U2623 (N_2623,N_2490,N_2319);
and U2624 (N_2624,N_1261,N_2287);
nor U2625 (N_2625,N_2423,N_2064);
and U2626 (N_2626,N_2065,N_1503);
nand U2627 (N_2627,N_2358,N_2138);
xor U2628 (N_2628,N_2387,N_1589);
nand U2629 (N_2629,N_2351,N_2283);
nand U2630 (N_2630,N_1971,N_1721);
nand U2631 (N_2631,N_2428,N_2060);
nor U2632 (N_2632,N_2329,N_1449);
or U2633 (N_2633,N_1815,N_2080);
and U2634 (N_2634,N_1510,N_2053);
nor U2635 (N_2635,N_1412,N_1476);
nand U2636 (N_2636,N_2436,N_2288);
nor U2637 (N_2637,N_1668,N_1486);
nand U2638 (N_2638,N_1375,N_1974);
nor U2639 (N_2639,N_2286,N_2061);
nor U2640 (N_2640,N_2314,N_2442);
or U2641 (N_2641,N_1661,N_1718);
nor U2642 (N_2642,N_2259,N_1559);
and U2643 (N_2643,N_2361,N_2204);
or U2644 (N_2644,N_1282,N_1553);
and U2645 (N_2645,N_2462,N_1937);
and U2646 (N_2646,N_1717,N_1710);
xnor U2647 (N_2647,N_2279,N_1986);
xnor U2648 (N_2648,N_1447,N_2008);
nand U2649 (N_2649,N_1907,N_2201);
xor U2650 (N_2650,N_2251,N_1859);
xor U2651 (N_2651,N_1742,N_1541);
and U2652 (N_2652,N_1292,N_1332);
nor U2653 (N_2653,N_2218,N_1366);
nand U2654 (N_2654,N_1764,N_2059);
nand U2655 (N_2655,N_1690,N_1965);
nor U2656 (N_2656,N_1659,N_1387);
nor U2657 (N_2657,N_1873,N_1356);
xor U2658 (N_2658,N_2117,N_2374);
xor U2659 (N_2659,N_1470,N_1933);
nor U2660 (N_2660,N_1293,N_1613);
nand U2661 (N_2661,N_1484,N_2466);
or U2662 (N_2662,N_2197,N_1490);
nor U2663 (N_2663,N_2125,N_1446);
nor U2664 (N_2664,N_1720,N_2317);
xor U2665 (N_2665,N_2231,N_2146);
xnor U2666 (N_2666,N_2224,N_2458);
xnor U2667 (N_2667,N_1919,N_1451);
or U2668 (N_2668,N_1539,N_1641);
or U2669 (N_2669,N_1567,N_2200);
or U2670 (N_2670,N_2236,N_1689);
or U2671 (N_2671,N_1517,N_1341);
xnor U2672 (N_2672,N_1266,N_1970);
xnor U2673 (N_2673,N_1653,N_2017);
or U2674 (N_2674,N_1429,N_1543);
nand U2675 (N_2675,N_1991,N_1702);
nor U2676 (N_2676,N_2071,N_1487);
and U2677 (N_2677,N_1973,N_2301);
or U2678 (N_2678,N_2069,N_1716);
and U2679 (N_2679,N_2097,N_1481);
nor U2680 (N_2680,N_1264,N_2042);
and U2681 (N_2681,N_2380,N_2293);
nand U2682 (N_2682,N_2184,N_1739);
and U2683 (N_2683,N_1331,N_2431);
xor U2684 (N_2684,N_1850,N_2232);
xor U2685 (N_2685,N_2384,N_2444);
or U2686 (N_2686,N_1315,N_2223);
or U2687 (N_2687,N_2048,N_2257);
or U2688 (N_2688,N_1333,N_1509);
nor U2689 (N_2689,N_1999,N_2073);
and U2690 (N_2690,N_1478,N_1912);
nand U2691 (N_2691,N_2349,N_1950);
or U2692 (N_2692,N_2179,N_2093);
and U2693 (N_2693,N_1833,N_2284);
nor U2694 (N_2694,N_1790,N_2476);
and U2695 (N_2695,N_2306,N_2497);
nor U2696 (N_2696,N_1817,N_1640);
nand U2697 (N_2697,N_1442,N_1458);
nor U2698 (N_2698,N_1308,N_2312);
and U2699 (N_2699,N_1631,N_1799);
or U2700 (N_2700,N_1952,N_1425);
or U2701 (N_2701,N_1497,N_1797);
nor U2702 (N_2702,N_1875,N_1976);
nand U2703 (N_2703,N_2254,N_1707);
nor U2704 (N_2704,N_2429,N_2268);
or U2705 (N_2705,N_2115,N_1418);
xnor U2706 (N_2706,N_1749,N_1964);
nor U2707 (N_2707,N_1432,N_2114);
xnor U2708 (N_2708,N_2424,N_1732);
or U2709 (N_2709,N_2496,N_1940);
and U2710 (N_2710,N_1754,N_2432);
and U2711 (N_2711,N_2481,N_1575);
or U2712 (N_2712,N_2303,N_2104);
nor U2713 (N_2713,N_2239,N_2499);
and U2714 (N_2714,N_1511,N_1772);
xor U2715 (N_2715,N_1993,N_1337);
and U2716 (N_2716,N_2352,N_1944);
and U2717 (N_2717,N_2324,N_1820);
xnor U2718 (N_2718,N_1812,N_1343);
nand U2719 (N_2719,N_2468,N_2249);
nand U2720 (N_2720,N_2402,N_1830);
xor U2721 (N_2721,N_2075,N_2007);
or U2722 (N_2722,N_2193,N_1252);
and U2723 (N_2723,N_1459,N_1419);
nor U2724 (N_2724,N_2336,N_1876);
nand U2725 (N_2725,N_1818,N_1796);
nor U2726 (N_2726,N_2145,N_2126);
and U2727 (N_2727,N_1474,N_2397);
or U2728 (N_2728,N_1453,N_1305);
xnor U2729 (N_2729,N_2426,N_2350);
and U2730 (N_2730,N_2137,N_1946);
nand U2731 (N_2731,N_2482,N_2182);
or U2732 (N_2732,N_1967,N_1355);
or U2733 (N_2733,N_1440,N_2261);
or U2734 (N_2734,N_1395,N_1892);
nor U2735 (N_2735,N_2241,N_1521);
xor U2736 (N_2736,N_1615,N_2129);
or U2737 (N_2737,N_1584,N_1639);
nand U2738 (N_2738,N_1393,N_2414);
and U2739 (N_2739,N_2029,N_1525);
or U2740 (N_2740,N_2021,N_1595);
nand U2741 (N_2741,N_1855,N_2139);
nand U2742 (N_2742,N_2398,N_1406);
xor U2743 (N_2743,N_1268,N_2020);
or U2744 (N_2744,N_1839,N_1520);
or U2745 (N_2745,N_1620,N_2074);
xor U2746 (N_2746,N_1834,N_1726);
nand U2747 (N_2747,N_1396,N_1887);
and U2748 (N_2748,N_1673,N_2152);
nor U2749 (N_2749,N_1776,N_1670);
or U2750 (N_2750,N_1862,N_2144);
nor U2751 (N_2751,N_2422,N_1909);
and U2752 (N_2752,N_1686,N_2471);
or U2753 (N_2753,N_1897,N_2298);
nor U2754 (N_2754,N_2392,N_1628);
xnor U2755 (N_2755,N_2247,N_2485);
nor U2756 (N_2756,N_2066,N_2149);
nor U2757 (N_2757,N_1400,N_1706);
and U2758 (N_2758,N_1302,N_2101);
and U2759 (N_2759,N_1598,N_1599);
or U2760 (N_2760,N_1379,N_1531);
xor U2761 (N_2761,N_2122,N_2216);
or U2762 (N_2762,N_1787,N_1295);
xor U2763 (N_2763,N_1901,N_1806);
nand U2764 (N_2764,N_2208,N_1587);
xor U2765 (N_2765,N_2211,N_1391);
nand U2766 (N_2766,N_1811,N_2416);
nand U2767 (N_2767,N_2016,N_2000);
xnor U2768 (N_2768,N_2209,N_1680);
nand U2769 (N_2769,N_1903,N_1652);
or U2770 (N_2770,N_1788,N_2281);
nand U2771 (N_2771,N_1258,N_1617);
xnor U2772 (N_2772,N_2375,N_1325);
nand U2773 (N_2773,N_1989,N_1832);
nand U2774 (N_2774,N_2457,N_2153);
xnor U2775 (N_2775,N_1498,N_1883);
xor U2776 (N_2776,N_2199,N_1401);
and U2777 (N_2777,N_1829,N_2168);
nand U2778 (N_2778,N_2187,N_1607);
nor U2779 (N_2779,N_1385,N_1995);
nor U2780 (N_2780,N_1947,N_1512);
or U2781 (N_2781,N_1358,N_2202);
nor U2782 (N_2782,N_1849,N_2467);
and U2783 (N_2783,N_1398,N_1262);
or U2784 (N_2784,N_2379,N_1462);
and U2785 (N_2785,N_2049,N_2320);
or U2786 (N_2786,N_1318,N_1761);
and U2787 (N_2787,N_2366,N_1938);
or U2788 (N_2788,N_2015,N_1951);
nand U2789 (N_2789,N_1624,N_1715);
nor U2790 (N_2790,N_2127,N_1255);
nand U2791 (N_2791,N_1775,N_1762);
and U2792 (N_2792,N_1612,N_2309);
or U2793 (N_2793,N_1314,N_2443);
and U2794 (N_2794,N_1957,N_1421);
and U2795 (N_2795,N_2041,N_2141);
and U2796 (N_2796,N_2226,N_2308);
nand U2797 (N_2797,N_2230,N_1700);
nand U2798 (N_2798,N_2253,N_1479);
nor U2799 (N_2799,N_2296,N_1920);
or U2800 (N_2800,N_2420,N_1848);
nor U2801 (N_2801,N_1692,N_2435);
and U2802 (N_2802,N_1552,N_1536);
xnor U2803 (N_2803,N_1253,N_1735);
or U2804 (N_2804,N_1979,N_2217);
nor U2805 (N_2805,N_1955,N_1869);
and U2806 (N_2806,N_2194,N_1751);
nand U2807 (N_2807,N_1745,N_1545);
nand U2808 (N_2808,N_1320,N_1913);
and U2809 (N_2809,N_1825,N_2390);
nand U2810 (N_2810,N_2151,N_2450);
and U2811 (N_2811,N_1380,N_1507);
and U2812 (N_2812,N_1256,N_1729);
and U2813 (N_2813,N_2134,N_2480);
and U2814 (N_2814,N_2313,N_2096);
nor U2815 (N_2815,N_1771,N_1564);
nor U2816 (N_2816,N_1382,N_2235);
and U2817 (N_2817,N_2234,N_2108);
and U2818 (N_2818,N_1286,N_2132);
or U2819 (N_2819,N_2070,N_1257);
or U2820 (N_2820,N_1345,N_2357);
xor U2821 (N_2821,N_1572,N_2340);
xnor U2822 (N_2822,N_2419,N_2272);
xor U2823 (N_2823,N_1687,N_1898);
or U2824 (N_2824,N_2353,N_1455);
nor U2825 (N_2825,N_1727,N_1397);
or U2826 (N_2826,N_1696,N_2393);
nand U2827 (N_2827,N_2189,N_1388);
and U2828 (N_2828,N_1603,N_1576);
nor U2829 (N_2829,N_1889,N_1853);
xor U2830 (N_2830,N_2203,N_2058);
or U2831 (N_2831,N_2348,N_2136);
or U2832 (N_2832,N_2381,N_1565);
and U2833 (N_2833,N_2124,N_1791);
xor U2834 (N_2834,N_2322,N_2086);
or U2835 (N_2835,N_1346,N_1568);
and U2836 (N_2836,N_1983,N_1968);
nand U2837 (N_2837,N_2470,N_2491);
nor U2838 (N_2838,N_1638,N_2386);
nand U2839 (N_2839,N_2297,N_1585);
nand U2840 (N_2840,N_2242,N_1334);
xor U2841 (N_2841,N_1596,N_2291);
nand U2842 (N_2842,N_1533,N_1778);
nor U2843 (N_2843,N_2119,N_1304);
nand U2844 (N_2844,N_2027,N_1277);
xnor U2845 (N_2845,N_2110,N_2460);
xor U2846 (N_2846,N_2477,N_2250);
and U2847 (N_2847,N_2159,N_2451);
xor U2848 (N_2848,N_1780,N_1942);
or U2849 (N_2849,N_1987,N_1621);
and U2850 (N_2850,N_1381,N_2292);
and U2851 (N_2851,N_2295,N_1538);
nand U2852 (N_2852,N_1998,N_1409);
nand U2853 (N_2853,N_1688,N_2328);
or U2854 (N_2854,N_2116,N_2043);
xnor U2855 (N_2855,N_2395,N_2181);
nand U2856 (N_2856,N_1527,N_1312);
nor U2857 (N_2857,N_2161,N_1808);
xnor U2858 (N_2858,N_2107,N_1684);
nand U2859 (N_2859,N_1701,N_1656);
or U2860 (N_2860,N_1428,N_1354);
nor U2861 (N_2861,N_1363,N_2207);
nor U2862 (N_2862,N_1943,N_1868);
nand U2863 (N_2863,N_1573,N_2372);
and U2864 (N_2864,N_2326,N_1475);
or U2865 (N_2865,N_1313,N_1969);
nor U2866 (N_2866,N_2221,N_2360);
and U2867 (N_2867,N_2140,N_1609);
and U2868 (N_2868,N_1551,N_1269);
nand U2869 (N_2869,N_1777,N_2245);
nand U2870 (N_2870,N_2373,N_1703);
xnor U2871 (N_2871,N_2098,N_1644);
nand U2872 (N_2872,N_2365,N_2031);
xor U2873 (N_2873,N_1386,N_1443);
nor U2874 (N_2874,N_1298,N_1714);
and U2875 (N_2875,N_1583,N_1349);
or U2876 (N_2876,N_2083,N_2213);
or U2877 (N_2877,N_2004,N_2025);
xnor U2878 (N_2878,N_2430,N_1931);
nand U2879 (N_2879,N_1317,N_1423);
nand U2880 (N_2880,N_1956,N_2359);
or U2881 (N_2881,N_1941,N_2258);
xnor U2882 (N_2882,N_1768,N_1272);
or U2883 (N_2883,N_2441,N_1779);
nand U2884 (N_2884,N_1633,N_1373);
nand U2885 (N_2885,N_1630,N_1767);
or U2886 (N_2886,N_2363,N_1279);
and U2887 (N_2887,N_2391,N_2331);
or U2888 (N_2888,N_1992,N_1939);
nand U2889 (N_2889,N_2023,N_1636);
or U2890 (N_2890,N_1737,N_2463);
or U2891 (N_2891,N_2333,N_1427);
nand U2892 (N_2892,N_1846,N_1795);
nor U2893 (N_2893,N_1563,N_1394);
or U2894 (N_2894,N_1571,N_2278);
nor U2895 (N_2895,N_2346,N_2323);
xor U2896 (N_2896,N_2370,N_1554);
or U2897 (N_2897,N_1274,N_1669);
nand U2898 (N_2898,N_1693,N_1766);
nand U2899 (N_2899,N_2033,N_2417);
nor U2900 (N_2900,N_2192,N_1792);
nand U2901 (N_2901,N_1860,N_2014);
xnor U2902 (N_2902,N_1329,N_2316);
xor U2903 (N_2903,N_1880,N_1683);
and U2904 (N_2904,N_1763,N_1891);
xnor U2905 (N_2905,N_1723,N_2269);
nand U2906 (N_2906,N_2454,N_1866);
xor U2907 (N_2907,N_1863,N_2210);
and U2908 (N_2908,N_1619,N_2248);
xor U2909 (N_2909,N_2332,N_2032);
nor U2910 (N_2910,N_1736,N_1996);
nor U2911 (N_2911,N_2050,N_1813);
nor U2912 (N_2912,N_1441,N_1606);
and U2913 (N_2913,N_1390,N_1783);
and U2914 (N_2914,N_1985,N_2040);
xnor U2915 (N_2915,N_2406,N_2009);
nor U2916 (N_2916,N_2133,N_1376);
nand U2917 (N_2917,N_1713,N_1649);
nor U2918 (N_2918,N_1301,N_1709);
xnor U2919 (N_2919,N_1691,N_2068);
xnor U2920 (N_2920,N_1600,N_2131);
nor U2921 (N_2921,N_1961,N_2212);
xnor U2922 (N_2922,N_2164,N_2165);
and U2923 (N_2923,N_1959,N_2160);
nand U2924 (N_2924,N_1467,N_1650);
nor U2925 (N_2925,N_1904,N_1984);
and U2926 (N_2926,N_1506,N_1353);
or U2927 (N_2927,N_2087,N_1878);
xor U2928 (N_2928,N_1962,N_1285);
or U2929 (N_2929,N_1885,N_2439);
and U2930 (N_2930,N_1283,N_1915);
nor U2931 (N_2931,N_1291,N_1637);
xor U2932 (N_2932,N_1537,N_2369);
nand U2933 (N_2933,N_2495,N_1288);
or U2934 (N_2934,N_1990,N_2228);
nor U2935 (N_2935,N_2091,N_1327);
or U2936 (N_2936,N_2438,N_2342);
xnor U2937 (N_2937,N_1408,N_1948);
or U2938 (N_2938,N_1578,N_1765);
xnor U2939 (N_2939,N_1874,N_1697);
nand U2940 (N_2940,N_2469,N_2196);
or U2941 (N_2941,N_1529,N_1558);
or U2942 (N_2942,N_1582,N_1359);
or U2943 (N_2943,N_1456,N_1518);
xor U2944 (N_2944,N_2166,N_1870);
xnor U2945 (N_2945,N_1900,N_1415);
nor U2946 (N_2946,N_1917,N_2112);
xnor U2947 (N_2947,N_2367,N_2325);
nand U2948 (N_2948,N_1647,N_2150);
nor U2949 (N_2949,N_2280,N_2282);
nor U2950 (N_2950,N_2255,N_1665);
and U2951 (N_2951,N_1340,N_1960);
xnor U2952 (N_2952,N_1671,N_1695);
nor U2953 (N_2953,N_2355,N_2002);
nor U2954 (N_2954,N_1823,N_2076);
xnor U2955 (N_2955,N_1438,N_2175);
nor U2956 (N_2956,N_2244,N_1774);
nand U2957 (N_2957,N_2085,N_1557);
nand U2958 (N_2958,N_1740,N_1667);
nor U2959 (N_2959,N_2425,N_1499);
and U2960 (N_2960,N_2154,N_2178);
nor U2961 (N_2961,N_1618,N_1932);
nand U2962 (N_2962,N_1259,N_1434);
and U2963 (N_2963,N_1845,N_1835);
nand U2964 (N_2964,N_1893,N_2267);
nor U2965 (N_2965,N_1294,N_1360);
or U2966 (N_2966,N_1857,N_1678);
nand U2967 (N_2967,N_2289,N_1581);
xnor U2968 (N_2968,N_1827,N_1750);
nand U2969 (N_2969,N_2300,N_2378);
xor U2970 (N_2970,N_1321,N_1819);
or U2971 (N_2971,N_2005,N_2155);
nor U2972 (N_2972,N_1471,N_2270);
xnor U2973 (N_2973,N_2413,N_2177);
nand U2974 (N_2974,N_2162,N_1297);
and U2975 (N_2975,N_1542,N_2345);
and U2976 (N_2976,N_1336,N_1728);
xor U2977 (N_2977,N_2487,N_1648);
xnor U2978 (N_2978,N_2089,N_2484);
xor U2979 (N_2979,N_1275,N_1374);
xor U2980 (N_2980,N_2079,N_1495);
and U2981 (N_2981,N_1828,N_1660);
and U2982 (N_2982,N_1523,N_1793);
nand U2983 (N_2983,N_2400,N_2294);
or U2984 (N_2984,N_1679,N_1923);
and U2985 (N_2985,N_2311,N_1437);
or U2986 (N_2986,N_1682,N_2176);
or U2987 (N_2987,N_2273,N_1954);
or U2988 (N_2988,N_1861,N_2028);
xnor U2989 (N_2989,N_2227,N_1342);
or U2990 (N_2990,N_1263,N_1924);
and U2991 (N_2991,N_1906,N_1594);
or U2992 (N_2992,N_1676,N_1770);
nand U2993 (N_2993,N_1747,N_1514);
and U2994 (N_2994,N_2389,N_2039);
or U2995 (N_2995,N_2385,N_1287);
and U2996 (N_2996,N_1841,N_2163);
nor U2997 (N_2997,N_1515,N_1271);
or U2998 (N_2998,N_1879,N_1335);
or U2999 (N_2999,N_1367,N_2220);
nand U3000 (N_3000,N_2018,N_1929);
nor U3001 (N_3001,N_1755,N_2299);
nand U3002 (N_3002,N_1890,N_1972);
nor U3003 (N_3003,N_2453,N_2052);
and U3004 (N_3004,N_1577,N_1416);
and U3005 (N_3005,N_1250,N_2243);
nor U3006 (N_3006,N_2318,N_1978);
xor U3007 (N_3007,N_2135,N_2265);
nand U3008 (N_3008,N_1579,N_1550);
nor U3009 (N_3009,N_2147,N_1601);
or U3010 (N_3010,N_1324,N_2240);
nor U3011 (N_3011,N_2148,N_2465);
nor U3012 (N_3012,N_1953,N_1556);
xnor U3013 (N_3013,N_1494,N_2315);
and U3014 (N_3014,N_2305,N_2022);
and U3015 (N_3015,N_2062,N_1608);
nor U3016 (N_3016,N_2158,N_2030);
nor U3017 (N_3017,N_1362,N_1402);
nand U3018 (N_3018,N_1368,N_1756);
nor U3019 (N_3019,N_2330,N_2038);
or U3020 (N_3020,N_1426,N_2082);
xnor U3021 (N_3021,N_1807,N_1311);
nor U3022 (N_3022,N_1548,N_1936);
nand U3023 (N_3023,N_1674,N_2405);
or U3024 (N_3024,N_2335,N_1886);
and U3025 (N_3025,N_1921,N_1328);
and U3026 (N_3026,N_2377,N_1782);
or U3027 (N_3027,N_1758,N_2290);
xnor U3028 (N_3028,N_1300,N_2246);
or U3029 (N_3029,N_2347,N_2121);
xnor U3030 (N_3030,N_1604,N_1645);
nand U3031 (N_3031,N_1698,N_2167);
or U3032 (N_3032,N_1963,N_2113);
nor U3033 (N_3033,N_2170,N_1384);
xor U3034 (N_3034,N_2304,N_2225);
and U3035 (N_3035,N_2063,N_2266);
or U3036 (N_3036,N_2409,N_1699);
xor U3037 (N_3037,N_1433,N_2475);
xnor U3038 (N_3038,N_1546,N_2498);
nand U3039 (N_3039,N_1303,N_2421);
or U3040 (N_3040,N_2446,N_1549);
and U3041 (N_3041,N_1842,N_1365);
or U3042 (N_3042,N_1642,N_1854);
xor U3043 (N_3043,N_1675,N_1593);
and U3044 (N_3044,N_1980,N_1574);
nand U3045 (N_3045,N_1672,N_1975);
xor U3046 (N_3046,N_1802,N_2077);
nor U3047 (N_3047,N_1881,N_1810);
or U3048 (N_3048,N_1508,N_1352);
nand U3049 (N_3049,N_1290,N_1580);
nor U3050 (N_3050,N_1934,N_1966);
nor U3051 (N_3051,N_1865,N_1605);
nor U3052 (N_3052,N_1420,N_1836);
or U3053 (N_3053,N_2339,N_2307);
and U3054 (N_3054,N_1847,N_1323);
nand U3055 (N_3055,N_1296,N_1306);
xnor U3056 (N_3056,N_1945,N_2118);
or U3057 (N_3057,N_2034,N_1896);
xnor U3058 (N_3058,N_2488,N_1908);
and U3059 (N_3059,N_1616,N_1591);
or U3060 (N_3060,N_1623,N_1460);
xor U3061 (N_3061,N_2099,N_2440);
nand U3062 (N_3062,N_1871,N_2026);
nand U3063 (N_3063,N_1431,N_1657);
nor U3064 (N_3064,N_1547,N_1491);
and U3065 (N_3065,N_1319,N_1781);
or U3066 (N_3066,N_1289,N_2215);
nand U3067 (N_3067,N_1597,N_1677);
nor U3068 (N_3068,N_2072,N_1798);
xor U3069 (N_3069,N_2473,N_1643);
nor U3070 (N_3070,N_1445,N_1658);
xor U3071 (N_3071,N_1528,N_2277);
xor U3072 (N_3072,N_2092,N_1614);
nand U3073 (N_3073,N_1655,N_1351);
nor U3074 (N_3074,N_1254,N_1666);
xor U3075 (N_3075,N_2011,N_1852);
nor U3076 (N_3076,N_1322,N_1602);
or U3077 (N_3077,N_2472,N_1473);
nand U3078 (N_3078,N_1372,N_2109);
xnor U3079 (N_3079,N_1634,N_1712);
nand U3080 (N_3080,N_2403,N_2260);
xnor U3081 (N_3081,N_1786,N_2205);
nand U3082 (N_3082,N_2051,N_2237);
nand U3083 (N_3083,N_1611,N_2399);
nand U3084 (N_3084,N_1759,N_1399);
and U3085 (N_3085,N_2344,N_1705);
or U3086 (N_3086,N_1725,N_1404);
and U3087 (N_3087,N_2362,N_2327);
and U3088 (N_3088,N_2036,N_2461);
xor U3089 (N_3089,N_2095,N_1544);
and U3090 (N_3090,N_1524,N_1821);
xor U3091 (N_3091,N_2415,N_1744);
or U3092 (N_3092,N_2056,N_1730);
and U3093 (N_3093,N_1627,N_1662);
nand U3094 (N_3094,N_2388,N_2106);
or U3095 (N_3095,N_1532,N_1925);
xor U3096 (N_3096,N_1251,N_1988);
nand U3097 (N_3097,N_1469,N_2123);
nor U3098 (N_3098,N_1831,N_1273);
or U3099 (N_3099,N_1731,N_2411);
xnor U3100 (N_3100,N_1570,N_1803);
xnor U3101 (N_3101,N_2174,N_2185);
nor U3102 (N_3102,N_2338,N_1502);
nand U3103 (N_3103,N_2128,N_2455);
and U3104 (N_3104,N_1914,N_1561);
nor U3105 (N_3105,N_2084,N_1801);
and U3106 (N_3106,N_1392,N_1926);
or U3107 (N_3107,N_2408,N_1260);
xor U3108 (N_3108,N_1378,N_1369);
nand U3109 (N_3109,N_1310,N_1822);
nor U3110 (N_3110,N_1461,N_1483);
and U3111 (N_3111,N_2046,N_1414);
or U3112 (N_3112,N_1773,N_1278);
or U3113 (N_3113,N_1694,N_2003);
and U3114 (N_3114,N_1330,N_2001);
nand U3115 (N_3115,N_2111,N_1918);
nor U3116 (N_3116,N_2173,N_1411);
and U3117 (N_3117,N_2437,N_1477);
or U3118 (N_3118,N_2013,N_2343);
or U3119 (N_3119,N_1704,N_1902);
nand U3120 (N_3120,N_1816,N_1757);
or U3121 (N_3121,N_2057,N_2045);
xor U3122 (N_3122,N_1800,N_1350);
and U3123 (N_3123,N_2010,N_2156);
xor U3124 (N_3124,N_1377,N_1265);
nand U3125 (N_3125,N_2042,N_2408);
nor U3126 (N_3126,N_1496,N_2337);
and U3127 (N_3127,N_1429,N_1520);
or U3128 (N_3128,N_1498,N_2310);
nand U3129 (N_3129,N_1773,N_1435);
nor U3130 (N_3130,N_1510,N_1477);
nor U3131 (N_3131,N_1441,N_2254);
nand U3132 (N_3132,N_2118,N_2212);
nand U3133 (N_3133,N_2321,N_1481);
and U3134 (N_3134,N_2243,N_1924);
xor U3135 (N_3135,N_1373,N_1974);
or U3136 (N_3136,N_2450,N_2399);
nand U3137 (N_3137,N_1321,N_1871);
nand U3138 (N_3138,N_2471,N_1350);
or U3139 (N_3139,N_1953,N_1840);
nand U3140 (N_3140,N_2169,N_1699);
or U3141 (N_3141,N_1919,N_2297);
and U3142 (N_3142,N_2273,N_2132);
xnor U3143 (N_3143,N_1927,N_2351);
nand U3144 (N_3144,N_1649,N_2405);
nand U3145 (N_3145,N_2065,N_2351);
xnor U3146 (N_3146,N_2317,N_1446);
or U3147 (N_3147,N_1762,N_2417);
or U3148 (N_3148,N_2064,N_2241);
nor U3149 (N_3149,N_1927,N_1810);
nor U3150 (N_3150,N_1346,N_1838);
or U3151 (N_3151,N_1421,N_1476);
nor U3152 (N_3152,N_1810,N_2065);
or U3153 (N_3153,N_2177,N_1607);
nor U3154 (N_3154,N_2136,N_2417);
or U3155 (N_3155,N_2484,N_2103);
nor U3156 (N_3156,N_1616,N_2269);
nor U3157 (N_3157,N_1929,N_1761);
or U3158 (N_3158,N_2464,N_1799);
and U3159 (N_3159,N_2147,N_1435);
xnor U3160 (N_3160,N_1462,N_2253);
xor U3161 (N_3161,N_2229,N_1607);
nor U3162 (N_3162,N_1423,N_1267);
or U3163 (N_3163,N_2343,N_1474);
or U3164 (N_3164,N_2420,N_1322);
and U3165 (N_3165,N_1722,N_1462);
and U3166 (N_3166,N_2150,N_1557);
nand U3167 (N_3167,N_1836,N_1940);
and U3168 (N_3168,N_2065,N_1251);
nand U3169 (N_3169,N_2025,N_1593);
xnor U3170 (N_3170,N_1707,N_2114);
nand U3171 (N_3171,N_1501,N_1333);
nor U3172 (N_3172,N_1617,N_1432);
nor U3173 (N_3173,N_2216,N_1862);
xnor U3174 (N_3174,N_2004,N_1414);
and U3175 (N_3175,N_1477,N_1698);
or U3176 (N_3176,N_1775,N_2150);
nand U3177 (N_3177,N_1704,N_1734);
and U3178 (N_3178,N_1848,N_1594);
or U3179 (N_3179,N_2204,N_1459);
nor U3180 (N_3180,N_2412,N_1442);
and U3181 (N_3181,N_1571,N_1858);
and U3182 (N_3182,N_2151,N_1487);
or U3183 (N_3183,N_2085,N_2030);
and U3184 (N_3184,N_1532,N_2498);
nand U3185 (N_3185,N_2403,N_2458);
and U3186 (N_3186,N_2015,N_1803);
nor U3187 (N_3187,N_2158,N_1287);
and U3188 (N_3188,N_1789,N_2178);
or U3189 (N_3189,N_1442,N_2431);
xnor U3190 (N_3190,N_1428,N_1491);
nand U3191 (N_3191,N_1528,N_1775);
nand U3192 (N_3192,N_2310,N_2391);
xnor U3193 (N_3193,N_2340,N_1457);
or U3194 (N_3194,N_1555,N_1421);
xnor U3195 (N_3195,N_2081,N_1362);
or U3196 (N_3196,N_1790,N_1970);
nor U3197 (N_3197,N_1292,N_2404);
nor U3198 (N_3198,N_1642,N_1941);
nand U3199 (N_3199,N_2394,N_2498);
or U3200 (N_3200,N_2368,N_2259);
and U3201 (N_3201,N_1375,N_2273);
nor U3202 (N_3202,N_2273,N_1903);
and U3203 (N_3203,N_1998,N_1524);
or U3204 (N_3204,N_2112,N_1814);
xor U3205 (N_3205,N_2019,N_1650);
nor U3206 (N_3206,N_1350,N_1804);
and U3207 (N_3207,N_2436,N_2367);
nand U3208 (N_3208,N_1344,N_1943);
and U3209 (N_3209,N_2186,N_1552);
and U3210 (N_3210,N_1601,N_1615);
and U3211 (N_3211,N_1502,N_1974);
and U3212 (N_3212,N_1778,N_1780);
nor U3213 (N_3213,N_1898,N_1631);
nor U3214 (N_3214,N_2459,N_1739);
xnor U3215 (N_3215,N_1577,N_2229);
xor U3216 (N_3216,N_1534,N_1887);
or U3217 (N_3217,N_1262,N_2189);
nor U3218 (N_3218,N_2391,N_2368);
xor U3219 (N_3219,N_2014,N_2330);
nand U3220 (N_3220,N_1297,N_1491);
xor U3221 (N_3221,N_1509,N_1950);
and U3222 (N_3222,N_1724,N_1531);
and U3223 (N_3223,N_2221,N_1544);
nand U3224 (N_3224,N_1368,N_2008);
xor U3225 (N_3225,N_1728,N_2105);
or U3226 (N_3226,N_2413,N_1287);
nand U3227 (N_3227,N_2207,N_1398);
xnor U3228 (N_3228,N_1517,N_1724);
nand U3229 (N_3229,N_2036,N_1255);
nor U3230 (N_3230,N_1948,N_2306);
or U3231 (N_3231,N_2134,N_1720);
xnor U3232 (N_3232,N_1852,N_2235);
xor U3233 (N_3233,N_1294,N_2003);
and U3234 (N_3234,N_1436,N_1704);
nand U3235 (N_3235,N_1301,N_2250);
nor U3236 (N_3236,N_1838,N_2151);
xor U3237 (N_3237,N_1518,N_1838);
nor U3238 (N_3238,N_1311,N_1810);
xnor U3239 (N_3239,N_1520,N_2087);
xnor U3240 (N_3240,N_1852,N_2389);
nand U3241 (N_3241,N_1935,N_1993);
xnor U3242 (N_3242,N_2269,N_2128);
nand U3243 (N_3243,N_1567,N_2022);
nor U3244 (N_3244,N_1775,N_2395);
and U3245 (N_3245,N_2351,N_1621);
nor U3246 (N_3246,N_1652,N_1894);
nand U3247 (N_3247,N_2229,N_2304);
and U3248 (N_3248,N_2353,N_1526);
or U3249 (N_3249,N_1254,N_1557);
nor U3250 (N_3250,N_2118,N_1496);
or U3251 (N_3251,N_1679,N_1447);
nand U3252 (N_3252,N_2196,N_2374);
and U3253 (N_3253,N_2499,N_1290);
xnor U3254 (N_3254,N_1738,N_2225);
or U3255 (N_3255,N_1862,N_2197);
xor U3256 (N_3256,N_1978,N_2313);
nand U3257 (N_3257,N_1383,N_1462);
nor U3258 (N_3258,N_2063,N_2201);
or U3259 (N_3259,N_1369,N_2036);
or U3260 (N_3260,N_1898,N_1346);
and U3261 (N_3261,N_2492,N_2399);
or U3262 (N_3262,N_1291,N_1691);
or U3263 (N_3263,N_2311,N_2063);
xnor U3264 (N_3264,N_2082,N_1827);
xnor U3265 (N_3265,N_2383,N_2055);
xnor U3266 (N_3266,N_2364,N_1562);
xor U3267 (N_3267,N_2327,N_2283);
nor U3268 (N_3268,N_1563,N_1601);
xnor U3269 (N_3269,N_1472,N_1958);
nor U3270 (N_3270,N_1271,N_2180);
and U3271 (N_3271,N_1880,N_1279);
nand U3272 (N_3272,N_2110,N_1430);
nor U3273 (N_3273,N_1395,N_1783);
xor U3274 (N_3274,N_1853,N_2292);
nand U3275 (N_3275,N_1308,N_1557);
nor U3276 (N_3276,N_1543,N_2309);
nand U3277 (N_3277,N_2446,N_2063);
nor U3278 (N_3278,N_1929,N_2250);
nor U3279 (N_3279,N_1840,N_1575);
and U3280 (N_3280,N_2156,N_1309);
and U3281 (N_3281,N_2038,N_1716);
or U3282 (N_3282,N_1382,N_2362);
and U3283 (N_3283,N_2492,N_2268);
or U3284 (N_3284,N_1806,N_1898);
nor U3285 (N_3285,N_1443,N_1834);
nor U3286 (N_3286,N_1609,N_1955);
and U3287 (N_3287,N_2155,N_1730);
or U3288 (N_3288,N_1887,N_1441);
xor U3289 (N_3289,N_1728,N_1640);
nor U3290 (N_3290,N_2012,N_1408);
or U3291 (N_3291,N_2441,N_1301);
or U3292 (N_3292,N_1669,N_2360);
nor U3293 (N_3293,N_1592,N_1849);
nor U3294 (N_3294,N_2323,N_2324);
nor U3295 (N_3295,N_1643,N_2025);
or U3296 (N_3296,N_1857,N_2308);
xnor U3297 (N_3297,N_2176,N_1693);
nand U3298 (N_3298,N_1529,N_1640);
nor U3299 (N_3299,N_2256,N_2078);
or U3300 (N_3300,N_1522,N_1253);
nor U3301 (N_3301,N_2219,N_2320);
nor U3302 (N_3302,N_1253,N_2151);
nand U3303 (N_3303,N_1960,N_2270);
xor U3304 (N_3304,N_1990,N_1939);
nand U3305 (N_3305,N_1811,N_2205);
xor U3306 (N_3306,N_1558,N_1956);
xor U3307 (N_3307,N_2168,N_1328);
xor U3308 (N_3308,N_1687,N_2116);
and U3309 (N_3309,N_1284,N_1321);
xnor U3310 (N_3310,N_1388,N_1523);
and U3311 (N_3311,N_2075,N_1511);
or U3312 (N_3312,N_2335,N_1389);
and U3313 (N_3313,N_2175,N_2420);
and U3314 (N_3314,N_2061,N_2308);
xnor U3315 (N_3315,N_2170,N_2011);
nor U3316 (N_3316,N_2278,N_1862);
and U3317 (N_3317,N_2157,N_2198);
nor U3318 (N_3318,N_2265,N_2446);
xor U3319 (N_3319,N_2100,N_1934);
xor U3320 (N_3320,N_1839,N_1335);
nor U3321 (N_3321,N_1338,N_2324);
and U3322 (N_3322,N_1508,N_1304);
and U3323 (N_3323,N_1904,N_1497);
and U3324 (N_3324,N_1466,N_2146);
nor U3325 (N_3325,N_1819,N_1599);
and U3326 (N_3326,N_2365,N_1513);
nand U3327 (N_3327,N_2054,N_1963);
xnor U3328 (N_3328,N_1634,N_2174);
or U3329 (N_3329,N_2381,N_1315);
and U3330 (N_3330,N_1606,N_1795);
nor U3331 (N_3331,N_1613,N_2251);
nand U3332 (N_3332,N_2065,N_2486);
or U3333 (N_3333,N_1369,N_1636);
or U3334 (N_3334,N_2049,N_2035);
or U3335 (N_3335,N_1958,N_1260);
xor U3336 (N_3336,N_2284,N_1947);
or U3337 (N_3337,N_2415,N_1422);
xor U3338 (N_3338,N_1898,N_1809);
nand U3339 (N_3339,N_2150,N_1434);
nor U3340 (N_3340,N_1692,N_2470);
and U3341 (N_3341,N_1423,N_2208);
nand U3342 (N_3342,N_2025,N_2357);
nor U3343 (N_3343,N_1476,N_1835);
or U3344 (N_3344,N_2187,N_1988);
and U3345 (N_3345,N_1903,N_1841);
and U3346 (N_3346,N_1526,N_1666);
or U3347 (N_3347,N_2200,N_1685);
and U3348 (N_3348,N_1958,N_1465);
nand U3349 (N_3349,N_2298,N_2171);
and U3350 (N_3350,N_2245,N_1260);
nor U3351 (N_3351,N_1717,N_2391);
nor U3352 (N_3352,N_1326,N_2144);
xor U3353 (N_3353,N_2370,N_1358);
nand U3354 (N_3354,N_2095,N_1462);
nand U3355 (N_3355,N_2131,N_2497);
nand U3356 (N_3356,N_1784,N_2311);
xnor U3357 (N_3357,N_1897,N_1312);
xor U3358 (N_3358,N_2262,N_1480);
and U3359 (N_3359,N_1742,N_1889);
nor U3360 (N_3360,N_2333,N_1440);
nand U3361 (N_3361,N_1302,N_1378);
nand U3362 (N_3362,N_2345,N_1816);
and U3363 (N_3363,N_2213,N_1901);
or U3364 (N_3364,N_1684,N_1251);
nor U3365 (N_3365,N_2179,N_1673);
xnor U3366 (N_3366,N_2322,N_1851);
or U3367 (N_3367,N_1268,N_1684);
and U3368 (N_3368,N_1541,N_2346);
nand U3369 (N_3369,N_1834,N_2130);
or U3370 (N_3370,N_2012,N_2332);
or U3371 (N_3371,N_1549,N_2296);
nor U3372 (N_3372,N_1551,N_1407);
or U3373 (N_3373,N_1783,N_1549);
nand U3374 (N_3374,N_1363,N_2480);
nand U3375 (N_3375,N_1623,N_1294);
nand U3376 (N_3376,N_1318,N_2222);
and U3377 (N_3377,N_1534,N_1971);
or U3378 (N_3378,N_1682,N_2273);
or U3379 (N_3379,N_1524,N_2185);
xor U3380 (N_3380,N_1631,N_2349);
nor U3381 (N_3381,N_1420,N_1903);
and U3382 (N_3382,N_2486,N_2373);
nor U3383 (N_3383,N_2363,N_2462);
xor U3384 (N_3384,N_1843,N_2071);
and U3385 (N_3385,N_1953,N_1904);
xor U3386 (N_3386,N_2471,N_2107);
nand U3387 (N_3387,N_2499,N_1689);
xnor U3388 (N_3388,N_1785,N_1804);
xor U3389 (N_3389,N_2315,N_1741);
and U3390 (N_3390,N_1671,N_1890);
nor U3391 (N_3391,N_2110,N_1739);
or U3392 (N_3392,N_2174,N_2194);
nor U3393 (N_3393,N_2491,N_2458);
nand U3394 (N_3394,N_1361,N_2122);
and U3395 (N_3395,N_1291,N_1928);
nor U3396 (N_3396,N_1815,N_1530);
or U3397 (N_3397,N_1993,N_1571);
or U3398 (N_3398,N_2361,N_1764);
nand U3399 (N_3399,N_1753,N_1411);
and U3400 (N_3400,N_2478,N_1314);
and U3401 (N_3401,N_2105,N_2218);
and U3402 (N_3402,N_1707,N_2119);
and U3403 (N_3403,N_2217,N_1735);
xnor U3404 (N_3404,N_2288,N_2150);
nand U3405 (N_3405,N_1928,N_1584);
and U3406 (N_3406,N_2172,N_1777);
nor U3407 (N_3407,N_1821,N_2278);
nor U3408 (N_3408,N_1855,N_2381);
xor U3409 (N_3409,N_1461,N_1812);
xnor U3410 (N_3410,N_1683,N_1679);
and U3411 (N_3411,N_1626,N_2453);
and U3412 (N_3412,N_1592,N_1771);
and U3413 (N_3413,N_2283,N_2005);
nor U3414 (N_3414,N_2442,N_2211);
nand U3415 (N_3415,N_1380,N_2120);
nor U3416 (N_3416,N_2067,N_1287);
nand U3417 (N_3417,N_2238,N_1401);
nor U3418 (N_3418,N_1727,N_1706);
nand U3419 (N_3419,N_2470,N_1900);
nand U3420 (N_3420,N_2078,N_1629);
and U3421 (N_3421,N_1577,N_1566);
nand U3422 (N_3422,N_1747,N_1960);
or U3423 (N_3423,N_1891,N_2116);
xnor U3424 (N_3424,N_2089,N_1705);
nor U3425 (N_3425,N_1515,N_1716);
nor U3426 (N_3426,N_2330,N_2206);
or U3427 (N_3427,N_2488,N_1745);
nand U3428 (N_3428,N_1464,N_1733);
and U3429 (N_3429,N_2419,N_1945);
nand U3430 (N_3430,N_2249,N_1988);
and U3431 (N_3431,N_1811,N_1474);
nand U3432 (N_3432,N_1834,N_2491);
and U3433 (N_3433,N_2277,N_1283);
nand U3434 (N_3434,N_1518,N_2336);
or U3435 (N_3435,N_1359,N_2211);
nor U3436 (N_3436,N_2290,N_2321);
and U3437 (N_3437,N_2454,N_2055);
nor U3438 (N_3438,N_2087,N_2245);
nor U3439 (N_3439,N_1723,N_2168);
nand U3440 (N_3440,N_2015,N_1489);
nor U3441 (N_3441,N_1464,N_2465);
xor U3442 (N_3442,N_1298,N_2199);
nand U3443 (N_3443,N_1312,N_1776);
or U3444 (N_3444,N_1968,N_2239);
xor U3445 (N_3445,N_1846,N_2426);
nand U3446 (N_3446,N_1804,N_1929);
xor U3447 (N_3447,N_2166,N_2413);
nor U3448 (N_3448,N_1687,N_1451);
or U3449 (N_3449,N_1388,N_2029);
nor U3450 (N_3450,N_2284,N_2164);
nand U3451 (N_3451,N_1443,N_2053);
nor U3452 (N_3452,N_1293,N_1727);
and U3453 (N_3453,N_2153,N_2243);
nand U3454 (N_3454,N_1695,N_2355);
xor U3455 (N_3455,N_2087,N_1456);
and U3456 (N_3456,N_2036,N_2264);
or U3457 (N_3457,N_2040,N_1362);
or U3458 (N_3458,N_1535,N_2451);
nor U3459 (N_3459,N_1767,N_2340);
nor U3460 (N_3460,N_2411,N_2176);
or U3461 (N_3461,N_1647,N_1704);
and U3462 (N_3462,N_1267,N_1577);
xor U3463 (N_3463,N_1763,N_2121);
xor U3464 (N_3464,N_1761,N_2268);
nor U3465 (N_3465,N_1324,N_2147);
nand U3466 (N_3466,N_2344,N_1476);
xnor U3467 (N_3467,N_1983,N_1790);
nor U3468 (N_3468,N_2412,N_2408);
nand U3469 (N_3469,N_1676,N_2188);
xor U3470 (N_3470,N_2269,N_1705);
nand U3471 (N_3471,N_1919,N_1624);
and U3472 (N_3472,N_1894,N_2430);
or U3473 (N_3473,N_2463,N_1354);
xnor U3474 (N_3474,N_2101,N_1506);
nor U3475 (N_3475,N_2127,N_1537);
xnor U3476 (N_3476,N_2341,N_2345);
nor U3477 (N_3477,N_1347,N_1967);
and U3478 (N_3478,N_1853,N_1795);
and U3479 (N_3479,N_2091,N_2460);
xnor U3480 (N_3480,N_1844,N_2096);
nand U3481 (N_3481,N_1360,N_2069);
xor U3482 (N_3482,N_2414,N_1703);
xor U3483 (N_3483,N_1511,N_2303);
nand U3484 (N_3484,N_2029,N_1982);
or U3485 (N_3485,N_2012,N_1339);
xnor U3486 (N_3486,N_2186,N_2138);
nand U3487 (N_3487,N_1554,N_2161);
or U3488 (N_3488,N_1287,N_2494);
and U3489 (N_3489,N_2177,N_1619);
nor U3490 (N_3490,N_2412,N_1395);
nor U3491 (N_3491,N_2449,N_1988);
or U3492 (N_3492,N_1324,N_1728);
nor U3493 (N_3493,N_1874,N_1792);
nand U3494 (N_3494,N_1487,N_2006);
or U3495 (N_3495,N_2233,N_1694);
and U3496 (N_3496,N_1521,N_2201);
nor U3497 (N_3497,N_2405,N_1848);
and U3498 (N_3498,N_1516,N_2019);
nand U3499 (N_3499,N_1685,N_2096);
nor U3500 (N_3500,N_2226,N_2373);
and U3501 (N_3501,N_2413,N_1625);
nand U3502 (N_3502,N_1516,N_1894);
nand U3503 (N_3503,N_1421,N_2124);
nand U3504 (N_3504,N_2357,N_1312);
nor U3505 (N_3505,N_1890,N_2279);
nand U3506 (N_3506,N_1388,N_2458);
nor U3507 (N_3507,N_1872,N_1941);
or U3508 (N_3508,N_2399,N_2113);
and U3509 (N_3509,N_2418,N_2376);
or U3510 (N_3510,N_2156,N_2498);
xor U3511 (N_3511,N_1395,N_2225);
xor U3512 (N_3512,N_1519,N_1633);
xor U3513 (N_3513,N_2118,N_1928);
or U3514 (N_3514,N_2026,N_1797);
and U3515 (N_3515,N_2221,N_1636);
nor U3516 (N_3516,N_1898,N_2089);
nand U3517 (N_3517,N_1461,N_1888);
or U3518 (N_3518,N_1275,N_1819);
nor U3519 (N_3519,N_1634,N_2405);
or U3520 (N_3520,N_2421,N_1852);
and U3521 (N_3521,N_1423,N_2378);
nand U3522 (N_3522,N_1577,N_1620);
or U3523 (N_3523,N_1834,N_1944);
or U3524 (N_3524,N_1661,N_1881);
nor U3525 (N_3525,N_2474,N_1957);
and U3526 (N_3526,N_1662,N_1309);
nor U3527 (N_3527,N_1402,N_1749);
and U3528 (N_3528,N_1266,N_2175);
or U3529 (N_3529,N_2037,N_1390);
xnor U3530 (N_3530,N_1689,N_2116);
nand U3531 (N_3531,N_2460,N_1712);
nand U3532 (N_3532,N_2377,N_2444);
and U3533 (N_3533,N_1857,N_2108);
xor U3534 (N_3534,N_1802,N_1469);
or U3535 (N_3535,N_1507,N_2364);
and U3536 (N_3536,N_1860,N_1355);
nand U3537 (N_3537,N_1433,N_2221);
and U3538 (N_3538,N_1407,N_2272);
nand U3539 (N_3539,N_1559,N_2237);
and U3540 (N_3540,N_1613,N_2158);
and U3541 (N_3541,N_2050,N_1419);
and U3542 (N_3542,N_2133,N_1659);
nand U3543 (N_3543,N_2270,N_2107);
or U3544 (N_3544,N_1807,N_2214);
or U3545 (N_3545,N_1579,N_1452);
nor U3546 (N_3546,N_2208,N_1283);
nor U3547 (N_3547,N_2165,N_2183);
and U3548 (N_3548,N_1398,N_2034);
and U3549 (N_3549,N_1272,N_1390);
and U3550 (N_3550,N_1529,N_1998);
or U3551 (N_3551,N_1540,N_2061);
nor U3552 (N_3552,N_1360,N_1409);
or U3553 (N_3553,N_1393,N_2198);
and U3554 (N_3554,N_1359,N_2424);
and U3555 (N_3555,N_1295,N_2153);
or U3556 (N_3556,N_1415,N_1961);
nand U3557 (N_3557,N_1494,N_1476);
xnor U3558 (N_3558,N_1393,N_2205);
xor U3559 (N_3559,N_2300,N_1563);
xnor U3560 (N_3560,N_2373,N_1913);
nor U3561 (N_3561,N_1300,N_1685);
nor U3562 (N_3562,N_2490,N_2130);
nor U3563 (N_3563,N_2224,N_2231);
nand U3564 (N_3564,N_1818,N_1431);
nor U3565 (N_3565,N_1341,N_1719);
nand U3566 (N_3566,N_1341,N_1361);
or U3567 (N_3567,N_1659,N_2019);
nor U3568 (N_3568,N_1858,N_2211);
and U3569 (N_3569,N_2210,N_2033);
nand U3570 (N_3570,N_1581,N_2363);
or U3571 (N_3571,N_2279,N_1563);
and U3572 (N_3572,N_1980,N_2128);
xor U3573 (N_3573,N_1696,N_2001);
xor U3574 (N_3574,N_1410,N_2466);
and U3575 (N_3575,N_2090,N_1551);
xor U3576 (N_3576,N_1739,N_1434);
or U3577 (N_3577,N_2185,N_1366);
nor U3578 (N_3578,N_1302,N_1459);
and U3579 (N_3579,N_1841,N_2361);
and U3580 (N_3580,N_1905,N_1659);
or U3581 (N_3581,N_1254,N_2175);
nor U3582 (N_3582,N_2262,N_2171);
and U3583 (N_3583,N_2176,N_1264);
xor U3584 (N_3584,N_2086,N_1270);
or U3585 (N_3585,N_1914,N_2285);
nor U3586 (N_3586,N_2155,N_1431);
and U3587 (N_3587,N_1410,N_1591);
nand U3588 (N_3588,N_1927,N_1803);
or U3589 (N_3589,N_1477,N_2015);
and U3590 (N_3590,N_1678,N_1396);
nor U3591 (N_3591,N_1676,N_1502);
nand U3592 (N_3592,N_1375,N_1499);
and U3593 (N_3593,N_2447,N_2008);
nor U3594 (N_3594,N_2294,N_2000);
nor U3595 (N_3595,N_2357,N_1419);
or U3596 (N_3596,N_1684,N_2008);
or U3597 (N_3597,N_1705,N_1840);
nand U3598 (N_3598,N_2244,N_2301);
or U3599 (N_3599,N_1721,N_1263);
and U3600 (N_3600,N_2164,N_1503);
and U3601 (N_3601,N_1646,N_1958);
and U3602 (N_3602,N_1885,N_1723);
nor U3603 (N_3603,N_1472,N_2241);
nor U3604 (N_3604,N_1255,N_2244);
nand U3605 (N_3605,N_1262,N_1565);
nand U3606 (N_3606,N_2457,N_1568);
or U3607 (N_3607,N_1302,N_1559);
nor U3608 (N_3608,N_2019,N_2175);
or U3609 (N_3609,N_1933,N_1606);
nor U3610 (N_3610,N_2235,N_2224);
and U3611 (N_3611,N_1353,N_1624);
and U3612 (N_3612,N_2079,N_2471);
xnor U3613 (N_3613,N_1575,N_1920);
nand U3614 (N_3614,N_1789,N_2332);
nor U3615 (N_3615,N_2253,N_2131);
xnor U3616 (N_3616,N_2240,N_1731);
and U3617 (N_3617,N_1571,N_2103);
xnor U3618 (N_3618,N_1468,N_2369);
and U3619 (N_3619,N_1968,N_2467);
xnor U3620 (N_3620,N_2129,N_1278);
or U3621 (N_3621,N_1962,N_1287);
or U3622 (N_3622,N_2062,N_1505);
xor U3623 (N_3623,N_2077,N_1486);
or U3624 (N_3624,N_1557,N_1332);
xor U3625 (N_3625,N_2210,N_2031);
nor U3626 (N_3626,N_2289,N_2245);
nor U3627 (N_3627,N_1837,N_1502);
nor U3628 (N_3628,N_1843,N_1410);
or U3629 (N_3629,N_2214,N_1875);
or U3630 (N_3630,N_2077,N_2465);
xnor U3631 (N_3631,N_1508,N_1591);
xnor U3632 (N_3632,N_2400,N_1988);
nand U3633 (N_3633,N_1686,N_2217);
nand U3634 (N_3634,N_1349,N_2358);
nor U3635 (N_3635,N_1843,N_2379);
xnor U3636 (N_3636,N_1529,N_1806);
or U3637 (N_3637,N_1535,N_2241);
nor U3638 (N_3638,N_1953,N_2095);
or U3639 (N_3639,N_1862,N_2182);
or U3640 (N_3640,N_1593,N_1806);
or U3641 (N_3641,N_1508,N_2316);
nand U3642 (N_3642,N_1262,N_2337);
nand U3643 (N_3643,N_1393,N_1962);
xnor U3644 (N_3644,N_1719,N_1708);
or U3645 (N_3645,N_2236,N_2117);
nand U3646 (N_3646,N_1818,N_2041);
nand U3647 (N_3647,N_1576,N_1738);
nand U3648 (N_3648,N_1892,N_1482);
nor U3649 (N_3649,N_1602,N_1403);
nor U3650 (N_3650,N_2423,N_2077);
nand U3651 (N_3651,N_1503,N_1882);
nand U3652 (N_3652,N_1697,N_1820);
nor U3653 (N_3653,N_1507,N_1395);
nand U3654 (N_3654,N_2302,N_2202);
nand U3655 (N_3655,N_1438,N_2335);
nand U3656 (N_3656,N_1365,N_1645);
nand U3657 (N_3657,N_1816,N_1937);
or U3658 (N_3658,N_2362,N_2284);
or U3659 (N_3659,N_2225,N_2423);
nor U3660 (N_3660,N_1457,N_1382);
nor U3661 (N_3661,N_2029,N_2402);
and U3662 (N_3662,N_2394,N_1574);
and U3663 (N_3663,N_2304,N_2008);
or U3664 (N_3664,N_1952,N_2255);
and U3665 (N_3665,N_2030,N_1671);
nand U3666 (N_3666,N_1752,N_2314);
nor U3667 (N_3667,N_1982,N_1268);
xnor U3668 (N_3668,N_1335,N_2067);
or U3669 (N_3669,N_1520,N_1997);
xnor U3670 (N_3670,N_1366,N_1363);
and U3671 (N_3671,N_2102,N_1999);
nor U3672 (N_3672,N_2443,N_1608);
or U3673 (N_3673,N_1792,N_2012);
and U3674 (N_3674,N_1394,N_1914);
nand U3675 (N_3675,N_1834,N_1354);
and U3676 (N_3676,N_1924,N_1252);
and U3677 (N_3677,N_1572,N_1827);
nor U3678 (N_3678,N_1575,N_2005);
xor U3679 (N_3679,N_2183,N_2434);
nand U3680 (N_3680,N_2359,N_1479);
xor U3681 (N_3681,N_1871,N_1418);
or U3682 (N_3682,N_2147,N_2299);
nand U3683 (N_3683,N_2208,N_2347);
nand U3684 (N_3684,N_2318,N_1720);
nand U3685 (N_3685,N_1742,N_1428);
or U3686 (N_3686,N_1559,N_2401);
xor U3687 (N_3687,N_2250,N_1412);
xnor U3688 (N_3688,N_2047,N_2394);
and U3689 (N_3689,N_1789,N_2080);
nand U3690 (N_3690,N_2210,N_2008);
and U3691 (N_3691,N_1281,N_1830);
or U3692 (N_3692,N_1706,N_1738);
nand U3693 (N_3693,N_1860,N_1698);
nor U3694 (N_3694,N_1965,N_1562);
or U3695 (N_3695,N_1518,N_1918);
xor U3696 (N_3696,N_1992,N_1262);
nand U3697 (N_3697,N_1873,N_2467);
nor U3698 (N_3698,N_2490,N_2013);
xor U3699 (N_3699,N_2056,N_2455);
xnor U3700 (N_3700,N_2432,N_1286);
or U3701 (N_3701,N_2300,N_2185);
and U3702 (N_3702,N_1857,N_1358);
nor U3703 (N_3703,N_1391,N_1372);
or U3704 (N_3704,N_1660,N_1478);
and U3705 (N_3705,N_1625,N_2192);
and U3706 (N_3706,N_2249,N_1394);
and U3707 (N_3707,N_1812,N_1752);
xnor U3708 (N_3708,N_2125,N_1675);
and U3709 (N_3709,N_1411,N_1919);
and U3710 (N_3710,N_2085,N_1276);
and U3711 (N_3711,N_2006,N_1386);
nand U3712 (N_3712,N_1881,N_1578);
nor U3713 (N_3713,N_2400,N_2373);
xnor U3714 (N_3714,N_2352,N_1713);
and U3715 (N_3715,N_1438,N_1455);
or U3716 (N_3716,N_1675,N_2040);
xnor U3717 (N_3717,N_1375,N_2440);
and U3718 (N_3718,N_1896,N_2406);
and U3719 (N_3719,N_1402,N_2314);
or U3720 (N_3720,N_1729,N_1351);
xnor U3721 (N_3721,N_1524,N_1798);
xor U3722 (N_3722,N_1526,N_1882);
or U3723 (N_3723,N_2023,N_1705);
or U3724 (N_3724,N_1821,N_1933);
xnor U3725 (N_3725,N_1758,N_2475);
xnor U3726 (N_3726,N_2108,N_2013);
nand U3727 (N_3727,N_1446,N_1497);
nand U3728 (N_3728,N_2426,N_1721);
and U3729 (N_3729,N_1810,N_1587);
nor U3730 (N_3730,N_1750,N_2388);
nand U3731 (N_3731,N_1352,N_1463);
and U3732 (N_3732,N_1391,N_1563);
and U3733 (N_3733,N_1824,N_1796);
nor U3734 (N_3734,N_1575,N_1568);
nor U3735 (N_3735,N_2441,N_1647);
or U3736 (N_3736,N_1698,N_1675);
and U3737 (N_3737,N_1496,N_1982);
nor U3738 (N_3738,N_2197,N_2173);
nor U3739 (N_3739,N_2420,N_1885);
nand U3740 (N_3740,N_1887,N_2463);
or U3741 (N_3741,N_2154,N_1949);
and U3742 (N_3742,N_1946,N_1331);
nor U3743 (N_3743,N_2452,N_1732);
nor U3744 (N_3744,N_2293,N_2237);
nor U3745 (N_3745,N_2378,N_1517);
xnor U3746 (N_3746,N_1508,N_1984);
or U3747 (N_3747,N_1822,N_1317);
nand U3748 (N_3748,N_1621,N_1444);
xor U3749 (N_3749,N_1401,N_2265);
nand U3750 (N_3750,N_2633,N_2984);
nor U3751 (N_3751,N_3624,N_2954);
nand U3752 (N_3752,N_2779,N_3697);
xor U3753 (N_3753,N_3371,N_3366);
or U3754 (N_3754,N_3210,N_3200);
and U3755 (N_3755,N_2591,N_2587);
and U3756 (N_3756,N_2694,N_3498);
and U3757 (N_3757,N_2829,N_3150);
or U3758 (N_3758,N_2827,N_2579);
or U3759 (N_3759,N_3402,N_3543);
nor U3760 (N_3760,N_2558,N_3289);
nor U3761 (N_3761,N_2836,N_2793);
nand U3762 (N_3762,N_3483,N_3456);
nor U3763 (N_3763,N_3255,N_3516);
or U3764 (N_3764,N_2666,N_3709);
and U3765 (N_3765,N_2759,N_3530);
and U3766 (N_3766,N_3021,N_2537);
or U3767 (N_3767,N_3023,N_3390);
nand U3768 (N_3768,N_2649,N_3217);
and U3769 (N_3769,N_3142,N_3558);
nor U3770 (N_3770,N_3644,N_3610);
nand U3771 (N_3771,N_3097,N_2795);
nor U3772 (N_3772,N_3221,N_3435);
xnor U3773 (N_3773,N_2609,N_2832);
and U3774 (N_3774,N_3723,N_2523);
nand U3775 (N_3775,N_3261,N_2664);
xnor U3776 (N_3776,N_2583,N_2862);
nand U3777 (N_3777,N_2782,N_3005);
xor U3778 (N_3778,N_3096,N_2699);
nand U3779 (N_3779,N_3242,N_2912);
or U3780 (N_3780,N_2627,N_3314);
or U3781 (N_3781,N_3631,N_2930);
or U3782 (N_3782,N_3646,N_3484);
and U3783 (N_3783,N_2527,N_2962);
nand U3784 (N_3784,N_2593,N_2828);
nand U3785 (N_3785,N_3545,N_3002);
or U3786 (N_3786,N_3111,N_3172);
nor U3787 (N_3787,N_2908,N_3547);
or U3788 (N_3788,N_3502,N_2612);
nor U3789 (N_3789,N_3017,N_2769);
and U3790 (N_3790,N_3469,N_2854);
or U3791 (N_3791,N_3313,N_2635);
xor U3792 (N_3792,N_3662,N_2853);
and U3793 (N_3793,N_3279,N_2598);
nor U3794 (N_3794,N_2777,N_2670);
or U3795 (N_3795,N_2837,N_3715);
nand U3796 (N_3796,N_3244,N_3676);
and U3797 (N_3797,N_3416,N_3716);
or U3798 (N_3798,N_2669,N_3088);
or U3799 (N_3799,N_2511,N_2760);
nand U3800 (N_3800,N_2608,N_3064);
and U3801 (N_3801,N_2820,N_2870);
and U3802 (N_3802,N_3344,N_2851);
or U3803 (N_3803,N_3085,N_3518);
xor U3804 (N_3804,N_3378,N_3041);
xor U3805 (N_3805,N_2657,N_2747);
xnor U3806 (N_3806,N_3609,N_2735);
and U3807 (N_3807,N_3372,N_3568);
nand U3808 (N_3808,N_2823,N_2926);
nand U3809 (N_3809,N_2811,N_3592);
xor U3810 (N_3810,N_2911,N_2840);
nand U3811 (N_3811,N_2951,N_3347);
or U3812 (N_3812,N_2695,N_2925);
and U3813 (N_3813,N_3431,N_3496);
and U3814 (N_3814,N_3690,N_2794);
xnor U3815 (N_3815,N_3499,N_3162);
nand U3816 (N_3816,N_2860,N_2973);
or U3817 (N_3817,N_3091,N_2617);
nand U3818 (N_3818,N_3247,N_2614);
or U3819 (N_3819,N_2597,N_3351);
or U3820 (N_3820,N_3109,N_3493);
xor U3821 (N_3821,N_3205,N_3550);
nor U3822 (N_3822,N_2894,N_2904);
xnor U3823 (N_3823,N_3497,N_3011);
or U3824 (N_3824,N_3309,N_3458);
or U3825 (N_3825,N_3546,N_3621);
xnor U3826 (N_3826,N_3278,N_2896);
and U3827 (N_3827,N_3001,N_3742);
or U3828 (N_3828,N_2529,N_2738);
and U3829 (N_3829,N_3448,N_2866);
xnor U3830 (N_3830,N_3039,N_2875);
nor U3831 (N_3831,N_3138,N_3196);
and U3832 (N_3832,N_3356,N_2819);
xnor U3833 (N_3833,N_3439,N_3016);
nor U3834 (N_3834,N_3026,N_2702);
nor U3835 (N_3835,N_3663,N_3674);
nand U3836 (N_3836,N_3419,N_2830);
xor U3837 (N_3837,N_3744,N_3301);
nor U3838 (N_3838,N_3513,N_3563);
or U3839 (N_3839,N_3033,N_3381);
nand U3840 (N_3840,N_3659,N_3077);
nand U3841 (N_3841,N_2736,N_2733);
nand U3842 (N_3842,N_3682,N_3565);
xnor U3843 (N_3843,N_3282,N_2570);
nand U3844 (N_3844,N_3086,N_2776);
xor U3845 (N_3845,N_2721,N_2920);
and U3846 (N_3846,N_3123,N_3102);
or U3847 (N_3847,N_3348,N_3280);
nand U3848 (N_3848,N_3046,N_2731);
nor U3849 (N_3849,N_2789,N_2900);
and U3850 (N_3850,N_3517,N_2620);
nor U3851 (N_3851,N_3334,N_3254);
and U3852 (N_3852,N_3534,N_2817);
nor U3853 (N_3853,N_3745,N_2661);
nand U3854 (N_3854,N_3283,N_3010);
or U3855 (N_3855,N_2895,N_2691);
xor U3856 (N_3856,N_3480,N_3081);
xor U3857 (N_3857,N_3043,N_2624);
xor U3858 (N_3858,N_3581,N_3163);
or U3859 (N_3859,N_3154,N_3367);
xnor U3860 (N_3860,N_2765,N_3125);
xor U3861 (N_3861,N_3616,N_3192);
and U3862 (N_3862,N_3685,N_3594);
and U3863 (N_3863,N_3595,N_2931);
nand U3864 (N_3864,N_3459,N_2578);
nor U3865 (N_3865,N_2816,N_3655);
nor U3866 (N_3866,N_3615,N_3054);
nand U3867 (N_3867,N_2883,N_2599);
nor U3868 (N_3868,N_3432,N_3074);
nor U3869 (N_3869,N_3423,N_2800);
and U3870 (N_3870,N_3350,N_3519);
nor U3871 (N_3871,N_2596,N_3444);
and U3872 (N_3872,N_2745,N_3134);
xnor U3873 (N_3873,N_3038,N_3443);
nand U3874 (N_3874,N_3104,N_3362);
xor U3875 (N_3875,N_3028,N_2772);
or U3876 (N_3876,N_3590,N_3322);
nor U3877 (N_3877,N_2799,N_3467);
xor U3878 (N_3878,N_3141,N_3706);
nand U3879 (N_3879,N_2713,N_3401);
nor U3880 (N_3880,N_3441,N_3298);
nand U3881 (N_3881,N_2671,N_2730);
nand U3882 (N_3882,N_3470,N_2863);
nor U3883 (N_3883,N_3571,N_3252);
nand U3884 (N_3884,N_3190,N_2964);
and U3885 (N_3885,N_2672,N_3073);
or U3886 (N_3886,N_2906,N_2775);
or U3887 (N_3887,N_2932,N_3640);
nor U3888 (N_3888,N_3494,N_2815);
or U3889 (N_3889,N_3276,N_3335);
and U3890 (N_3890,N_3100,N_3698);
nor U3891 (N_3891,N_3705,N_3666);
nor U3892 (N_3892,N_2982,N_2905);
xnor U3893 (N_3893,N_3364,N_2709);
and U3894 (N_3894,N_2554,N_3067);
xnor U3895 (N_3895,N_3230,N_2801);
xor U3896 (N_3896,N_3562,N_3434);
and U3897 (N_3897,N_2513,N_3520);
or U3898 (N_3898,N_3414,N_3528);
nand U3899 (N_3899,N_3338,N_3537);
and U3900 (N_3900,N_3159,N_2567);
and U3901 (N_3901,N_3526,N_3725);
nor U3902 (N_3902,N_3570,N_3525);
xnor U3903 (N_3903,N_2636,N_3296);
nor U3904 (N_3904,N_2571,N_3184);
and U3905 (N_3905,N_2923,N_2580);
and U3906 (N_3906,N_3233,N_3042);
nor U3907 (N_3907,N_2734,N_3256);
and U3908 (N_3908,N_2653,N_2590);
nand U3909 (N_3909,N_3397,N_2956);
or U3910 (N_3910,N_3675,N_3567);
and U3911 (N_3911,N_3266,N_2989);
and U3912 (N_3912,N_2739,N_2880);
nand U3913 (N_3913,N_3087,N_2850);
or U3914 (N_3914,N_2656,N_2654);
and U3915 (N_3915,N_3457,N_2879);
nand U3916 (N_3916,N_3564,N_3211);
xor U3917 (N_3917,N_3668,N_3034);
nor U3918 (N_3918,N_3552,N_3639);
or U3919 (N_3919,N_3695,N_2665);
and U3920 (N_3920,N_2771,N_3551);
xnor U3921 (N_3921,N_2958,N_3079);
xor U3922 (N_3922,N_3536,N_3454);
xnor U3923 (N_3923,N_2986,N_3169);
xnor U3924 (N_3924,N_3427,N_3689);
and U3925 (N_3925,N_3410,N_2886);
nor U3926 (N_3926,N_3116,N_3664);
nand U3927 (N_3927,N_3415,N_3625);
nor U3928 (N_3928,N_3599,N_2564);
and U3929 (N_3929,N_3170,N_3007);
nor U3930 (N_3930,N_3243,N_2980);
nand U3931 (N_3931,N_3503,N_2897);
or U3932 (N_3932,N_3103,N_2963);
and U3933 (N_3933,N_3556,N_3311);
and U3934 (N_3934,N_2676,N_3185);
and U3935 (N_3935,N_2533,N_2544);
nand U3936 (N_3936,N_2839,N_2700);
nand U3937 (N_3937,N_3144,N_3549);
and U3938 (N_3938,N_3653,N_3129);
xnor U3939 (N_3939,N_3369,N_3747);
xor U3940 (N_3940,N_3288,N_3627);
xnor U3941 (N_3941,N_2998,N_3587);
nand U3942 (N_3942,N_3234,N_2822);
or U3943 (N_3943,N_3460,N_3337);
xor U3944 (N_3944,N_3475,N_2647);
nor U3945 (N_3945,N_2502,N_2899);
nand U3946 (N_3946,N_3388,N_3020);
and U3947 (N_3947,N_3405,N_2844);
nor U3948 (N_3948,N_3323,N_3593);
and U3949 (N_3949,N_3466,N_3115);
or U3950 (N_3950,N_2887,N_2503);
nand U3951 (N_3951,N_2500,N_3476);
xor U3952 (N_3952,N_3683,N_3677);
nand U3953 (N_3953,N_3209,N_3608);
nor U3954 (N_3954,N_3361,N_2660);
and U3955 (N_3955,N_2845,N_3089);
nand U3956 (N_3956,N_2961,N_2915);
nor U3957 (N_3957,N_2907,N_3522);
xor U3958 (N_3958,N_3094,N_3710);
xor U3959 (N_3959,N_2808,N_2868);
xnor U3960 (N_3960,N_3749,N_2551);
xor U3961 (N_3961,N_3486,N_3511);
or U3962 (N_3962,N_2611,N_2871);
nor U3963 (N_3963,N_3275,N_3130);
nor U3964 (N_3964,N_3058,N_3611);
nor U3965 (N_3965,N_3739,N_2948);
or U3966 (N_3966,N_2773,N_3228);
nand U3967 (N_3967,N_3317,N_3557);
xnor U3968 (N_3968,N_2914,N_2634);
nor U3969 (N_3969,N_2568,N_2509);
or U3970 (N_3970,N_2615,N_3354);
and U3971 (N_3971,N_2806,N_3613);
or U3972 (N_3972,N_3665,N_3436);
nor U3973 (N_3973,N_3704,N_3168);
nand U3974 (N_3974,N_3320,N_3569);
or U3975 (N_3975,N_3580,N_3307);
and U3976 (N_3976,N_3012,N_3693);
xor U3977 (N_3977,N_2791,N_2877);
or U3978 (N_3978,N_2976,N_2530);
nor U3979 (N_3979,N_3137,N_3684);
and U3980 (N_3980,N_3355,N_2909);
nand U3981 (N_3981,N_3147,N_2938);
nand U3982 (N_3982,N_2701,N_2574);
or U3983 (N_3983,N_2852,N_3535);
or U3984 (N_3984,N_3294,N_3128);
xor U3985 (N_3985,N_3143,N_3738);
nor U3986 (N_3986,N_3368,N_3040);
and U3987 (N_3987,N_2835,N_2687);
and U3988 (N_3988,N_2507,N_2628);
or U3989 (N_3989,N_2746,N_3304);
nand U3990 (N_3990,N_2719,N_3579);
nor U3991 (N_3991,N_2994,N_2869);
nand U3992 (N_3992,N_3022,N_2737);
or U3993 (N_3993,N_2514,N_2553);
and U3994 (N_3994,N_3452,N_2622);
or U3995 (N_3995,N_3648,N_3741);
or U3996 (N_3996,N_2752,N_2662);
nand U3997 (N_3997,N_3117,N_2740);
nand U3998 (N_3998,N_3490,N_2546);
xnor U3999 (N_3999,N_2913,N_2833);
xnor U4000 (N_4000,N_3037,N_3281);
nor U4001 (N_4001,N_2588,N_2601);
nor U4002 (N_4002,N_2902,N_3602);
xor U4003 (N_4003,N_2517,N_2838);
nor U4004 (N_4004,N_2910,N_2903);
nor U4005 (N_4005,N_3406,N_3057);
xnor U4006 (N_4006,N_3413,N_3018);
xnor U4007 (N_4007,N_3321,N_2566);
or U4008 (N_4008,N_2841,N_3092);
or U4009 (N_4009,N_3412,N_2798);
or U4010 (N_4010,N_2510,N_2781);
nor U4011 (N_4011,N_3131,N_2924);
xor U4012 (N_4012,N_3177,N_2890);
nor U4013 (N_4013,N_3035,N_2878);
and U4014 (N_4014,N_2983,N_2764);
and U4015 (N_4015,N_3702,N_3612);
or U4016 (N_4016,N_3474,N_2623);
xnor U4017 (N_4017,N_2990,N_3214);
and U4018 (N_4018,N_3342,N_3400);
nor U4019 (N_4019,N_3030,N_3420);
nand U4020 (N_4020,N_3036,N_3465);
or U4021 (N_4021,N_2917,N_3329);
nand U4022 (N_4022,N_3249,N_3136);
or U4023 (N_4023,N_2802,N_3634);
and U4024 (N_4024,N_2565,N_2710);
or U4025 (N_4025,N_3736,N_3241);
or U4026 (N_4026,N_2645,N_2945);
or U4027 (N_4027,N_3195,N_2748);
nand U4028 (N_4028,N_3687,N_2981);
nor U4029 (N_4029,N_3272,N_2643);
xnor U4030 (N_4030,N_3376,N_3575);
or U4031 (N_4031,N_2720,N_3636);
nand U4032 (N_4032,N_3740,N_2606);
and U4033 (N_4033,N_2655,N_3188);
xnor U4034 (N_4034,N_3628,N_2508);
nand U4035 (N_4035,N_3186,N_3070);
or U4036 (N_4036,N_3409,N_3287);
nand U4037 (N_4037,N_3515,N_2563);
xnor U4038 (N_4038,N_3076,N_2992);
nand U4039 (N_4039,N_3544,N_2761);
nand U4040 (N_4040,N_3353,N_3157);
and U4041 (N_4041,N_3245,N_2979);
nor U4042 (N_4042,N_2526,N_3645);
nand U4043 (N_4043,N_3201,N_3250);
nor U4044 (N_4044,N_3669,N_3377);
xor U4045 (N_4045,N_3121,N_3422);
xnor U4046 (N_4046,N_3090,N_3622);
nand U4047 (N_4047,N_2921,N_3541);
nand U4048 (N_4048,N_3048,N_3025);
xnor U4049 (N_4049,N_3671,N_2814);
and U4050 (N_4050,N_3227,N_2936);
or U4051 (N_4051,N_3286,N_2667);
and U4052 (N_4052,N_3160,N_2684);
or U4053 (N_4053,N_2753,N_2757);
or U4054 (N_4054,N_3449,N_3181);
nor U4055 (N_4055,N_3632,N_3626);
nand U4056 (N_4056,N_2785,N_3438);
nand U4057 (N_4057,N_3061,N_3491);
xor U4058 (N_4058,N_2569,N_2703);
nor U4059 (N_4059,N_3722,N_3508);
and U4060 (N_4060,N_2847,N_2749);
xor U4061 (N_4061,N_3492,N_3204);
xor U4062 (N_4062,N_2967,N_3174);
nand U4063 (N_4063,N_3461,N_3696);
nor U4064 (N_4064,N_2638,N_3315);
nor U4065 (N_4065,N_3446,N_3734);
nand U4066 (N_4066,N_2605,N_2812);
nand U4067 (N_4067,N_2725,N_3198);
nand U4068 (N_4068,N_2901,N_3468);
nor U4069 (N_4069,N_2690,N_3265);
xor U4070 (N_4070,N_3729,N_3505);
xor U4071 (N_4071,N_3225,N_3614);
or U4072 (N_4072,N_3207,N_3000);
or U4073 (N_4073,N_2625,N_3728);
or U4074 (N_4074,N_3336,N_3328);
and U4075 (N_4075,N_2673,N_3641);
and U4076 (N_4076,N_3084,N_2631);
nor U4077 (N_4077,N_3330,N_3219);
or U4078 (N_4078,N_2648,N_2646);
nor U4079 (N_4079,N_3193,N_3426);
xor U4080 (N_4080,N_3013,N_3395);
xnor U4081 (N_4081,N_2572,N_2797);
and U4082 (N_4082,N_2918,N_3643);
and U4083 (N_4083,N_2521,N_3507);
nor U4084 (N_4084,N_3360,N_3319);
and U4085 (N_4085,N_2679,N_3327);
or U4086 (N_4086,N_3232,N_3029);
and U4087 (N_4087,N_2744,N_3657);
nand U4088 (N_4088,N_2966,N_3008);
nand U4089 (N_4089,N_2552,N_3450);
and U4090 (N_4090,N_2663,N_2864);
nor U4091 (N_4091,N_2621,N_2941);
or U4092 (N_4092,N_3386,N_2518);
nor U4093 (N_4093,N_2865,N_2585);
xor U4094 (N_4094,N_3711,N_3686);
nand U4095 (N_4095,N_3447,N_2548);
or U4096 (N_4096,N_2849,N_3075);
nor U4097 (N_4097,N_3727,N_2882);
and U4098 (N_4098,N_3127,N_3268);
or U4099 (N_4099,N_3239,N_2592);
and U4100 (N_4100,N_2950,N_2610);
or U4101 (N_4101,N_2715,N_2780);
nand U4102 (N_4102,N_3384,N_3485);
nor U4103 (N_4103,N_2639,N_3718);
or U4104 (N_4104,N_2652,N_3099);
xnor U4105 (N_4105,N_3730,N_3072);
and U4106 (N_4106,N_2573,N_3066);
nand U4107 (N_4107,N_2547,N_3681);
nor U4108 (N_4108,N_3310,N_3477);
nand U4109 (N_4109,N_2618,N_3661);
and U4110 (N_4110,N_3270,N_2867);
nand U4111 (N_4111,N_3118,N_3672);
or U4112 (N_4112,N_2534,N_2751);
nand U4113 (N_4113,N_2602,N_3688);
xnor U4114 (N_4114,N_2506,N_2589);
xor U4115 (N_4115,N_2804,N_3318);
or U4116 (N_4116,N_3290,N_3324);
and U4117 (N_4117,N_2978,N_3560);
nand U4118 (N_4118,N_2540,N_3071);
or U4119 (N_4119,N_3357,N_3240);
nor U4120 (N_4120,N_2784,N_2557);
nand U4121 (N_4121,N_3095,N_3737);
and U4122 (N_4122,N_3654,N_3218);
nand U4123 (N_4123,N_3743,N_2697);
nand U4124 (N_4124,N_2810,N_2803);
and U4125 (N_4125,N_3396,N_3500);
nand U4126 (N_4126,N_3065,N_3540);
xor U4127 (N_4127,N_3308,N_2825);
nor U4128 (N_4128,N_3341,N_2937);
and U4129 (N_4129,N_3047,N_2708);
nor U4130 (N_4130,N_3429,N_2532);
and U4131 (N_4131,N_3649,N_3638);
or U4132 (N_4132,N_3604,N_3044);
nor U4133 (N_4133,N_3052,N_2857);
nor U4134 (N_4134,N_3373,N_2504);
nor U4135 (N_4135,N_3586,N_3206);
and U4136 (N_4136,N_2619,N_3049);
and U4137 (N_4137,N_3605,N_2616);
nand U4138 (N_4138,N_2520,N_2650);
xnor U4139 (N_4139,N_3146,N_2724);
and U4140 (N_4140,N_2524,N_3126);
nand U4141 (N_4141,N_3292,N_2774);
xnor U4142 (N_4142,N_2675,N_3006);
xnor U4143 (N_4143,N_3591,N_3455);
or U4144 (N_4144,N_2988,N_3488);
nand U4145 (N_4145,N_3300,N_3692);
xnor U4146 (N_4146,N_2728,N_2995);
nor U4147 (N_4147,N_3365,N_3180);
nor U4148 (N_4148,N_3251,N_3291);
nor U4149 (N_4149,N_2550,N_3231);
xnor U4150 (N_4150,N_3343,N_3445);
and U4151 (N_4151,N_2792,N_2522);
xor U4152 (N_4152,N_3375,N_3119);
nand U4153 (N_4153,N_3331,N_3374);
or U4154 (N_4154,N_2756,N_3277);
and U4155 (N_4155,N_3236,N_3701);
nand U4156 (N_4156,N_2696,N_3179);
nand U4157 (N_4157,N_2898,N_2516);
xnor U4158 (N_4158,N_2556,N_2581);
or U4159 (N_4159,N_2916,N_3597);
and U4160 (N_4160,N_3027,N_2818);
nand U4161 (N_4161,N_3700,N_2668);
or U4162 (N_4162,N_2965,N_3358);
nand U4163 (N_4163,N_2584,N_3559);
nand U4164 (N_4164,N_3167,N_3582);
nand U4165 (N_4165,N_2939,N_2873);
nand U4166 (N_4166,N_3216,N_2767);
nor U4167 (N_4167,N_2974,N_2706);
and U4168 (N_4168,N_3194,N_3050);
or U4169 (N_4169,N_2575,N_3726);
or U4170 (N_4170,N_2999,N_3238);
nand U4171 (N_4171,N_3398,N_3418);
xnor U4172 (N_4172,N_3083,N_2968);
nand U4173 (N_4173,N_3471,N_3585);
or U4174 (N_4174,N_3258,N_3062);
or U4175 (N_4175,N_3472,N_2613);
xnor U4176 (N_4176,N_3260,N_3603);
or U4177 (N_4177,N_3312,N_2848);
nand U4178 (N_4178,N_3158,N_2885);
or U4179 (N_4179,N_3407,N_2977);
and U4180 (N_4180,N_3098,N_3403);
nor U4181 (N_4181,N_2519,N_3656);
or U4182 (N_4182,N_3506,N_2874);
xor U4183 (N_4183,N_3731,N_2722);
nand U4184 (N_4184,N_2600,N_3155);
xnor U4185 (N_4185,N_3139,N_3339);
and U4186 (N_4186,N_2778,N_3617);
xor U4187 (N_4187,N_3630,N_2985);
xnor U4188 (N_4188,N_2718,N_2834);
or U4189 (N_4189,N_2603,N_3382);
or U4190 (N_4190,N_3417,N_3340);
xor U4191 (N_4191,N_3433,N_3584);
nor U4192 (N_4192,N_3349,N_3712);
xnor U4193 (N_4193,N_3093,N_3151);
or U4194 (N_4194,N_3060,N_3153);
and U4195 (N_4195,N_3229,N_3113);
xor U4196 (N_4196,N_2543,N_3735);
nor U4197 (N_4197,N_3667,N_2641);
nor U4198 (N_4198,N_3208,N_3120);
and U4199 (N_4199,N_2766,N_3724);
xor U4200 (N_4200,N_3024,N_3080);
and U4201 (N_4201,N_2528,N_2549);
and U4202 (N_4202,N_3110,N_2682);
nor U4203 (N_4203,N_2934,N_2861);
xor U4204 (N_4204,N_2831,N_3202);
or U4205 (N_4205,N_2842,N_3014);
or U4206 (N_4206,N_3363,N_2594);
xnor U4207 (N_4207,N_3133,N_2658);
and U4208 (N_4208,N_3352,N_2927);
and U4209 (N_4209,N_3680,N_3389);
or U4210 (N_4210,N_3583,N_3269);
nor U4211 (N_4211,N_3577,N_2630);
nor U4212 (N_4212,N_3713,N_3411);
xnor U4213 (N_4213,N_2762,N_3316);
nand U4214 (N_4214,N_2884,N_2889);
or U4215 (N_4215,N_2933,N_2993);
nand U4216 (N_4216,N_2881,N_2512);
nand U4217 (N_4217,N_3056,N_2971);
and U4218 (N_4218,N_3391,N_3679);
nor U4219 (N_4219,N_2683,N_3453);
and U4220 (N_4220,N_2876,N_3345);
or U4221 (N_4221,N_3618,N_3482);
nand U4222 (N_4222,N_3148,N_2640);
nand U4223 (N_4223,N_3512,N_3222);
and U4224 (N_4224,N_2692,N_3542);
nand U4225 (N_4225,N_3473,N_3370);
or U4226 (N_4226,N_3464,N_3380);
and U4227 (N_4227,N_2629,N_2712);
xnor U4228 (N_4228,N_2758,N_2763);
nand U4229 (N_4229,N_2813,N_3107);
xor U4230 (N_4230,N_3660,N_2729);
xor U4231 (N_4231,N_3257,N_2940);
xor U4232 (N_4232,N_3699,N_2531);
or U4233 (N_4233,N_2846,N_3189);
and U4234 (N_4234,N_2535,N_3068);
nand U4235 (N_4235,N_3297,N_2659);
xor U4236 (N_4236,N_3504,N_2770);
xnor U4237 (N_4237,N_3514,N_2525);
nand U4238 (N_4238,N_3521,N_2946);
nor U4239 (N_4239,N_3285,N_2826);
xnor U4240 (N_4240,N_2577,N_3478);
or U4241 (N_4241,N_3019,N_2996);
nor U4242 (N_4242,N_2807,N_3399);
and U4243 (N_4243,N_3105,N_2949);
nor U4244 (N_4244,N_2714,N_2505);
nor U4245 (N_4245,N_2970,N_3430);
nor U4246 (N_4246,N_3732,N_3108);
nand U4247 (N_4247,N_3305,N_3199);
xnor U4248 (N_4248,N_3529,N_2542);
nand U4249 (N_4249,N_3428,N_2576);
nor U4250 (N_4250,N_2677,N_3387);
xor U4251 (N_4251,N_3051,N_3176);
or U4252 (N_4252,N_2893,N_3721);
xor U4253 (N_4253,N_3031,N_3302);
xnor U4254 (N_4254,N_3203,N_2872);
xnor U4255 (N_4255,N_2607,N_2859);
and U4256 (N_4256,N_3122,N_2536);
xnor U4257 (N_4257,N_2929,N_2858);
and U4258 (N_4258,N_3442,N_3523);
and U4259 (N_4259,N_3145,N_3299);
nor U4260 (N_4260,N_3694,N_2582);
nand U4261 (N_4261,N_2680,N_3132);
nand U4262 (N_4262,N_2821,N_2693);
and U4263 (N_4263,N_2626,N_3220);
and U4264 (N_4264,N_3578,N_3248);
or U4265 (N_4265,N_3424,N_2942);
xor U4266 (N_4266,N_3589,N_3533);
xnor U4267 (N_4267,N_3212,N_3596);
nand U4268 (N_4268,N_3332,N_3509);
nor U4269 (N_4269,N_3259,N_3015);
nor U4270 (N_4270,N_3273,N_3003);
or U4271 (N_4271,N_3101,N_3263);
nor U4272 (N_4272,N_3032,N_3566);
or U4273 (N_4273,N_3235,N_2997);
and U4274 (N_4274,N_2783,N_3246);
and U4275 (N_4275,N_3479,N_3156);
and U4276 (N_4276,N_3703,N_3532);
xnor U4277 (N_4277,N_3404,N_2959);
nor U4278 (N_4278,N_2919,N_3264);
xnor U4279 (N_4279,N_3173,N_3325);
or U4280 (N_4280,N_3633,N_3670);
xnor U4281 (N_4281,N_3262,N_2560);
nor U4282 (N_4282,N_3393,N_3237);
nor U4283 (N_4283,N_2539,N_2698);
and U4284 (N_4284,N_2928,N_3481);
nor U4285 (N_4285,N_3106,N_3553);
and U4286 (N_4286,N_3383,N_3379);
xnor U4287 (N_4287,N_2644,N_2943);
nand U4288 (N_4288,N_2991,N_3600);
nand U4289 (N_4289,N_2790,N_2726);
or U4290 (N_4290,N_3607,N_3191);
nor U4291 (N_4291,N_3573,N_3495);
or U4292 (N_4292,N_3748,N_3708);
and U4293 (N_4293,N_2855,N_3187);
xnor U4294 (N_4294,N_3063,N_3619);
nor U4295 (N_4295,N_3501,N_3326);
or U4296 (N_4296,N_3149,N_2796);
xor U4297 (N_4297,N_3009,N_2786);
or U4298 (N_4298,N_2960,N_2711);
nand U4299 (N_4299,N_3719,N_3053);
xnor U4300 (N_4300,N_2545,N_3746);
xnor U4301 (N_4301,N_2559,N_3548);
or U4302 (N_4302,N_2856,N_3114);
nor U4303 (N_4303,N_3510,N_2892);
nor U4304 (N_4304,N_2562,N_3333);
and U4305 (N_4305,N_2741,N_3175);
and U4306 (N_4306,N_3165,N_3425);
nor U4307 (N_4307,N_3647,N_3135);
or U4308 (N_4308,N_2805,N_2538);
nand U4309 (N_4309,N_3178,N_3124);
or U4310 (N_4310,N_3171,N_2716);
and U4311 (N_4311,N_3306,N_3487);
and U4312 (N_4312,N_3720,N_3539);
xor U4313 (N_4313,N_2843,N_2743);
nor U4314 (N_4314,N_3462,N_2637);
nor U4315 (N_4315,N_3652,N_3651);
nand U4316 (N_4316,N_3714,N_3223);
or U4317 (N_4317,N_3554,N_3678);
nand U4318 (N_4318,N_3691,N_2947);
xnor U4319 (N_4319,N_3055,N_3524);
and U4320 (N_4320,N_2969,N_3140);
and U4321 (N_4321,N_2561,N_3623);
and U4322 (N_4322,N_3274,N_3650);
nand U4323 (N_4323,N_2788,N_3197);
nand U4324 (N_4324,N_3166,N_3451);
xnor U4325 (N_4325,N_3213,N_3161);
and U4326 (N_4326,N_2952,N_2975);
or U4327 (N_4327,N_3658,N_3673);
or U4328 (N_4328,N_2681,N_2555);
nand U4329 (N_4329,N_2922,N_2955);
or U4330 (N_4330,N_3527,N_2754);
or U4331 (N_4331,N_3082,N_3112);
and U4332 (N_4332,N_3295,N_2586);
and U4333 (N_4333,N_2642,N_3293);
or U4334 (N_4334,N_2723,N_3271);
xnor U4335 (N_4335,N_3284,N_2888);
nor U4336 (N_4336,N_3045,N_2935);
nand U4337 (N_4337,N_3437,N_2689);
nor U4338 (N_4338,N_3267,N_2824);
and U4339 (N_4339,N_3394,N_2632);
nor U4340 (N_4340,N_3606,N_2674);
or U4341 (N_4341,N_2595,N_3572);
xnor U4342 (N_4342,N_3152,N_2707);
nand U4343 (N_4343,N_2953,N_3642);
nand U4344 (N_4344,N_3059,N_2541);
or U4345 (N_4345,N_2972,N_3538);
nand U4346 (N_4346,N_2678,N_3182);
and U4347 (N_4347,N_2957,N_3561);
xor U4348 (N_4348,N_3489,N_2809);
xor U4349 (N_4349,N_3215,N_2768);
and U4350 (N_4350,N_2515,N_3598);
and U4351 (N_4351,N_2688,N_3555);
or U4352 (N_4352,N_2944,N_3707);
nand U4353 (N_4353,N_2686,N_3601);
nor U4354 (N_4354,N_3440,N_3303);
and U4355 (N_4355,N_3635,N_2755);
xnor U4356 (N_4356,N_3629,N_3620);
nand U4357 (N_4357,N_3463,N_3253);
or U4358 (N_4358,N_3531,N_2685);
or U4359 (N_4359,N_2727,N_3078);
or U4360 (N_4360,N_3421,N_2651);
or U4361 (N_4361,N_3576,N_2705);
xnor U4362 (N_4362,N_2891,N_2704);
and U4363 (N_4363,N_2501,N_3637);
nand U4364 (N_4364,N_2987,N_2742);
nor U4365 (N_4365,N_3392,N_2787);
nand U4366 (N_4366,N_2732,N_3164);
nor U4367 (N_4367,N_3069,N_3574);
and U4368 (N_4368,N_3346,N_3226);
nand U4369 (N_4369,N_3183,N_3717);
xor U4370 (N_4370,N_2717,N_3385);
xnor U4371 (N_4371,N_3359,N_3224);
nor U4372 (N_4372,N_2750,N_3408);
and U4373 (N_4373,N_3733,N_3588);
nor U4374 (N_4374,N_2604,N_3004);
xor U4375 (N_4375,N_2595,N_2829);
or U4376 (N_4376,N_2739,N_3434);
and U4377 (N_4377,N_3053,N_3179);
and U4378 (N_4378,N_2907,N_3017);
xor U4379 (N_4379,N_2826,N_3089);
nor U4380 (N_4380,N_3019,N_2851);
or U4381 (N_4381,N_2610,N_3495);
xor U4382 (N_4382,N_3532,N_2802);
and U4383 (N_4383,N_2643,N_3030);
nand U4384 (N_4384,N_3385,N_2989);
and U4385 (N_4385,N_2509,N_2828);
nand U4386 (N_4386,N_3465,N_3583);
nand U4387 (N_4387,N_2817,N_3153);
and U4388 (N_4388,N_3477,N_3721);
and U4389 (N_4389,N_2517,N_3561);
or U4390 (N_4390,N_2767,N_2645);
nor U4391 (N_4391,N_3166,N_3742);
nand U4392 (N_4392,N_3293,N_3017);
nand U4393 (N_4393,N_2635,N_2770);
and U4394 (N_4394,N_3507,N_3305);
nand U4395 (N_4395,N_3124,N_3033);
xnor U4396 (N_4396,N_2923,N_3698);
nor U4397 (N_4397,N_3527,N_3081);
nand U4398 (N_4398,N_2719,N_3656);
nor U4399 (N_4399,N_2817,N_3388);
and U4400 (N_4400,N_3186,N_3408);
and U4401 (N_4401,N_3385,N_3185);
or U4402 (N_4402,N_3709,N_3242);
xnor U4403 (N_4403,N_2778,N_3556);
or U4404 (N_4404,N_3438,N_2520);
nor U4405 (N_4405,N_3454,N_3234);
xor U4406 (N_4406,N_3092,N_2506);
or U4407 (N_4407,N_3726,N_2925);
nor U4408 (N_4408,N_3042,N_3401);
nand U4409 (N_4409,N_2579,N_3031);
nor U4410 (N_4410,N_3243,N_3578);
nor U4411 (N_4411,N_3429,N_3634);
xnor U4412 (N_4412,N_2860,N_3519);
and U4413 (N_4413,N_2835,N_3234);
nand U4414 (N_4414,N_3086,N_3520);
xor U4415 (N_4415,N_2576,N_3257);
xor U4416 (N_4416,N_2987,N_3398);
nand U4417 (N_4417,N_3653,N_3595);
nand U4418 (N_4418,N_3191,N_2662);
or U4419 (N_4419,N_3236,N_3325);
xnor U4420 (N_4420,N_3168,N_2618);
nor U4421 (N_4421,N_3566,N_2680);
nor U4422 (N_4422,N_2740,N_2881);
nor U4423 (N_4423,N_3346,N_3224);
nor U4424 (N_4424,N_3458,N_2943);
xnor U4425 (N_4425,N_2655,N_2589);
xor U4426 (N_4426,N_2983,N_3382);
and U4427 (N_4427,N_3574,N_3707);
xnor U4428 (N_4428,N_3491,N_2603);
nand U4429 (N_4429,N_2905,N_2956);
xor U4430 (N_4430,N_3441,N_2785);
nand U4431 (N_4431,N_3335,N_2520);
or U4432 (N_4432,N_3483,N_3346);
and U4433 (N_4433,N_3745,N_2704);
nor U4434 (N_4434,N_3081,N_2568);
nand U4435 (N_4435,N_3067,N_2624);
or U4436 (N_4436,N_3431,N_2521);
and U4437 (N_4437,N_2643,N_3525);
nand U4438 (N_4438,N_2629,N_2836);
xnor U4439 (N_4439,N_2837,N_3385);
xnor U4440 (N_4440,N_3488,N_2873);
or U4441 (N_4441,N_3634,N_3405);
and U4442 (N_4442,N_3573,N_3140);
xnor U4443 (N_4443,N_2796,N_3296);
and U4444 (N_4444,N_2687,N_2512);
nor U4445 (N_4445,N_3345,N_3660);
and U4446 (N_4446,N_3024,N_2732);
and U4447 (N_4447,N_2704,N_3366);
xor U4448 (N_4448,N_3161,N_3277);
nor U4449 (N_4449,N_3652,N_2577);
xnor U4450 (N_4450,N_3418,N_2702);
nand U4451 (N_4451,N_3114,N_3342);
nor U4452 (N_4452,N_3696,N_2973);
xor U4453 (N_4453,N_3071,N_2812);
nand U4454 (N_4454,N_3169,N_2824);
nor U4455 (N_4455,N_3449,N_3261);
and U4456 (N_4456,N_3184,N_2641);
or U4457 (N_4457,N_2808,N_3510);
nand U4458 (N_4458,N_2664,N_2633);
or U4459 (N_4459,N_3329,N_2748);
and U4460 (N_4460,N_2991,N_3644);
or U4461 (N_4461,N_3558,N_3396);
or U4462 (N_4462,N_2668,N_3504);
or U4463 (N_4463,N_3228,N_3214);
nand U4464 (N_4464,N_2618,N_2773);
nand U4465 (N_4465,N_2527,N_3142);
or U4466 (N_4466,N_3051,N_3066);
xor U4467 (N_4467,N_3745,N_3343);
nand U4468 (N_4468,N_2879,N_2641);
xor U4469 (N_4469,N_3034,N_2634);
xnor U4470 (N_4470,N_3333,N_2680);
nand U4471 (N_4471,N_3199,N_3119);
and U4472 (N_4472,N_2559,N_2851);
or U4473 (N_4473,N_2847,N_2923);
nand U4474 (N_4474,N_2716,N_2816);
or U4475 (N_4475,N_3007,N_3199);
nor U4476 (N_4476,N_3143,N_3614);
or U4477 (N_4477,N_2661,N_3411);
nor U4478 (N_4478,N_3706,N_3151);
xnor U4479 (N_4479,N_2739,N_3061);
and U4480 (N_4480,N_2533,N_3234);
and U4481 (N_4481,N_2654,N_3282);
nand U4482 (N_4482,N_2943,N_3097);
nor U4483 (N_4483,N_2844,N_2804);
nor U4484 (N_4484,N_3714,N_2726);
xor U4485 (N_4485,N_2637,N_3407);
xnor U4486 (N_4486,N_3109,N_3727);
and U4487 (N_4487,N_2578,N_2882);
xor U4488 (N_4488,N_2550,N_2775);
or U4489 (N_4489,N_3055,N_2667);
or U4490 (N_4490,N_3604,N_3627);
xnor U4491 (N_4491,N_2977,N_2846);
and U4492 (N_4492,N_3194,N_3207);
xnor U4493 (N_4493,N_3200,N_3395);
and U4494 (N_4494,N_3273,N_3617);
xnor U4495 (N_4495,N_2925,N_3156);
or U4496 (N_4496,N_3703,N_3167);
and U4497 (N_4497,N_2802,N_2896);
nor U4498 (N_4498,N_3483,N_3568);
nor U4499 (N_4499,N_2615,N_3254);
nor U4500 (N_4500,N_2614,N_3046);
nor U4501 (N_4501,N_2560,N_2733);
and U4502 (N_4502,N_2699,N_3305);
and U4503 (N_4503,N_2810,N_3401);
nor U4504 (N_4504,N_2611,N_2717);
or U4505 (N_4505,N_2855,N_3098);
or U4506 (N_4506,N_3625,N_3199);
or U4507 (N_4507,N_2752,N_3663);
nand U4508 (N_4508,N_3538,N_3320);
and U4509 (N_4509,N_2568,N_3600);
and U4510 (N_4510,N_3252,N_3366);
nor U4511 (N_4511,N_3332,N_2566);
nor U4512 (N_4512,N_2883,N_3253);
or U4513 (N_4513,N_2599,N_3393);
or U4514 (N_4514,N_3426,N_3018);
or U4515 (N_4515,N_2688,N_2710);
nor U4516 (N_4516,N_3120,N_3532);
xnor U4517 (N_4517,N_3117,N_3466);
nor U4518 (N_4518,N_2629,N_2692);
or U4519 (N_4519,N_3700,N_3129);
or U4520 (N_4520,N_3511,N_2546);
nand U4521 (N_4521,N_3461,N_2971);
or U4522 (N_4522,N_3341,N_3602);
nor U4523 (N_4523,N_3704,N_3211);
and U4524 (N_4524,N_3220,N_2743);
or U4525 (N_4525,N_3688,N_3308);
and U4526 (N_4526,N_2971,N_2766);
xnor U4527 (N_4527,N_2760,N_3667);
and U4528 (N_4528,N_3734,N_2852);
or U4529 (N_4529,N_3253,N_3491);
and U4530 (N_4530,N_2909,N_3557);
nand U4531 (N_4531,N_3131,N_2524);
xor U4532 (N_4532,N_3246,N_2712);
nand U4533 (N_4533,N_3513,N_3491);
nand U4534 (N_4534,N_2654,N_3623);
or U4535 (N_4535,N_3191,N_3083);
or U4536 (N_4536,N_3259,N_2662);
nor U4537 (N_4537,N_3038,N_2773);
xnor U4538 (N_4538,N_3734,N_3237);
xnor U4539 (N_4539,N_2983,N_3735);
nand U4540 (N_4540,N_2567,N_2602);
nand U4541 (N_4541,N_3052,N_3604);
xor U4542 (N_4542,N_2901,N_3105);
nand U4543 (N_4543,N_2992,N_3715);
nand U4544 (N_4544,N_3214,N_3134);
xnor U4545 (N_4545,N_2767,N_3439);
and U4546 (N_4546,N_2905,N_3183);
nand U4547 (N_4547,N_2856,N_2520);
and U4548 (N_4548,N_3087,N_2700);
nand U4549 (N_4549,N_3033,N_2720);
or U4550 (N_4550,N_3119,N_3243);
nor U4551 (N_4551,N_3653,N_2927);
nor U4552 (N_4552,N_3478,N_3726);
nand U4553 (N_4553,N_3275,N_3715);
and U4554 (N_4554,N_2552,N_2592);
and U4555 (N_4555,N_3523,N_2684);
nor U4556 (N_4556,N_3202,N_3418);
nand U4557 (N_4557,N_3135,N_3673);
nand U4558 (N_4558,N_2569,N_3675);
nor U4559 (N_4559,N_3006,N_3373);
xnor U4560 (N_4560,N_2638,N_2977);
xnor U4561 (N_4561,N_3669,N_2817);
and U4562 (N_4562,N_2529,N_3741);
nand U4563 (N_4563,N_3259,N_2782);
xnor U4564 (N_4564,N_3372,N_2523);
nand U4565 (N_4565,N_2527,N_3024);
and U4566 (N_4566,N_3261,N_2616);
and U4567 (N_4567,N_3392,N_3475);
nand U4568 (N_4568,N_3487,N_2953);
and U4569 (N_4569,N_3727,N_2782);
nor U4570 (N_4570,N_3061,N_2588);
nand U4571 (N_4571,N_3416,N_2607);
xnor U4572 (N_4572,N_3075,N_3420);
and U4573 (N_4573,N_3297,N_3709);
and U4574 (N_4574,N_3058,N_2868);
nand U4575 (N_4575,N_3699,N_2921);
and U4576 (N_4576,N_2751,N_3718);
nand U4577 (N_4577,N_2592,N_3698);
or U4578 (N_4578,N_3195,N_3272);
xor U4579 (N_4579,N_3039,N_3388);
xor U4580 (N_4580,N_3027,N_3418);
and U4581 (N_4581,N_2682,N_2864);
xnor U4582 (N_4582,N_2562,N_3362);
xnor U4583 (N_4583,N_3725,N_2555);
and U4584 (N_4584,N_2734,N_2761);
nor U4585 (N_4585,N_3672,N_3548);
nor U4586 (N_4586,N_3504,N_2994);
nand U4587 (N_4587,N_3439,N_2811);
nand U4588 (N_4588,N_3536,N_2816);
or U4589 (N_4589,N_2615,N_3676);
and U4590 (N_4590,N_3397,N_2833);
xor U4591 (N_4591,N_3310,N_2828);
or U4592 (N_4592,N_2979,N_3385);
or U4593 (N_4593,N_3597,N_2674);
and U4594 (N_4594,N_3022,N_2843);
xor U4595 (N_4595,N_3009,N_3164);
or U4596 (N_4596,N_2676,N_2809);
or U4597 (N_4597,N_2585,N_2532);
nor U4598 (N_4598,N_2501,N_3153);
nor U4599 (N_4599,N_3619,N_3657);
or U4600 (N_4600,N_2844,N_3740);
and U4601 (N_4601,N_3498,N_3090);
xnor U4602 (N_4602,N_3358,N_3410);
or U4603 (N_4603,N_3001,N_3632);
xnor U4604 (N_4604,N_3576,N_3514);
and U4605 (N_4605,N_3279,N_2712);
and U4606 (N_4606,N_3257,N_3371);
nor U4607 (N_4607,N_3333,N_3491);
nor U4608 (N_4608,N_3393,N_3424);
or U4609 (N_4609,N_2963,N_3128);
and U4610 (N_4610,N_3451,N_3694);
nor U4611 (N_4611,N_3476,N_3024);
xor U4612 (N_4612,N_2990,N_2887);
nand U4613 (N_4613,N_3199,N_3198);
nand U4614 (N_4614,N_3742,N_2961);
or U4615 (N_4615,N_2609,N_3425);
nand U4616 (N_4616,N_2623,N_2731);
or U4617 (N_4617,N_2788,N_2785);
and U4618 (N_4618,N_3288,N_2648);
xnor U4619 (N_4619,N_3660,N_2857);
xor U4620 (N_4620,N_3409,N_3456);
or U4621 (N_4621,N_3353,N_3587);
and U4622 (N_4622,N_3336,N_2802);
nor U4623 (N_4623,N_3401,N_2705);
and U4624 (N_4624,N_3139,N_2850);
nor U4625 (N_4625,N_2712,N_3646);
nand U4626 (N_4626,N_3226,N_3164);
nor U4627 (N_4627,N_2535,N_3373);
nand U4628 (N_4628,N_3435,N_2800);
or U4629 (N_4629,N_3649,N_2537);
or U4630 (N_4630,N_2825,N_3083);
nand U4631 (N_4631,N_3186,N_3599);
nand U4632 (N_4632,N_2979,N_3279);
nand U4633 (N_4633,N_3477,N_3466);
nand U4634 (N_4634,N_2893,N_3562);
nand U4635 (N_4635,N_2742,N_3650);
or U4636 (N_4636,N_2764,N_3315);
and U4637 (N_4637,N_3444,N_3308);
or U4638 (N_4638,N_3026,N_2936);
nand U4639 (N_4639,N_3480,N_3063);
nor U4640 (N_4640,N_2620,N_3594);
nand U4641 (N_4641,N_3708,N_2665);
xor U4642 (N_4642,N_3190,N_2832);
nand U4643 (N_4643,N_2787,N_3721);
nand U4644 (N_4644,N_3419,N_3101);
xnor U4645 (N_4645,N_2756,N_3502);
or U4646 (N_4646,N_3043,N_3222);
nand U4647 (N_4647,N_3442,N_3279);
nor U4648 (N_4648,N_2806,N_3144);
or U4649 (N_4649,N_3549,N_2846);
or U4650 (N_4650,N_2972,N_3383);
nand U4651 (N_4651,N_3634,N_2621);
nor U4652 (N_4652,N_2681,N_3719);
xnor U4653 (N_4653,N_3145,N_3473);
nor U4654 (N_4654,N_2961,N_3388);
nor U4655 (N_4655,N_3542,N_3539);
or U4656 (N_4656,N_2629,N_2779);
nand U4657 (N_4657,N_2970,N_3188);
and U4658 (N_4658,N_3614,N_3484);
and U4659 (N_4659,N_3313,N_2630);
nand U4660 (N_4660,N_2851,N_3301);
and U4661 (N_4661,N_2723,N_2618);
nand U4662 (N_4662,N_2938,N_2949);
xor U4663 (N_4663,N_2734,N_2612);
nor U4664 (N_4664,N_3219,N_3374);
and U4665 (N_4665,N_2628,N_3562);
xnor U4666 (N_4666,N_3735,N_2874);
and U4667 (N_4667,N_3002,N_2700);
or U4668 (N_4668,N_3504,N_3643);
xnor U4669 (N_4669,N_3025,N_3530);
nand U4670 (N_4670,N_3520,N_2566);
or U4671 (N_4671,N_2754,N_2704);
nor U4672 (N_4672,N_3041,N_3121);
nand U4673 (N_4673,N_2844,N_2613);
or U4674 (N_4674,N_3381,N_3670);
or U4675 (N_4675,N_3076,N_2611);
nor U4676 (N_4676,N_2734,N_3260);
nor U4677 (N_4677,N_2606,N_2717);
nor U4678 (N_4678,N_3223,N_2648);
and U4679 (N_4679,N_3113,N_2524);
and U4680 (N_4680,N_2523,N_3690);
xnor U4681 (N_4681,N_3273,N_3637);
or U4682 (N_4682,N_2826,N_2793);
and U4683 (N_4683,N_3166,N_3084);
nand U4684 (N_4684,N_2933,N_3622);
and U4685 (N_4685,N_3271,N_3462);
nand U4686 (N_4686,N_3591,N_3140);
and U4687 (N_4687,N_3528,N_2738);
nor U4688 (N_4688,N_3488,N_2638);
or U4689 (N_4689,N_2971,N_3422);
or U4690 (N_4690,N_3640,N_2622);
and U4691 (N_4691,N_2801,N_2642);
or U4692 (N_4692,N_2741,N_3490);
xor U4693 (N_4693,N_3657,N_3233);
or U4694 (N_4694,N_2890,N_3658);
nand U4695 (N_4695,N_3442,N_3482);
or U4696 (N_4696,N_2874,N_2905);
and U4697 (N_4697,N_2981,N_3378);
or U4698 (N_4698,N_3513,N_3373);
xnor U4699 (N_4699,N_3115,N_3471);
nand U4700 (N_4700,N_3057,N_2990);
nand U4701 (N_4701,N_2526,N_3191);
nand U4702 (N_4702,N_3157,N_3000);
or U4703 (N_4703,N_2736,N_3707);
or U4704 (N_4704,N_3325,N_3504);
nand U4705 (N_4705,N_3544,N_2686);
or U4706 (N_4706,N_3456,N_3052);
nand U4707 (N_4707,N_2984,N_3460);
nor U4708 (N_4708,N_3285,N_3557);
xnor U4709 (N_4709,N_3151,N_3470);
nand U4710 (N_4710,N_3619,N_3555);
or U4711 (N_4711,N_3725,N_3193);
nor U4712 (N_4712,N_3607,N_3223);
or U4713 (N_4713,N_3148,N_3275);
nor U4714 (N_4714,N_3648,N_2629);
or U4715 (N_4715,N_2724,N_3326);
nand U4716 (N_4716,N_3166,N_3306);
xor U4717 (N_4717,N_2580,N_3144);
nand U4718 (N_4718,N_2942,N_3355);
xnor U4719 (N_4719,N_2897,N_2747);
xnor U4720 (N_4720,N_3482,N_3596);
nor U4721 (N_4721,N_2614,N_2955);
xor U4722 (N_4722,N_3396,N_3137);
and U4723 (N_4723,N_3301,N_3026);
or U4724 (N_4724,N_3618,N_2622);
xor U4725 (N_4725,N_3205,N_2762);
and U4726 (N_4726,N_3395,N_3637);
or U4727 (N_4727,N_2574,N_2587);
nand U4728 (N_4728,N_3252,N_3678);
and U4729 (N_4729,N_3164,N_2988);
xor U4730 (N_4730,N_3124,N_3699);
nand U4731 (N_4731,N_2569,N_3473);
and U4732 (N_4732,N_3689,N_2571);
nor U4733 (N_4733,N_3353,N_3746);
nand U4734 (N_4734,N_2728,N_3393);
nor U4735 (N_4735,N_2546,N_2944);
xnor U4736 (N_4736,N_3421,N_2919);
nand U4737 (N_4737,N_3344,N_2965);
or U4738 (N_4738,N_3629,N_2934);
xnor U4739 (N_4739,N_2812,N_2691);
xor U4740 (N_4740,N_3467,N_2601);
nand U4741 (N_4741,N_2724,N_3714);
nand U4742 (N_4742,N_3521,N_2743);
nor U4743 (N_4743,N_2584,N_3409);
nand U4744 (N_4744,N_3184,N_2892);
xor U4745 (N_4745,N_3632,N_3009);
or U4746 (N_4746,N_3360,N_2570);
xnor U4747 (N_4747,N_2625,N_3207);
nand U4748 (N_4748,N_2588,N_2850);
nand U4749 (N_4749,N_3165,N_3547);
nand U4750 (N_4750,N_2832,N_3694);
nor U4751 (N_4751,N_3399,N_2773);
nor U4752 (N_4752,N_2577,N_2930);
nand U4753 (N_4753,N_3375,N_3214);
nor U4754 (N_4754,N_2813,N_3026);
or U4755 (N_4755,N_2719,N_2530);
or U4756 (N_4756,N_2854,N_3414);
or U4757 (N_4757,N_3572,N_3732);
nand U4758 (N_4758,N_3405,N_2592);
and U4759 (N_4759,N_2522,N_3667);
nand U4760 (N_4760,N_3319,N_2820);
and U4761 (N_4761,N_2827,N_3524);
nor U4762 (N_4762,N_3309,N_3376);
nor U4763 (N_4763,N_3071,N_3555);
nand U4764 (N_4764,N_2587,N_3293);
and U4765 (N_4765,N_3370,N_2920);
nor U4766 (N_4766,N_3608,N_3577);
and U4767 (N_4767,N_3691,N_2634);
or U4768 (N_4768,N_2548,N_3015);
nor U4769 (N_4769,N_3435,N_3427);
xor U4770 (N_4770,N_3193,N_3688);
or U4771 (N_4771,N_2525,N_3078);
nand U4772 (N_4772,N_2959,N_3418);
or U4773 (N_4773,N_2976,N_3091);
xnor U4774 (N_4774,N_2708,N_2630);
nor U4775 (N_4775,N_3677,N_3115);
nor U4776 (N_4776,N_2737,N_2599);
xnor U4777 (N_4777,N_3504,N_3080);
xnor U4778 (N_4778,N_2979,N_2649);
nand U4779 (N_4779,N_3007,N_3009);
nand U4780 (N_4780,N_2820,N_3580);
nand U4781 (N_4781,N_3248,N_2942);
and U4782 (N_4782,N_2752,N_3249);
and U4783 (N_4783,N_2824,N_2983);
nor U4784 (N_4784,N_3181,N_3591);
nand U4785 (N_4785,N_2781,N_2795);
xnor U4786 (N_4786,N_2517,N_3489);
nor U4787 (N_4787,N_3452,N_2590);
nand U4788 (N_4788,N_3048,N_3322);
or U4789 (N_4789,N_2667,N_3397);
and U4790 (N_4790,N_3745,N_3447);
and U4791 (N_4791,N_2881,N_3316);
and U4792 (N_4792,N_3665,N_2848);
xor U4793 (N_4793,N_3670,N_2722);
nor U4794 (N_4794,N_3705,N_2854);
nand U4795 (N_4795,N_2691,N_3618);
xor U4796 (N_4796,N_2851,N_3702);
xor U4797 (N_4797,N_2604,N_2980);
nand U4798 (N_4798,N_3225,N_3376);
xor U4799 (N_4799,N_3199,N_2879);
and U4800 (N_4800,N_2708,N_3159);
nor U4801 (N_4801,N_3721,N_3339);
xnor U4802 (N_4802,N_3617,N_2834);
or U4803 (N_4803,N_2877,N_2800);
nor U4804 (N_4804,N_3016,N_2948);
and U4805 (N_4805,N_3428,N_3360);
nor U4806 (N_4806,N_3198,N_3125);
nor U4807 (N_4807,N_2892,N_3722);
or U4808 (N_4808,N_2578,N_2964);
and U4809 (N_4809,N_3360,N_2770);
nand U4810 (N_4810,N_3169,N_2907);
nand U4811 (N_4811,N_2931,N_2705);
or U4812 (N_4812,N_3169,N_3316);
or U4813 (N_4813,N_3172,N_2678);
xnor U4814 (N_4814,N_2805,N_2651);
and U4815 (N_4815,N_2617,N_3619);
and U4816 (N_4816,N_3623,N_2699);
and U4817 (N_4817,N_2585,N_3678);
xnor U4818 (N_4818,N_2864,N_3615);
nor U4819 (N_4819,N_3126,N_2906);
xnor U4820 (N_4820,N_2958,N_3315);
nor U4821 (N_4821,N_2564,N_3688);
and U4822 (N_4822,N_3376,N_2758);
nor U4823 (N_4823,N_3122,N_3145);
nor U4824 (N_4824,N_2947,N_3584);
nor U4825 (N_4825,N_2802,N_2860);
and U4826 (N_4826,N_3531,N_2556);
nor U4827 (N_4827,N_3539,N_2858);
xnor U4828 (N_4828,N_3515,N_3717);
nor U4829 (N_4829,N_2560,N_2617);
xor U4830 (N_4830,N_3727,N_2741);
and U4831 (N_4831,N_3438,N_2857);
or U4832 (N_4832,N_3709,N_3479);
nor U4833 (N_4833,N_3518,N_3641);
or U4834 (N_4834,N_2990,N_2670);
nor U4835 (N_4835,N_2539,N_2980);
nor U4836 (N_4836,N_3078,N_2788);
or U4837 (N_4837,N_3236,N_3180);
nor U4838 (N_4838,N_2616,N_2962);
nor U4839 (N_4839,N_3477,N_3297);
or U4840 (N_4840,N_3187,N_2745);
xor U4841 (N_4841,N_2609,N_3284);
xnor U4842 (N_4842,N_3290,N_3189);
nand U4843 (N_4843,N_3249,N_3002);
and U4844 (N_4844,N_2706,N_3368);
and U4845 (N_4845,N_2589,N_2995);
xor U4846 (N_4846,N_3121,N_3265);
or U4847 (N_4847,N_3638,N_3007);
xnor U4848 (N_4848,N_2788,N_2812);
nor U4849 (N_4849,N_2940,N_3524);
nand U4850 (N_4850,N_3709,N_3606);
or U4851 (N_4851,N_2860,N_2842);
xor U4852 (N_4852,N_2596,N_3116);
xnor U4853 (N_4853,N_3281,N_3149);
xnor U4854 (N_4854,N_2789,N_2653);
xor U4855 (N_4855,N_3478,N_3545);
nor U4856 (N_4856,N_3148,N_3338);
nand U4857 (N_4857,N_3340,N_2583);
and U4858 (N_4858,N_2745,N_3274);
xnor U4859 (N_4859,N_2863,N_3207);
or U4860 (N_4860,N_2557,N_2774);
or U4861 (N_4861,N_2619,N_3372);
nor U4862 (N_4862,N_2829,N_3266);
and U4863 (N_4863,N_3497,N_3127);
xor U4864 (N_4864,N_2993,N_2538);
xor U4865 (N_4865,N_3157,N_3065);
or U4866 (N_4866,N_3158,N_3522);
or U4867 (N_4867,N_3608,N_3535);
nor U4868 (N_4868,N_2949,N_3641);
nand U4869 (N_4869,N_3322,N_2536);
nand U4870 (N_4870,N_2827,N_3166);
and U4871 (N_4871,N_3465,N_3437);
nand U4872 (N_4872,N_2781,N_2979);
xnor U4873 (N_4873,N_2669,N_2964);
nand U4874 (N_4874,N_3319,N_3423);
xor U4875 (N_4875,N_2868,N_3575);
nor U4876 (N_4876,N_3529,N_2516);
xor U4877 (N_4877,N_3164,N_3408);
nand U4878 (N_4878,N_3597,N_3271);
or U4879 (N_4879,N_2771,N_2791);
nor U4880 (N_4880,N_3144,N_3497);
nand U4881 (N_4881,N_2665,N_2683);
nor U4882 (N_4882,N_3116,N_3350);
and U4883 (N_4883,N_3199,N_3529);
nor U4884 (N_4884,N_2784,N_2623);
or U4885 (N_4885,N_3240,N_3567);
and U4886 (N_4886,N_3706,N_2759);
nand U4887 (N_4887,N_3513,N_3586);
xnor U4888 (N_4888,N_3251,N_2666);
nor U4889 (N_4889,N_3515,N_3089);
nand U4890 (N_4890,N_2988,N_3539);
nor U4891 (N_4891,N_3593,N_3155);
nand U4892 (N_4892,N_2772,N_3125);
and U4893 (N_4893,N_2587,N_3023);
nand U4894 (N_4894,N_3619,N_3032);
and U4895 (N_4895,N_2680,N_2503);
or U4896 (N_4896,N_3707,N_3665);
or U4897 (N_4897,N_2945,N_3383);
nor U4898 (N_4898,N_2584,N_2936);
nand U4899 (N_4899,N_2942,N_2872);
xor U4900 (N_4900,N_2719,N_2604);
nand U4901 (N_4901,N_2639,N_3296);
xor U4902 (N_4902,N_2670,N_2786);
and U4903 (N_4903,N_3605,N_3488);
nand U4904 (N_4904,N_3280,N_3354);
and U4905 (N_4905,N_3112,N_2724);
and U4906 (N_4906,N_2960,N_3731);
nand U4907 (N_4907,N_3354,N_3014);
or U4908 (N_4908,N_3175,N_2844);
nor U4909 (N_4909,N_2896,N_3547);
and U4910 (N_4910,N_3634,N_3538);
nand U4911 (N_4911,N_2934,N_3000);
nand U4912 (N_4912,N_3726,N_3680);
nor U4913 (N_4913,N_2551,N_3423);
xor U4914 (N_4914,N_2986,N_3711);
xor U4915 (N_4915,N_3424,N_3167);
nor U4916 (N_4916,N_2645,N_3321);
and U4917 (N_4917,N_3590,N_2728);
xor U4918 (N_4918,N_3031,N_3417);
xor U4919 (N_4919,N_2570,N_2780);
nor U4920 (N_4920,N_3512,N_3559);
nand U4921 (N_4921,N_3375,N_3273);
nand U4922 (N_4922,N_3528,N_2867);
xor U4923 (N_4923,N_2802,N_3344);
and U4924 (N_4924,N_3565,N_2546);
and U4925 (N_4925,N_2796,N_3650);
and U4926 (N_4926,N_2680,N_2863);
nand U4927 (N_4927,N_3349,N_3548);
and U4928 (N_4928,N_2752,N_3445);
or U4929 (N_4929,N_3649,N_2697);
or U4930 (N_4930,N_2538,N_3735);
nor U4931 (N_4931,N_2737,N_3594);
or U4932 (N_4932,N_2822,N_2664);
nor U4933 (N_4933,N_2754,N_3300);
or U4934 (N_4934,N_2750,N_2580);
xnor U4935 (N_4935,N_3544,N_3334);
nand U4936 (N_4936,N_3248,N_3520);
nor U4937 (N_4937,N_3494,N_3380);
nand U4938 (N_4938,N_3306,N_2992);
and U4939 (N_4939,N_3472,N_3347);
and U4940 (N_4940,N_2871,N_3191);
nor U4941 (N_4941,N_2859,N_2809);
or U4942 (N_4942,N_2512,N_2887);
or U4943 (N_4943,N_3166,N_3077);
and U4944 (N_4944,N_3433,N_3308);
nor U4945 (N_4945,N_2772,N_3127);
xor U4946 (N_4946,N_3119,N_3093);
xor U4947 (N_4947,N_2691,N_3258);
or U4948 (N_4948,N_2858,N_3735);
nor U4949 (N_4949,N_2735,N_2581);
nor U4950 (N_4950,N_3708,N_2715);
nor U4951 (N_4951,N_3731,N_3342);
nand U4952 (N_4952,N_2851,N_3653);
and U4953 (N_4953,N_3351,N_2571);
xor U4954 (N_4954,N_3620,N_3668);
xor U4955 (N_4955,N_2851,N_2797);
nand U4956 (N_4956,N_3716,N_2510);
and U4957 (N_4957,N_3049,N_3221);
nor U4958 (N_4958,N_2785,N_3670);
or U4959 (N_4959,N_3021,N_3381);
nor U4960 (N_4960,N_2990,N_2932);
or U4961 (N_4961,N_3345,N_3640);
nor U4962 (N_4962,N_3279,N_2993);
or U4963 (N_4963,N_3042,N_2549);
nor U4964 (N_4964,N_3703,N_3172);
nor U4965 (N_4965,N_2811,N_2860);
and U4966 (N_4966,N_3572,N_3428);
and U4967 (N_4967,N_2599,N_2568);
and U4968 (N_4968,N_2704,N_3264);
and U4969 (N_4969,N_3563,N_2937);
and U4970 (N_4970,N_3432,N_3399);
xnor U4971 (N_4971,N_3308,N_2731);
nor U4972 (N_4972,N_3032,N_2905);
and U4973 (N_4973,N_2590,N_2987);
xor U4974 (N_4974,N_2547,N_2985);
xor U4975 (N_4975,N_2899,N_3691);
or U4976 (N_4976,N_2840,N_3635);
and U4977 (N_4977,N_3249,N_3523);
nand U4978 (N_4978,N_3489,N_3660);
xnor U4979 (N_4979,N_2915,N_2513);
and U4980 (N_4980,N_2753,N_3058);
nor U4981 (N_4981,N_2604,N_3065);
or U4982 (N_4982,N_2679,N_3249);
nand U4983 (N_4983,N_3637,N_3232);
nand U4984 (N_4984,N_2795,N_2977);
and U4985 (N_4985,N_3580,N_3330);
nor U4986 (N_4986,N_2997,N_3449);
nor U4987 (N_4987,N_2923,N_3258);
xnor U4988 (N_4988,N_3486,N_2596);
xnor U4989 (N_4989,N_3661,N_2693);
and U4990 (N_4990,N_3488,N_3420);
nor U4991 (N_4991,N_2939,N_3598);
or U4992 (N_4992,N_3657,N_2958);
nand U4993 (N_4993,N_3656,N_3504);
and U4994 (N_4994,N_3231,N_2663);
nand U4995 (N_4995,N_3104,N_3165);
xor U4996 (N_4996,N_2546,N_3140);
nor U4997 (N_4997,N_3488,N_3523);
and U4998 (N_4998,N_3154,N_3088);
nand U4999 (N_4999,N_2920,N_2812);
xnor U5000 (N_5000,N_4866,N_4565);
and U5001 (N_5001,N_4177,N_4399);
nand U5002 (N_5002,N_3831,N_4571);
xnor U5003 (N_5003,N_4311,N_4377);
nand U5004 (N_5004,N_4685,N_4484);
nor U5005 (N_5005,N_4445,N_4572);
nor U5006 (N_5006,N_4480,N_3773);
or U5007 (N_5007,N_4705,N_3941);
or U5008 (N_5008,N_3960,N_4440);
nand U5009 (N_5009,N_4890,N_4292);
xnor U5010 (N_5010,N_3842,N_4095);
nor U5011 (N_5011,N_4148,N_4842);
and U5012 (N_5012,N_4453,N_4619);
and U5013 (N_5013,N_4186,N_4670);
xnor U5014 (N_5014,N_4144,N_3926);
xor U5015 (N_5015,N_4225,N_4415);
xor U5016 (N_5016,N_4044,N_4644);
xnor U5017 (N_5017,N_3895,N_4636);
xnor U5018 (N_5018,N_3778,N_3966);
or U5019 (N_5019,N_4495,N_4403);
nor U5020 (N_5020,N_3907,N_4784);
nand U5021 (N_5021,N_4498,N_4859);
or U5022 (N_5022,N_4150,N_3997);
xnor U5023 (N_5023,N_4537,N_4991);
nand U5024 (N_5024,N_3770,N_4457);
nor U5025 (N_5025,N_4265,N_4492);
and U5026 (N_5026,N_4838,N_3756);
or U5027 (N_5027,N_3763,N_4740);
and U5028 (N_5028,N_4928,N_4826);
and U5029 (N_5029,N_4230,N_4205);
nor U5030 (N_5030,N_3987,N_3936);
nor U5031 (N_5031,N_4173,N_4601);
or U5032 (N_5032,N_4166,N_4902);
nor U5033 (N_5033,N_4794,N_4438);
and U5034 (N_5034,N_4620,N_4811);
or U5035 (N_5035,N_4764,N_4421);
and U5036 (N_5036,N_4692,N_4746);
nand U5037 (N_5037,N_4730,N_4924);
nor U5038 (N_5038,N_3788,N_4954);
or U5039 (N_5039,N_3802,N_4040);
nor U5040 (N_5040,N_3925,N_4960);
nand U5041 (N_5041,N_4101,N_4561);
and U5042 (N_5042,N_4455,N_4939);
nand U5043 (N_5043,N_4018,N_3977);
and U5044 (N_5044,N_4860,N_4391);
and U5045 (N_5045,N_4989,N_4988);
nor U5046 (N_5046,N_3912,N_4473);
xnor U5047 (N_5047,N_4791,N_4020);
nor U5048 (N_5048,N_4888,N_4809);
nand U5049 (N_5049,N_4726,N_4761);
or U5050 (N_5050,N_3794,N_4033);
and U5051 (N_5051,N_4518,N_4666);
nand U5052 (N_5052,N_3956,N_4779);
and U5053 (N_5053,N_4118,N_3806);
nand U5054 (N_5054,N_4376,N_3891);
nor U5055 (N_5055,N_4341,N_4560);
xor U5056 (N_5056,N_3863,N_3883);
xnor U5057 (N_5057,N_4734,N_3865);
or U5058 (N_5058,N_4822,N_3760);
nor U5059 (N_5059,N_3851,N_4886);
or U5060 (N_5060,N_4219,N_4336);
nand U5061 (N_5061,N_4626,N_4815);
xor U5062 (N_5062,N_4089,N_4743);
and U5063 (N_5063,N_4906,N_4994);
nand U5064 (N_5064,N_4270,N_4025);
and U5065 (N_5065,N_4060,N_4212);
nand U5066 (N_5066,N_3820,N_4789);
xor U5067 (N_5067,N_4370,N_4948);
nor U5068 (N_5068,N_4727,N_3896);
nand U5069 (N_5069,N_4539,N_4594);
xor U5070 (N_5070,N_4373,N_4675);
xor U5071 (N_5071,N_4722,N_4750);
nand U5072 (N_5072,N_4434,N_4963);
xnor U5073 (N_5073,N_4971,N_4299);
nor U5074 (N_5074,N_3877,N_4097);
nand U5075 (N_5075,N_3969,N_3939);
nor U5076 (N_5076,N_4679,N_4855);
and U5077 (N_5077,N_3971,N_4709);
nor U5078 (N_5078,N_4309,N_4523);
or U5079 (N_5079,N_3990,N_4153);
xor U5080 (N_5080,N_4072,N_4188);
or U5081 (N_5081,N_4303,N_4987);
nor U5082 (N_5082,N_4213,N_3991);
or U5083 (N_5083,N_3796,N_4437);
nor U5084 (N_5084,N_4057,N_3777);
nor U5085 (N_5085,N_4986,N_4277);
xor U5086 (N_5086,N_3949,N_4147);
nand U5087 (N_5087,N_4354,N_4613);
nor U5088 (N_5088,N_4725,N_4404);
xor U5089 (N_5089,N_4413,N_4853);
nor U5090 (N_5090,N_4375,N_4787);
and U5091 (N_5091,N_4946,N_4955);
nand U5092 (N_5092,N_4747,N_4306);
or U5093 (N_5093,N_4280,N_4107);
nand U5094 (N_5094,N_4231,N_4489);
xnor U5095 (N_5095,N_4351,N_4062);
nand U5096 (N_5096,N_4068,N_4580);
and U5097 (N_5097,N_4045,N_4076);
nor U5098 (N_5098,N_3935,N_4773);
or U5099 (N_5099,N_4202,N_4908);
or U5100 (N_5100,N_4331,N_4239);
xor U5101 (N_5101,N_4934,N_4801);
nor U5102 (N_5102,N_4246,N_4691);
or U5103 (N_5103,N_4003,N_4812);
xor U5104 (N_5104,N_3860,N_4783);
xor U5105 (N_5105,N_4884,N_4154);
xor U5106 (N_5106,N_4477,N_4897);
nor U5107 (N_5107,N_4481,N_4871);
nand U5108 (N_5108,N_4732,N_4925);
nand U5109 (N_5109,N_4968,N_4831);
nand U5110 (N_5110,N_4688,N_4632);
and U5111 (N_5111,N_4304,N_4417);
or U5112 (N_5112,N_3959,N_3767);
nor U5113 (N_5113,N_4138,N_4876);
or U5114 (N_5114,N_4329,N_3921);
nand U5115 (N_5115,N_4528,N_4942);
nor U5116 (N_5116,N_3750,N_4332);
xnor U5117 (N_5117,N_4302,N_4328);
nand U5118 (N_5118,N_4658,N_4111);
and U5119 (N_5119,N_4190,N_4360);
nand U5120 (N_5120,N_4568,N_4296);
xnor U5121 (N_5121,N_4476,N_4402);
nand U5122 (N_5122,N_4065,N_3849);
and U5123 (N_5123,N_3946,N_4012);
or U5124 (N_5124,N_4366,N_3898);
xnor U5125 (N_5125,N_4929,N_4651);
and U5126 (N_5126,N_4669,N_3948);
nor U5127 (N_5127,N_4913,N_3985);
or U5128 (N_5128,N_4979,N_4843);
nor U5129 (N_5129,N_4663,N_4485);
xor U5130 (N_5130,N_3902,N_4271);
or U5131 (N_5131,N_3759,N_4266);
nand U5132 (N_5132,N_4661,N_3850);
and U5133 (N_5133,N_4577,N_4869);
or U5134 (N_5134,N_4352,N_3869);
nor U5135 (N_5135,N_4662,N_4947);
and U5136 (N_5136,N_3995,N_4088);
nor U5137 (N_5137,N_4985,N_4878);
or U5138 (N_5138,N_3786,N_4597);
nand U5139 (N_5139,N_4185,N_4439);
nand U5140 (N_5140,N_4538,N_3817);
nand U5141 (N_5141,N_4106,N_3975);
and U5142 (N_5142,N_4610,N_4999);
xnor U5143 (N_5143,N_4034,N_4247);
nand U5144 (N_5144,N_3848,N_4255);
xor U5145 (N_5145,N_3903,N_4760);
xnor U5146 (N_5146,N_4983,N_3812);
xnor U5147 (N_5147,N_4562,N_4226);
and U5148 (N_5148,N_4140,N_3920);
xnor U5149 (N_5149,N_4972,N_4549);
nor U5150 (N_5150,N_4357,N_4788);
nor U5151 (N_5151,N_3847,N_4804);
or U5152 (N_5152,N_4317,N_4061);
nand U5153 (N_5153,N_4359,N_4011);
nand U5154 (N_5154,N_4193,N_4478);
nor U5155 (N_5155,N_4405,N_4083);
or U5156 (N_5156,N_4541,N_4700);
xnor U5157 (N_5157,N_4735,N_4608);
and U5158 (N_5158,N_4023,N_3843);
nand U5159 (N_5159,N_4390,N_3841);
or U5160 (N_5160,N_4507,N_4943);
and U5161 (N_5161,N_4337,N_4251);
or U5162 (N_5162,N_4527,N_4285);
or U5163 (N_5163,N_4508,N_3961);
xnor U5164 (N_5164,N_4338,N_4534);
nand U5165 (N_5165,N_4681,N_4981);
or U5166 (N_5166,N_4080,N_4487);
and U5167 (N_5167,N_4520,N_4069);
nor U5168 (N_5168,N_4491,N_4032);
nand U5169 (N_5169,N_3915,N_4459);
or U5170 (N_5170,N_4151,N_4005);
or U5171 (N_5171,N_4660,N_4475);
nand U5172 (N_5172,N_4930,N_4852);
or U5173 (N_5173,N_4659,N_3758);
nor U5174 (N_5174,N_3938,N_3889);
xnor U5175 (N_5175,N_4633,N_4813);
or U5176 (N_5176,N_4241,N_3928);
or U5177 (N_5177,N_4990,N_4259);
or U5178 (N_5178,N_4711,N_4575);
xnor U5179 (N_5179,N_4396,N_4622);
nand U5180 (N_5180,N_4428,N_4035);
xnor U5181 (N_5181,N_3774,N_4261);
xor U5182 (N_5182,N_4139,N_4053);
or U5183 (N_5183,N_3771,N_4300);
nor U5184 (N_5184,N_4919,N_4217);
and U5185 (N_5185,N_4710,N_4087);
nor U5186 (N_5186,N_4365,N_4828);
nand U5187 (N_5187,N_4287,N_3866);
or U5188 (N_5188,N_3810,N_4098);
nor U5189 (N_5189,N_4494,N_4236);
or U5190 (N_5190,N_4056,N_4599);
xor U5191 (N_5191,N_3840,N_4614);
xor U5192 (N_5192,N_4353,N_4808);
xnor U5193 (N_5193,N_3828,N_3862);
and U5194 (N_5194,N_4641,N_3798);
nand U5195 (N_5195,N_4016,N_4105);
xor U5196 (N_5196,N_4524,N_3845);
nand U5197 (N_5197,N_4100,N_4596);
xor U5198 (N_5198,N_4041,N_4310);
or U5199 (N_5199,N_4321,N_4368);
or U5200 (N_5200,N_4503,N_4689);
xnor U5201 (N_5201,N_4774,N_3830);
xor U5202 (N_5202,N_4465,N_4698);
xnor U5203 (N_5203,N_3881,N_4133);
xor U5204 (N_5204,N_4708,N_4081);
nand U5205 (N_5205,N_4501,N_4279);
and U5206 (N_5206,N_4850,N_4701);
or U5207 (N_5207,N_4249,N_4120);
or U5208 (N_5208,N_3807,N_4163);
and U5209 (N_5209,N_4851,N_4687);
nand U5210 (N_5210,N_3892,N_4298);
or U5211 (N_5211,N_4112,N_3854);
or U5212 (N_5212,N_4319,N_4218);
nor U5213 (N_5213,N_4274,N_4461);
nand U5214 (N_5214,N_4469,N_4532);
and U5215 (N_5215,N_4047,N_4414);
nor U5216 (N_5216,N_4637,N_3782);
and U5217 (N_5217,N_4579,N_4430);
nand U5218 (N_5218,N_4315,N_3914);
and U5219 (N_5219,N_4322,N_4993);
nor U5220 (N_5220,N_4982,N_4770);
nor U5221 (N_5221,N_4115,N_4778);
nor U5222 (N_5222,N_4880,N_4182);
or U5223 (N_5223,N_4733,N_4466);
and U5224 (N_5224,N_4731,N_4738);
or U5225 (N_5225,N_4326,N_4119);
or U5226 (N_5226,N_3870,N_4785);
nor U5227 (N_5227,N_3973,N_4482);
and U5228 (N_5228,N_4891,N_3775);
nand U5229 (N_5229,N_4867,N_4678);
and U5230 (N_5230,N_4936,N_4829);
nand U5231 (N_5231,N_4706,N_4776);
and U5232 (N_5232,N_4612,N_4167);
xor U5233 (N_5233,N_4894,N_4531);
nand U5234 (N_5234,N_4702,N_4171);
and U5235 (N_5235,N_4384,N_4806);
or U5236 (N_5236,N_3893,N_4419);
and U5237 (N_5237,N_4029,N_4195);
nor U5238 (N_5238,N_3876,N_4748);
nor U5239 (N_5239,N_4635,N_4209);
nand U5240 (N_5240,N_4868,N_4067);
nor U5241 (N_5241,N_4420,N_4237);
or U5242 (N_5242,N_4969,N_3814);
nor U5243 (N_5243,N_3999,N_3937);
nor U5244 (N_5244,N_4054,N_4912);
and U5245 (N_5245,N_4854,N_3924);
nand U5246 (N_5246,N_4515,N_3856);
nand U5247 (N_5247,N_4327,N_4961);
nor U5248 (N_5248,N_3943,N_4564);
or U5249 (N_5249,N_4937,N_4093);
xnor U5250 (N_5250,N_4559,N_4388);
xor U5251 (N_5251,N_4174,N_3931);
and U5252 (N_5252,N_4416,N_4634);
and U5253 (N_5253,N_4703,N_3789);
nor U5254 (N_5254,N_4526,N_4695);
or U5255 (N_5255,N_3779,N_3989);
nand U5256 (N_5256,N_4052,N_4940);
nand U5257 (N_5257,N_4381,N_4574);
or U5258 (N_5258,N_4629,N_4717);
or U5259 (N_5259,N_4668,N_4625);
nand U5260 (N_5260,N_4825,N_4066);
and U5261 (N_5261,N_3962,N_4452);
nor U5262 (N_5262,N_4566,N_4435);
nor U5263 (N_5263,N_4245,N_4471);
or U5264 (N_5264,N_3955,N_4349);
nand U5265 (N_5265,N_3905,N_4131);
and U5266 (N_5266,N_4109,N_4051);
nor U5267 (N_5267,N_4116,N_4429);
xor U5268 (N_5268,N_3981,N_4155);
xnor U5269 (N_5269,N_4922,N_4953);
and U5270 (N_5270,N_4649,N_4000);
xnor U5271 (N_5271,N_4143,N_4974);
nor U5272 (N_5272,N_4042,N_4938);
and U5273 (N_5273,N_4652,N_4552);
nor U5274 (N_5274,N_4578,N_4207);
nor U5275 (N_5275,N_4462,N_4673);
xnor U5276 (N_5276,N_4721,N_4158);
xor U5277 (N_5277,N_4753,N_4238);
or U5278 (N_5278,N_3769,N_3826);
or U5279 (N_5279,N_4345,N_3824);
nand U5280 (N_5280,N_4984,N_4858);
or U5281 (N_5281,N_3970,N_4426);
and U5282 (N_5282,N_3894,N_4078);
xnor U5283 (N_5283,N_4017,N_4130);
nand U5284 (N_5284,N_4911,N_4645);
nand U5285 (N_5285,N_4175,N_4995);
or U5286 (N_5286,N_4227,N_4063);
xnor U5287 (N_5287,N_4600,N_4903);
nor U5288 (N_5288,N_4224,N_4550);
nor U5289 (N_5289,N_3976,N_4581);
nor U5290 (N_5290,N_4313,N_3761);
or U5291 (N_5291,N_4113,N_4398);
or U5292 (N_5292,N_4022,N_4777);
and U5293 (N_5293,N_3916,N_3988);
nor U5294 (N_5294,N_4915,N_4917);
nor U5295 (N_5295,N_4514,N_4926);
and U5296 (N_5296,N_3954,N_4164);
xor U5297 (N_5297,N_4604,N_4046);
and U5298 (N_5298,N_3913,N_4099);
xnor U5299 (N_5299,N_4286,N_3986);
xor U5300 (N_5300,N_4257,N_4959);
and U5301 (N_5301,N_4921,N_4551);
xor U5302 (N_5302,N_4293,N_3792);
nor U5303 (N_5303,N_4425,N_4754);
or U5304 (N_5304,N_3901,N_4680);
nand U5305 (N_5305,N_4208,N_4244);
nor U5306 (N_5306,N_4933,N_4883);
and U5307 (N_5307,N_4820,N_4800);
nor U5308 (N_5308,N_4793,N_3780);
and U5309 (N_5309,N_4071,N_4281);
or U5310 (N_5310,N_4646,N_4607);
and U5311 (N_5311,N_4275,N_4010);
nand U5312 (N_5312,N_4588,N_3801);
or U5313 (N_5313,N_3952,N_4529);
or U5314 (N_5314,N_4656,N_4200);
nand U5315 (N_5315,N_4262,N_3923);
nand U5316 (N_5316,N_4104,N_4348);
and U5317 (N_5317,N_4795,N_3958);
or U5318 (N_5318,N_4102,N_4432);
xnor U5319 (N_5319,N_3996,N_3757);
or U5320 (N_5320,N_4611,N_4533);
xor U5321 (N_5321,N_4769,N_3839);
and U5322 (N_5322,N_4817,N_4371);
xnor U5323 (N_5323,N_4672,N_3776);
or U5324 (N_5324,N_4905,N_4001);
nor U5325 (N_5325,N_4665,N_4335);
xor U5326 (N_5326,N_4864,N_4179);
nor U5327 (N_5327,N_4519,N_4161);
or U5328 (N_5328,N_4240,N_4639);
nor U5329 (N_5329,N_3879,N_4308);
nand U5330 (N_5330,N_4235,N_4627);
nand U5331 (N_5331,N_4316,N_3787);
or U5332 (N_5332,N_3993,N_4768);
nor U5333 (N_5333,N_4856,N_4932);
xnor U5334 (N_5334,N_4904,N_4970);
nor U5335 (N_5335,N_4320,N_4254);
xor U5336 (N_5336,N_4467,N_4334);
xor U5337 (N_5337,N_4555,N_4406);
nor U5338 (N_5338,N_4058,N_4638);
nor U5339 (N_5339,N_4749,N_4759);
and U5340 (N_5340,N_4916,N_3852);
nor U5341 (N_5341,N_3880,N_4587);
xnor U5342 (N_5342,N_4879,N_4542);
nand U5343 (N_5343,N_3793,N_4616);
xnor U5344 (N_5344,N_4720,N_4422);
and U5345 (N_5345,N_4479,N_4499);
nor U5346 (N_5346,N_4350,N_4470);
and U5347 (N_5347,N_4301,N_3846);
nor U5348 (N_5348,N_4766,N_4818);
xnor U5349 (N_5349,N_4424,N_4497);
or U5350 (N_5350,N_4950,N_4075);
xor U5351 (N_5351,N_4729,N_4704);
and U5352 (N_5352,N_4008,N_4289);
or U5353 (N_5353,N_4372,N_3816);
nor U5354 (N_5354,N_3945,N_4914);
nor U5355 (N_5355,N_4126,N_4771);
or U5356 (N_5356,N_4603,N_4050);
nand U5357 (N_5357,N_4004,N_4447);
xnor U5358 (N_5358,N_4535,N_3844);
nand U5359 (N_5359,N_4039,N_4964);
and U5360 (N_5360,N_4136,N_4650);
nand U5361 (N_5361,N_3800,N_4229);
and U5362 (N_5362,N_4975,N_4870);
xor U5363 (N_5363,N_4623,N_4324);
and U5364 (N_5364,N_4840,N_3822);
nand U5365 (N_5365,N_4211,N_4845);
and U5366 (N_5366,N_4282,N_4263);
nand U5367 (N_5367,N_4194,N_4456);
nand U5368 (N_5368,N_4253,N_3900);
or U5369 (N_5369,N_4090,N_4250);
and U5370 (N_5370,N_4583,N_4573);
or U5371 (N_5371,N_4189,N_3835);
xor U5372 (N_5372,N_4248,N_4128);
or U5373 (N_5373,N_4506,N_3825);
nand U5374 (N_5374,N_4693,N_4796);
nand U5375 (N_5375,N_3884,N_4183);
nor U5376 (N_5376,N_4418,N_4141);
nand U5377 (N_5377,N_4206,N_4899);
nand U5378 (N_5378,N_4944,N_4677);
nor U5379 (N_5379,N_3833,N_4595);
or U5380 (N_5380,N_4220,N_4460);
nand U5381 (N_5381,N_4443,N_4618);
or U5382 (N_5382,N_4885,N_3963);
nand U5383 (N_5383,N_3932,N_4361);
or U5384 (N_5384,N_4187,N_4997);
nand U5385 (N_5385,N_4221,N_4387);
or U5386 (N_5386,N_4273,N_4493);
nand U5387 (N_5387,N_4841,N_4043);
or U5388 (N_5388,N_4745,N_4865);
nand U5389 (N_5389,N_4333,N_4536);
nand U5390 (N_5390,N_4889,N_3772);
xnor U5391 (N_5391,N_4135,N_4294);
nand U5392 (N_5392,N_4874,N_4123);
xor U5393 (N_5393,N_4742,N_4160);
xor U5394 (N_5394,N_3911,N_3868);
nor U5395 (N_5395,N_3836,N_3904);
or U5396 (N_5396,N_3957,N_4516);
xor U5397 (N_5397,N_3875,N_4631);
nand U5398 (N_5398,N_3783,N_3813);
and U5399 (N_5399,N_3853,N_4048);
and U5400 (N_5400,N_4228,N_4875);
or U5401 (N_5401,N_4821,N_4762);
nor U5402 (N_5402,N_3878,N_4472);
nor U5403 (N_5403,N_4395,N_4367);
and U5404 (N_5404,N_3818,N_4307);
xor U5405 (N_5405,N_4980,N_4602);
nor U5406 (N_5406,N_3858,N_4628);
or U5407 (N_5407,N_4483,N_4243);
or U5408 (N_5408,N_3934,N_4512);
xnor U5409 (N_5409,N_4122,N_4682);
and U5410 (N_5410,N_4409,N_4802);
nand U5411 (N_5411,N_4664,N_4252);
nor U5412 (N_5412,N_4496,N_3834);
and U5413 (N_5413,N_4260,N_4444);
nor U5414 (N_5414,N_3927,N_4965);
xor U5415 (N_5415,N_3910,N_3809);
nand U5416 (N_5416,N_4397,N_4347);
nor U5417 (N_5417,N_4923,N_4276);
and U5418 (N_5418,N_4657,N_4323);
and U5419 (N_5419,N_4810,N_4737);
nand U5420 (N_5420,N_4697,N_4149);
or U5421 (N_5421,N_4269,N_4676);
nand U5422 (N_5422,N_4803,N_4907);
or U5423 (N_5423,N_4077,N_3765);
and U5424 (N_5424,N_4168,N_4379);
nand U5425 (N_5425,N_4758,N_4952);
or U5426 (N_5426,N_4807,N_4554);
nand U5427 (N_5427,N_4699,N_3753);
nand U5428 (N_5428,N_4198,N_4385);
or U5429 (N_5429,N_3811,N_4756);
or U5430 (N_5430,N_4744,N_4543);
and U5431 (N_5431,N_4007,N_4900);
nand U5432 (N_5432,N_4978,N_4103);
and U5433 (N_5433,N_4223,N_4145);
nor U5434 (N_5434,N_4584,N_4707);
nand U5435 (N_5435,N_4896,N_4451);
xnor U5436 (N_5436,N_4127,N_3887);
or U5437 (N_5437,N_3909,N_3947);
nand U5438 (N_5438,N_3754,N_4517);
xnor U5439 (N_5439,N_4191,N_3791);
xor U5440 (N_5440,N_4216,N_3980);
and U5441 (N_5441,N_4752,N_4192);
or U5442 (N_5442,N_3766,N_4958);
and U5443 (N_5443,N_4775,N_4522);
nand U5444 (N_5444,N_4165,N_4449);
xnor U5445 (N_5445,N_3953,N_4169);
and U5446 (N_5446,N_3908,N_4442);
nand U5447 (N_5447,N_3781,N_4598);
nand U5448 (N_5448,N_4159,N_4291);
nor U5449 (N_5449,N_4945,N_4129);
xnor U5450 (N_5450,N_4197,N_4064);
nor U5451 (N_5451,N_4640,N_4343);
xor U5452 (N_5452,N_4935,N_4015);
and U5453 (N_5453,N_4458,N_4872);
nand U5454 (N_5454,N_3872,N_4410);
or U5455 (N_5455,N_4002,N_4839);
and U5456 (N_5456,N_4655,N_4196);
nand U5457 (N_5457,N_4346,N_4992);
nor U5458 (N_5458,N_4427,N_4400);
and U5459 (N_5459,N_4910,N_4976);
nand U5460 (N_5460,N_4272,N_4079);
nor U5461 (N_5461,N_4530,N_4297);
xor U5462 (N_5462,N_4407,N_4038);
and U5463 (N_5463,N_4835,N_3982);
or U5464 (N_5464,N_4464,N_4757);
xor U5465 (N_5465,N_4718,N_3804);
nand U5466 (N_5466,N_4355,N_4998);
and U5467 (N_5467,N_3972,N_4833);
nand U5468 (N_5468,N_3944,N_4278);
nor U5469 (N_5469,N_4392,N_4436);
nor U5470 (N_5470,N_3967,N_4027);
nand U5471 (N_5471,N_4070,N_4049);
and U5472 (N_5472,N_4741,N_4882);
xnor U5473 (N_5473,N_4214,N_4755);
nor U5474 (N_5474,N_4210,N_4178);
nor U5475 (N_5475,N_3864,N_4152);
xor U5476 (N_5476,N_4956,N_3940);
xnor U5477 (N_5477,N_4096,N_3874);
and U5478 (N_5478,N_3838,N_4605);
or U5479 (N_5479,N_4569,N_4967);
nor U5480 (N_5480,N_4340,N_4585);
nor U5481 (N_5481,N_4823,N_4411);
xnor U5482 (N_5482,N_3998,N_3861);
nor U5483 (N_5483,N_4792,N_4268);
nand U5484 (N_5484,N_4026,N_4454);
or U5485 (N_5485,N_4146,N_4790);
nor U5486 (N_5486,N_4124,N_4949);
xnor U5487 (N_5487,N_4132,N_4318);
and U5488 (N_5488,N_4763,N_3917);
and U5489 (N_5489,N_4389,N_4684);
nor U5490 (N_5490,N_4504,N_4648);
xnor U5491 (N_5491,N_4203,N_3823);
nor U5492 (N_5492,N_4862,N_4846);
and U5493 (N_5493,N_3983,N_4814);
xnor U5494 (N_5494,N_3837,N_4877);
nand U5495 (N_5495,N_3829,N_4920);
or U5496 (N_5496,N_4547,N_4617);
or U5497 (N_5497,N_4591,N_4125);
nand U5498 (N_5498,N_4030,N_4448);
nor U5499 (N_5499,N_4401,N_4881);
xnor U5500 (N_5500,N_4713,N_3968);
xnor U5501 (N_5501,N_4824,N_4288);
or U5502 (N_5502,N_4085,N_3890);
nand U5503 (N_5503,N_3764,N_4582);
nor U5504 (N_5504,N_4314,N_4006);
xor U5505 (N_5505,N_4009,N_3797);
nor U5506 (N_5506,N_4798,N_4450);
and U5507 (N_5507,N_3951,N_3964);
xnor U5508 (N_5508,N_3942,N_3768);
nor U5509 (N_5509,N_4486,N_4715);
and U5510 (N_5510,N_4117,N_4844);
nor U5511 (N_5511,N_4511,N_4363);
and U5512 (N_5512,N_4525,N_4267);
or U5513 (N_5513,N_3873,N_4290);
and U5514 (N_5514,N_4739,N_4819);
and U5515 (N_5515,N_3979,N_4234);
nand U5516 (N_5516,N_4654,N_3974);
nand U5517 (N_5517,N_4201,N_4909);
nor U5518 (N_5518,N_4502,N_3808);
or U5519 (N_5519,N_4037,N_4674);
or U5520 (N_5520,N_4157,N_4723);
xor U5521 (N_5521,N_4284,N_4686);
xor U5522 (N_5522,N_4446,N_3751);
nand U5523 (N_5523,N_4513,N_4642);
or U5524 (N_5524,N_4545,N_4780);
or U5525 (N_5525,N_4567,N_4393);
nand U5526 (N_5526,N_4181,N_4505);
xnor U5527 (N_5527,N_4683,N_4358);
xor U5528 (N_5528,N_4394,N_4094);
nor U5529 (N_5529,N_3984,N_4898);
nor U5530 (N_5530,N_4772,N_4339);
and U5531 (N_5531,N_4589,N_4172);
nand U5532 (N_5532,N_4383,N_4615);
and U5533 (N_5533,N_3785,N_4962);
xnor U5534 (N_5534,N_4719,N_4816);
xnor U5535 (N_5535,N_4609,N_4647);
or U5536 (N_5536,N_4957,N_4378);
or U5537 (N_5537,N_4441,N_4621);
nand U5538 (N_5538,N_4423,N_4863);
nand U5539 (N_5539,N_3855,N_4356);
xor U5540 (N_5540,N_4295,N_4055);
and U5541 (N_5541,N_4861,N_4108);
and U5542 (N_5542,N_4592,N_4586);
or U5543 (N_5543,N_4176,N_4086);
xor U5544 (N_5544,N_3799,N_4857);
nand U5545 (N_5545,N_4204,N_4199);
nor U5546 (N_5546,N_4724,N_4031);
xnor U5547 (N_5547,N_4362,N_4074);
and U5548 (N_5548,N_4966,N_3922);
nor U5549 (N_5549,N_4563,N_3950);
and U5550 (N_5550,N_4590,N_3859);
or U5551 (N_5551,N_4797,N_4408);
or U5552 (N_5552,N_4593,N_4728);
nand U5553 (N_5553,N_4510,N_4073);
and U5554 (N_5554,N_4887,N_4156);
nor U5555 (N_5555,N_3994,N_4059);
nand U5556 (N_5556,N_4028,N_4781);
nor U5557 (N_5557,N_4142,N_4170);
or U5558 (N_5558,N_4036,N_4500);
or U5559 (N_5559,N_4712,N_3918);
and U5560 (N_5560,N_4330,N_3857);
xnor U5561 (N_5561,N_4488,N_4019);
or U5562 (N_5562,N_4941,N_4834);
nor U5563 (N_5563,N_4873,N_4233);
and U5564 (N_5564,N_3886,N_4468);
or U5565 (N_5565,N_4630,N_3867);
and U5566 (N_5566,N_4973,N_4386);
xor U5567 (N_5567,N_3784,N_4977);
nor U5568 (N_5568,N_4024,N_4463);
xnor U5569 (N_5569,N_4380,N_4256);
xor U5570 (N_5570,N_4714,N_3882);
nor U5571 (N_5571,N_4767,N_4222);
nor U5572 (N_5572,N_4895,N_4624);
nor U5573 (N_5573,N_4013,N_4548);
and U5574 (N_5574,N_3978,N_4474);
xor U5575 (N_5575,N_4557,N_3871);
xnor U5576 (N_5576,N_4325,N_4558);
xnor U5577 (N_5577,N_4431,N_4927);
or U5578 (N_5578,N_4110,N_4951);
nand U5579 (N_5579,N_4799,N_4344);
nand U5580 (N_5580,N_4232,N_3805);
nor U5581 (N_5581,N_4137,N_4892);
and U5582 (N_5582,N_4342,N_4751);
nor U5583 (N_5583,N_4509,N_4305);
nor U5584 (N_5584,N_4258,N_3897);
nor U5585 (N_5585,N_3755,N_4283);
and U5586 (N_5586,N_3815,N_4805);
nor U5587 (N_5587,N_4082,N_4671);
nand U5588 (N_5588,N_3885,N_4832);
nor U5589 (N_5589,N_4643,N_3899);
and U5590 (N_5590,N_4836,N_3832);
or U5591 (N_5591,N_4716,N_4134);
nor U5592 (N_5592,N_4848,N_4931);
xor U5593 (N_5593,N_4736,N_3821);
xor U5594 (N_5594,N_4606,N_4570);
or U5595 (N_5595,N_4765,N_4546);
nor U5596 (N_5596,N_4369,N_4184);
or U5597 (N_5597,N_4690,N_3752);
nand U5598 (N_5598,N_4215,N_4312);
and U5599 (N_5599,N_4382,N_3919);
xnor U5600 (N_5600,N_4242,N_4830);
and U5601 (N_5601,N_4162,N_4553);
and U5602 (N_5602,N_4786,N_4490);
or U5603 (N_5603,N_4918,N_4782);
or U5604 (N_5604,N_4540,N_3930);
and U5605 (N_5605,N_4901,N_3888);
xor U5606 (N_5606,N_4653,N_4180);
nor U5607 (N_5607,N_4667,N_4014);
nand U5608 (N_5608,N_3819,N_3827);
nor U5609 (N_5609,N_4412,N_3906);
nor U5610 (N_5610,N_3790,N_3965);
nor U5611 (N_5611,N_4556,N_4374);
nor U5612 (N_5612,N_4084,N_4433);
nand U5613 (N_5613,N_4837,N_4121);
or U5614 (N_5614,N_3762,N_4893);
and U5615 (N_5615,N_4264,N_4827);
or U5616 (N_5616,N_4996,N_4849);
or U5617 (N_5617,N_4521,N_3929);
or U5618 (N_5618,N_4696,N_4092);
or U5619 (N_5619,N_3933,N_4091);
xnor U5620 (N_5620,N_4364,N_4114);
or U5621 (N_5621,N_3795,N_4694);
nand U5622 (N_5622,N_4847,N_3803);
nor U5623 (N_5623,N_4021,N_4576);
or U5624 (N_5624,N_3992,N_4544);
nor U5625 (N_5625,N_4013,N_3936);
and U5626 (N_5626,N_4432,N_4072);
and U5627 (N_5627,N_4831,N_4589);
nand U5628 (N_5628,N_4489,N_3904);
nor U5629 (N_5629,N_4954,N_4085);
nand U5630 (N_5630,N_4459,N_4604);
and U5631 (N_5631,N_4873,N_4184);
or U5632 (N_5632,N_3906,N_4254);
nand U5633 (N_5633,N_3983,N_4047);
xor U5634 (N_5634,N_4005,N_4596);
nor U5635 (N_5635,N_4971,N_4564);
or U5636 (N_5636,N_4816,N_4856);
nand U5637 (N_5637,N_3874,N_4199);
nor U5638 (N_5638,N_4735,N_4597);
nand U5639 (N_5639,N_4590,N_4524);
and U5640 (N_5640,N_4816,N_3977);
nor U5641 (N_5641,N_4624,N_4348);
or U5642 (N_5642,N_4372,N_4324);
nand U5643 (N_5643,N_4427,N_4918);
nor U5644 (N_5644,N_4417,N_3829);
and U5645 (N_5645,N_4201,N_4106);
nor U5646 (N_5646,N_4353,N_4682);
nand U5647 (N_5647,N_4664,N_4295);
and U5648 (N_5648,N_4121,N_4762);
or U5649 (N_5649,N_4995,N_4327);
nand U5650 (N_5650,N_4061,N_4470);
and U5651 (N_5651,N_4396,N_4595);
and U5652 (N_5652,N_4207,N_3767);
xnor U5653 (N_5653,N_4642,N_4240);
nor U5654 (N_5654,N_4794,N_4947);
nand U5655 (N_5655,N_4879,N_4236);
nor U5656 (N_5656,N_4203,N_4011);
or U5657 (N_5657,N_4428,N_4165);
and U5658 (N_5658,N_4841,N_3921);
nor U5659 (N_5659,N_4894,N_4076);
nor U5660 (N_5660,N_4678,N_4025);
nor U5661 (N_5661,N_4789,N_4609);
nand U5662 (N_5662,N_4572,N_4585);
or U5663 (N_5663,N_3772,N_3977);
xnor U5664 (N_5664,N_4296,N_3949);
xnor U5665 (N_5665,N_4417,N_4832);
or U5666 (N_5666,N_3956,N_4504);
nor U5667 (N_5667,N_4612,N_4834);
and U5668 (N_5668,N_3759,N_4745);
xnor U5669 (N_5669,N_4587,N_4972);
and U5670 (N_5670,N_4770,N_4812);
or U5671 (N_5671,N_3907,N_3980);
nand U5672 (N_5672,N_4238,N_4130);
or U5673 (N_5673,N_4627,N_4900);
nor U5674 (N_5674,N_4082,N_4958);
xor U5675 (N_5675,N_4593,N_4912);
nor U5676 (N_5676,N_4042,N_4959);
or U5677 (N_5677,N_4926,N_4245);
or U5678 (N_5678,N_4509,N_4838);
nor U5679 (N_5679,N_4469,N_4926);
nor U5680 (N_5680,N_4654,N_4651);
nand U5681 (N_5681,N_4655,N_3879);
or U5682 (N_5682,N_4426,N_3961);
and U5683 (N_5683,N_4921,N_4043);
or U5684 (N_5684,N_3892,N_4210);
xor U5685 (N_5685,N_4821,N_4891);
or U5686 (N_5686,N_3947,N_4153);
nand U5687 (N_5687,N_4913,N_4403);
nor U5688 (N_5688,N_4795,N_3890);
nand U5689 (N_5689,N_4556,N_4489);
or U5690 (N_5690,N_4643,N_3836);
nand U5691 (N_5691,N_3773,N_4599);
nor U5692 (N_5692,N_4139,N_3922);
and U5693 (N_5693,N_3997,N_4664);
or U5694 (N_5694,N_4110,N_4611);
nor U5695 (N_5695,N_4175,N_4041);
nand U5696 (N_5696,N_4688,N_3784);
or U5697 (N_5697,N_3796,N_4512);
or U5698 (N_5698,N_4447,N_4304);
xnor U5699 (N_5699,N_4934,N_4220);
nor U5700 (N_5700,N_4248,N_4515);
nor U5701 (N_5701,N_4970,N_4155);
nand U5702 (N_5702,N_4362,N_4680);
xor U5703 (N_5703,N_3771,N_4638);
nor U5704 (N_5704,N_4259,N_4134);
nor U5705 (N_5705,N_4545,N_4868);
nor U5706 (N_5706,N_4509,N_4920);
or U5707 (N_5707,N_4512,N_4230);
xor U5708 (N_5708,N_4428,N_4096);
xnor U5709 (N_5709,N_3778,N_4547);
or U5710 (N_5710,N_4314,N_4330);
xor U5711 (N_5711,N_4652,N_4141);
nand U5712 (N_5712,N_3754,N_4401);
and U5713 (N_5713,N_4521,N_4768);
xor U5714 (N_5714,N_4053,N_4003);
and U5715 (N_5715,N_4339,N_4139);
nor U5716 (N_5716,N_4242,N_3907);
xor U5717 (N_5717,N_4932,N_4060);
or U5718 (N_5718,N_4887,N_3994);
or U5719 (N_5719,N_4343,N_4189);
or U5720 (N_5720,N_4781,N_4931);
xor U5721 (N_5721,N_4377,N_4033);
nor U5722 (N_5722,N_4390,N_4110);
nor U5723 (N_5723,N_3907,N_4371);
nor U5724 (N_5724,N_4304,N_4710);
and U5725 (N_5725,N_4852,N_4776);
xor U5726 (N_5726,N_4872,N_4928);
and U5727 (N_5727,N_4761,N_4357);
or U5728 (N_5728,N_4062,N_4931);
nand U5729 (N_5729,N_4342,N_4053);
or U5730 (N_5730,N_4217,N_4110);
nor U5731 (N_5731,N_4307,N_3762);
nand U5732 (N_5732,N_3909,N_4607);
xor U5733 (N_5733,N_4988,N_4470);
nor U5734 (N_5734,N_4965,N_4750);
nand U5735 (N_5735,N_4765,N_4897);
nand U5736 (N_5736,N_4259,N_4064);
nand U5737 (N_5737,N_4851,N_4309);
and U5738 (N_5738,N_3926,N_4908);
or U5739 (N_5739,N_4627,N_4130);
and U5740 (N_5740,N_3797,N_4536);
nor U5741 (N_5741,N_4764,N_4806);
xnor U5742 (N_5742,N_4576,N_4085);
xnor U5743 (N_5743,N_4734,N_4735);
xor U5744 (N_5744,N_3820,N_4912);
nand U5745 (N_5745,N_3975,N_4265);
and U5746 (N_5746,N_4428,N_4587);
or U5747 (N_5747,N_4147,N_4928);
xnor U5748 (N_5748,N_4851,N_4046);
nor U5749 (N_5749,N_4657,N_4603);
xor U5750 (N_5750,N_4912,N_4505);
xor U5751 (N_5751,N_4431,N_3888);
nor U5752 (N_5752,N_4149,N_4365);
or U5753 (N_5753,N_4645,N_4048);
xor U5754 (N_5754,N_3802,N_4778);
or U5755 (N_5755,N_4543,N_4800);
and U5756 (N_5756,N_4685,N_4409);
nand U5757 (N_5757,N_4054,N_4869);
nand U5758 (N_5758,N_4604,N_4661);
nand U5759 (N_5759,N_3892,N_4918);
nor U5760 (N_5760,N_4140,N_3963);
xnor U5761 (N_5761,N_4623,N_4069);
nor U5762 (N_5762,N_4079,N_4736);
and U5763 (N_5763,N_4321,N_4086);
nand U5764 (N_5764,N_4985,N_4788);
nor U5765 (N_5765,N_4191,N_4952);
nor U5766 (N_5766,N_4458,N_4807);
xnor U5767 (N_5767,N_4161,N_3851);
and U5768 (N_5768,N_4155,N_4513);
xor U5769 (N_5769,N_4979,N_4903);
or U5770 (N_5770,N_4288,N_3827);
xor U5771 (N_5771,N_4388,N_4631);
xor U5772 (N_5772,N_3980,N_4784);
xor U5773 (N_5773,N_3814,N_4898);
and U5774 (N_5774,N_4373,N_4354);
and U5775 (N_5775,N_4574,N_3845);
or U5776 (N_5776,N_3828,N_4955);
and U5777 (N_5777,N_3870,N_4426);
xnor U5778 (N_5778,N_4361,N_3799);
and U5779 (N_5779,N_4027,N_4719);
nor U5780 (N_5780,N_3788,N_3948);
nor U5781 (N_5781,N_4545,N_4069);
and U5782 (N_5782,N_4588,N_3885);
or U5783 (N_5783,N_4353,N_4062);
and U5784 (N_5784,N_4262,N_4457);
xnor U5785 (N_5785,N_4270,N_4680);
nor U5786 (N_5786,N_4249,N_4973);
nor U5787 (N_5787,N_4573,N_4179);
nor U5788 (N_5788,N_4922,N_4517);
nand U5789 (N_5789,N_4872,N_4582);
nand U5790 (N_5790,N_4844,N_4578);
nand U5791 (N_5791,N_3890,N_3896);
or U5792 (N_5792,N_4896,N_4467);
xnor U5793 (N_5793,N_4989,N_4827);
or U5794 (N_5794,N_4192,N_4621);
and U5795 (N_5795,N_4200,N_4519);
and U5796 (N_5796,N_4072,N_4993);
nor U5797 (N_5797,N_4085,N_3776);
nor U5798 (N_5798,N_4426,N_3843);
xor U5799 (N_5799,N_4996,N_4323);
xnor U5800 (N_5800,N_4188,N_4393);
and U5801 (N_5801,N_4159,N_4626);
nor U5802 (N_5802,N_4350,N_4577);
or U5803 (N_5803,N_4842,N_4787);
xor U5804 (N_5804,N_4331,N_4447);
nand U5805 (N_5805,N_3904,N_4497);
nand U5806 (N_5806,N_4038,N_3831);
nand U5807 (N_5807,N_4250,N_3938);
xnor U5808 (N_5808,N_4326,N_4105);
xor U5809 (N_5809,N_4514,N_4043);
xnor U5810 (N_5810,N_3851,N_4608);
and U5811 (N_5811,N_4718,N_4304);
nor U5812 (N_5812,N_4830,N_4917);
or U5813 (N_5813,N_4136,N_4769);
nand U5814 (N_5814,N_4812,N_4057);
nand U5815 (N_5815,N_3813,N_4715);
nand U5816 (N_5816,N_4342,N_4586);
and U5817 (N_5817,N_3888,N_4760);
nor U5818 (N_5818,N_4040,N_4523);
nand U5819 (N_5819,N_3967,N_3957);
or U5820 (N_5820,N_4588,N_3922);
nand U5821 (N_5821,N_4277,N_4300);
and U5822 (N_5822,N_4751,N_4650);
nor U5823 (N_5823,N_4074,N_3881);
nand U5824 (N_5824,N_4612,N_4760);
or U5825 (N_5825,N_4957,N_4936);
nor U5826 (N_5826,N_3947,N_4266);
xnor U5827 (N_5827,N_4253,N_4621);
and U5828 (N_5828,N_3806,N_3998);
and U5829 (N_5829,N_4406,N_4354);
xor U5830 (N_5830,N_3947,N_4423);
or U5831 (N_5831,N_4609,N_4166);
nor U5832 (N_5832,N_4719,N_4708);
nor U5833 (N_5833,N_4278,N_4347);
nand U5834 (N_5834,N_4615,N_4488);
nor U5835 (N_5835,N_4767,N_4087);
nor U5836 (N_5836,N_4101,N_4517);
or U5837 (N_5837,N_3833,N_4041);
xor U5838 (N_5838,N_4660,N_4935);
xor U5839 (N_5839,N_4170,N_4398);
or U5840 (N_5840,N_4952,N_4638);
nor U5841 (N_5841,N_4996,N_4034);
xor U5842 (N_5842,N_4838,N_4621);
nor U5843 (N_5843,N_4792,N_4235);
or U5844 (N_5844,N_4932,N_4273);
xnor U5845 (N_5845,N_4274,N_3971);
xor U5846 (N_5846,N_4029,N_4863);
and U5847 (N_5847,N_3925,N_4572);
and U5848 (N_5848,N_3922,N_4383);
and U5849 (N_5849,N_4060,N_4405);
and U5850 (N_5850,N_4343,N_3924);
xor U5851 (N_5851,N_4035,N_4957);
xor U5852 (N_5852,N_3937,N_4613);
and U5853 (N_5853,N_4818,N_3959);
and U5854 (N_5854,N_4804,N_4215);
nor U5855 (N_5855,N_3774,N_4205);
and U5856 (N_5856,N_4143,N_4457);
and U5857 (N_5857,N_4703,N_4295);
nor U5858 (N_5858,N_4438,N_4692);
and U5859 (N_5859,N_4065,N_3975);
xor U5860 (N_5860,N_3862,N_4759);
nor U5861 (N_5861,N_4396,N_3813);
nand U5862 (N_5862,N_4888,N_4474);
xnor U5863 (N_5863,N_4475,N_4265);
and U5864 (N_5864,N_4183,N_4467);
nand U5865 (N_5865,N_4805,N_4232);
or U5866 (N_5866,N_4875,N_4587);
or U5867 (N_5867,N_4060,N_4656);
nor U5868 (N_5868,N_3882,N_4355);
and U5869 (N_5869,N_4074,N_4581);
nor U5870 (N_5870,N_4764,N_4395);
xnor U5871 (N_5871,N_3757,N_4380);
nor U5872 (N_5872,N_3978,N_4914);
and U5873 (N_5873,N_3810,N_4107);
nor U5874 (N_5874,N_4106,N_4087);
xnor U5875 (N_5875,N_4125,N_4876);
or U5876 (N_5876,N_3864,N_4494);
nor U5877 (N_5877,N_4798,N_4528);
xor U5878 (N_5878,N_4320,N_4430);
xor U5879 (N_5879,N_4225,N_4467);
xor U5880 (N_5880,N_4364,N_4600);
and U5881 (N_5881,N_4203,N_4613);
and U5882 (N_5882,N_4682,N_4841);
nor U5883 (N_5883,N_4507,N_4327);
and U5884 (N_5884,N_3803,N_4232);
or U5885 (N_5885,N_4595,N_3829);
nand U5886 (N_5886,N_4093,N_4430);
nor U5887 (N_5887,N_4836,N_3876);
and U5888 (N_5888,N_4336,N_4043);
nor U5889 (N_5889,N_4988,N_4100);
or U5890 (N_5890,N_4271,N_4784);
xnor U5891 (N_5891,N_4668,N_4565);
and U5892 (N_5892,N_4943,N_4773);
nor U5893 (N_5893,N_4649,N_3842);
nor U5894 (N_5894,N_4071,N_4864);
xor U5895 (N_5895,N_3976,N_4535);
nor U5896 (N_5896,N_4880,N_4945);
xor U5897 (N_5897,N_4922,N_4518);
xor U5898 (N_5898,N_3865,N_3919);
and U5899 (N_5899,N_4938,N_4559);
or U5900 (N_5900,N_4067,N_3895);
or U5901 (N_5901,N_4317,N_4886);
xor U5902 (N_5902,N_4903,N_4974);
xnor U5903 (N_5903,N_4101,N_4294);
or U5904 (N_5904,N_4270,N_4740);
nor U5905 (N_5905,N_4132,N_4718);
nand U5906 (N_5906,N_4786,N_4279);
and U5907 (N_5907,N_3883,N_4861);
nor U5908 (N_5908,N_4827,N_4188);
nor U5909 (N_5909,N_4552,N_4895);
nand U5910 (N_5910,N_4835,N_4971);
nand U5911 (N_5911,N_3785,N_3949);
nand U5912 (N_5912,N_3952,N_4969);
and U5913 (N_5913,N_3872,N_4919);
xor U5914 (N_5914,N_4941,N_3942);
xor U5915 (N_5915,N_4514,N_4137);
and U5916 (N_5916,N_3951,N_4247);
nor U5917 (N_5917,N_4174,N_4238);
and U5918 (N_5918,N_4541,N_4874);
and U5919 (N_5919,N_4612,N_4114);
nand U5920 (N_5920,N_3807,N_3981);
or U5921 (N_5921,N_4134,N_4658);
xnor U5922 (N_5922,N_4382,N_4078);
nand U5923 (N_5923,N_3994,N_4265);
xor U5924 (N_5924,N_4160,N_4981);
nand U5925 (N_5925,N_4619,N_4662);
nor U5926 (N_5926,N_4677,N_4670);
nand U5927 (N_5927,N_4085,N_4966);
and U5928 (N_5928,N_4017,N_4337);
nand U5929 (N_5929,N_3765,N_4464);
nor U5930 (N_5930,N_4254,N_3901);
nand U5931 (N_5931,N_4580,N_4959);
nand U5932 (N_5932,N_4428,N_4553);
nand U5933 (N_5933,N_4387,N_4755);
and U5934 (N_5934,N_4599,N_4936);
nand U5935 (N_5935,N_3941,N_4578);
and U5936 (N_5936,N_4475,N_4665);
or U5937 (N_5937,N_3785,N_4538);
and U5938 (N_5938,N_4347,N_4915);
nor U5939 (N_5939,N_4114,N_4047);
and U5940 (N_5940,N_3947,N_4771);
xnor U5941 (N_5941,N_4071,N_4773);
and U5942 (N_5942,N_4422,N_4573);
nand U5943 (N_5943,N_4900,N_4358);
nand U5944 (N_5944,N_3886,N_4481);
or U5945 (N_5945,N_4849,N_4555);
nor U5946 (N_5946,N_4045,N_4493);
nor U5947 (N_5947,N_4160,N_3837);
and U5948 (N_5948,N_4312,N_4616);
and U5949 (N_5949,N_4770,N_4768);
nor U5950 (N_5950,N_4098,N_4792);
nor U5951 (N_5951,N_4412,N_3974);
and U5952 (N_5952,N_3856,N_4432);
nor U5953 (N_5953,N_4510,N_4477);
and U5954 (N_5954,N_3896,N_4018);
xnor U5955 (N_5955,N_4892,N_4724);
nand U5956 (N_5956,N_3928,N_3787);
or U5957 (N_5957,N_4861,N_4251);
or U5958 (N_5958,N_4828,N_4952);
nor U5959 (N_5959,N_4067,N_4583);
and U5960 (N_5960,N_3802,N_3954);
nor U5961 (N_5961,N_4054,N_4135);
xor U5962 (N_5962,N_4071,N_4453);
and U5963 (N_5963,N_3758,N_4734);
nor U5964 (N_5964,N_4773,N_4702);
and U5965 (N_5965,N_4471,N_4134);
nand U5966 (N_5966,N_4160,N_4997);
nand U5967 (N_5967,N_4223,N_4462);
nor U5968 (N_5968,N_3767,N_4395);
nand U5969 (N_5969,N_4298,N_4351);
xor U5970 (N_5970,N_4615,N_4343);
or U5971 (N_5971,N_4481,N_4319);
nand U5972 (N_5972,N_4061,N_4920);
or U5973 (N_5973,N_4208,N_4508);
or U5974 (N_5974,N_4099,N_4529);
or U5975 (N_5975,N_4536,N_3773);
nor U5976 (N_5976,N_4718,N_4459);
or U5977 (N_5977,N_3922,N_4461);
and U5978 (N_5978,N_3851,N_4930);
nand U5979 (N_5979,N_4533,N_4479);
nand U5980 (N_5980,N_3946,N_4482);
nand U5981 (N_5981,N_4268,N_4953);
or U5982 (N_5982,N_4452,N_4285);
and U5983 (N_5983,N_4303,N_4691);
or U5984 (N_5984,N_4584,N_4237);
nand U5985 (N_5985,N_4035,N_3774);
xnor U5986 (N_5986,N_4126,N_4283);
nor U5987 (N_5987,N_3768,N_3895);
xnor U5988 (N_5988,N_4386,N_4151);
and U5989 (N_5989,N_4096,N_4366);
nor U5990 (N_5990,N_4512,N_3899);
and U5991 (N_5991,N_4104,N_4323);
xnor U5992 (N_5992,N_3833,N_4696);
and U5993 (N_5993,N_4136,N_4580);
xor U5994 (N_5994,N_3967,N_4152);
nand U5995 (N_5995,N_4815,N_4259);
and U5996 (N_5996,N_3879,N_4186);
nand U5997 (N_5997,N_4647,N_3832);
nand U5998 (N_5998,N_4414,N_4328);
xnor U5999 (N_5999,N_4155,N_4981);
or U6000 (N_6000,N_4371,N_4742);
nand U6001 (N_6001,N_4867,N_4375);
xnor U6002 (N_6002,N_4336,N_3777);
nor U6003 (N_6003,N_4275,N_4988);
nor U6004 (N_6004,N_4350,N_4649);
or U6005 (N_6005,N_4383,N_4827);
nor U6006 (N_6006,N_4318,N_3962);
nor U6007 (N_6007,N_3945,N_4613);
or U6008 (N_6008,N_4187,N_4260);
xor U6009 (N_6009,N_3837,N_4319);
xnor U6010 (N_6010,N_4695,N_4277);
and U6011 (N_6011,N_4592,N_3753);
or U6012 (N_6012,N_4726,N_4486);
or U6013 (N_6013,N_3797,N_4810);
xor U6014 (N_6014,N_3807,N_4672);
xnor U6015 (N_6015,N_3949,N_4318);
xnor U6016 (N_6016,N_4558,N_4229);
xor U6017 (N_6017,N_4839,N_4711);
xnor U6018 (N_6018,N_4307,N_4193);
nor U6019 (N_6019,N_3806,N_3993);
nand U6020 (N_6020,N_3877,N_4985);
xor U6021 (N_6021,N_4288,N_4721);
nor U6022 (N_6022,N_4134,N_4081);
and U6023 (N_6023,N_4473,N_4006);
or U6024 (N_6024,N_4052,N_3763);
nand U6025 (N_6025,N_4854,N_3875);
and U6026 (N_6026,N_4035,N_4181);
nor U6027 (N_6027,N_4798,N_4726);
and U6028 (N_6028,N_3866,N_4674);
nor U6029 (N_6029,N_3893,N_4546);
or U6030 (N_6030,N_4350,N_4778);
or U6031 (N_6031,N_3971,N_4476);
xor U6032 (N_6032,N_4855,N_4211);
nor U6033 (N_6033,N_3993,N_4526);
and U6034 (N_6034,N_4704,N_4770);
or U6035 (N_6035,N_4929,N_3957);
xnor U6036 (N_6036,N_4117,N_4923);
nor U6037 (N_6037,N_4104,N_4532);
or U6038 (N_6038,N_4928,N_4878);
nor U6039 (N_6039,N_4561,N_4741);
nor U6040 (N_6040,N_4561,N_4992);
nor U6041 (N_6041,N_4492,N_4866);
nor U6042 (N_6042,N_4117,N_4354);
nor U6043 (N_6043,N_3947,N_4106);
nor U6044 (N_6044,N_4314,N_4320);
nor U6045 (N_6045,N_3925,N_4371);
and U6046 (N_6046,N_4680,N_4702);
nand U6047 (N_6047,N_3967,N_4592);
nand U6048 (N_6048,N_4697,N_4653);
nor U6049 (N_6049,N_4250,N_4060);
or U6050 (N_6050,N_4741,N_3822);
nor U6051 (N_6051,N_4635,N_4741);
xor U6052 (N_6052,N_4284,N_3915);
nand U6053 (N_6053,N_4429,N_4682);
nand U6054 (N_6054,N_4678,N_4389);
or U6055 (N_6055,N_4558,N_3902);
nand U6056 (N_6056,N_4365,N_3856);
nand U6057 (N_6057,N_4185,N_4138);
and U6058 (N_6058,N_4879,N_3862);
or U6059 (N_6059,N_4050,N_4453);
xor U6060 (N_6060,N_4097,N_4312);
nor U6061 (N_6061,N_4009,N_4904);
nor U6062 (N_6062,N_4332,N_4920);
nor U6063 (N_6063,N_4654,N_4488);
nand U6064 (N_6064,N_3767,N_4391);
xnor U6065 (N_6065,N_4844,N_4396);
nor U6066 (N_6066,N_4623,N_4802);
and U6067 (N_6067,N_4544,N_3883);
nand U6068 (N_6068,N_4984,N_4516);
xor U6069 (N_6069,N_4389,N_4500);
xnor U6070 (N_6070,N_4252,N_4052);
nor U6071 (N_6071,N_3982,N_4659);
nor U6072 (N_6072,N_4572,N_4806);
xor U6073 (N_6073,N_4894,N_3968);
xnor U6074 (N_6074,N_4521,N_3944);
xor U6075 (N_6075,N_4450,N_4790);
nand U6076 (N_6076,N_4365,N_4927);
nand U6077 (N_6077,N_4188,N_4475);
nor U6078 (N_6078,N_3999,N_3799);
and U6079 (N_6079,N_4250,N_4129);
and U6080 (N_6080,N_3998,N_4139);
nand U6081 (N_6081,N_4575,N_4439);
nand U6082 (N_6082,N_4005,N_3802);
nor U6083 (N_6083,N_4860,N_4124);
or U6084 (N_6084,N_3981,N_4697);
nor U6085 (N_6085,N_4394,N_4994);
nand U6086 (N_6086,N_4976,N_4626);
and U6087 (N_6087,N_4336,N_4318);
nand U6088 (N_6088,N_4999,N_4632);
nand U6089 (N_6089,N_4151,N_4040);
or U6090 (N_6090,N_4831,N_4996);
xnor U6091 (N_6091,N_4092,N_4850);
and U6092 (N_6092,N_4856,N_4287);
or U6093 (N_6093,N_4016,N_4413);
or U6094 (N_6094,N_4236,N_4775);
nand U6095 (N_6095,N_4561,N_4226);
xor U6096 (N_6096,N_4570,N_4097);
or U6097 (N_6097,N_4595,N_4910);
or U6098 (N_6098,N_4123,N_4549);
and U6099 (N_6099,N_4335,N_4076);
or U6100 (N_6100,N_4632,N_4200);
or U6101 (N_6101,N_4331,N_3936);
or U6102 (N_6102,N_3981,N_4063);
and U6103 (N_6103,N_3760,N_4179);
or U6104 (N_6104,N_4881,N_4721);
xnor U6105 (N_6105,N_4593,N_3900);
and U6106 (N_6106,N_3840,N_4081);
nor U6107 (N_6107,N_4535,N_3951);
and U6108 (N_6108,N_3788,N_4746);
or U6109 (N_6109,N_3793,N_4176);
and U6110 (N_6110,N_3982,N_4613);
xor U6111 (N_6111,N_4075,N_3948);
nor U6112 (N_6112,N_4341,N_4116);
xor U6113 (N_6113,N_3969,N_3750);
nor U6114 (N_6114,N_4836,N_4565);
nor U6115 (N_6115,N_4450,N_4710);
xnor U6116 (N_6116,N_3818,N_4347);
nor U6117 (N_6117,N_3892,N_4004);
xnor U6118 (N_6118,N_4963,N_4940);
or U6119 (N_6119,N_4260,N_4901);
xnor U6120 (N_6120,N_4812,N_4754);
and U6121 (N_6121,N_4417,N_4536);
xnor U6122 (N_6122,N_4324,N_4314);
xnor U6123 (N_6123,N_4580,N_4329);
xnor U6124 (N_6124,N_4250,N_4239);
or U6125 (N_6125,N_4666,N_4067);
and U6126 (N_6126,N_4926,N_4933);
or U6127 (N_6127,N_3996,N_4581);
nor U6128 (N_6128,N_4245,N_4750);
nor U6129 (N_6129,N_4440,N_4384);
nand U6130 (N_6130,N_3830,N_4363);
xor U6131 (N_6131,N_4993,N_4704);
and U6132 (N_6132,N_4746,N_4921);
and U6133 (N_6133,N_4136,N_3754);
nand U6134 (N_6134,N_4518,N_3953);
and U6135 (N_6135,N_4007,N_4604);
and U6136 (N_6136,N_4643,N_4897);
nor U6137 (N_6137,N_3966,N_4352);
nand U6138 (N_6138,N_4979,N_3913);
or U6139 (N_6139,N_4002,N_4084);
xnor U6140 (N_6140,N_4677,N_4860);
xor U6141 (N_6141,N_3845,N_4834);
and U6142 (N_6142,N_4461,N_4727);
nand U6143 (N_6143,N_3760,N_3830);
or U6144 (N_6144,N_3991,N_3822);
xnor U6145 (N_6145,N_4228,N_4494);
and U6146 (N_6146,N_4545,N_4273);
nand U6147 (N_6147,N_4521,N_4418);
nor U6148 (N_6148,N_4887,N_4013);
nor U6149 (N_6149,N_4468,N_3978);
xor U6150 (N_6150,N_4031,N_3935);
or U6151 (N_6151,N_4833,N_4367);
nor U6152 (N_6152,N_3831,N_4271);
and U6153 (N_6153,N_4944,N_4703);
nand U6154 (N_6154,N_4233,N_3827);
xor U6155 (N_6155,N_4259,N_4151);
or U6156 (N_6156,N_4903,N_4031);
and U6157 (N_6157,N_4689,N_4232);
or U6158 (N_6158,N_4667,N_3862);
and U6159 (N_6159,N_4351,N_4313);
nor U6160 (N_6160,N_3826,N_4297);
and U6161 (N_6161,N_4054,N_4319);
and U6162 (N_6162,N_4707,N_4943);
or U6163 (N_6163,N_4154,N_4492);
nor U6164 (N_6164,N_4573,N_4977);
nand U6165 (N_6165,N_3844,N_4497);
and U6166 (N_6166,N_4354,N_4463);
or U6167 (N_6167,N_4472,N_4209);
xnor U6168 (N_6168,N_4054,N_4183);
and U6169 (N_6169,N_4915,N_4344);
or U6170 (N_6170,N_4889,N_4265);
and U6171 (N_6171,N_4510,N_4237);
xnor U6172 (N_6172,N_4815,N_4990);
and U6173 (N_6173,N_4628,N_4730);
nor U6174 (N_6174,N_4391,N_4553);
or U6175 (N_6175,N_4640,N_4832);
nor U6176 (N_6176,N_4485,N_4180);
nor U6177 (N_6177,N_4865,N_3823);
or U6178 (N_6178,N_4688,N_4390);
nor U6179 (N_6179,N_3966,N_4324);
nor U6180 (N_6180,N_4900,N_4815);
or U6181 (N_6181,N_3859,N_4305);
or U6182 (N_6182,N_4268,N_4718);
or U6183 (N_6183,N_3909,N_3840);
and U6184 (N_6184,N_4643,N_4116);
or U6185 (N_6185,N_4825,N_3984);
xor U6186 (N_6186,N_4879,N_4677);
or U6187 (N_6187,N_4941,N_3994);
and U6188 (N_6188,N_4008,N_3861);
and U6189 (N_6189,N_4675,N_4746);
xnor U6190 (N_6190,N_4924,N_4706);
xnor U6191 (N_6191,N_4616,N_4723);
and U6192 (N_6192,N_4892,N_4046);
or U6193 (N_6193,N_4936,N_4225);
xor U6194 (N_6194,N_4399,N_4847);
nor U6195 (N_6195,N_3818,N_3858);
and U6196 (N_6196,N_4311,N_4571);
xor U6197 (N_6197,N_3886,N_4924);
or U6198 (N_6198,N_4786,N_4788);
xnor U6199 (N_6199,N_4398,N_3870);
xnor U6200 (N_6200,N_4349,N_4567);
or U6201 (N_6201,N_4162,N_4779);
xnor U6202 (N_6202,N_4309,N_4655);
or U6203 (N_6203,N_4270,N_4045);
or U6204 (N_6204,N_4607,N_4564);
xor U6205 (N_6205,N_4595,N_4457);
or U6206 (N_6206,N_3987,N_3848);
or U6207 (N_6207,N_4474,N_3903);
nand U6208 (N_6208,N_4850,N_4218);
nor U6209 (N_6209,N_4205,N_4103);
xnor U6210 (N_6210,N_4591,N_4981);
and U6211 (N_6211,N_4159,N_4492);
nand U6212 (N_6212,N_4464,N_4094);
and U6213 (N_6213,N_4525,N_4304);
or U6214 (N_6214,N_4032,N_4220);
or U6215 (N_6215,N_4619,N_4714);
xor U6216 (N_6216,N_4471,N_4364);
and U6217 (N_6217,N_4123,N_4987);
nor U6218 (N_6218,N_3889,N_4996);
or U6219 (N_6219,N_3861,N_4764);
or U6220 (N_6220,N_3842,N_4196);
and U6221 (N_6221,N_4002,N_3977);
and U6222 (N_6222,N_3979,N_4665);
nand U6223 (N_6223,N_4532,N_4112);
xnor U6224 (N_6224,N_4271,N_4738);
nor U6225 (N_6225,N_4119,N_3785);
or U6226 (N_6226,N_4371,N_4550);
nor U6227 (N_6227,N_4538,N_4456);
xnor U6228 (N_6228,N_4061,N_4296);
nor U6229 (N_6229,N_4041,N_4728);
and U6230 (N_6230,N_4268,N_4036);
xor U6231 (N_6231,N_4294,N_4649);
xnor U6232 (N_6232,N_3759,N_4552);
nand U6233 (N_6233,N_4712,N_4732);
xor U6234 (N_6234,N_4436,N_4595);
nand U6235 (N_6235,N_4379,N_4607);
and U6236 (N_6236,N_3765,N_4909);
nor U6237 (N_6237,N_3846,N_4337);
or U6238 (N_6238,N_3878,N_4266);
nor U6239 (N_6239,N_4378,N_4603);
nor U6240 (N_6240,N_4841,N_3777);
and U6241 (N_6241,N_4853,N_4755);
nand U6242 (N_6242,N_4381,N_4883);
and U6243 (N_6243,N_4034,N_4262);
xor U6244 (N_6244,N_4413,N_4512);
nor U6245 (N_6245,N_4042,N_4691);
nor U6246 (N_6246,N_4452,N_3948);
nand U6247 (N_6247,N_4045,N_4039);
xnor U6248 (N_6248,N_4345,N_4515);
and U6249 (N_6249,N_4876,N_3820);
and U6250 (N_6250,N_5523,N_5287);
nor U6251 (N_6251,N_5850,N_5646);
and U6252 (N_6252,N_6122,N_6120);
xor U6253 (N_6253,N_5012,N_5201);
nor U6254 (N_6254,N_5694,N_5993);
nor U6255 (N_6255,N_5574,N_5038);
or U6256 (N_6256,N_5578,N_6226);
nand U6257 (N_6257,N_5693,N_5063);
or U6258 (N_6258,N_6072,N_5653);
nor U6259 (N_6259,N_6092,N_5582);
and U6260 (N_6260,N_5099,N_5974);
nor U6261 (N_6261,N_5129,N_6210);
and U6262 (N_6262,N_5948,N_5704);
and U6263 (N_6263,N_5103,N_5042);
nand U6264 (N_6264,N_5961,N_5673);
nor U6265 (N_6265,N_5313,N_5527);
and U6266 (N_6266,N_5194,N_6194);
or U6267 (N_6267,N_5290,N_5700);
nand U6268 (N_6268,N_5973,N_5713);
and U6269 (N_6269,N_5421,N_5737);
nand U6270 (N_6270,N_5598,N_5772);
nand U6271 (N_6271,N_5108,N_5798);
or U6272 (N_6272,N_5849,N_5390);
and U6273 (N_6273,N_6112,N_5327);
nor U6274 (N_6274,N_5599,N_5770);
xnor U6275 (N_6275,N_5956,N_5371);
xnor U6276 (N_6276,N_5433,N_5138);
nand U6277 (N_6277,N_5116,N_5286);
and U6278 (N_6278,N_6055,N_5724);
or U6279 (N_6279,N_6063,N_5660);
nor U6280 (N_6280,N_6191,N_5796);
or U6281 (N_6281,N_6236,N_6169);
or U6282 (N_6282,N_5469,N_5615);
nand U6283 (N_6283,N_5228,N_5324);
xnor U6284 (N_6284,N_5592,N_5377);
nand U6285 (N_6285,N_5905,N_5268);
xnor U6286 (N_6286,N_5087,N_5546);
xor U6287 (N_6287,N_6244,N_5271);
or U6288 (N_6288,N_6080,N_5786);
and U6289 (N_6289,N_5581,N_5213);
xor U6290 (N_6290,N_5586,N_5720);
or U6291 (N_6291,N_5912,N_5818);
nor U6292 (N_6292,N_5101,N_5497);
or U6293 (N_6293,N_5998,N_5435);
xor U6294 (N_6294,N_5193,N_5519);
nand U6295 (N_6295,N_5965,N_6139);
xor U6296 (N_6296,N_6059,N_5983);
or U6297 (N_6297,N_5662,N_6104);
or U6298 (N_6298,N_5924,N_5621);
nor U6299 (N_6299,N_5488,N_5867);
and U6300 (N_6300,N_5507,N_5580);
nor U6301 (N_6301,N_5367,N_5057);
or U6302 (N_6302,N_6167,N_5024);
nor U6303 (N_6303,N_5452,N_5455);
or U6304 (N_6304,N_5141,N_5957);
xor U6305 (N_6305,N_5337,N_5557);
and U6306 (N_6306,N_5828,N_5872);
or U6307 (N_6307,N_6188,N_5757);
and U6308 (N_6308,N_5127,N_6027);
xor U6309 (N_6309,N_5902,N_5645);
nand U6310 (N_6310,N_5603,N_5449);
or U6311 (N_6311,N_5280,N_5665);
nand U6312 (N_6312,N_5445,N_5172);
nand U6313 (N_6313,N_5352,N_6213);
and U6314 (N_6314,N_5545,N_5035);
and U6315 (N_6315,N_5089,N_5827);
xor U6316 (N_6316,N_5779,N_5190);
and U6317 (N_6317,N_5356,N_5289);
nor U6318 (N_6318,N_5782,N_6121);
xor U6319 (N_6319,N_5636,N_5878);
or U6320 (N_6320,N_5418,N_5602);
and U6321 (N_6321,N_5230,N_5282);
nand U6322 (N_6322,N_6000,N_5382);
nor U6323 (N_6323,N_5078,N_5852);
nand U6324 (N_6324,N_5162,N_6175);
or U6325 (N_6325,N_5503,N_5526);
and U6326 (N_6326,N_6118,N_5404);
and U6327 (N_6327,N_5016,N_5717);
nand U6328 (N_6328,N_6046,N_5736);
nor U6329 (N_6329,N_5262,N_6102);
or U6330 (N_6330,N_6200,N_5837);
or U6331 (N_6331,N_6076,N_5628);
nor U6332 (N_6332,N_5409,N_6119);
or U6333 (N_6333,N_6151,N_5699);
and U6334 (N_6334,N_6128,N_5734);
nor U6335 (N_6335,N_5088,N_5184);
and U6336 (N_6336,N_5284,N_5774);
xnor U6337 (N_6337,N_5761,N_5627);
xnor U6338 (N_6338,N_5319,N_5363);
or U6339 (N_6339,N_6212,N_5590);
nor U6340 (N_6340,N_5408,N_5933);
xnor U6341 (N_6341,N_5113,N_5369);
xnor U6342 (N_6342,N_5744,N_6068);
nand U6343 (N_6343,N_6029,N_5906);
nand U6344 (N_6344,N_5611,N_5056);
xor U6345 (N_6345,N_6131,N_5986);
and U6346 (N_6346,N_5053,N_6089);
nand U6347 (N_6347,N_5679,N_5111);
xor U6348 (N_6348,N_5964,N_5972);
nor U6349 (N_6349,N_5270,N_5345);
and U6350 (N_6350,N_5820,N_5259);
and U6351 (N_6351,N_5773,N_5996);
or U6352 (N_6352,N_5960,N_5624);
and U6353 (N_6353,N_5335,N_6126);
or U6354 (N_6354,N_5305,N_5067);
nand U6355 (N_6355,N_6082,N_5894);
xor U6356 (N_6356,N_5385,N_5727);
nand U6357 (N_6357,N_5414,N_5552);
and U6358 (N_6358,N_5712,N_6032);
nor U6359 (N_6359,N_5068,N_5076);
and U6360 (N_6360,N_5953,N_5043);
nor U6361 (N_6361,N_5496,N_6084);
nand U6362 (N_6362,N_5539,N_5186);
nor U6363 (N_6363,N_5039,N_5183);
xor U6364 (N_6364,N_5466,N_6061);
nand U6365 (N_6365,N_5821,N_5913);
nand U6366 (N_6366,N_5220,N_5465);
and U6367 (N_6367,N_5946,N_5984);
nor U6368 (N_6368,N_5672,N_6222);
and U6369 (N_6369,N_5656,N_5588);
nor U6370 (N_6370,N_6058,N_5637);
nor U6371 (N_6371,N_6117,N_6196);
or U6372 (N_6372,N_5529,N_5781);
xor U6373 (N_6373,N_6217,N_5294);
xor U6374 (N_6374,N_6006,N_6001);
nand U6375 (N_6375,N_5364,N_5224);
nor U6376 (N_6376,N_5187,N_6004);
and U6377 (N_6377,N_5929,N_5413);
xnor U6378 (N_6378,N_5124,N_5571);
nor U6379 (N_6379,N_5533,N_5778);
and U6380 (N_6380,N_5267,N_5178);
nor U6381 (N_6381,N_5301,N_5733);
or U6382 (N_6382,N_6144,N_5154);
nand U6383 (N_6383,N_6241,N_5416);
or U6384 (N_6384,N_5304,N_5399);
or U6385 (N_6385,N_5968,N_5297);
nor U6386 (N_6386,N_5623,N_5292);
xor U6387 (N_6387,N_5419,N_5380);
and U6388 (N_6388,N_5198,N_5521);
and U6389 (N_6389,N_5942,N_5444);
nand U6390 (N_6390,N_5118,N_5311);
xor U6391 (N_6391,N_5943,N_5215);
xor U6392 (N_6392,N_5810,N_5987);
nand U6393 (N_6393,N_5797,N_5988);
nor U6394 (N_6394,N_5793,N_6164);
nor U6395 (N_6395,N_5572,N_5075);
or U6396 (N_6396,N_5668,N_6028);
nor U6397 (N_6397,N_5216,N_5403);
nand U6398 (N_6398,N_6024,N_5688);
nor U6399 (N_6399,N_6242,N_5205);
or U6400 (N_6400,N_6043,N_5877);
and U6401 (N_6401,N_5897,N_5844);
and U6402 (N_6402,N_5875,N_5083);
or U6403 (N_6403,N_5179,N_5966);
and U6404 (N_6404,N_5246,N_5510);
or U6405 (N_6405,N_5567,N_5936);
nor U6406 (N_6406,N_5130,N_5204);
and U6407 (N_6407,N_5888,N_5368);
nand U6408 (N_6408,N_5619,N_6240);
nand U6409 (N_6409,N_6176,N_6127);
and U6410 (N_6410,N_6160,N_5633);
nor U6411 (N_6411,N_5429,N_5298);
and U6412 (N_6412,N_5746,N_5989);
nor U6413 (N_6413,N_5247,N_6037);
xor U6414 (N_6414,N_5155,N_5642);
or U6415 (N_6415,N_5066,N_5890);
nor U6416 (N_6416,N_6054,N_5378);
xor U6417 (N_6417,N_5254,N_5440);
nor U6418 (N_6418,N_5165,N_5175);
or U6419 (N_6419,N_5861,N_6173);
xor U6420 (N_6420,N_5532,N_6197);
and U6421 (N_6421,N_5438,N_6181);
xnor U6422 (N_6422,N_5344,N_6039);
nand U6423 (N_6423,N_5979,N_5841);
xor U6424 (N_6424,N_5019,N_5383);
or U6425 (N_6425,N_5881,N_6180);
and U6426 (N_6426,N_5226,N_6035);
nand U6427 (N_6427,N_5857,N_5027);
nand U6428 (N_6428,N_5070,N_5730);
or U6429 (N_6429,N_5657,N_5077);
or U6430 (N_6430,N_6022,N_5769);
or U6431 (N_6431,N_5457,N_5361);
xnor U6432 (N_6432,N_5343,N_5762);
or U6433 (N_6433,N_5710,N_5949);
nor U6434 (N_6434,N_5119,N_5015);
xor U6435 (N_6435,N_5499,N_6062);
and U6436 (N_6436,N_5425,N_5095);
xor U6437 (N_6437,N_6235,N_5609);
or U6438 (N_6438,N_5397,N_6225);
nand U6439 (N_6439,N_6227,N_5823);
or U6440 (N_6440,N_5062,N_5522);
nor U6441 (N_6441,N_6165,N_6049);
or U6442 (N_6442,N_5826,N_5302);
and U6443 (N_6443,N_5051,N_5145);
or U6444 (N_6444,N_5775,N_6232);
and U6445 (N_6445,N_5631,N_5255);
nor U6446 (N_6446,N_5033,N_5629);
and U6447 (N_6447,N_5923,N_5227);
xnor U6448 (N_6448,N_5928,N_5136);
nor U6449 (N_6449,N_5675,N_5670);
nor U6450 (N_6450,N_5703,N_6234);
nand U6451 (N_6451,N_5046,N_5091);
xor U6452 (N_6452,N_6243,N_5235);
xor U6453 (N_6453,N_5954,N_5054);
or U6454 (N_6454,N_6184,N_5125);
xnor U6455 (N_6455,N_5269,N_5030);
nor U6456 (N_6456,N_5721,N_5803);
xor U6457 (N_6457,N_5517,N_6183);
nor U6458 (N_6458,N_6141,N_5667);
or U6459 (N_6459,N_5719,N_5277);
nor U6460 (N_6460,N_5505,N_5150);
nand U6461 (N_6461,N_5855,N_5909);
and U6462 (N_6462,N_5807,N_5738);
xnor U6463 (N_6463,N_6033,N_6093);
xnor U6464 (N_6464,N_5661,N_5384);
xor U6465 (N_6465,N_5501,N_6145);
nand U6466 (N_6466,N_6150,N_5472);
or U6467 (N_6467,N_5221,N_5718);
nor U6468 (N_6468,N_6067,N_5579);
or U6469 (N_6469,N_6186,N_5635);
and U6470 (N_6470,N_6245,N_6171);
nor U6471 (N_6471,N_5654,N_5180);
xor U6472 (N_6472,N_6203,N_5819);
and U6473 (N_6473,N_5439,N_5847);
and U6474 (N_6474,N_6090,N_6237);
nand U6475 (N_6475,N_5239,N_5182);
nor U6476 (N_6476,N_5174,N_5899);
nor U6477 (N_6477,N_5211,N_5809);
and U6478 (N_6478,N_5504,N_5799);
or U6479 (N_6479,N_5028,N_5478);
xor U6480 (N_6480,N_5214,N_5664);
xor U6481 (N_6481,N_5423,N_6132);
and U6482 (N_6482,N_5453,N_6130);
and U6483 (N_6483,N_5682,N_5045);
and U6484 (N_6484,N_5585,N_5766);
and U6485 (N_6485,N_5307,N_6110);
and U6486 (N_6486,N_5134,N_5569);
xor U6487 (N_6487,N_5584,N_6052);
xnor U6488 (N_6488,N_5490,N_5749);
nand U6489 (N_6489,N_5471,N_5206);
nand U6490 (N_6490,N_5346,N_5832);
nor U6491 (N_6491,N_6034,N_5272);
nor U6492 (N_6492,N_6157,N_5728);
and U6493 (N_6493,N_5997,N_5651);
nand U6494 (N_6494,N_5641,N_5374);
xor U6495 (N_6495,N_6073,N_5559);
xor U6496 (N_6496,N_5107,N_5926);
nor U6497 (N_6497,N_6168,N_5350);
nor U6498 (N_6498,N_6010,N_5649);
or U6499 (N_6499,N_5040,N_5197);
nand U6500 (N_6500,N_6185,N_5243);
or U6501 (N_6501,N_5595,N_5537);
or U6502 (N_6502,N_5223,N_5308);
nor U6503 (N_6503,N_6099,N_5244);
or U6504 (N_6504,N_5941,N_5322);
nand U6505 (N_6505,N_5907,N_5242);
and U6506 (N_6506,N_6195,N_5241);
nand U6507 (N_6507,N_5555,N_5003);
or U6508 (N_6508,N_5225,N_6097);
and U6509 (N_6509,N_5426,N_5591);
and U6510 (N_6510,N_5353,N_6041);
xnor U6511 (N_6511,N_5880,N_5340);
or U6512 (N_6512,N_5001,N_5562);
and U6513 (N_6513,N_5306,N_5032);
nand U6514 (N_6514,N_5073,N_5741);
or U6515 (N_6515,N_6088,N_5316);
nand U6516 (N_6516,N_5658,N_5952);
or U6517 (N_6517,N_5854,N_6106);
and U6518 (N_6518,N_6045,N_5879);
xnor U6519 (N_6519,N_6030,N_5678);
or U6520 (N_6520,N_5671,N_6163);
xnor U6521 (N_6521,N_5731,N_5436);
nor U6522 (N_6522,N_5299,N_5376);
nand U6523 (N_6523,N_5825,N_5959);
or U6524 (N_6524,N_5348,N_6153);
nand U6525 (N_6525,N_5093,N_6026);
nand U6526 (N_6526,N_5838,N_5549);
nor U6527 (N_6527,N_5222,N_5686);
nand U6528 (N_6528,N_5474,N_6162);
nand U6529 (N_6529,N_6040,N_5123);
or U6530 (N_6530,N_6075,N_5771);
and U6531 (N_6531,N_5594,N_5883);
xor U6532 (N_6532,N_6048,N_5314);
nor U6533 (N_6533,N_5696,N_5085);
nor U6534 (N_6534,N_5434,N_5231);
and U6535 (N_6535,N_6060,N_5164);
xor U6536 (N_6536,N_5437,N_5945);
nand U6537 (N_6537,N_6214,N_5655);
xor U6538 (N_6538,N_5084,N_5566);
and U6539 (N_6539,N_5617,N_5812);
and U6540 (N_6540,N_5424,N_5804);
or U6541 (N_6541,N_5233,N_5695);
xnor U6542 (N_6542,N_5596,N_5309);
nand U6543 (N_6543,N_5919,N_5753);
and U6544 (N_6544,N_5393,N_5994);
or U6545 (N_6545,N_5120,N_5709);
nor U6546 (N_6546,N_5169,N_5776);
and U6547 (N_6547,N_5331,N_5064);
nand U6548 (N_6548,N_5568,N_5940);
or U6549 (N_6549,N_5310,N_5652);
and U6550 (N_6550,N_5958,N_5515);
xor U6551 (N_6551,N_5431,N_5132);
or U6552 (N_6552,N_5139,N_5944);
and U6553 (N_6553,N_5342,N_5339);
xnor U6554 (N_6554,N_5274,N_5153);
nor U6555 (N_6555,N_6193,N_6123);
xnor U6556 (N_6556,N_6051,N_5498);
xnor U6557 (N_6557,N_5163,N_6115);
xnor U6558 (N_6558,N_5447,N_6015);
nand U6559 (N_6559,N_5927,N_5092);
and U6560 (N_6560,N_5105,N_5104);
or U6561 (N_6561,N_5885,N_5379);
nand U6562 (N_6562,N_5583,N_5514);
nor U6563 (N_6563,N_5554,N_5052);
nor U6564 (N_6564,N_5612,N_6125);
or U6565 (N_6565,N_5604,N_5813);
or U6566 (N_6566,N_5536,N_6154);
xor U6567 (N_6567,N_5842,N_5748);
nand U6568 (N_6568,N_5041,N_5112);
and U6569 (N_6569,N_5542,N_5422);
or U6570 (N_6570,N_6019,N_5874);
nor U6571 (N_6571,N_5570,N_5920);
nor U6572 (N_6572,N_6229,N_5010);
nand U6573 (N_6573,N_5530,N_5630);
or U6574 (N_6574,N_5253,N_5764);
nand U6575 (N_6575,N_5754,N_5939);
xnor U6576 (N_6576,N_5824,N_5442);
nor U6577 (N_6577,N_6057,N_5896);
or U6578 (N_6578,N_5690,N_5715);
xnor U6579 (N_6579,N_5428,N_5765);
and U6580 (N_6580,N_5538,N_5427);
nor U6581 (N_6581,N_5683,N_5577);
nand U6582 (N_6582,N_5281,N_5295);
or U6583 (N_6583,N_5788,N_5975);
or U6584 (N_6584,N_6220,N_6149);
xnor U6585 (N_6585,N_5341,N_5816);
nand U6586 (N_6586,N_6129,N_6158);
or U6587 (N_6587,N_5918,N_6247);
nor U6588 (N_6588,N_5362,N_5315);
nand U6589 (N_6589,N_5669,N_5689);
and U6590 (N_6590,N_5049,N_5021);
or U6591 (N_6591,N_5937,N_6142);
or U6592 (N_6592,N_5140,N_5934);
and U6593 (N_6593,N_5389,N_5014);
or U6594 (N_6594,N_5144,N_5462);
nand U6595 (N_6595,N_5476,N_5209);
xnor U6596 (N_6596,N_5412,N_5848);
xor U6597 (N_6597,N_5777,N_5701);
and U6598 (N_6598,N_5464,N_5865);
or U6599 (N_6599,N_5258,N_6053);
xnor U6600 (N_6600,N_5170,N_5707);
or U6601 (N_6601,N_5691,N_5454);
or U6602 (N_6602,N_5017,N_6233);
xnor U6603 (N_6603,N_6155,N_6042);
or U6604 (N_6604,N_5148,N_5513);
or U6605 (N_6605,N_5394,N_5047);
nand U6606 (N_6606,N_5747,N_5547);
nand U6607 (N_6607,N_5279,N_6206);
nand U6608 (N_6608,N_5659,N_5240);
or U6609 (N_6609,N_5976,N_6025);
or U6610 (N_6610,N_5026,N_6170);
nand U6611 (N_6611,N_6103,N_5483);
and U6612 (N_6612,N_5999,N_5893);
or U6613 (N_6613,N_5373,N_5589);
xnor U6614 (N_6614,N_5330,N_5025);
and U6615 (N_6615,N_5296,N_5648);
and U6616 (N_6616,N_5106,N_5978);
nand U6617 (N_6617,N_5729,N_5058);
and U6618 (N_6618,N_5795,N_5917);
xnor U6619 (N_6619,N_6177,N_6178);
xor U6620 (N_6620,N_5991,N_5685);
nand U6621 (N_6621,N_5705,N_5548);
and U6622 (N_6622,N_5189,N_5980);
xor U6623 (N_6623,N_5236,N_6207);
nand U6624 (N_6624,N_5234,N_5856);
or U6625 (N_6625,N_5317,N_5614);
nand U6626 (N_6626,N_6079,N_5891);
xor U6627 (N_6627,N_6036,N_5288);
nor U6628 (N_6628,N_5723,N_6136);
nor U6629 (N_6629,N_5525,N_5050);
xor U6630 (N_6630,N_5732,N_6116);
and U6631 (N_6631,N_5059,N_5491);
or U6632 (N_6632,N_5535,N_5805);
nand U6633 (N_6633,N_6134,N_5925);
and U6634 (N_6634,N_5843,N_5963);
or U6635 (N_6635,N_5470,N_5808);
nand U6636 (N_6636,N_5610,N_6101);
xnor U6637 (N_6637,N_6108,N_5556);
nor U6638 (N_6638,N_5458,N_5887);
xor U6639 (N_6639,N_5202,N_5763);
and U6640 (N_6640,N_5131,N_5420);
xor U6641 (N_6641,N_5698,N_6248);
xor U6642 (N_6642,N_6018,N_6017);
nand U6643 (N_6643,N_5261,N_6107);
and U6644 (N_6644,N_5372,N_5787);
nor U6645 (N_6645,N_5702,N_6211);
or U6646 (N_6646,N_5607,N_5643);
xor U6647 (N_6647,N_5512,N_5173);
and U6648 (N_6648,N_5250,N_5600);
or U6649 (N_6649,N_5575,N_5485);
nor U6650 (N_6650,N_5831,N_6198);
and U6651 (N_6651,N_5351,N_6013);
nor U6652 (N_6652,N_5484,N_6147);
nand U6653 (N_6653,N_6113,N_5932);
nand U6654 (N_6654,N_5325,N_6050);
and U6655 (N_6655,N_5320,N_6064);
or U6656 (N_6656,N_5200,N_5060);
or U6657 (N_6657,N_5009,N_5995);
nand U6658 (N_6658,N_5487,N_5029);
nor U6659 (N_6659,N_5275,N_5725);
nand U6660 (N_6660,N_5410,N_5480);
xor U6661 (N_6661,N_6124,N_5392);
nand U6662 (N_6662,N_5739,N_5540);
or U6663 (N_6663,N_5072,N_5677);
nand U6664 (N_6664,N_5981,N_5801);
xnor U6665 (N_6665,N_5830,N_5862);
or U6666 (N_6666,N_5871,N_5573);
nand U6667 (N_6667,N_5044,N_5520);
xor U6668 (N_6668,N_5868,N_5811);
or U6669 (N_6669,N_5620,N_5264);
nand U6670 (N_6670,N_6215,N_5212);
xor U6671 (N_6671,N_6140,N_5606);
nand U6672 (N_6672,N_5473,N_5516);
nor U6673 (N_6673,N_5935,N_5869);
and U6674 (N_6674,N_5502,N_5097);
xor U6675 (N_6675,N_5743,N_6109);
or U6676 (N_6676,N_5597,N_5931);
nor U6677 (N_6677,N_5098,N_6077);
nand U6678 (N_6678,N_6005,N_6135);
nand U6679 (N_6679,N_6078,N_5370);
or U6680 (N_6680,N_5185,N_5156);
nand U6681 (N_6681,N_5493,N_5143);
xor U6682 (N_6682,N_5817,N_5355);
or U6683 (N_6683,N_5219,N_5835);
and U6684 (N_6684,N_5790,N_6096);
nor U6685 (N_6685,N_5767,N_5815);
nand U6686 (N_6686,N_5333,N_5110);
or U6687 (N_6687,N_5278,N_5004);
nor U6688 (N_6688,N_5866,N_5357);
nand U6689 (N_6689,N_6209,N_5950);
xor U6690 (N_6690,N_5158,N_5405);
nand U6691 (N_6691,N_5759,N_6230);
and U6692 (N_6692,N_6066,N_5524);
xnor U6693 (N_6693,N_5347,N_5086);
or U6694 (N_6694,N_6228,N_5632);
nand U6695 (N_6695,N_5181,N_6083);
nand U6696 (N_6696,N_5265,N_5252);
nand U6697 (N_6697,N_5318,N_5128);
and U6698 (N_6698,N_5133,N_5388);
nand U6699 (N_6699,N_5889,N_5531);
nand U6700 (N_6700,N_5587,N_5726);
xnor U6701 (N_6701,N_5663,N_5676);
xnor U6702 (N_6702,N_5323,N_5916);
nand U6703 (N_6703,N_6238,N_5443);
nor U6704 (N_6704,N_5366,N_5400);
and U6705 (N_6705,N_5199,N_5495);
or U6706 (N_6706,N_5249,N_5121);
xnor U6707 (N_6707,N_5463,N_5303);
xor U6708 (N_6708,N_5257,N_5802);
and U6709 (N_6709,N_5716,N_5626);
and U6710 (N_6710,N_6086,N_6095);
and U6711 (N_6711,N_5845,N_5500);
nand U6712 (N_6712,N_5638,N_5750);
and U6713 (N_6713,N_6148,N_5055);
nor U6714 (N_6714,N_5432,N_6065);
xnor U6715 (N_6715,N_5446,N_5232);
nor U6716 (N_6716,N_5489,N_5011);
xnor U6717 (N_6717,N_5951,N_5081);
xor U6718 (N_6718,N_5161,N_6249);
xnor U6719 (N_6719,N_6182,N_5780);
nor U6720 (N_6720,N_5650,N_5708);
or U6721 (N_6721,N_6187,N_5647);
nor U6722 (N_6722,N_5002,N_5518);
and U6723 (N_6723,N_5210,N_5985);
or U6724 (N_6724,N_5938,N_5398);
nor U6725 (N_6725,N_5031,N_6199);
nand U6726 (N_6726,N_5565,N_5114);
nor U6727 (N_6727,N_5982,N_6189);
nand U6728 (N_6728,N_5171,N_5450);
xor U6729 (N_6729,N_5895,N_5365);
and U6730 (N_6730,N_5137,N_5618);
nor U6731 (N_6731,N_5904,N_6098);
or U6732 (N_6732,N_6085,N_5740);
or U6733 (N_6733,N_5544,N_5094);
xor U6734 (N_6734,N_5395,N_5622);
and U6735 (N_6735,N_5967,N_5840);
nand U6736 (N_6736,N_5147,N_5177);
nand U6737 (N_6737,N_5460,N_5564);
and U6738 (N_6738,N_5751,N_5321);
nor U6739 (N_6739,N_6205,N_6208);
and U6740 (N_6740,N_5349,N_5018);
nor U6741 (N_6741,N_5601,N_5007);
or U6742 (N_6742,N_5921,N_5149);
nor U6743 (N_6743,N_6239,N_5005);
and U6744 (N_6744,N_5706,N_5992);
and U6745 (N_6745,N_6172,N_6221);
xor U6746 (N_6746,N_5901,N_5401);
and U6747 (N_6747,N_5506,N_5534);
or U6748 (N_6748,N_5191,N_5300);
and U6749 (N_6749,N_5386,N_5245);
xnor U6750 (N_6750,N_5238,N_5494);
and U6751 (N_6751,N_6003,N_5013);
xor U6752 (N_6752,N_5160,N_5692);
xor U6753 (N_6753,N_6071,N_6216);
or U6754 (N_6754,N_5608,N_6074);
or U6755 (N_6755,N_6105,N_5375);
or U6756 (N_6756,N_5508,N_5285);
nor U6757 (N_6757,N_5406,N_5276);
or U6758 (N_6758,N_5448,N_5468);
or U6759 (N_6759,N_5755,N_5217);
nor U6760 (N_6760,N_5644,N_5910);
nor U6761 (N_6761,N_6070,N_5151);
or U6762 (N_6762,N_6021,N_6016);
nor U6763 (N_6763,N_5674,N_5860);
and U6764 (N_6764,N_5846,N_5441);
and U6765 (N_6765,N_5312,N_5882);
xor U6766 (N_6766,N_5758,N_5605);
or U6767 (N_6767,N_5248,N_6023);
or U6768 (N_6768,N_5157,N_5511);
nor U6769 (N_6769,N_5541,N_6204);
xnor U6770 (N_6770,N_5543,N_5756);
and U6771 (N_6771,N_5794,N_5970);
and U6772 (N_6772,N_5022,N_5332);
nand U6773 (N_6773,N_5911,N_5260);
xor U6774 (N_6774,N_5834,N_5459);
and U6775 (N_6775,N_5218,N_5354);
nand U6776 (N_6776,N_5036,N_5908);
and U6777 (N_6777,N_5176,N_5687);
or U6778 (N_6778,N_5188,N_5415);
nor U6779 (N_6779,N_5971,N_5625);
or U6780 (N_6780,N_5486,N_6166);
nor U6781 (N_6781,N_6031,N_5955);
nand U6782 (N_6782,N_5836,N_5814);
or U6783 (N_6783,N_5266,N_5822);
nor U6784 (N_6784,N_6156,N_5806);
or U6785 (N_6785,N_5876,N_5760);
or U6786 (N_6786,N_5742,N_6219);
or U6787 (N_6787,N_5873,N_5467);
and U6788 (N_6788,N_5071,N_5791);
and U6789 (N_6789,N_5962,N_6047);
or U6790 (N_6790,N_5338,N_5680);
nor U6791 (N_6791,N_6008,N_5195);
and U6792 (N_6792,N_5558,N_5407);
nor U6793 (N_6793,N_5451,N_5560);
and U6794 (N_6794,N_5329,N_6011);
nor U6795 (N_6795,N_5152,N_5864);
nand U6796 (N_6796,N_6114,N_5851);
nor U6797 (N_6797,N_5977,N_6069);
nor U6798 (N_6798,N_5168,N_5100);
nor U6799 (N_6799,N_5482,N_5898);
or U6800 (N_6800,N_5142,N_6014);
xor U6801 (N_6801,N_5023,N_5892);
nand U6802 (N_6802,N_6002,N_6192);
nand U6803 (N_6803,N_6218,N_5528);
and U6804 (N_6804,N_5922,N_5359);
or U6805 (N_6805,N_5020,N_5461);
nand U6806 (N_6806,N_5553,N_5800);
nand U6807 (N_6807,N_6246,N_5117);
and U6808 (N_6808,N_5251,N_5593);
xnor U6809 (N_6809,N_5000,N_5697);
nor U6810 (N_6810,N_5914,N_6044);
and U6811 (N_6811,N_6038,N_5237);
or U6812 (N_6812,N_5069,N_5203);
xor U6813 (N_6813,N_5639,N_5858);
or U6814 (N_6814,N_5477,N_5037);
and U6815 (N_6815,N_5196,N_5789);
or U6816 (N_6816,N_5402,N_5745);
nor U6817 (N_6817,N_5783,N_5034);
or U6818 (N_6818,N_6224,N_5256);
nor U6819 (N_6819,N_5391,N_5109);
and U6820 (N_6820,N_5291,N_5634);
and U6821 (N_6821,N_6159,N_5159);
or U6822 (N_6822,N_5456,N_5561);
nand U6823 (N_6823,N_5870,N_5768);
nand U6824 (N_6824,N_5411,N_5616);
and U6825 (N_6825,N_6143,N_5681);
nor U6826 (N_6826,N_5475,N_5930);
or U6827 (N_6827,N_5509,N_5492);
nand U6828 (N_6828,N_6231,N_6111);
nor U6829 (N_6829,N_5396,N_5784);
nand U6830 (N_6830,N_6133,N_5102);
nor U6831 (N_6831,N_6179,N_5551);
and U6832 (N_6832,N_5903,N_5192);
nand U6833 (N_6833,N_5479,N_5065);
or U6834 (N_6834,N_5666,N_5135);
or U6835 (N_6835,N_5283,N_5900);
nor U6836 (N_6836,N_5711,N_5074);
or U6837 (N_6837,N_5722,N_6202);
and U6838 (N_6838,N_5969,N_5061);
and U6839 (N_6839,N_6094,N_6152);
and U6840 (N_6840,N_5122,N_6081);
nand U6841 (N_6841,N_5166,N_6174);
xnor U6842 (N_6842,N_6056,N_5853);
and U6843 (N_6843,N_5481,N_5126);
nand U6844 (N_6844,N_5863,N_5096);
or U6845 (N_6845,N_6223,N_5293);
xnor U6846 (N_6846,N_6190,N_5326);
nand U6847 (N_6847,N_5080,N_6012);
nor U6848 (N_6848,N_5785,N_5417);
and U6849 (N_6849,N_5886,N_6087);
nand U6850 (N_6850,N_6138,N_5358);
or U6851 (N_6851,N_5990,N_5563);
nand U6852 (N_6852,N_5381,N_5387);
nand U6853 (N_6853,N_5208,N_5328);
nor U6854 (N_6854,N_5048,N_6009);
and U6855 (N_6855,N_6007,N_5833);
and U6856 (N_6856,N_5273,N_6020);
or U6857 (N_6857,N_5915,N_5146);
nand U6858 (N_6858,N_6201,N_5684);
nand U6859 (N_6859,N_5115,N_5550);
nand U6860 (N_6860,N_5336,N_5829);
and U6861 (N_6861,N_5884,N_5360);
or U6862 (N_6862,N_5207,N_5576);
and U6863 (N_6863,N_5752,N_5792);
nor U6864 (N_6864,N_5613,N_5735);
xor U6865 (N_6865,N_5263,N_5008);
or U6866 (N_6866,N_5839,N_5079);
or U6867 (N_6867,N_5640,N_6146);
nor U6868 (N_6868,N_5947,N_5006);
and U6869 (N_6869,N_6100,N_6091);
xnor U6870 (N_6870,N_5430,N_5334);
xor U6871 (N_6871,N_6161,N_5229);
or U6872 (N_6872,N_5859,N_5167);
nor U6873 (N_6873,N_5714,N_6137);
and U6874 (N_6874,N_5082,N_5090);
nand U6875 (N_6875,N_5154,N_5902);
and U6876 (N_6876,N_6209,N_5972);
or U6877 (N_6877,N_5914,N_5418);
or U6878 (N_6878,N_5817,N_6241);
nand U6879 (N_6879,N_5164,N_6079);
nand U6880 (N_6880,N_5643,N_5383);
or U6881 (N_6881,N_5871,N_5768);
xor U6882 (N_6882,N_5470,N_5142);
and U6883 (N_6883,N_5723,N_5429);
and U6884 (N_6884,N_5149,N_5308);
and U6885 (N_6885,N_6109,N_5489);
xnor U6886 (N_6886,N_6157,N_5493);
or U6887 (N_6887,N_6178,N_6012);
xor U6888 (N_6888,N_5247,N_6043);
or U6889 (N_6889,N_6160,N_5868);
xnor U6890 (N_6890,N_5228,N_6226);
xor U6891 (N_6891,N_5459,N_5448);
nor U6892 (N_6892,N_6102,N_5629);
xor U6893 (N_6893,N_5315,N_5807);
or U6894 (N_6894,N_5877,N_5345);
and U6895 (N_6895,N_5295,N_5859);
and U6896 (N_6896,N_6191,N_5545);
nand U6897 (N_6897,N_5361,N_5881);
xor U6898 (N_6898,N_5834,N_5677);
or U6899 (N_6899,N_5076,N_5446);
and U6900 (N_6900,N_5771,N_5992);
xor U6901 (N_6901,N_5967,N_5718);
xor U6902 (N_6902,N_5652,N_5435);
nor U6903 (N_6903,N_5111,N_5840);
xor U6904 (N_6904,N_5301,N_5514);
or U6905 (N_6905,N_5933,N_5558);
nor U6906 (N_6906,N_5661,N_5458);
nand U6907 (N_6907,N_5562,N_6061);
or U6908 (N_6908,N_5997,N_5220);
xnor U6909 (N_6909,N_5120,N_5653);
and U6910 (N_6910,N_5993,N_5310);
and U6911 (N_6911,N_5773,N_5701);
and U6912 (N_6912,N_5722,N_5785);
xor U6913 (N_6913,N_5949,N_5057);
or U6914 (N_6914,N_5177,N_5144);
or U6915 (N_6915,N_5887,N_5929);
nand U6916 (N_6916,N_5667,N_5727);
or U6917 (N_6917,N_6023,N_5333);
xor U6918 (N_6918,N_5391,N_6164);
nor U6919 (N_6919,N_5851,N_6207);
or U6920 (N_6920,N_5923,N_5041);
nor U6921 (N_6921,N_5629,N_6177);
xnor U6922 (N_6922,N_6097,N_5837);
xor U6923 (N_6923,N_5165,N_5709);
nand U6924 (N_6924,N_5843,N_5933);
xor U6925 (N_6925,N_6054,N_5525);
or U6926 (N_6926,N_5983,N_5320);
and U6927 (N_6927,N_6200,N_6204);
xor U6928 (N_6928,N_5026,N_5762);
and U6929 (N_6929,N_6128,N_5589);
or U6930 (N_6930,N_6191,N_6156);
and U6931 (N_6931,N_6034,N_5605);
nor U6932 (N_6932,N_5683,N_5446);
and U6933 (N_6933,N_5978,N_5604);
xor U6934 (N_6934,N_5961,N_5081);
nor U6935 (N_6935,N_5027,N_5635);
or U6936 (N_6936,N_5526,N_5371);
xor U6937 (N_6937,N_5883,N_5038);
and U6938 (N_6938,N_5490,N_5282);
or U6939 (N_6939,N_5918,N_5153);
nor U6940 (N_6940,N_5606,N_5156);
xor U6941 (N_6941,N_5096,N_5117);
or U6942 (N_6942,N_5471,N_6226);
nand U6943 (N_6943,N_6007,N_5205);
or U6944 (N_6944,N_5389,N_5471);
nand U6945 (N_6945,N_6187,N_5811);
nand U6946 (N_6946,N_6134,N_5793);
nand U6947 (N_6947,N_5559,N_5963);
or U6948 (N_6948,N_6043,N_6246);
xnor U6949 (N_6949,N_5443,N_5995);
or U6950 (N_6950,N_5567,N_5519);
nor U6951 (N_6951,N_5662,N_5267);
nor U6952 (N_6952,N_5265,N_5804);
nor U6953 (N_6953,N_5292,N_5754);
and U6954 (N_6954,N_5566,N_5246);
and U6955 (N_6955,N_5374,N_5548);
and U6956 (N_6956,N_5135,N_6124);
nand U6957 (N_6957,N_5204,N_5060);
or U6958 (N_6958,N_5346,N_6027);
nor U6959 (N_6959,N_5868,N_5553);
and U6960 (N_6960,N_5286,N_5850);
and U6961 (N_6961,N_5247,N_5433);
and U6962 (N_6962,N_6172,N_5604);
nand U6963 (N_6963,N_5092,N_5634);
nand U6964 (N_6964,N_5690,N_5148);
or U6965 (N_6965,N_5645,N_6021);
nor U6966 (N_6966,N_5752,N_5901);
nor U6967 (N_6967,N_5540,N_5996);
nor U6968 (N_6968,N_5504,N_6094);
nand U6969 (N_6969,N_5545,N_5308);
xnor U6970 (N_6970,N_6112,N_5132);
xnor U6971 (N_6971,N_5725,N_5583);
xnor U6972 (N_6972,N_5594,N_6102);
nand U6973 (N_6973,N_6076,N_5830);
xor U6974 (N_6974,N_5790,N_5350);
or U6975 (N_6975,N_5066,N_5753);
nand U6976 (N_6976,N_5329,N_5104);
and U6977 (N_6977,N_6160,N_5836);
nor U6978 (N_6978,N_5128,N_5518);
and U6979 (N_6979,N_5034,N_5749);
or U6980 (N_6980,N_5299,N_5310);
xor U6981 (N_6981,N_6113,N_5508);
xnor U6982 (N_6982,N_5744,N_6247);
or U6983 (N_6983,N_5850,N_5604);
xor U6984 (N_6984,N_5907,N_5663);
and U6985 (N_6985,N_5474,N_5558);
nor U6986 (N_6986,N_5125,N_5777);
nand U6987 (N_6987,N_5879,N_5312);
or U6988 (N_6988,N_5997,N_6239);
and U6989 (N_6989,N_5613,N_5185);
and U6990 (N_6990,N_5818,N_5891);
or U6991 (N_6991,N_6142,N_6122);
xor U6992 (N_6992,N_5436,N_5258);
nor U6993 (N_6993,N_5989,N_5829);
nand U6994 (N_6994,N_5725,N_5141);
nor U6995 (N_6995,N_6180,N_5578);
nand U6996 (N_6996,N_5117,N_6225);
nor U6997 (N_6997,N_5801,N_5540);
xnor U6998 (N_6998,N_5443,N_5125);
nor U6999 (N_6999,N_5801,N_5013);
or U7000 (N_7000,N_5164,N_5257);
nand U7001 (N_7001,N_5618,N_5492);
nand U7002 (N_7002,N_5698,N_5082);
nor U7003 (N_7003,N_5808,N_5028);
or U7004 (N_7004,N_5120,N_5402);
nor U7005 (N_7005,N_5215,N_5470);
or U7006 (N_7006,N_5669,N_5953);
xnor U7007 (N_7007,N_5443,N_5144);
and U7008 (N_7008,N_5368,N_5613);
xnor U7009 (N_7009,N_5898,N_5197);
xor U7010 (N_7010,N_5777,N_5902);
or U7011 (N_7011,N_5916,N_5591);
xnor U7012 (N_7012,N_6192,N_6092);
nand U7013 (N_7013,N_5339,N_5967);
or U7014 (N_7014,N_5201,N_5412);
or U7015 (N_7015,N_5184,N_5481);
and U7016 (N_7016,N_5647,N_5998);
or U7017 (N_7017,N_5425,N_5188);
and U7018 (N_7018,N_5971,N_5849);
xor U7019 (N_7019,N_5704,N_6003);
nand U7020 (N_7020,N_5546,N_5795);
nand U7021 (N_7021,N_5633,N_5504);
or U7022 (N_7022,N_5328,N_6107);
nand U7023 (N_7023,N_5373,N_5842);
and U7024 (N_7024,N_5997,N_5394);
xor U7025 (N_7025,N_5941,N_6173);
nand U7026 (N_7026,N_5644,N_6222);
nand U7027 (N_7027,N_6136,N_5275);
xor U7028 (N_7028,N_6009,N_5065);
nand U7029 (N_7029,N_6017,N_6080);
nand U7030 (N_7030,N_5017,N_5805);
or U7031 (N_7031,N_5371,N_5129);
nor U7032 (N_7032,N_5130,N_5659);
nand U7033 (N_7033,N_5520,N_5807);
nand U7034 (N_7034,N_5539,N_5579);
nand U7035 (N_7035,N_5290,N_5472);
nand U7036 (N_7036,N_6096,N_6084);
xor U7037 (N_7037,N_5059,N_5940);
or U7038 (N_7038,N_5049,N_5415);
and U7039 (N_7039,N_5129,N_5876);
or U7040 (N_7040,N_5615,N_5045);
nor U7041 (N_7041,N_5529,N_5278);
nand U7042 (N_7042,N_6111,N_5042);
nor U7043 (N_7043,N_5018,N_5973);
and U7044 (N_7044,N_5365,N_5724);
nor U7045 (N_7045,N_5605,N_5301);
nor U7046 (N_7046,N_5303,N_6093);
and U7047 (N_7047,N_5031,N_6010);
nand U7048 (N_7048,N_5120,N_6136);
xor U7049 (N_7049,N_5160,N_5780);
nor U7050 (N_7050,N_5119,N_5056);
and U7051 (N_7051,N_5795,N_5632);
nand U7052 (N_7052,N_5669,N_5794);
nand U7053 (N_7053,N_5848,N_5240);
xor U7054 (N_7054,N_5877,N_5124);
and U7055 (N_7055,N_5372,N_5547);
and U7056 (N_7056,N_6012,N_6014);
xnor U7057 (N_7057,N_5578,N_5833);
and U7058 (N_7058,N_6219,N_5224);
xnor U7059 (N_7059,N_5144,N_5678);
or U7060 (N_7060,N_5623,N_6048);
xnor U7061 (N_7061,N_5605,N_6068);
and U7062 (N_7062,N_5502,N_5468);
nor U7063 (N_7063,N_5807,N_5627);
or U7064 (N_7064,N_5078,N_5871);
or U7065 (N_7065,N_5193,N_5229);
or U7066 (N_7066,N_5729,N_5022);
nor U7067 (N_7067,N_6122,N_5354);
and U7068 (N_7068,N_5291,N_6029);
nand U7069 (N_7069,N_5129,N_5823);
nor U7070 (N_7070,N_5964,N_5119);
or U7071 (N_7071,N_5012,N_5329);
nor U7072 (N_7072,N_5582,N_5386);
xnor U7073 (N_7073,N_5291,N_5384);
nor U7074 (N_7074,N_5382,N_5365);
nor U7075 (N_7075,N_5463,N_5721);
or U7076 (N_7076,N_5834,N_6155);
xor U7077 (N_7077,N_6074,N_5574);
nand U7078 (N_7078,N_5445,N_5081);
nor U7079 (N_7079,N_6238,N_5140);
xor U7080 (N_7080,N_5288,N_5318);
nand U7081 (N_7081,N_6159,N_5099);
nor U7082 (N_7082,N_5169,N_6035);
xnor U7083 (N_7083,N_5144,N_6059);
nor U7084 (N_7084,N_6169,N_5692);
and U7085 (N_7085,N_5107,N_5719);
or U7086 (N_7086,N_5446,N_5823);
and U7087 (N_7087,N_5250,N_5258);
xor U7088 (N_7088,N_5439,N_5058);
and U7089 (N_7089,N_5172,N_5485);
or U7090 (N_7090,N_5591,N_5606);
nor U7091 (N_7091,N_6029,N_5251);
or U7092 (N_7092,N_5179,N_5948);
nor U7093 (N_7093,N_6198,N_6090);
and U7094 (N_7094,N_5571,N_5760);
nand U7095 (N_7095,N_5951,N_5921);
nor U7096 (N_7096,N_5315,N_5518);
or U7097 (N_7097,N_5359,N_5684);
or U7098 (N_7098,N_5331,N_5722);
or U7099 (N_7099,N_5367,N_6203);
nor U7100 (N_7100,N_5992,N_5664);
and U7101 (N_7101,N_6115,N_5699);
xor U7102 (N_7102,N_5966,N_6030);
or U7103 (N_7103,N_5664,N_5814);
nand U7104 (N_7104,N_6149,N_5310);
or U7105 (N_7105,N_6193,N_5204);
nand U7106 (N_7106,N_6186,N_5560);
xor U7107 (N_7107,N_6248,N_5380);
nor U7108 (N_7108,N_5192,N_5164);
xnor U7109 (N_7109,N_5178,N_6090);
xnor U7110 (N_7110,N_6205,N_5482);
or U7111 (N_7111,N_5822,N_5727);
nand U7112 (N_7112,N_6102,N_6157);
nor U7113 (N_7113,N_5899,N_5040);
xor U7114 (N_7114,N_6160,N_5983);
nand U7115 (N_7115,N_5902,N_5756);
xnor U7116 (N_7116,N_5603,N_5958);
and U7117 (N_7117,N_5480,N_6146);
xnor U7118 (N_7118,N_5703,N_6126);
and U7119 (N_7119,N_5737,N_6000);
nand U7120 (N_7120,N_5205,N_5010);
or U7121 (N_7121,N_5468,N_5832);
or U7122 (N_7122,N_5975,N_5974);
and U7123 (N_7123,N_5082,N_5256);
nand U7124 (N_7124,N_5666,N_5347);
nand U7125 (N_7125,N_6147,N_5021);
nand U7126 (N_7126,N_5569,N_5519);
nand U7127 (N_7127,N_5545,N_5788);
nand U7128 (N_7128,N_6040,N_5043);
or U7129 (N_7129,N_5181,N_5699);
and U7130 (N_7130,N_5342,N_6109);
nor U7131 (N_7131,N_5762,N_5294);
nor U7132 (N_7132,N_5626,N_5526);
xor U7133 (N_7133,N_6091,N_5557);
nor U7134 (N_7134,N_5834,N_5047);
nand U7135 (N_7135,N_5984,N_5101);
and U7136 (N_7136,N_5077,N_5904);
nand U7137 (N_7137,N_5589,N_5689);
or U7138 (N_7138,N_5739,N_5285);
or U7139 (N_7139,N_5461,N_5679);
nor U7140 (N_7140,N_5640,N_5540);
or U7141 (N_7141,N_5066,N_5341);
and U7142 (N_7142,N_5248,N_5420);
and U7143 (N_7143,N_5326,N_5293);
and U7144 (N_7144,N_5559,N_6185);
and U7145 (N_7145,N_5386,N_5905);
or U7146 (N_7146,N_5532,N_5505);
or U7147 (N_7147,N_5641,N_6010);
or U7148 (N_7148,N_6201,N_5626);
nor U7149 (N_7149,N_5475,N_6018);
nor U7150 (N_7150,N_5103,N_5659);
nor U7151 (N_7151,N_5019,N_6041);
or U7152 (N_7152,N_6031,N_5720);
nor U7153 (N_7153,N_6022,N_5304);
nand U7154 (N_7154,N_5592,N_5068);
nor U7155 (N_7155,N_6188,N_6107);
nor U7156 (N_7156,N_5169,N_5058);
xor U7157 (N_7157,N_6103,N_5655);
and U7158 (N_7158,N_6086,N_5405);
and U7159 (N_7159,N_5614,N_5380);
and U7160 (N_7160,N_6039,N_5198);
nand U7161 (N_7161,N_5829,N_5091);
and U7162 (N_7162,N_5464,N_5830);
nor U7163 (N_7163,N_5858,N_6225);
xor U7164 (N_7164,N_5186,N_5056);
xnor U7165 (N_7165,N_5659,N_5928);
or U7166 (N_7166,N_5467,N_5855);
xnor U7167 (N_7167,N_5036,N_6104);
nor U7168 (N_7168,N_6057,N_6003);
and U7169 (N_7169,N_5654,N_5016);
xor U7170 (N_7170,N_6178,N_5918);
nand U7171 (N_7171,N_5371,N_5553);
and U7172 (N_7172,N_6081,N_6109);
or U7173 (N_7173,N_6133,N_5833);
nand U7174 (N_7174,N_6019,N_6225);
nand U7175 (N_7175,N_5155,N_5105);
and U7176 (N_7176,N_5821,N_5572);
nand U7177 (N_7177,N_5130,N_6200);
or U7178 (N_7178,N_5916,N_5001);
nor U7179 (N_7179,N_6106,N_5076);
nor U7180 (N_7180,N_5730,N_5074);
nand U7181 (N_7181,N_5424,N_5218);
xor U7182 (N_7182,N_5644,N_5006);
or U7183 (N_7183,N_5946,N_5504);
nor U7184 (N_7184,N_5392,N_5900);
nand U7185 (N_7185,N_6051,N_5396);
or U7186 (N_7186,N_5495,N_5452);
xor U7187 (N_7187,N_5053,N_5949);
or U7188 (N_7188,N_6216,N_6195);
xor U7189 (N_7189,N_5300,N_5380);
nor U7190 (N_7190,N_6049,N_5880);
nand U7191 (N_7191,N_5059,N_5052);
nand U7192 (N_7192,N_5945,N_5612);
nor U7193 (N_7193,N_5928,N_5082);
nor U7194 (N_7194,N_5400,N_5717);
xnor U7195 (N_7195,N_5236,N_5395);
xnor U7196 (N_7196,N_5207,N_5473);
and U7197 (N_7197,N_5638,N_6018);
and U7198 (N_7198,N_5169,N_6128);
or U7199 (N_7199,N_6120,N_6186);
xor U7200 (N_7200,N_6104,N_6042);
nand U7201 (N_7201,N_6193,N_5325);
xor U7202 (N_7202,N_5269,N_5093);
and U7203 (N_7203,N_5715,N_6043);
nand U7204 (N_7204,N_5422,N_5515);
and U7205 (N_7205,N_5906,N_5347);
and U7206 (N_7206,N_5698,N_6034);
xnor U7207 (N_7207,N_5714,N_5330);
or U7208 (N_7208,N_5914,N_5171);
xnor U7209 (N_7209,N_5760,N_5706);
xnor U7210 (N_7210,N_5643,N_5355);
or U7211 (N_7211,N_5227,N_5342);
nand U7212 (N_7212,N_5646,N_5899);
nor U7213 (N_7213,N_5452,N_5150);
or U7214 (N_7214,N_5194,N_5004);
or U7215 (N_7215,N_5485,N_5605);
and U7216 (N_7216,N_5493,N_5395);
and U7217 (N_7217,N_6003,N_5403);
or U7218 (N_7218,N_5830,N_6058);
nand U7219 (N_7219,N_5983,N_6129);
nand U7220 (N_7220,N_5517,N_5352);
nand U7221 (N_7221,N_6057,N_6137);
xnor U7222 (N_7222,N_5304,N_6096);
nor U7223 (N_7223,N_5603,N_5345);
nand U7224 (N_7224,N_5335,N_6122);
nand U7225 (N_7225,N_5823,N_5944);
nand U7226 (N_7226,N_6208,N_5169);
nor U7227 (N_7227,N_5476,N_5105);
or U7228 (N_7228,N_5182,N_5306);
xor U7229 (N_7229,N_5505,N_6217);
or U7230 (N_7230,N_6216,N_6093);
nand U7231 (N_7231,N_5253,N_5785);
and U7232 (N_7232,N_5078,N_5599);
nor U7233 (N_7233,N_5789,N_5744);
nor U7234 (N_7234,N_6229,N_5533);
nand U7235 (N_7235,N_5075,N_5843);
and U7236 (N_7236,N_5869,N_5568);
and U7237 (N_7237,N_5112,N_5315);
xnor U7238 (N_7238,N_5477,N_5549);
nand U7239 (N_7239,N_5932,N_5376);
xor U7240 (N_7240,N_6192,N_5881);
and U7241 (N_7241,N_6172,N_5447);
xor U7242 (N_7242,N_5644,N_5081);
nand U7243 (N_7243,N_5752,N_6163);
and U7244 (N_7244,N_5403,N_6108);
or U7245 (N_7245,N_5026,N_5232);
and U7246 (N_7246,N_5862,N_5383);
nand U7247 (N_7247,N_5540,N_5707);
nand U7248 (N_7248,N_5994,N_5316);
and U7249 (N_7249,N_5816,N_5117);
nand U7250 (N_7250,N_5947,N_5525);
xnor U7251 (N_7251,N_5978,N_5935);
nand U7252 (N_7252,N_6000,N_5240);
and U7253 (N_7253,N_5989,N_5204);
and U7254 (N_7254,N_5101,N_5015);
or U7255 (N_7255,N_5311,N_6056);
or U7256 (N_7256,N_5785,N_5779);
nor U7257 (N_7257,N_5981,N_5446);
nand U7258 (N_7258,N_5034,N_6195);
or U7259 (N_7259,N_5897,N_6003);
xnor U7260 (N_7260,N_5216,N_5257);
nand U7261 (N_7261,N_5042,N_5027);
nor U7262 (N_7262,N_6111,N_5875);
nor U7263 (N_7263,N_6149,N_5087);
and U7264 (N_7264,N_5587,N_5706);
nand U7265 (N_7265,N_5945,N_5774);
or U7266 (N_7266,N_6153,N_5543);
xnor U7267 (N_7267,N_6139,N_5177);
nor U7268 (N_7268,N_5231,N_5041);
or U7269 (N_7269,N_5975,N_6139);
nand U7270 (N_7270,N_5747,N_5128);
nor U7271 (N_7271,N_5571,N_5317);
and U7272 (N_7272,N_6146,N_5448);
or U7273 (N_7273,N_5910,N_5311);
nor U7274 (N_7274,N_5153,N_5217);
and U7275 (N_7275,N_5957,N_5002);
xor U7276 (N_7276,N_5979,N_5693);
and U7277 (N_7277,N_5948,N_5886);
xnor U7278 (N_7278,N_5517,N_5689);
nor U7279 (N_7279,N_5231,N_5955);
or U7280 (N_7280,N_6246,N_5931);
nor U7281 (N_7281,N_5633,N_5542);
or U7282 (N_7282,N_5018,N_5704);
xor U7283 (N_7283,N_5267,N_5112);
or U7284 (N_7284,N_5944,N_5688);
and U7285 (N_7285,N_5893,N_5500);
nor U7286 (N_7286,N_5464,N_5611);
nand U7287 (N_7287,N_6023,N_5024);
nor U7288 (N_7288,N_5671,N_5395);
xnor U7289 (N_7289,N_6131,N_5929);
nor U7290 (N_7290,N_5688,N_5831);
and U7291 (N_7291,N_5930,N_5221);
or U7292 (N_7292,N_5210,N_6012);
and U7293 (N_7293,N_5403,N_5605);
and U7294 (N_7294,N_5532,N_5263);
and U7295 (N_7295,N_5419,N_5073);
and U7296 (N_7296,N_6248,N_5370);
and U7297 (N_7297,N_5329,N_6067);
or U7298 (N_7298,N_5538,N_5420);
or U7299 (N_7299,N_5102,N_5625);
and U7300 (N_7300,N_5135,N_5093);
or U7301 (N_7301,N_5635,N_5132);
nor U7302 (N_7302,N_6047,N_5389);
nor U7303 (N_7303,N_5431,N_5921);
or U7304 (N_7304,N_5370,N_5272);
xnor U7305 (N_7305,N_5306,N_6158);
xnor U7306 (N_7306,N_5254,N_5721);
xor U7307 (N_7307,N_5955,N_5523);
nand U7308 (N_7308,N_5623,N_5874);
or U7309 (N_7309,N_6038,N_5048);
or U7310 (N_7310,N_5552,N_5976);
or U7311 (N_7311,N_5494,N_5517);
or U7312 (N_7312,N_5050,N_5330);
xor U7313 (N_7313,N_5227,N_5358);
nor U7314 (N_7314,N_6014,N_5481);
or U7315 (N_7315,N_6065,N_5594);
xor U7316 (N_7316,N_5142,N_5050);
nor U7317 (N_7317,N_5353,N_5561);
nand U7318 (N_7318,N_5020,N_5341);
xor U7319 (N_7319,N_5289,N_5812);
nor U7320 (N_7320,N_5699,N_5453);
nand U7321 (N_7321,N_5854,N_6003);
and U7322 (N_7322,N_6135,N_5765);
or U7323 (N_7323,N_5687,N_5531);
nor U7324 (N_7324,N_5734,N_5694);
nand U7325 (N_7325,N_5697,N_5825);
xnor U7326 (N_7326,N_6228,N_5966);
nor U7327 (N_7327,N_5396,N_5257);
or U7328 (N_7328,N_5904,N_5923);
xor U7329 (N_7329,N_5870,N_5983);
xor U7330 (N_7330,N_5293,N_5248);
and U7331 (N_7331,N_6212,N_5538);
or U7332 (N_7332,N_5879,N_5095);
or U7333 (N_7333,N_6003,N_5201);
nor U7334 (N_7334,N_5989,N_5193);
or U7335 (N_7335,N_6218,N_5834);
nor U7336 (N_7336,N_5230,N_5521);
or U7337 (N_7337,N_5136,N_5924);
nand U7338 (N_7338,N_5431,N_5145);
nand U7339 (N_7339,N_5703,N_6115);
and U7340 (N_7340,N_5004,N_5078);
xor U7341 (N_7341,N_5000,N_6103);
nand U7342 (N_7342,N_5107,N_6000);
nand U7343 (N_7343,N_6192,N_5534);
nor U7344 (N_7344,N_5677,N_5785);
and U7345 (N_7345,N_5169,N_6120);
nor U7346 (N_7346,N_6217,N_5196);
nand U7347 (N_7347,N_5851,N_5406);
xnor U7348 (N_7348,N_5636,N_6079);
and U7349 (N_7349,N_5443,N_5976);
or U7350 (N_7350,N_5437,N_5316);
nand U7351 (N_7351,N_6216,N_6179);
and U7352 (N_7352,N_5937,N_5998);
and U7353 (N_7353,N_5060,N_5677);
nor U7354 (N_7354,N_5865,N_6243);
and U7355 (N_7355,N_5342,N_5455);
or U7356 (N_7356,N_5008,N_5793);
nor U7357 (N_7357,N_5893,N_6155);
xnor U7358 (N_7358,N_5988,N_5556);
xor U7359 (N_7359,N_6211,N_6225);
or U7360 (N_7360,N_6071,N_6044);
or U7361 (N_7361,N_6017,N_5506);
nand U7362 (N_7362,N_5554,N_6074);
xnor U7363 (N_7363,N_5960,N_5063);
nor U7364 (N_7364,N_5091,N_5857);
nand U7365 (N_7365,N_5964,N_5235);
and U7366 (N_7366,N_5535,N_6086);
or U7367 (N_7367,N_5646,N_5566);
or U7368 (N_7368,N_5194,N_5236);
or U7369 (N_7369,N_6113,N_5507);
nor U7370 (N_7370,N_6165,N_6154);
and U7371 (N_7371,N_5747,N_6074);
and U7372 (N_7372,N_5206,N_6169);
xnor U7373 (N_7373,N_5511,N_5221);
nor U7374 (N_7374,N_5092,N_5160);
nor U7375 (N_7375,N_6191,N_5466);
or U7376 (N_7376,N_5329,N_5615);
xnor U7377 (N_7377,N_5347,N_5832);
nor U7378 (N_7378,N_5687,N_5601);
nor U7379 (N_7379,N_5727,N_5710);
nor U7380 (N_7380,N_6129,N_5541);
and U7381 (N_7381,N_5464,N_6056);
xor U7382 (N_7382,N_5831,N_6163);
xnor U7383 (N_7383,N_5854,N_5065);
and U7384 (N_7384,N_5766,N_6113);
nand U7385 (N_7385,N_5835,N_5805);
or U7386 (N_7386,N_5304,N_5531);
or U7387 (N_7387,N_5252,N_5902);
or U7388 (N_7388,N_5479,N_6021);
nand U7389 (N_7389,N_5817,N_5796);
nor U7390 (N_7390,N_5036,N_5733);
nor U7391 (N_7391,N_5657,N_5562);
nand U7392 (N_7392,N_5641,N_5385);
nand U7393 (N_7393,N_5912,N_5082);
and U7394 (N_7394,N_6220,N_5776);
xor U7395 (N_7395,N_5722,N_5880);
nand U7396 (N_7396,N_5336,N_6232);
or U7397 (N_7397,N_5731,N_5341);
xor U7398 (N_7398,N_5180,N_5606);
or U7399 (N_7399,N_6093,N_5212);
or U7400 (N_7400,N_6238,N_5226);
and U7401 (N_7401,N_5779,N_5950);
and U7402 (N_7402,N_5368,N_5917);
and U7403 (N_7403,N_6089,N_5476);
xnor U7404 (N_7404,N_5845,N_5691);
xor U7405 (N_7405,N_5047,N_6239);
and U7406 (N_7406,N_5126,N_5834);
and U7407 (N_7407,N_5187,N_5795);
and U7408 (N_7408,N_5430,N_5344);
nor U7409 (N_7409,N_6048,N_6183);
and U7410 (N_7410,N_5719,N_5857);
nand U7411 (N_7411,N_5799,N_5858);
or U7412 (N_7412,N_5103,N_5566);
nand U7413 (N_7413,N_5365,N_6201);
nor U7414 (N_7414,N_6122,N_5220);
or U7415 (N_7415,N_5381,N_5948);
nand U7416 (N_7416,N_5715,N_5413);
or U7417 (N_7417,N_5086,N_5450);
nand U7418 (N_7418,N_5506,N_5268);
nand U7419 (N_7419,N_5751,N_5870);
nor U7420 (N_7420,N_5815,N_5332);
or U7421 (N_7421,N_5322,N_5527);
nand U7422 (N_7422,N_5142,N_5978);
nor U7423 (N_7423,N_5322,N_5055);
xor U7424 (N_7424,N_5022,N_5277);
and U7425 (N_7425,N_6069,N_5530);
xnor U7426 (N_7426,N_5726,N_5402);
xnor U7427 (N_7427,N_5709,N_5519);
xnor U7428 (N_7428,N_5004,N_5905);
and U7429 (N_7429,N_5493,N_5486);
and U7430 (N_7430,N_5741,N_5653);
or U7431 (N_7431,N_5634,N_5315);
nand U7432 (N_7432,N_5432,N_5066);
or U7433 (N_7433,N_5571,N_5819);
nor U7434 (N_7434,N_5468,N_5697);
xnor U7435 (N_7435,N_5052,N_5386);
and U7436 (N_7436,N_5002,N_5017);
nand U7437 (N_7437,N_5748,N_5443);
or U7438 (N_7438,N_5421,N_6195);
or U7439 (N_7439,N_5996,N_5718);
xnor U7440 (N_7440,N_5808,N_5461);
and U7441 (N_7441,N_5735,N_5156);
nor U7442 (N_7442,N_5953,N_6118);
xor U7443 (N_7443,N_5295,N_5492);
or U7444 (N_7444,N_5890,N_6196);
and U7445 (N_7445,N_5350,N_5634);
and U7446 (N_7446,N_5713,N_5638);
and U7447 (N_7447,N_5461,N_5591);
nor U7448 (N_7448,N_5265,N_5624);
nand U7449 (N_7449,N_5243,N_5356);
or U7450 (N_7450,N_5576,N_5029);
nor U7451 (N_7451,N_5478,N_6163);
nor U7452 (N_7452,N_5304,N_5106);
xor U7453 (N_7453,N_5606,N_5568);
nor U7454 (N_7454,N_5409,N_5616);
or U7455 (N_7455,N_5056,N_5488);
or U7456 (N_7456,N_5295,N_5228);
xnor U7457 (N_7457,N_5217,N_5367);
nor U7458 (N_7458,N_6042,N_6209);
nand U7459 (N_7459,N_5913,N_5846);
or U7460 (N_7460,N_5706,N_5054);
or U7461 (N_7461,N_5948,N_5655);
or U7462 (N_7462,N_5627,N_6032);
and U7463 (N_7463,N_6212,N_6205);
or U7464 (N_7464,N_5722,N_6238);
nand U7465 (N_7465,N_5517,N_5701);
or U7466 (N_7466,N_5621,N_5109);
xor U7467 (N_7467,N_5715,N_6188);
nor U7468 (N_7468,N_5738,N_5897);
and U7469 (N_7469,N_5535,N_5721);
nand U7470 (N_7470,N_6206,N_5497);
xnor U7471 (N_7471,N_5873,N_5108);
or U7472 (N_7472,N_6056,N_5031);
and U7473 (N_7473,N_5403,N_5057);
nor U7474 (N_7474,N_5474,N_5089);
nor U7475 (N_7475,N_5300,N_6011);
and U7476 (N_7476,N_6215,N_5414);
nand U7477 (N_7477,N_5462,N_5517);
nor U7478 (N_7478,N_6106,N_6124);
or U7479 (N_7479,N_5877,N_6076);
xor U7480 (N_7480,N_5808,N_5198);
nor U7481 (N_7481,N_6003,N_5823);
nor U7482 (N_7482,N_5493,N_6007);
nand U7483 (N_7483,N_5717,N_5593);
xor U7484 (N_7484,N_5347,N_5543);
nand U7485 (N_7485,N_5524,N_5320);
nor U7486 (N_7486,N_5712,N_6176);
nor U7487 (N_7487,N_5341,N_5260);
nand U7488 (N_7488,N_5253,N_5340);
xnor U7489 (N_7489,N_5564,N_5405);
xnor U7490 (N_7490,N_5723,N_5300);
nand U7491 (N_7491,N_6223,N_5106);
xor U7492 (N_7492,N_5294,N_5808);
or U7493 (N_7493,N_5643,N_6023);
nor U7494 (N_7494,N_6096,N_5468);
and U7495 (N_7495,N_5981,N_6101);
and U7496 (N_7496,N_5713,N_5992);
xnor U7497 (N_7497,N_5637,N_6002);
xnor U7498 (N_7498,N_6092,N_5564);
and U7499 (N_7499,N_5427,N_6044);
nor U7500 (N_7500,N_7279,N_6992);
nand U7501 (N_7501,N_7393,N_6943);
nor U7502 (N_7502,N_6469,N_6779);
or U7503 (N_7503,N_7210,N_7420);
nand U7504 (N_7504,N_7088,N_6482);
nand U7505 (N_7505,N_6912,N_6823);
and U7506 (N_7506,N_6502,N_6840);
nand U7507 (N_7507,N_7077,N_7196);
or U7508 (N_7508,N_6807,N_6980);
and U7509 (N_7509,N_7058,N_6302);
xor U7510 (N_7510,N_6820,N_7296);
or U7511 (N_7511,N_6527,N_7485);
nor U7512 (N_7512,N_6568,N_6949);
nor U7513 (N_7513,N_7273,N_6917);
xnor U7514 (N_7514,N_6539,N_6273);
and U7515 (N_7515,N_7452,N_6562);
xnor U7516 (N_7516,N_6853,N_6848);
nand U7517 (N_7517,N_6261,N_6587);
or U7518 (N_7518,N_6269,N_6277);
and U7519 (N_7519,N_6579,N_6691);
nand U7520 (N_7520,N_7321,N_6835);
or U7521 (N_7521,N_7234,N_6343);
or U7522 (N_7522,N_6530,N_7072);
nand U7523 (N_7523,N_6485,N_6729);
and U7524 (N_7524,N_7075,N_6792);
nor U7525 (N_7525,N_7397,N_7489);
and U7526 (N_7526,N_6793,N_6958);
and U7527 (N_7527,N_6459,N_7112);
and U7528 (N_7528,N_6726,N_7410);
and U7529 (N_7529,N_7288,N_6760);
nand U7530 (N_7530,N_7154,N_6250);
and U7531 (N_7531,N_6412,N_6311);
or U7532 (N_7532,N_7428,N_7053);
or U7533 (N_7533,N_6493,N_7156);
nand U7534 (N_7534,N_6800,N_6531);
xor U7535 (N_7535,N_7046,N_7498);
nor U7536 (N_7536,N_6518,N_6836);
and U7537 (N_7537,N_6329,N_7435);
nand U7538 (N_7538,N_6733,N_6477);
nand U7539 (N_7539,N_7318,N_7097);
nor U7540 (N_7540,N_6395,N_7176);
and U7541 (N_7541,N_7221,N_6722);
nand U7542 (N_7542,N_6920,N_6745);
or U7543 (N_7543,N_7301,N_7206);
nor U7544 (N_7544,N_7125,N_7089);
nor U7545 (N_7545,N_6418,N_7385);
nor U7546 (N_7546,N_6400,N_6725);
or U7547 (N_7547,N_7329,N_6950);
xor U7548 (N_7548,N_7354,N_7023);
xor U7549 (N_7549,N_6609,N_6638);
and U7550 (N_7550,N_7025,N_6580);
or U7551 (N_7551,N_7412,N_6782);
and U7552 (N_7552,N_6285,N_6647);
nor U7553 (N_7553,N_6289,N_6936);
and U7554 (N_7554,N_6666,N_7267);
nand U7555 (N_7555,N_7158,N_6746);
nand U7556 (N_7556,N_6721,N_7457);
xnor U7557 (N_7557,N_6299,N_6708);
nor U7558 (N_7558,N_7306,N_6436);
nor U7559 (N_7559,N_6762,N_6690);
and U7560 (N_7560,N_7418,N_7143);
or U7561 (N_7561,N_7099,N_7050);
and U7562 (N_7562,N_6942,N_7269);
nand U7563 (N_7563,N_6463,N_6780);
xor U7564 (N_7564,N_6737,N_6611);
and U7565 (N_7565,N_6319,N_7432);
nor U7566 (N_7566,N_6529,N_7482);
nand U7567 (N_7567,N_7049,N_6614);
nor U7568 (N_7568,N_6607,N_7363);
or U7569 (N_7569,N_6781,N_6264);
or U7570 (N_7570,N_6565,N_7274);
and U7571 (N_7571,N_6447,N_6973);
or U7572 (N_7572,N_6382,N_7038);
nor U7573 (N_7573,N_6483,N_6589);
nor U7574 (N_7574,N_7396,N_6754);
or U7575 (N_7575,N_6694,N_7226);
nor U7576 (N_7576,N_7126,N_6918);
xor U7577 (N_7577,N_6724,N_7483);
and U7578 (N_7578,N_6506,N_6255);
nor U7579 (N_7579,N_7240,N_7365);
nand U7580 (N_7580,N_6718,N_7350);
nor U7581 (N_7581,N_6643,N_6528);
or U7582 (N_7582,N_6897,N_7081);
nor U7583 (N_7583,N_6676,N_6372);
or U7584 (N_7584,N_6898,N_6639);
xnor U7585 (N_7585,N_6636,N_6685);
nand U7586 (N_7586,N_7106,N_6444);
nand U7587 (N_7587,N_6271,N_7451);
nand U7588 (N_7588,N_7445,N_6838);
and U7589 (N_7589,N_7473,N_7317);
xor U7590 (N_7590,N_6410,N_6542);
nor U7591 (N_7591,N_6773,N_7007);
nand U7592 (N_7592,N_7311,N_6703);
xor U7593 (N_7593,N_7183,N_6561);
and U7594 (N_7594,N_7228,N_6866);
or U7595 (N_7595,N_6660,N_7233);
nand U7596 (N_7596,N_7337,N_6262);
nand U7597 (N_7597,N_7167,N_7446);
or U7598 (N_7598,N_7031,N_7387);
or U7599 (N_7599,N_7402,N_6507);
nor U7600 (N_7600,N_7111,N_6964);
or U7601 (N_7601,N_6550,N_7254);
and U7602 (N_7602,N_6769,N_6628);
or U7603 (N_7603,N_6486,N_6505);
xnor U7604 (N_7604,N_6736,N_7180);
xnor U7605 (N_7605,N_7212,N_7359);
nor U7606 (N_7606,N_6925,N_7448);
or U7607 (N_7607,N_6849,N_6668);
nor U7608 (N_7608,N_6496,N_7235);
nor U7609 (N_7609,N_6605,N_6368);
and U7610 (N_7610,N_7048,N_6409);
nand U7611 (N_7611,N_7401,N_7458);
xor U7612 (N_7612,N_6624,N_6476);
nor U7613 (N_7613,N_6998,N_6837);
nand U7614 (N_7614,N_6543,N_6442);
or U7615 (N_7615,N_7471,N_6545);
and U7616 (N_7616,N_7065,N_7142);
or U7617 (N_7617,N_7360,N_6510);
nor U7618 (N_7618,N_7144,N_6830);
nor U7619 (N_7619,N_6306,N_7199);
and U7620 (N_7620,N_7152,N_6832);
or U7621 (N_7621,N_6683,N_6880);
xnor U7622 (N_7622,N_7343,N_6675);
xor U7623 (N_7623,N_6581,N_7488);
nand U7624 (N_7624,N_6524,N_7316);
and U7625 (N_7625,N_6615,N_6604);
nand U7626 (N_7626,N_6622,N_7093);
nand U7627 (N_7627,N_7484,N_6821);
nor U7628 (N_7628,N_7164,N_6598);
xnor U7629 (N_7629,N_6787,N_6514);
nand U7630 (N_7630,N_7487,N_6327);
xnor U7631 (N_7631,N_6759,N_7377);
nor U7632 (N_7632,N_6602,N_6411);
nand U7633 (N_7633,N_6603,N_7021);
nand U7634 (N_7634,N_7422,N_6612);
or U7635 (N_7635,N_6620,N_7294);
nand U7636 (N_7636,N_6532,N_7364);
xor U7637 (N_7637,N_6574,N_6474);
xor U7638 (N_7638,N_7168,N_6549);
nand U7639 (N_7639,N_7309,N_7148);
xnor U7640 (N_7640,N_7016,N_7115);
or U7641 (N_7641,N_6886,N_6903);
or U7642 (N_7642,N_6921,N_7315);
nor U7643 (N_7643,N_7101,N_6297);
and U7644 (N_7644,N_6796,N_6361);
and U7645 (N_7645,N_7278,N_7000);
or U7646 (N_7646,N_7320,N_7474);
and U7647 (N_7647,N_6687,N_6259);
xor U7648 (N_7648,N_7389,N_6422);
xnor U7649 (N_7649,N_6872,N_6349);
or U7650 (N_7650,N_7182,N_6592);
or U7651 (N_7651,N_7208,N_7461);
or U7652 (N_7652,N_7314,N_6952);
or U7653 (N_7653,N_6630,N_7263);
and U7654 (N_7654,N_6583,N_6825);
and U7655 (N_7655,N_6446,N_6650);
xnor U7656 (N_7656,N_6460,N_7270);
nand U7657 (N_7657,N_6803,N_6670);
nor U7658 (N_7658,N_6572,N_6326);
nor U7659 (N_7659,N_6944,N_6540);
nor U7660 (N_7660,N_7127,N_6938);
xnor U7661 (N_7661,N_6352,N_6727);
and U7662 (N_7662,N_7004,N_7366);
xnor U7663 (N_7663,N_6342,N_7114);
xor U7664 (N_7664,N_6437,N_6286);
xor U7665 (N_7665,N_6279,N_6535);
and U7666 (N_7666,N_6818,N_7223);
xnor U7667 (N_7667,N_6929,N_7014);
or U7668 (N_7668,N_6902,N_6559);
nand U7669 (N_7669,N_6979,N_7486);
and U7670 (N_7670,N_7376,N_7430);
or U7671 (N_7671,N_6582,N_6257);
and U7672 (N_7672,N_6495,N_6310);
or U7673 (N_7673,N_7247,N_6619);
or U7674 (N_7674,N_7382,N_6627);
or U7675 (N_7675,N_6430,N_7424);
xnor U7676 (N_7676,N_7024,N_6516);
nor U7677 (N_7677,N_6906,N_7224);
nand U7678 (N_7678,N_7204,N_6993);
xor U7679 (N_7679,N_6435,N_7059);
xnor U7680 (N_7680,N_6616,N_6263);
nor U7681 (N_7681,N_7417,N_7078);
nand U7682 (N_7682,N_6290,N_6710);
and U7683 (N_7683,N_6308,N_6696);
or U7684 (N_7684,N_6366,N_6320);
nor U7685 (N_7685,N_6939,N_7032);
nor U7686 (N_7686,N_6995,N_6945);
and U7687 (N_7687,N_7439,N_6744);
nand U7688 (N_7688,N_6763,N_6864);
nand U7689 (N_7689,N_6909,N_6775);
nand U7690 (N_7690,N_7336,N_6393);
nand U7691 (N_7691,N_7478,N_6251);
or U7692 (N_7692,N_7444,N_7388);
nor U7693 (N_7693,N_6719,N_7197);
xor U7694 (N_7694,N_6371,N_6802);
or U7695 (N_7695,N_7098,N_6834);
nand U7696 (N_7696,N_6323,N_7022);
and U7697 (N_7697,N_6613,N_7283);
and U7698 (N_7698,N_7150,N_6546);
or U7699 (N_7699,N_6651,N_7241);
xnor U7700 (N_7700,N_6312,N_7145);
xnor U7701 (N_7701,N_6480,N_6623);
or U7702 (N_7702,N_6711,N_6738);
xnor U7703 (N_7703,N_7230,N_6552);
and U7704 (N_7704,N_6987,N_6573);
and U7705 (N_7705,N_6294,N_6978);
nand U7706 (N_7706,N_6369,N_7490);
nor U7707 (N_7707,N_6593,N_6862);
and U7708 (N_7708,N_7450,N_7379);
or U7709 (N_7709,N_6567,N_7341);
xnor U7710 (N_7710,N_6934,N_6896);
nor U7711 (N_7711,N_7459,N_7147);
or U7712 (N_7712,N_6791,N_7330);
nor U7713 (N_7713,N_7003,N_7431);
xor U7714 (N_7714,N_6337,N_7340);
or U7715 (N_7715,N_6827,N_6932);
or U7716 (N_7716,N_7352,N_7061);
xnor U7717 (N_7717,N_6901,N_7104);
nand U7718 (N_7718,N_6272,N_6481);
nand U7719 (N_7719,N_6700,N_6662);
nand U7720 (N_7720,N_6566,N_7079);
nor U7721 (N_7721,N_7013,N_6503);
and U7722 (N_7722,N_6307,N_6431);
nor U7723 (N_7723,N_7259,N_7463);
nor U7724 (N_7724,N_6657,N_7286);
or U7725 (N_7725,N_6874,N_6956);
xnor U7726 (N_7726,N_7056,N_6723);
and U7727 (N_7727,N_6734,N_6984);
xor U7728 (N_7728,N_6653,N_7066);
and U7729 (N_7729,N_6955,N_6692);
nand U7730 (N_7730,N_7429,N_6776);
or U7731 (N_7731,N_6799,N_6895);
or U7732 (N_7732,N_7277,N_6768);
nor U7733 (N_7733,N_6808,N_6801);
or U7734 (N_7734,N_7477,N_6680);
xor U7735 (N_7735,N_6714,N_6946);
xnor U7736 (N_7736,N_6771,N_7189);
and U7737 (N_7737,N_7476,N_7123);
xnor U7738 (N_7738,N_6288,N_6826);
and U7739 (N_7739,N_6487,N_6332);
or U7740 (N_7740,N_6293,N_6440);
or U7741 (N_7741,N_6421,N_6875);
and U7742 (N_7742,N_7047,N_6785);
xnor U7743 (N_7743,N_6961,N_7391);
and U7744 (N_7744,N_6538,N_6965);
nand U7745 (N_7745,N_6656,N_6515);
and U7746 (N_7746,N_7082,N_7120);
and U7747 (N_7747,N_6355,N_6570);
and U7748 (N_7748,N_7002,N_7102);
or U7749 (N_7749,N_6789,N_6260);
or U7750 (N_7750,N_7362,N_7149);
and U7751 (N_7751,N_6554,N_6595);
nor U7752 (N_7752,N_6816,N_6497);
xnor U7753 (N_7753,N_6797,N_7361);
nand U7754 (N_7754,N_6910,N_6625);
nand U7755 (N_7755,N_6673,N_6974);
xnor U7756 (N_7756,N_6633,N_6885);
or U7757 (N_7757,N_7438,N_6869);
or U7758 (N_7758,N_7260,N_6427);
xnor U7759 (N_7759,N_6686,N_6353);
xor U7760 (N_7760,N_6341,N_7371);
nor U7761 (N_7761,N_7403,N_6815);
nand U7762 (N_7762,N_6606,N_7172);
or U7763 (N_7763,N_6465,N_7261);
or U7764 (N_7764,N_6968,N_7338);
xor U7765 (N_7765,N_6387,N_7019);
xnor U7766 (N_7766,N_7119,N_7480);
or U7767 (N_7767,N_7054,N_6743);
or U7768 (N_7768,N_7243,N_6253);
xnor U7769 (N_7769,N_7117,N_7229);
or U7770 (N_7770,N_7236,N_6588);
xnor U7771 (N_7771,N_6907,N_6316);
or U7772 (N_7772,N_7005,N_6536);
xor U7773 (N_7773,N_6766,N_7174);
nand U7774 (N_7774,N_6520,N_6394);
nor U7775 (N_7775,N_7035,N_6985);
nand U7776 (N_7776,N_7033,N_7238);
nand U7777 (N_7777,N_6937,N_6865);
or U7778 (N_7778,N_6664,N_6585);
xnor U7779 (N_7779,N_7335,N_7372);
nand U7780 (N_7780,N_7251,N_7434);
or U7781 (N_7781,N_7185,N_6557);
and U7782 (N_7782,N_6809,N_6709);
xnor U7783 (N_7783,N_6911,N_7357);
xnor U7784 (N_7784,N_6900,N_7194);
and U7785 (N_7785,N_7384,N_6720);
and U7786 (N_7786,N_6892,N_6810);
nor U7787 (N_7787,N_7456,N_7497);
xnor U7788 (N_7788,N_6697,N_7460);
nor U7789 (N_7789,N_7297,N_7442);
and U7790 (N_7790,N_6578,N_7266);
xor U7791 (N_7791,N_7055,N_6863);
or U7792 (N_7792,N_7281,N_6357);
and U7793 (N_7793,N_6940,N_6432);
and U7794 (N_7794,N_6695,N_6661);
xnor U7795 (N_7795,N_7390,N_6850);
nor U7796 (N_7796,N_6547,N_6556);
nor U7797 (N_7797,N_6795,N_7249);
xor U7798 (N_7798,N_7063,N_7289);
and U7799 (N_7799,N_7245,N_7121);
and U7800 (N_7800,N_7256,N_7310);
or U7801 (N_7801,N_7303,N_6379);
or U7802 (N_7802,N_7153,N_6458);
nand U7803 (N_7803,N_6904,N_6915);
nand U7804 (N_7804,N_6812,N_6972);
and U7805 (N_7805,N_6464,N_7349);
or U7806 (N_7806,N_6999,N_6313);
nor U7807 (N_7807,N_6389,N_7400);
nor U7808 (N_7808,N_6391,N_6748);
nor U7809 (N_7809,N_6752,N_6635);
and U7810 (N_7810,N_7322,N_6504);
or U7811 (N_7811,N_7109,N_6989);
nand U7812 (N_7812,N_6742,N_7344);
xnor U7813 (N_7813,N_7227,N_6665);
xor U7814 (N_7814,N_7140,N_7200);
nand U7815 (N_7815,N_7324,N_6935);
nand U7816 (N_7816,N_7447,N_6363);
or U7817 (N_7817,N_6451,N_6479);
nor U7818 (N_7818,N_7203,N_6541);
nand U7819 (N_7819,N_6462,N_6854);
xor U7820 (N_7820,N_6916,N_6354);
or U7821 (N_7821,N_7380,N_6772);
nor U7822 (N_7822,N_6891,N_7348);
nand U7823 (N_7823,N_6908,N_7179);
nand U7824 (N_7824,N_6362,N_7220);
xor U7825 (N_7825,N_6969,N_6356);
or U7826 (N_7826,N_7437,N_6889);
xor U7827 (N_7827,N_6621,N_7239);
nor U7828 (N_7828,N_7202,N_6484);
and U7829 (N_7829,N_6649,N_7037);
and U7830 (N_7830,N_7181,N_6986);
xnor U7831 (N_7831,N_6684,N_7333);
nor U7832 (N_7832,N_7467,N_7201);
nor U7833 (N_7833,N_6674,N_6617);
xor U7834 (N_7834,N_6663,N_6367);
nor U7835 (N_7835,N_6383,N_6571);
nor U7836 (N_7836,N_6919,N_6870);
or U7837 (N_7837,N_6377,N_6677);
nor U7838 (N_7838,N_6632,N_7177);
xor U7839 (N_7839,N_7253,N_6804);
or U7840 (N_7840,N_7124,N_6735);
nor U7841 (N_7841,N_6267,N_6640);
or U7842 (N_7842,N_6659,N_6702);
xor U7843 (N_7843,N_7017,N_6478);
nor U7844 (N_7844,N_7421,N_6596);
nor U7845 (N_7845,N_6511,N_7345);
xor U7846 (N_7846,N_7096,N_7358);
or U7847 (N_7847,N_7195,N_7076);
nand U7848 (N_7848,N_6280,N_6879);
nor U7849 (N_7849,N_7231,N_7041);
or U7850 (N_7850,N_6758,N_7378);
nand U7851 (N_7851,N_6774,N_6433);
nand U7852 (N_7852,N_6948,N_7392);
or U7853 (N_7853,N_7155,N_6303);
xor U7854 (N_7854,N_6777,N_6330);
nor U7855 (N_7855,N_6334,N_7427);
nor U7856 (N_7856,N_6499,N_6378);
or U7857 (N_7857,N_6652,N_7469);
or U7858 (N_7858,N_7134,N_7009);
or U7859 (N_7859,N_7369,N_7129);
or U7860 (N_7860,N_7373,N_6519);
or U7861 (N_7861,N_6429,N_6441);
or U7862 (N_7862,N_6309,N_6689);
or U7863 (N_7863,N_6454,N_6407);
nand U7864 (N_7864,N_6388,N_7029);
or U7865 (N_7865,N_7415,N_6526);
xor U7866 (N_7866,N_7346,N_7113);
or U7867 (N_7867,N_6560,N_7067);
or U7868 (N_7868,N_7043,N_6851);
xor U7869 (N_7869,N_6404,N_6295);
xnor U7870 (N_7870,N_7295,N_6730);
xnor U7871 (N_7871,N_6301,N_6890);
nor U7872 (N_7872,N_6704,N_7213);
xor U7873 (N_7873,N_6646,N_6860);
or U7874 (N_7874,N_6600,N_7328);
and U7875 (N_7875,N_6765,N_6266);
and U7876 (N_7876,N_6951,N_7095);
xnor U7877 (N_7877,N_6913,N_6899);
and U7878 (N_7878,N_7108,N_6941);
xnor U7879 (N_7879,N_6894,N_6406);
or U7880 (N_7880,N_7250,N_6811);
nand U7881 (N_7881,N_6461,N_7219);
nor U7882 (N_7882,N_7215,N_6275);
nor U7883 (N_7883,N_6551,N_7441);
nor U7884 (N_7884,N_6281,N_6416);
xnor U7885 (N_7885,N_7091,N_6473);
and U7886 (N_7886,N_7170,N_7068);
xnor U7887 (N_7887,N_7064,N_6822);
nor U7888 (N_7888,N_7405,N_6601);
nand U7889 (N_7889,N_6284,N_6975);
xnor U7890 (N_7890,N_7028,N_6268);
nor U7891 (N_7891,N_6976,N_7280);
xor U7892 (N_7892,N_6732,N_7413);
nor U7893 (N_7893,N_6755,N_7375);
nor U7894 (N_7894,N_6492,N_6386);
xnor U7895 (N_7895,N_7175,N_6555);
or U7896 (N_7896,N_6424,N_6928);
nor U7897 (N_7897,N_7408,N_7087);
or U7898 (N_7898,N_7205,N_6877);
nand U7899 (N_7899,N_6428,N_7414);
xnor U7900 (N_7900,N_6390,N_6924);
or U7901 (N_7901,N_6591,N_7398);
or U7902 (N_7902,N_7299,N_6586);
nand U7903 (N_7903,N_7036,N_7313);
nand U7904 (N_7904,N_7130,N_7433);
nand U7905 (N_7905,N_7131,N_6346);
or U7906 (N_7906,N_6857,N_7479);
nand U7907 (N_7907,N_6831,N_6883);
xor U7908 (N_7908,N_6548,N_7464);
xor U7909 (N_7909,N_6788,N_6618);
and U7910 (N_7910,N_6882,N_6265);
xnor U7911 (N_7911,N_7045,N_6728);
or U7912 (N_7912,N_6876,N_7381);
nand U7913 (N_7913,N_6971,N_6402);
xnor U7914 (N_7914,N_6715,N_6576);
and U7915 (N_7915,N_7186,N_6868);
and U7916 (N_7916,N_6521,N_7449);
nand U7917 (N_7917,N_6648,N_6452);
nand U7918 (N_7918,N_6977,N_6914);
xor U7919 (N_7919,N_7207,N_7118);
nand U7920 (N_7920,N_7496,N_6384);
nand U7921 (N_7921,N_7105,N_7103);
nor U7922 (N_7922,N_7425,N_6450);
and U7923 (N_7923,N_6610,N_7347);
nand U7924 (N_7924,N_6375,N_7339);
nand U7925 (N_7925,N_7020,N_7436);
nor U7926 (N_7926,N_7018,N_6873);
xnor U7927 (N_7927,N_7242,N_6399);
nand U7928 (N_7928,N_6888,N_6923);
nand U7929 (N_7929,N_6324,N_7161);
xor U7930 (N_7930,N_7006,N_6360);
xor U7931 (N_7931,N_6962,N_6642);
xnor U7932 (N_7932,N_7304,N_7472);
nor U7933 (N_7933,N_7423,N_6842);
nor U7934 (N_7934,N_7248,N_6905);
nand U7935 (N_7935,N_7191,N_6339);
or U7936 (N_7936,N_7015,N_6833);
or U7937 (N_7937,N_7034,N_7374);
xor U7938 (N_7938,N_7198,N_6466);
nor U7939 (N_7939,N_6252,N_6654);
nor U7940 (N_7940,N_7331,N_6322);
and U7941 (N_7941,N_6373,N_6824);
xnor U7942 (N_7942,N_7368,N_7351);
nor U7943 (N_7943,N_6449,N_7494);
nand U7944 (N_7944,N_7030,N_6798);
xor U7945 (N_7945,N_6629,N_6359);
xor U7946 (N_7946,N_7443,N_6828);
and U7947 (N_7947,N_7305,N_6438);
nand U7948 (N_7948,N_7416,N_7169);
nor U7949 (N_7949,N_7468,N_6858);
or U7950 (N_7950,N_7308,N_6698);
nand U7951 (N_7951,N_6364,N_7367);
nor U7952 (N_7952,N_6403,N_7492);
and U7953 (N_7953,N_6300,N_6522);
or U7954 (N_7954,N_7291,N_6996);
nand U7955 (N_7955,N_6751,N_7052);
or U7956 (N_7956,N_6852,N_6374);
xor U7957 (N_7957,N_6445,N_7332);
xor U7958 (N_7958,N_7454,N_7342);
xor U7959 (N_7959,N_7455,N_7462);
or U7960 (N_7960,N_6739,N_6786);
or U7961 (N_7961,N_6381,N_7162);
xnor U7962 (N_7962,N_7298,N_7257);
nor U7963 (N_7963,N_7327,N_7166);
or U7964 (N_7964,N_6350,N_6489);
and U7965 (N_7965,N_7128,N_6455);
nand U7966 (N_7966,N_6867,N_6509);
nor U7967 (N_7967,N_6457,N_7107);
or U7968 (N_7968,N_6523,N_7264);
nand U7969 (N_7969,N_6966,N_7040);
nor U7970 (N_7970,N_7323,N_7453);
nor U7971 (N_7971,N_7491,N_6258);
or U7972 (N_7972,N_6292,N_6672);
xnor U7973 (N_7973,N_7136,N_6855);
and U7974 (N_7974,N_7062,N_6767);
nor U7975 (N_7975,N_7214,N_7302);
or U7976 (N_7976,N_6348,N_6844);
and U7977 (N_7977,N_7272,N_6778);
or U7978 (N_7978,N_6525,N_7151);
and U7979 (N_7979,N_6417,N_7039);
or U7980 (N_7980,N_6276,N_7057);
nor U7981 (N_7981,N_6317,N_7010);
nand U7982 (N_7982,N_6839,N_6365);
nor U7983 (N_7983,N_6960,N_6667);
and U7984 (N_7984,N_7353,N_7060);
nor U7985 (N_7985,N_6287,N_6380);
nand U7986 (N_7986,N_6553,N_6344);
and U7987 (N_7987,N_7285,N_6688);
xor U7988 (N_7988,N_7395,N_7409);
xnor U7989 (N_7989,N_7216,N_7426);
xnor U7990 (N_7990,N_6983,N_6770);
and U7991 (N_7991,N_6298,N_6376);
nor U7992 (N_7992,N_6405,N_7440);
or U7993 (N_7993,N_6753,N_6563);
nor U7994 (N_7994,N_6706,N_6385);
or U7995 (N_7995,N_7325,N_6594);
and U7996 (N_7996,N_6856,N_6731);
xnor U7997 (N_7997,N_6671,N_7159);
nand U7998 (N_7998,N_6413,N_6861);
nand U7999 (N_7999,N_7187,N_7051);
xor U8000 (N_8000,N_6254,N_6453);
nand U8001 (N_8001,N_7300,N_6681);
and U8002 (N_8002,N_7465,N_6717);
and U8003 (N_8003,N_6508,N_6947);
xnor U8004 (N_8004,N_6533,N_6783);
nand U8005 (N_8005,N_7481,N_6757);
xor U8006 (N_8006,N_6988,N_7334);
nand U8007 (N_8007,N_6333,N_6488);
and U8008 (N_8008,N_6847,N_6981);
nand U8009 (N_8009,N_6335,N_7122);
or U8010 (N_8010,N_6448,N_6475);
or U8011 (N_8011,N_6471,N_7190);
nor U8012 (N_8012,N_6881,N_7137);
xnor U8013 (N_8013,N_7284,N_7276);
and U8014 (N_8014,N_6470,N_6517);
and U8015 (N_8015,N_6713,N_6699);
nand U8016 (N_8016,N_6658,N_6845);
xnor U8017 (N_8017,N_7292,N_7470);
nor U8018 (N_8018,N_7133,N_6953);
nor U8019 (N_8019,N_6997,N_7406);
nand U8020 (N_8020,N_7282,N_6679);
nand U8021 (N_8021,N_6740,N_6701);
or U8022 (N_8022,N_6930,N_7042);
nor U8023 (N_8023,N_7287,N_6784);
and U8024 (N_8024,N_7084,N_6926);
nor U8025 (N_8025,N_7192,N_6278);
nor U8026 (N_8026,N_7157,N_7090);
nand U8027 (N_8027,N_6434,N_6922);
and U8028 (N_8028,N_6637,N_6443);
nand U8029 (N_8029,N_6871,N_7071);
or U8030 (N_8030,N_6814,N_6931);
and U8031 (N_8031,N_7086,N_7008);
and U8032 (N_8032,N_7394,N_6982);
nor U8033 (N_8033,N_7160,N_6305);
nand U8034 (N_8034,N_7184,N_7383);
or U8035 (N_8035,N_6817,N_6408);
nor U8036 (N_8036,N_6597,N_6599);
and U8037 (N_8037,N_6315,N_6283);
and U8038 (N_8038,N_7222,N_7044);
xor U8039 (N_8039,N_6318,N_6347);
and U8040 (N_8040,N_6716,N_7232);
or U8041 (N_8041,N_6584,N_6534);
nor U8042 (N_8042,N_7001,N_7139);
or U8043 (N_8043,N_7132,N_7356);
nor U8044 (N_8044,N_6819,N_6398);
nand U8045 (N_8045,N_7475,N_7252);
and U8046 (N_8046,N_7404,N_7074);
xor U8047 (N_8047,N_6500,N_7255);
nand U8048 (N_8048,N_6358,N_7244);
and U8049 (N_8049,N_7217,N_6396);
nor U8050 (N_8050,N_6959,N_7163);
nor U8051 (N_8051,N_6707,N_6741);
and U8052 (N_8052,N_7262,N_6415);
nor U8053 (N_8053,N_6841,N_7027);
nor U8054 (N_8054,N_6328,N_6512);
nand U8055 (N_8055,N_6790,N_7012);
nor U8056 (N_8056,N_6846,N_6878);
nand U8057 (N_8057,N_7326,N_6426);
and U8058 (N_8058,N_6655,N_6626);
xnor U8059 (N_8059,N_6419,N_7218);
nor U8060 (N_8060,N_6678,N_6761);
and U8061 (N_8061,N_6794,N_7110);
nand U8062 (N_8062,N_6756,N_6296);
nor U8063 (N_8063,N_6669,N_6954);
or U8064 (N_8064,N_6325,N_7312);
or U8065 (N_8065,N_7466,N_7116);
nand U8066 (N_8066,N_6843,N_7165);
nor U8067 (N_8067,N_6608,N_6933);
and U8068 (N_8068,N_7499,N_6631);
or U8069 (N_8069,N_6397,N_7193);
nand U8070 (N_8070,N_6577,N_6994);
or U8071 (N_8071,N_7100,N_6705);
nand U8072 (N_8072,N_6682,N_7135);
nor U8073 (N_8073,N_6747,N_6641);
nand U8074 (N_8074,N_6274,N_7085);
xor U8075 (N_8075,N_6401,N_7293);
xnor U8076 (N_8076,N_6644,N_6558);
nor U8077 (N_8077,N_7290,N_6693);
xor U8078 (N_8078,N_7370,N_6991);
and U8079 (N_8079,N_6338,N_6420);
nand U8080 (N_8080,N_6544,N_6392);
nand U8081 (N_8081,N_6256,N_6537);
and U8082 (N_8082,N_7493,N_7211);
or U8083 (N_8083,N_7173,N_6304);
nand U8084 (N_8084,N_7386,N_6414);
nor U8085 (N_8085,N_7094,N_7307);
or U8086 (N_8086,N_7399,N_6472);
or U8087 (N_8087,N_6963,N_7178);
xnor U8088 (N_8088,N_6806,N_6927);
and U8089 (N_8089,N_7246,N_7275);
nor U8090 (N_8090,N_6439,N_6282);
and U8091 (N_8091,N_6575,N_6564);
xnor U8092 (N_8092,N_6340,N_6494);
and U8093 (N_8093,N_6467,N_6970);
xor U8094 (N_8094,N_6490,N_6893);
or U8095 (N_8095,N_7138,N_6351);
xnor U8096 (N_8096,N_6967,N_6859);
nor U8097 (N_8097,N_6498,N_7092);
nand U8098 (N_8098,N_6645,N_6270);
or U8099 (N_8099,N_7171,N_7069);
and U8100 (N_8100,N_7225,N_6569);
or U8101 (N_8101,N_6425,N_6345);
or U8102 (N_8102,N_7407,N_7237);
nand U8103 (N_8103,N_7083,N_6764);
nor U8104 (N_8104,N_6501,N_7411);
and U8105 (N_8105,N_6590,N_6887);
nor U8106 (N_8106,N_6957,N_6829);
or U8107 (N_8107,N_6468,N_7419);
nor U8108 (N_8108,N_7026,N_7146);
or U8109 (N_8109,N_6749,N_7271);
nor U8110 (N_8110,N_6634,N_7080);
nand U8111 (N_8111,N_6750,N_7495);
and U8112 (N_8112,N_7209,N_6805);
nand U8113 (N_8113,N_6314,N_7188);
nand U8114 (N_8114,N_6884,N_6456);
and U8115 (N_8115,N_6331,N_6491);
and U8116 (N_8116,N_6321,N_6712);
or U8117 (N_8117,N_7258,N_7268);
or U8118 (N_8118,N_6336,N_7011);
xnor U8119 (N_8119,N_6370,N_7319);
and U8120 (N_8120,N_6423,N_6291);
and U8121 (N_8121,N_6990,N_6513);
nand U8122 (N_8122,N_7070,N_7073);
xnor U8123 (N_8123,N_7265,N_7141);
nor U8124 (N_8124,N_7355,N_6813);
and U8125 (N_8125,N_6750,N_6977);
nand U8126 (N_8126,N_6681,N_6290);
or U8127 (N_8127,N_7188,N_7358);
nand U8128 (N_8128,N_7141,N_7343);
nor U8129 (N_8129,N_6658,N_6575);
nand U8130 (N_8130,N_7302,N_7419);
xnor U8131 (N_8131,N_6735,N_6964);
or U8132 (N_8132,N_7420,N_6599);
and U8133 (N_8133,N_7348,N_6826);
xor U8134 (N_8134,N_6697,N_7035);
nor U8135 (N_8135,N_6633,N_6879);
nand U8136 (N_8136,N_6336,N_6803);
nor U8137 (N_8137,N_6682,N_6300);
or U8138 (N_8138,N_7371,N_7411);
nor U8139 (N_8139,N_6767,N_6984);
xnor U8140 (N_8140,N_6716,N_6593);
nand U8141 (N_8141,N_6471,N_6292);
nor U8142 (N_8142,N_6865,N_7193);
or U8143 (N_8143,N_7034,N_6647);
nor U8144 (N_8144,N_7425,N_7071);
xor U8145 (N_8145,N_7209,N_6506);
nor U8146 (N_8146,N_6674,N_7146);
and U8147 (N_8147,N_7119,N_6733);
xor U8148 (N_8148,N_6776,N_6584);
xor U8149 (N_8149,N_7174,N_7095);
nor U8150 (N_8150,N_6593,N_6725);
nor U8151 (N_8151,N_6873,N_6997);
xor U8152 (N_8152,N_7072,N_6967);
xor U8153 (N_8153,N_7272,N_7031);
nor U8154 (N_8154,N_6825,N_7049);
or U8155 (N_8155,N_7284,N_7383);
nor U8156 (N_8156,N_7173,N_6476);
or U8157 (N_8157,N_6367,N_7353);
nor U8158 (N_8158,N_6561,N_6451);
or U8159 (N_8159,N_7368,N_7207);
nor U8160 (N_8160,N_7144,N_7056);
or U8161 (N_8161,N_6829,N_7165);
and U8162 (N_8162,N_7439,N_7116);
nor U8163 (N_8163,N_6302,N_7274);
xor U8164 (N_8164,N_7277,N_7306);
and U8165 (N_8165,N_6689,N_6437);
and U8166 (N_8166,N_6318,N_6552);
nor U8167 (N_8167,N_6501,N_6638);
nor U8168 (N_8168,N_7050,N_7304);
xor U8169 (N_8169,N_7178,N_6506);
nand U8170 (N_8170,N_6995,N_7391);
nor U8171 (N_8171,N_6789,N_6270);
and U8172 (N_8172,N_7060,N_6864);
nand U8173 (N_8173,N_6576,N_6856);
or U8174 (N_8174,N_7308,N_7172);
or U8175 (N_8175,N_6629,N_7197);
xnor U8176 (N_8176,N_6524,N_6458);
or U8177 (N_8177,N_6993,N_7442);
nor U8178 (N_8178,N_7336,N_7005);
nand U8179 (N_8179,N_7376,N_7113);
nand U8180 (N_8180,N_6841,N_7151);
xnor U8181 (N_8181,N_7307,N_6811);
nand U8182 (N_8182,N_6803,N_6637);
xor U8183 (N_8183,N_6440,N_6821);
and U8184 (N_8184,N_6611,N_6522);
or U8185 (N_8185,N_6870,N_6262);
nor U8186 (N_8186,N_7275,N_6854);
and U8187 (N_8187,N_7118,N_6847);
nand U8188 (N_8188,N_6327,N_6491);
nand U8189 (N_8189,N_7250,N_6379);
nor U8190 (N_8190,N_7256,N_7094);
and U8191 (N_8191,N_6530,N_6940);
nand U8192 (N_8192,N_6905,N_6266);
and U8193 (N_8193,N_6931,N_6270);
nand U8194 (N_8194,N_7464,N_6781);
nand U8195 (N_8195,N_7411,N_7154);
nand U8196 (N_8196,N_7373,N_7147);
or U8197 (N_8197,N_6980,N_7104);
and U8198 (N_8198,N_6598,N_6392);
nor U8199 (N_8199,N_6682,N_6920);
or U8200 (N_8200,N_7386,N_7320);
nor U8201 (N_8201,N_6445,N_7093);
nand U8202 (N_8202,N_6739,N_6903);
xnor U8203 (N_8203,N_7169,N_7230);
and U8204 (N_8204,N_6976,N_6336);
nor U8205 (N_8205,N_7430,N_7297);
and U8206 (N_8206,N_7444,N_7080);
xnor U8207 (N_8207,N_7330,N_6677);
nor U8208 (N_8208,N_6881,N_6905);
and U8209 (N_8209,N_6870,N_6799);
nand U8210 (N_8210,N_7400,N_6550);
or U8211 (N_8211,N_6820,N_6358);
nor U8212 (N_8212,N_6821,N_6900);
nand U8213 (N_8213,N_6492,N_6439);
xnor U8214 (N_8214,N_6919,N_6797);
nand U8215 (N_8215,N_6969,N_7497);
xor U8216 (N_8216,N_6801,N_7260);
and U8217 (N_8217,N_6306,N_7421);
or U8218 (N_8218,N_6820,N_7457);
xnor U8219 (N_8219,N_6876,N_6821);
and U8220 (N_8220,N_6875,N_6863);
and U8221 (N_8221,N_6505,N_6450);
nor U8222 (N_8222,N_7144,N_7399);
xnor U8223 (N_8223,N_6346,N_6520);
nand U8224 (N_8224,N_6989,N_6251);
and U8225 (N_8225,N_7008,N_6472);
xor U8226 (N_8226,N_6532,N_7486);
xnor U8227 (N_8227,N_6395,N_6332);
and U8228 (N_8228,N_6898,N_7307);
nor U8229 (N_8229,N_7433,N_6462);
nor U8230 (N_8230,N_6361,N_6618);
nand U8231 (N_8231,N_7074,N_6449);
nor U8232 (N_8232,N_7394,N_7108);
xor U8233 (N_8233,N_6523,N_7139);
xor U8234 (N_8234,N_6710,N_6407);
nand U8235 (N_8235,N_7259,N_6489);
nor U8236 (N_8236,N_6271,N_6673);
xor U8237 (N_8237,N_6857,N_6280);
xor U8238 (N_8238,N_6820,N_6645);
nor U8239 (N_8239,N_7348,N_7404);
xor U8240 (N_8240,N_7085,N_6307);
nand U8241 (N_8241,N_7138,N_7285);
nand U8242 (N_8242,N_6575,N_7178);
or U8243 (N_8243,N_7040,N_6613);
xnor U8244 (N_8244,N_7497,N_7066);
xnor U8245 (N_8245,N_7007,N_7385);
xnor U8246 (N_8246,N_6625,N_6575);
nand U8247 (N_8247,N_6310,N_6500);
and U8248 (N_8248,N_7113,N_6788);
xnor U8249 (N_8249,N_7265,N_7277);
nand U8250 (N_8250,N_7242,N_7358);
or U8251 (N_8251,N_6992,N_6427);
or U8252 (N_8252,N_6609,N_7276);
and U8253 (N_8253,N_6715,N_6878);
or U8254 (N_8254,N_7359,N_6716);
nor U8255 (N_8255,N_6736,N_7028);
nor U8256 (N_8256,N_6419,N_7384);
nand U8257 (N_8257,N_7393,N_6815);
xor U8258 (N_8258,N_6581,N_7498);
or U8259 (N_8259,N_6779,N_6512);
nand U8260 (N_8260,N_6922,N_6508);
xnor U8261 (N_8261,N_6629,N_7401);
nand U8262 (N_8262,N_7465,N_6661);
nor U8263 (N_8263,N_7454,N_7032);
xnor U8264 (N_8264,N_6677,N_6864);
nand U8265 (N_8265,N_6578,N_7159);
nor U8266 (N_8266,N_7109,N_6494);
nand U8267 (N_8267,N_6631,N_6807);
nor U8268 (N_8268,N_7454,N_7305);
and U8269 (N_8269,N_6728,N_6337);
nor U8270 (N_8270,N_6669,N_6343);
nor U8271 (N_8271,N_7227,N_6594);
nand U8272 (N_8272,N_6896,N_6668);
or U8273 (N_8273,N_6831,N_7358);
or U8274 (N_8274,N_6358,N_7119);
or U8275 (N_8275,N_7168,N_6435);
or U8276 (N_8276,N_7274,N_7335);
and U8277 (N_8277,N_7051,N_6288);
and U8278 (N_8278,N_7392,N_7481);
and U8279 (N_8279,N_6514,N_6857);
and U8280 (N_8280,N_7352,N_6515);
nor U8281 (N_8281,N_7025,N_7109);
or U8282 (N_8282,N_6986,N_6868);
nand U8283 (N_8283,N_6410,N_7329);
and U8284 (N_8284,N_6973,N_6956);
xor U8285 (N_8285,N_6367,N_6814);
xnor U8286 (N_8286,N_6412,N_7377);
and U8287 (N_8287,N_7210,N_6303);
nor U8288 (N_8288,N_6588,N_6597);
nand U8289 (N_8289,N_7243,N_7326);
and U8290 (N_8290,N_7244,N_6792);
nor U8291 (N_8291,N_7153,N_7164);
or U8292 (N_8292,N_7473,N_7248);
nor U8293 (N_8293,N_7444,N_6483);
xor U8294 (N_8294,N_6752,N_6707);
nand U8295 (N_8295,N_6323,N_7390);
nor U8296 (N_8296,N_7450,N_7032);
nor U8297 (N_8297,N_6880,N_6263);
nor U8298 (N_8298,N_6587,N_6329);
nand U8299 (N_8299,N_7436,N_6414);
nand U8300 (N_8300,N_6268,N_6297);
nor U8301 (N_8301,N_7231,N_7099);
xnor U8302 (N_8302,N_7179,N_6737);
xor U8303 (N_8303,N_6347,N_6516);
nand U8304 (N_8304,N_6259,N_6479);
nand U8305 (N_8305,N_7373,N_6702);
nor U8306 (N_8306,N_7420,N_7324);
nand U8307 (N_8307,N_6706,N_6589);
and U8308 (N_8308,N_7069,N_7498);
xnor U8309 (N_8309,N_6957,N_7095);
xor U8310 (N_8310,N_6844,N_6302);
xnor U8311 (N_8311,N_7370,N_6943);
or U8312 (N_8312,N_7430,N_6961);
nand U8313 (N_8313,N_7432,N_6383);
and U8314 (N_8314,N_6408,N_7022);
and U8315 (N_8315,N_6478,N_7138);
xnor U8316 (N_8316,N_7315,N_6960);
xor U8317 (N_8317,N_6430,N_6516);
xor U8318 (N_8318,N_6257,N_6369);
xor U8319 (N_8319,N_7417,N_7463);
nor U8320 (N_8320,N_7217,N_6947);
nand U8321 (N_8321,N_6325,N_7140);
and U8322 (N_8322,N_7071,N_6449);
nand U8323 (N_8323,N_7007,N_7230);
xor U8324 (N_8324,N_7308,N_6730);
and U8325 (N_8325,N_6453,N_6560);
nand U8326 (N_8326,N_7449,N_7029);
or U8327 (N_8327,N_7304,N_7437);
or U8328 (N_8328,N_7333,N_6577);
nor U8329 (N_8329,N_6877,N_6825);
nand U8330 (N_8330,N_6324,N_6796);
or U8331 (N_8331,N_6655,N_6930);
xor U8332 (N_8332,N_6298,N_6317);
nand U8333 (N_8333,N_7108,N_7329);
nor U8334 (N_8334,N_7049,N_6269);
xor U8335 (N_8335,N_6623,N_6811);
nor U8336 (N_8336,N_7234,N_7488);
xnor U8337 (N_8337,N_6439,N_6524);
nand U8338 (N_8338,N_6563,N_6772);
and U8339 (N_8339,N_6930,N_6578);
nor U8340 (N_8340,N_7427,N_6822);
or U8341 (N_8341,N_6949,N_7013);
and U8342 (N_8342,N_6513,N_6434);
xnor U8343 (N_8343,N_6950,N_6591);
or U8344 (N_8344,N_7005,N_7087);
xor U8345 (N_8345,N_6812,N_7266);
and U8346 (N_8346,N_7123,N_6362);
nor U8347 (N_8347,N_6350,N_7023);
nand U8348 (N_8348,N_7010,N_7011);
nand U8349 (N_8349,N_6398,N_6627);
and U8350 (N_8350,N_7227,N_7082);
xnor U8351 (N_8351,N_6784,N_6319);
nand U8352 (N_8352,N_6650,N_7130);
and U8353 (N_8353,N_6971,N_6629);
nand U8354 (N_8354,N_6834,N_6806);
or U8355 (N_8355,N_6941,N_6955);
nand U8356 (N_8356,N_6254,N_6456);
nor U8357 (N_8357,N_7352,N_7261);
nand U8358 (N_8358,N_7161,N_7156);
and U8359 (N_8359,N_7335,N_7422);
xnor U8360 (N_8360,N_7056,N_6534);
and U8361 (N_8361,N_6822,N_6359);
or U8362 (N_8362,N_6266,N_6443);
nand U8363 (N_8363,N_7301,N_7223);
and U8364 (N_8364,N_6597,N_7447);
nor U8365 (N_8365,N_7106,N_6920);
nand U8366 (N_8366,N_7214,N_6771);
nand U8367 (N_8367,N_7135,N_6616);
nand U8368 (N_8368,N_6542,N_6426);
or U8369 (N_8369,N_6357,N_6964);
xor U8370 (N_8370,N_7035,N_6682);
nor U8371 (N_8371,N_6585,N_6677);
or U8372 (N_8372,N_7489,N_6747);
and U8373 (N_8373,N_6807,N_6782);
nor U8374 (N_8374,N_7485,N_6477);
or U8375 (N_8375,N_7357,N_7163);
or U8376 (N_8376,N_6339,N_6465);
xor U8377 (N_8377,N_6971,N_6561);
xnor U8378 (N_8378,N_7405,N_6931);
and U8379 (N_8379,N_7195,N_6375);
and U8380 (N_8380,N_6713,N_6811);
or U8381 (N_8381,N_6882,N_7218);
and U8382 (N_8382,N_7427,N_6556);
nand U8383 (N_8383,N_6614,N_6584);
nor U8384 (N_8384,N_6545,N_6445);
or U8385 (N_8385,N_6821,N_7185);
or U8386 (N_8386,N_7246,N_7290);
and U8387 (N_8387,N_7093,N_7218);
nand U8388 (N_8388,N_7396,N_6939);
nand U8389 (N_8389,N_6875,N_6387);
and U8390 (N_8390,N_7282,N_7086);
nor U8391 (N_8391,N_6639,N_6585);
nor U8392 (N_8392,N_7428,N_6660);
nor U8393 (N_8393,N_6823,N_6634);
xnor U8394 (N_8394,N_6780,N_7011);
and U8395 (N_8395,N_6391,N_6996);
nor U8396 (N_8396,N_6775,N_6318);
or U8397 (N_8397,N_7255,N_7429);
or U8398 (N_8398,N_6608,N_7250);
or U8399 (N_8399,N_6922,N_6782);
and U8400 (N_8400,N_7297,N_6583);
or U8401 (N_8401,N_7141,N_6560);
nand U8402 (N_8402,N_6497,N_6598);
nor U8403 (N_8403,N_7185,N_6558);
or U8404 (N_8404,N_6713,N_7171);
nor U8405 (N_8405,N_6794,N_6719);
nand U8406 (N_8406,N_7337,N_6609);
or U8407 (N_8407,N_7131,N_6482);
nor U8408 (N_8408,N_6325,N_6504);
or U8409 (N_8409,N_6983,N_7188);
nand U8410 (N_8410,N_7211,N_7127);
and U8411 (N_8411,N_7286,N_7345);
or U8412 (N_8412,N_7085,N_7472);
and U8413 (N_8413,N_6933,N_7258);
and U8414 (N_8414,N_6787,N_7485);
xor U8415 (N_8415,N_7460,N_6891);
and U8416 (N_8416,N_7115,N_6583);
or U8417 (N_8417,N_6617,N_6576);
or U8418 (N_8418,N_6465,N_7451);
nand U8419 (N_8419,N_6911,N_6487);
or U8420 (N_8420,N_6870,N_6329);
nand U8421 (N_8421,N_6351,N_7172);
nor U8422 (N_8422,N_7173,N_7442);
nor U8423 (N_8423,N_6824,N_6558);
xnor U8424 (N_8424,N_7436,N_6635);
xor U8425 (N_8425,N_6876,N_6815);
xor U8426 (N_8426,N_7449,N_6656);
and U8427 (N_8427,N_7210,N_6384);
and U8428 (N_8428,N_7320,N_6346);
nand U8429 (N_8429,N_7473,N_6320);
nand U8430 (N_8430,N_6684,N_6283);
xor U8431 (N_8431,N_7335,N_6315);
and U8432 (N_8432,N_6977,N_6645);
nand U8433 (N_8433,N_6320,N_6311);
nand U8434 (N_8434,N_7492,N_7142);
xor U8435 (N_8435,N_7439,N_6667);
xnor U8436 (N_8436,N_6250,N_6569);
or U8437 (N_8437,N_7414,N_6814);
xor U8438 (N_8438,N_6510,N_7346);
nand U8439 (N_8439,N_7099,N_6686);
and U8440 (N_8440,N_6266,N_6999);
nand U8441 (N_8441,N_6747,N_6263);
xor U8442 (N_8442,N_6672,N_6679);
xnor U8443 (N_8443,N_6400,N_6908);
nand U8444 (N_8444,N_6380,N_7142);
or U8445 (N_8445,N_6449,N_6262);
or U8446 (N_8446,N_6822,N_7372);
or U8447 (N_8447,N_7417,N_7088);
and U8448 (N_8448,N_7475,N_6918);
or U8449 (N_8449,N_7322,N_6909);
and U8450 (N_8450,N_6371,N_7088);
nor U8451 (N_8451,N_7136,N_7012);
nand U8452 (N_8452,N_6913,N_6707);
and U8453 (N_8453,N_6412,N_6906);
nand U8454 (N_8454,N_7340,N_6720);
and U8455 (N_8455,N_7478,N_7291);
or U8456 (N_8456,N_6873,N_6321);
nand U8457 (N_8457,N_7493,N_7235);
nand U8458 (N_8458,N_7305,N_6690);
nand U8459 (N_8459,N_6960,N_7489);
nor U8460 (N_8460,N_6781,N_7209);
or U8461 (N_8461,N_6966,N_6478);
nand U8462 (N_8462,N_7288,N_7443);
nand U8463 (N_8463,N_6961,N_7296);
and U8464 (N_8464,N_6585,N_6423);
nand U8465 (N_8465,N_6855,N_7215);
xor U8466 (N_8466,N_6904,N_6866);
xor U8467 (N_8467,N_7497,N_6734);
nand U8468 (N_8468,N_7259,N_6715);
nand U8469 (N_8469,N_6663,N_6288);
or U8470 (N_8470,N_6976,N_7230);
nand U8471 (N_8471,N_7271,N_7477);
and U8472 (N_8472,N_7371,N_6511);
and U8473 (N_8473,N_7352,N_7263);
xnor U8474 (N_8474,N_6354,N_6872);
and U8475 (N_8475,N_7375,N_6684);
and U8476 (N_8476,N_7342,N_7330);
xnor U8477 (N_8477,N_6483,N_7034);
nand U8478 (N_8478,N_7481,N_6678);
xnor U8479 (N_8479,N_6853,N_7160);
xnor U8480 (N_8480,N_7211,N_7015);
nand U8481 (N_8481,N_7430,N_7109);
xor U8482 (N_8482,N_6808,N_6481);
xor U8483 (N_8483,N_6459,N_7128);
nand U8484 (N_8484,N_6824,N_6332);
nand U8485 (N_8485,N_6313,N_7184);
nor U8486 (N_8486,N_6253,N_6637);
and U8487 (N_8487,N_6921,N_7193);
xnor U8488 (N_8488,N_6977,N_6354);
xor U8489 (N_8489,N_7381,N_6913);
xnor U8490 (N_8490,N_6270,N_6669);
nor U8491 (N_8491,N_7077,N_6627);
nor U8492 (N_8492,N_6482,N_6513);
xnor U8493 (N_8493,N_7276,N_6410);
xnor U8494 (N_8494,N_6282,N_7396);
nor U8495 (N_8495,N_6299,N_6370);
nor U8496 (N_8496,N_7480,N_6852);
and U8497 (N_8497,N_7016,N_6716);
xor U8498 (N_8498,N_7235,N_7096);
or U8499 (N_8499,N_6384,N_6544);
xor U8500 (N_8500,N_7180,N_6350);
or U8501 (N_8501,N_6452,N_6975);
nor U8502 (N_8502,N_6629,N_6546);
or U8503 (N_8503,N_6554,N_7295);
nor U8504 (N_8504,N_7129,N_6447);
xnor U8505 (N_8505,N_7136,N_7437);
xor U8506 (N_8506,N_6765,N_7382);
or U8507 (N_8507,N_7272,N_7394);
nand U8508 (N_8508,N_6831,N_6879);
nand U8509 (N_8509,N_7237,N_6501);
nor U8510 (N_8510,N_6596,N_6846);
and U8511 (N_8511,N_7319,N_6341);
xor U8512 (N_8512,N_6900,N_6867);
and U8513 (N_8513,N_6387,N_7182);
xnor U8514 (N_8514,N_6280,N_7433);
nand U8515 (N_8515,N_7426,N_6792);
nor U8516 (N_8516,N_7344,N_7095);
xor U8517 (N_8517,N_7438,N_7043);
and U8518 (N_8518,N_7422,N_6344);
and U8519 (N_8519,N_7254,N_6428);
and U8520 (N_8520,N_6636,N_6442);
nor U8521 (N_8521,N_7291,N_6772);
nor U8522 (N_8522,N_7333,N_6410);
or U8523 (N_8523,N_6739,N_7480);
nand U8524 (N_8524,N_6840,N_6836);
or U8525 (N_8525,N_6342,N_6429);
nand U8526 (N_8526,N_7385,N_6882);
or U8527 (N_8527,N_6611,N_6745);
and U8528 (N_8528,N_6277,N_7444);
or U8529 (N_8529,N_6452,N_6346);
or U8530 (N_8530,N_6681,N_6631);
nor U8531 (N_8531,N_7195,N_6527);
or U8532 (N_8532,N_6524,N_7245);
and U8533 (N_8533,N_6627,N_7349);
and U8534 (N_8534,N_6747,N_6969);
nand U8535 (N_8535,N_6619,N_7040);
and U8536 (N_8536,N_6645,N_6255);
and U8537 (N_8537,N_7132,N_6305);
xnor U8538 (N_8538,N_7222,N_6575);
nor U8539 (N_8539,N_7453,N_7272);
nor U8540 (N_8540,N_6636,N_6264);
xor U8541 (N_8541,N_6334,N_7084);
nor U8542 (N_8542,N_6686,N_7086);
and U8543 (N_8543,N_7405,N_7393);
nor U8544 (N_8544,N_7013,N_7192);
nand U8545 (N_8545,N_6482,N_6344);
xor U8546 (N_8546,N_7419,N_6955);
nor U8547 (N_8547,N_7287,N_7152);
nor U8548 (N_8548,N_6950,N_7047);
nor U8549 (N_8549,N_6805,N_6488);
nor U8550 (N_8550,N_6358,N_7061);
or U8551 (N_8551,N_7354,N_7424);
xor U8552 (N_8552,N_6933,N_6429);
and U8553 (N_8553,N_6720,N_6625);
nand U8554 (N_8554,N_7292,N_7119);
xnor U8555 (N_8555,N_7088,N_6624);
nand U8556 (N_8556,N_6813,N_6307);
or U8557 (N_8557,N_6710,N_6615);
or U8558 (N_8558,N_6606,N_6265);
and U8559 (N_8559,N_6871,N_6919);
nand U8560 (N_8560,N_6377,N_6375);
or U8561 (N_8561,N_7361,N_6276);
nor U8562 (N_8562,N_6520,N_6576);
and U8563 (N_8563,N_6918,N_7373);
nand U8564 (N_8564,N_6981,N_7085);
nand U8565 (N_8565,N_6261,N_6548);
xnor U8566 (N_8566,N_6480,N_6489);
xor U8567 (N_8567,N_6516,N_7069);
nand U8568 (N_8568,N_6844,N_7144);
nor U8569 (N_8569,N_7171,N_7084);
nor U8570 (N_8570,N_6570,N_7106);
nor U8571 (N_8571,N_6889,N_7147);
nor U8572 (N_8572,N_7384,N_6540);
or U8573 (N_8573,N_6291,N_6388);
nand U8574 (N_8574,N_6303,N_6430);
nand U8575 (N_8575,N_7247,N_6488);
or U8576 (N_8576,N_6776,N_6693);
and U8577 (N_8577,N_7038,N_6861);
or U8578 (N_8578,N_6432,N_6370);
or U8579 (N_8579,N_7384,N_6314);
nand U8580 (N_8580,N_6941,N_6629);
xor U8581 (N_8581,N_6627,N_6774);
and U8582 (N_8582,N_6693,N_6763);
and U8583 (N_8583,N_6843,N_6651);
nor U8584 (N_8584,N_7447,N_6846);
and U8585 (N_8585,N_7285,N_7490);
xor U8586 (N_8586,N_6662,N_7112);
or U8587 (N_8587,N_6349,N_7065);
nor U8588 (N_8588,N_7243,N_6754);
xnor U8589 (N_8589,N_6475,N_7022);
or U8590 (N_8590,N_6722,N_6922);
or U8591 (N_8591,N_7470,N_6592);
nor U8592 (N_8592,N_7067,N_6904);
xor U8593 (N_8593,N_6572,N_7167);
xnor U8594 (N_8594,N_7432,N_7185);
nor U8595 (N_8595,N_7011,N_6272);
xnor U8596 (N_8596,N_6832,N_6955);
xor U8597 (N_8597,N_7119,N_6762);
nand U8598 (N_8598,N_7162,N_7421);
or U8599 (N_8599,N_6310,N_6585);
and U8600 (N_8600,N_7242,N_6888);
xnor U8601 (N_8601,N_6543,N_7450);
or U8602 (N_8602,N_6418,N_7480);
xor U8603 (N_8603,N_6607,N_6992);
nor U8604 (N_8604,N_6410,N_7142);
or U8605 (N_8605,N_6367,N_6264);
xor U8606 (N_8606,N_7452,N_6691);
or U8607 (N_8607,N_6667,N_6959);
nor U8608 (N_8608,N_7084,N_6309);
xor U8609 (N_8609,N_7201,N_7473);
nor U8610 (N_8610,N_7405,N_6517);
and U8611 (N_8611,N_6319,N_6660);
or U8612 (N_8612,N_7461,N_7017);
or U8613 (N_8613,N_6797,N_7347);
nand U8614 (N_8614,N_6976,N_6281);
nand U8615 (N_8615,N_6782,N_7295);
and U8616 (N_8616,N_7180,N_7337);
nor U8617 (N_8617,N_6257,N_6388);
and U8618 (N_8618,N_6688,N_7010);
and U8619 (N_8619,N_7166,N_6378);
or U8620 (N_8620,N_6808,N_7427);
or U8621 (N_8621,N_7409,N_6501);
or U8622 (N_8622,N_7439,N_6845);
or U8623 (N_8623,N_6685,N_6409);
nor U8624 (N_8624,N_6482,N_6529);
nand U8625 (N_8625,N_6371,N_7060);
nor U8626 (N_8626,N_7367,N_6526);
or U8627 (N_8627,N_7201,N_7310);
xnor U8628 (N_8628,N_6336,N_6583);
or U8629 (N_8629,N_6511,N_6569);
and U8630 (N_8630,N_7436,N_7058);
and U8631 (N_8631,N_7153,N_7370);
or U8632 (N_8632,N_7480,N_7243);
nand U8633 (N_8633,N_6610,N_7173);
or U8634 (N_8634,N_6989,N_6740);
or U8635 (N_8635,N_6722,N_7080);
nand U8636 (N_8636,N_6598,N_6737);
or U8637 (N_8637,N_6833,N_6526);
nand U8638 (N_8638,N_6762,N_7443);
or U8639 (N_8639,N_7055,N_7291);
xor U8640 (N_8640,N_6757,N_6716);
nand U8641 (N_8641,N_7219,N_6594);
nor U8642 (N_8642,N_6587,N_6489);
xor U8643 (N_8643,N_7302,N_6961);
nor U8644 (N_8644,N_6729,N_6497);
or U8645 (N_8645,N_6875,N_6801);
or U8646 (N_8646,N_7453,N_6514);
xor U8647 (N_8647,N_6962,N_7145);
and U8648 (N_8648,N_6421,N_6498);
nand U8649 (N_8649,N_7442,N_6531);
and U8650 (N_8650,N_7329,N_6399);
nor U8651 (N_8651,N_6845,N_7330);
and U8652 (N_8652,N_6783,N_6558);
nand U8653 (N_8653,N_7159,N_6680);
and U8654 (N_8654,N_6635,N_7373);
and U8655 (N_8655,N_6569,N_6464);
and U8656 (N_8656,N_6826,N_7360);
xor U8657 (N_8657,N_7150,N_7030);
xnor U8658 (N_8658,N_7005,N_6794);
nand U8659 (N_8659,N_6277,N_6260);
xnor U8660 (N_8660,N_6331,N_6412);
and U8661 (N_8661,N_6630,N_6836);
nor U8662 (N_8662,N_7083,N_7220);
xor U8663 (N_8663,N_6708,N_6385);
xor U8664 (N_8664,N_6945,N_6703);
nor U8665 (N_8665,N_6710,N_6498);
nand U8666 (N_8666,N_7350,N_6827);
xnor U8667 (N_8667,N_6739,N_7031);
and U8668 (N_8668,N_7072,N_6952);
xnor U8669 (N_8669,N_6663,N_6462);
xnor U8670 (N_8670,N_6899,N_6451);
xnor U8671 (N_8671,N_6725,N_6302);
or U8672 (N_8672,N_6758,N_6778);
nand U8673 (N_8673,N_6947,N_6583);
xnor U8674 (N_8674,N_7250,N_7189);
and U8675 (N_8675,N_6284,N_6268);
nand U8676 (N_8676,N_7413,N_6469);
and U8677 (N_8677,N_6396,N_6651);
xor U8678 (N_8678,N_7312,N_6307);
and U8679 (N_8679,N_6998,N_6742);
and U8680 (N_8680,N_7186,N_6520);
xnor U8681 (N_8681,N_6664,N_6768);
nand U8682 (N_8682,N_7287,N_6309);
xnor U8683 (N_8683,N_7485,N_7237);
nand U8684 (N_8684,N_7187,N_6399);
nand U8685 (N_8685,N_7036,N_6911);
nor U8686 (N_8686,N_7164,N_6351);
nand U8687 (N_8687,N_6722,N_7226);
or U8688 (N_8688,N_7251,N_6606);
and U8689 (N_8689,N_6797,N_7255);
nor U8690 (N_8690,N_6956,N_7329);
nand U8691 (N_8691,N_6838,N_7065);
xnor U8692 (N_8692,N_7038,N_7037);
nand U8693 (N_8693,N_7059,N_7108);
nor U8694 (N_8694,N_6649,N_6403);
xor U8695 (N_8695,N_7123,N_7201);
or U8696 (N_8696,N_6488,N_6407);
nand U8697 (N_8697,N_7446,N_6709);
and U8698 (N_8698,N_7248,N_6647);
or U8699 (N_8699,N_6996,N_6900);
nor U8700 (N_8700,N_7185,N_6279);
nor U8701 (N_8701,N_6958,N_6448);
or U8702 (N_8702,N_6673,N_7460);
nor U8703 (N_8703,N_7277,N_6707);
xnor U8704 (N_8704,N_7236,N_6805);
xnor U8705 (N_8705,N_6253,N_7372);
or U8706 (N_8706,N_7133,N_7096);
xnor U8707 (N_8707,N_6918,N_6318);
nand U8708 (N_8708,N_6394,N_6930);
nand U8709 (N_8709,N_6712,N_6594);
and U8710 (N_8710,N_6707,N_6603);
nand U8711 (N_8711,N_6402,N_6644);
and U8712 (N_8712,N_6547,N_6435);
nor U8713 (N_8713,N_7181,N_6705);
and U8714 (N_8714,N_7385,N_7300);
or U8715 (N_8715,N_6285,N_6723);
nand U8716 (N_8716,N_6272,N_6973);
nor U8717 (N_8717,N_7118,N_7194);
or U8718 (N_8718,N_6315,N_7201);
and U8719 (N_8719,N_7092,N_6928);
or U8720 (N_8720,N_7437,N_7392);
xor U8721 (N_8721,N_7456,N_7068);
xor U8722 (N_8722,N_7315,N_6988);
or U8723 (N_8723,N_6704,N_6990);
and U8724 (N_8724,N_6810,N_7434);
or U8725 (N_8725,N_7183,N_6672);
and U8726 (N_8726,N_7160,N_6881);
nor U8727 (N_8727,N_6649,N_6391);
xnor U8728 (N_8728,N_7056,N_6732);
nor U8729 (N_8729,N_7106,N_6448);
or U8730 (N_8730,N_7324,N_6554);
nand U8731 (N_8731,N_6390,N_6996);
nand U8732 (N_8732,N_6948,N_6664);
and U8733 (N_8733,N_7272,N_7105);
nor U8734 (N_8734,N_7338,N_6253);
xor U8735 (N_8735,N_6410,N_6867);
nor U8736 (N_8736,N_6577,N_6953);
xnor U8737 (N_8737,N_6805,N_6495);
nand U8738 (N_8738,N_6445,N_7312);
nand U8739 (N_8739,N_6608,N_6821);
nor U8740 (N_8740,N_7026,N_7309);
or U8741 (N_8741,N_7381,N_6938);
nor U8742 (N_8742,N_6278,N_6577);
and U8743 (N_8743,N_7036,N_6470);
and U8744 (N_8744,N_7134,N_6327);
and U8745 (N_8745,N_6979,N_6915);
or U8746 (N_8746,N_6580,N_6711);
nor U8747 (N_8747,N_7461,N_6863);
nor U8748 (N_8748,N_7461,N_6569);
nor U8749 (N_8749,N_7052,N_7251);
xnor U8750 (N_8750,N_8159,N_7975);
nor U8751 (N_8751,N_7822,N_8172);
xnor U8752 (N_8752,N_8713,N_8135);
or U8753 (N_8753,N_8346,N_7512);
nor U8754 (N_8754,N_8710,N_7768);
nand U8755 (N_8755,N_7885,N_8484);
nor U8756 (N_8756,N_8513,N_7775);
or U8757 (N_8757,N_8546,N_7749);
or U8758 (N_8758,N_7525,N_8017);
or U8759 (N_8759,N_8120,N_8072);
or U8760 (N_8760,N_8586,N_8089);
or U8761 (N_8761,N_8523,N_8048);
or U8762 (N_8762,N_7794,N_8291);
nand U8763 (N_8763,N_8499,N_7659);
or U8764 (N_8764,N_8412,N_8070);
nor U8765 (N_8765,N_8243,N_8659);
nand U8766 (N_8766,N_8099,N_7691);
nand U8767 (N_8767,N_8162,N_8347);
nor U8768 (N_8768,N_8229,N_8000);
nor U8769 (N_8769,N_8724,N_8644);
nor U8770 (N_8770,N_7937,N_7529);
or U8771 (N_8771,N_7619,N_8675);
nand U8772 (N_8772,N_7579,N_8485);
or U8773 (N_8773,N_8511,N_8578);
and U8774 (N_8774,N_8080,N_7983);
and U8775 (N_8775,N_8205,N_7653);
nor U8776 (N_8776,N_8280,N_7916);
or U8777 (N_8777,N_7564,N_8394);
nand U8778 (N_8778,N_8627,N_7900);
xor U8779 (N_8779,N_7896,N_7969);
nand U8780 (N_8780,N_8401,N_8130);
or U8781 (N_8781,N_8373,N_8340);
or U8782 (N_8782,N_8518,N_8443);
nor U8783 (N_8783,N_8093,N_8730);
xnor U8784 (N_8784,N_8196,N_8605);
nand U8785 (N_8785,N_8136,N_8163);
nand U8786 (N_8786,N_7608,N_8661);
xnor U8787 (N_8787,N_8043,N_7733);
nand U8788 (N_8788,N_7607,N_8472);
or U8789 (N_8789,N_8282,N_7962);
xnor U8790 (N_8790,N_8720,N_8144);
nor U8791 (N_8791,N_7957,N_8001);
nand U8792 (N_8792,N_8180,N_7845);
xor U8793 (N_8793,N_8300,N_7755);
or U8794 (N_8794,N_7924,N_8168);
nand U8795 (N_8795,N_8193,N_8454);
nand U8796 (N_8796,N_8446,N_7816);
or U8797 (N_8797,N_7996,N_7663);
and U8798 (N_8798,N_8474,N_8557);
xor U8799 (N_8799,N_7920,N_8747);
xor U8800 (N_8800,N_8704,N_8034);
xor U8801 (N_8801,N_7696,N_7578);
or U8802 (N_8802,N_7649,N_7847);
xnor U8803 (N_8803,N_7734,N_8061);
and U8804 (N_8804,N_7912,N_7868);
xor U8805 (N_8805,N_7753,N_8363);
nand U8806 (N_8806,N_8224,N_8177);
and U8807 (N_8807,N_7621,N_8512);
and U8808 (N_8808,N_8678,N_7821);
or U8809 (N_8809,N_7859,N_8569);
nor U8810 (N_8810,N_7708,N_7567);
and U8811 (N_8811,N_7810,N_8744);
and U8812 (N_8812,N_8580,N_8515);
or U8813 (N_8813,N_8725,N_8258);
nor U8814 (N_8814,N_8077,N_8129);
xor U8815 (N_8815,N_7875,N_7940);
nand U8816 (N_8816,N_7844,N_7718);
nand U8817 (N_8817,N_8413,N_7568);
or U8818 (N_8818,N_8082,N_8425);
or U8819 (N_8819,N_8111,N_7672);
and U8820 (N_8820,N_8471,N_7577);
xnor U8821 (N_8821,N_8279,N_7848);
and U8822 (N_8822,N_8548,N_8406);
nor U8823 (N_8823,N_8619,N_7784);
and U8824 (N_8824,N_7800,N_8391);
nor U8825 (N_8825,N_8343,N_7706);
or U8826 (N_8826,N_8012,N_7640);
and U8827 (N_8827,N_8235,N_8429);
and U8828 (N_8828,N_7767,N_7692);
and U8829 (N_8829,N_8231,N_8433);
or U8830 (N_8830,N_8360,N_7552);
xor U8831 (N_8831,N_8132,N_8620);
nand U8832 (N_8832,N_7815,N_8721);
nand U8833 (N_8833,N_7772,N_8478);
or U8834 (N_8834,N_7520,N_8590);
xnor U8835 (N_8835,N_7785,N_7790);
and U8836 (N_8836,N_8101,N_7536);
and U8837 (N_8837,N_7903,N_7908);
xnor U8838 (N_8838,N_8265,N_7628);
or U8839 (N_8839,N_8648,N_7919);
and U8840 (N_8840,N_8727,N_8598);
xor U8841 (N_8841,N_7952,N_8189);
nand U8842 (N_8842,N_7732,N_8260);
and U8843 (N_8843,N_7931,N_8726);
nor U8844 (N_8844,N_8537,N_8158);
nand U8845 (N_8845,N_7562,N_8524);
nand U8846 (N_8846,N_7752,N_8284);
nor U8847 (N_8847,N_8103,N_7667);
and U8848 (N_8848,N_7994,N_7570);
nand U8849 (N_8849,N_8083,N_7933);
nor U8850 (N_8850,N_8091,N_8121);
xnor U8851 (N_8851,N_7740,N_8079);
nand U8852 (N_8852,N_8187,N_8175);
nand U8853 (N_8853,N_8161,N_7674);
xor U8854 (N_8854,N_7700,N_8044);
or U8855 (N_8855,N_8213,N_8336);
xor U8856 (N_8856,N_7850,N_8358);
or U8857 (N_8857,N_7910,N_7584);
xnor U8858 (N_8858,N_8587,N_8325);
nand U8859 (N_8859,N_8409,N_7995);
xnor U8860 (N_8860,N_8497,N_8221);
and U8861 (N_8861,N_7730,N_8050);
xor U8862 (N_8862,N_8496,N_7725);
xor U8863 (N_8863,N_7554,N_8021);
nor U8864 (N_8864,N_7647,N_8564);
nor U8865 (N_8865,N_7992,N_8475);
nand U8866 (N_8866,N_8232,N_7532);
and U8867 (N_8867,N_7863,N_8278);
and U8868 (N_8868,N_8608,N_8313);
nand U8869 (N_8869,N_8692,N_7798);
nand U8870 (N_8870,N_7825,N_8712);
and U8871 (N_8871,N_8290,N_8481);
and U8872 (N_8872,N_8319,N_7813);
xnor U8873 (N_8873,N_7958,N_8003);
nor U8874 (N_8874,N_8098,N_8669);
xor U8875 (N_8875,N_8603,N_8549);
nor U8876 (N_8876,N_7549,N_7664);
and U8877 (N_8877,N_8301,N_8310);
or U8878 (N_8878,N_8223,N_8328);
or U8879 (N_8879,N_8657,N_8124);
nor U8880 (N_8880,N_8480,N_8390);
xnor U8881 (N_8881,N_8440,N_8057);
nand U8882 (N_8882,N_8702,N_7606);
nor U8883 (N_8883,N_8560,N_7826);
or U8884 (N_8884,N_8731,N_7551);
or U8885 (N_8885,N_7820,N_8222);
and U8886 (N_8886,N_7872,N_7781);
or U8887 (N_8887,N_7698,N_8010);
xor U8888 (N_8888,N_8227,N_8027);
or U8889 (N_8889,N_8025,N_7635);
or U8890 (N_8890,N_8366,N_7571);
or U8891 (N_8891,N_8670,N_8625);
xor U8892 (N_8892,N_8385,N_8426);
and U8893 (N_8893,N_8439,N_8029);
nand U8894 (N_8894,N_8635,N_7737);
nand U8895 (N_8895,N_8249,N_8420);
nand U8896 (N_8896,N_8531,N_8684);
or U8897 (N_8897,N_8638,N_8453);
or U8898 (N_8898,N_8656,N_8115);
xor U8899 (N_8899,N_8622,N_8194);
nand U8900 (N_8900,N_8059,N_8544);
nand U8901 (N_8901,N_7693,N_7843);
nand U8902 (N_8902,N_8517,N_8428);
xor U8903 (N_8903,N_8287,N_8508);
or U8904 (N_8904,N_7811,N_7831);
or U8905 (N_8905,N_8460,N_7889);
or U8906 (N_8906,N_7757,N_8173);
or U8907 (N_8907,N_7837,N_7716);
or U8908 (N_8908,N_8152,N_7906);
nand U8909 (N_8909,N_7864,N_7651);
nor U8910 (N_8910,N_7964,N_7522);
and U8911 (N_8911,N_8673,N_7505);
nand U8912 (N_8912,N_7793,N_8672);
xnor U8913 (N_8913,N_8255,N_8149);
xnor U8914 (N_8914,N_8477,N_8397);
or U8915 (N_8915,N_7963,N_8032);
xor U8916 (N_8916,N_8049,N_7712);
and U8917 (N_8917,N_8198,N_8388);
and U8918 (N_8918,N_7892,N_7704);
xnor U8919 (N_8919,N_8634,N_8606);
and U8920 (N_8920,N_8455,N_8691);
and U8921 (N_8921,N_8253,N_7661);
nand U8922 (N_8922,N_8600,N_8112);
nor U8923 (N_8923,N_7719,N_7699);
or U8924 (N_8924,N_8631,N_8465);
nor U8925 (N_8925,N_8199,N_7928);
and U8926 (N_8926,N_7675,N_8538);
xnor U8927 (N_8927,N_8674,N_8362);
nand U8928 (N_8928,N_8005,N_8555);
or U8929 (N_8929,N_8131,N_7839);
nand U8930 (N_8930,N_7555,N_7803);
nand U8931 (N_8931,N_7759,N_8554);
xnor U8932 (N_8932,N_8090,N_8382);
nand U8933 (N_8933,N_7600,N_7987);
xnor U8934 (N_8934,N_8682,N_8601);
xor U8935 (N_8935,N_7893,N_7644);
nor U8936 (N_8936,N_8327,N_7656);
nand U8937 (N_8937,N_8410,N_8550);
nand U8938 (N_8938,N_8617,N_7846);
nand U8939 (N_8939,N_7801,N_8652);
xnor U8940 (N_8940,N_7882,N_7819);
and U8941 (N_8941,N_7531,N_8259);
nand U8942 (N_8942,N_8214,N_8685);
or U8943 (N_8943,N_8191,N_7538);
or U8944 (N_8944,N_7954,N_8654);
xor U8945 (N_8945,N_8493,N_8233);
and U8946 (N_8946,N_8246,N_8312);
and U8947 (N_8947,N_8637,N_8289);
or U8948 (N_8948,N_8256,N_8491);
and U8949 (N_8949,N_8107,N_8626);
nand U8950 (N_8950,N_8170,N_8039);
or U8951 (N_8951,N_8295,N_8540);
and U8952 (N_8952,N_7535,N_8195);
and U8953 (N_8953,N_7685,N_8505);
and U8954 (N_8954,N_8597,N_7799);
xnor U8955 (N_8955,N_7633,N_8370);
and U8956 (N_8956,N_7573,N_8140);
and U8957 (N_8957,N_7824,N_7603);
nor U8958 (N_8958,N_8054,N_8671);
nand U8959 (N_8959,N_8697,N_8357);
xor U8960 (N_8960,N_7860,N_7743);
or U8961 (N_8961,N_8060,N_7509);
nor U8962 (N_8962,N_7955,N_8324);
and U8963 (N_8963,N_8745,N_8009);
nand U8964 (N_8964,N_8589,N_7673);
xor U8965 (N_8965,N_7662,N_8404);
and U8966 (N_8966,N_8640,N_7738);
nor U8967 (N_8967,N_8658,N_7899);
nand U8968 (N_8968,N_8562,N_7714);
or U8969 (N_8969,N_8237,N_7769);
nand U8970 (N_8970,N_8040,N_7841);
or U8971 (N_8971,N_8240,N_7722);
nor U8972 (N_8972,N_7881,N_8514);
nor U8973 (N_8973,N_8575,N_8705);
nor U8974 (N_8974,N_7947,N_7973);
nor U8975 (N_8975,N_8424,N_7695);
xnor U8976 (N_8976,N_7866,N_7537);
and U8977 (N_8977,N_7516,N_7938);
nor U8978 (N_8978,N_8679,N_7823);
nand U8979 (N_8979,N_7533,N_8273);
nand U8980 (N_8980,N_7990,N_7745);
or U8981 (N_8981,N_8529,N_8616);
or U8982 (N_8982,N_8178,N_7944);
or U8983 (N_8983,N_7658,N_7741);
xnor U8984 (N_8984,N_7923,N_8206);
nor U8985 (N_8985,N_8449,N_7984);
nand U8986 (N_8986,N_7982,N_7879);
nor U8987 (N_8987,N_7681,N_8667);
or U8988 (N_8988,N_7932,N_7670);
nand U8989 (N_8989,N_7548,N_7508);
nand U8990 (N_8990,N_8242,N_8568);
nand U8991 (N_8991,N_8146,N_8094);
or U8992 (N_8992,N_7833,N_8128);
nor U8993 (N_8993,N_8160,N_7526);
nand U8994 (N_8994,N_7774,N_8086);
xor U8995 (N_8995,N_7852,N_7974);
or U8996 (N_8996,N_7678,N_8486);
xor U8997 (N_8997,N_7805,N_7540);
nand U8998 (N_8998,N_7762,N_8567);
nand U8999 (N_8999,N_8071,N_7814);
nand U9000 (N_9000,N_7626,N_8592);
and U9001 (N_9001,N_8650,N_8542);
and U9002 (N_9002,N_7773,N_8165);
nor U9003 (N_9003,N_8134,N_8105);
nor U9004 (N_9004,N_7941,N_7849);
xnor U9005 (N_9005,N_8274,N_8201);
and U9006 (N_9006,N_8607,N_8572);
xor U9007 (N_9007,N_8349,N_7746);
nor U9008 (N_9008,N_8452,N_7666);
nor U9009 (N_9009,N_7998,N_8075);
nor U9010 (N_9010,N_8041,N_8645);
nor U9011 (N_9011,N_8408,N_8078);
nand U9012 (N_9012,N_7586,N_8266);
nor U9013 (N_9013,N_8076,N_8058);
and U9014 (N_9014,N_8378,N_8148);
nor U9015 (N_9015,N_8615,N_8746);
nor U9016 (N_9016,N_8294,N_7976);
xnor U9017 (N_9017,N_8585,N_8577);
nand U9018 (N_9018,N_7542,N_8293);
or U9019 (N_9019,N_8329,N_7715);
or U9020 (N_9020,N_8104,N_8431);
or U9021 (N_9021,N_8387,N_8063);
xor U9022 (N_9022,N_7970,N_7927);
nand U9023 (N_9023,N_8488,N_8686);
and U9024 (N_9024,N_8599,N_7583);
or U9025 (N_9025,N_8226,N_8641);
nand U9026 (N_9026,N_8338,N_8383);
nand U9027 (N_9027,N_7953,N_8056);
xnor U9028 (N_9028,N_8516,N_8444);
or U9029 (N_9029,N_7575,N_8393);
and U9030 (N_9030,N_8594,N_7630);
nor U9031 (N_9031,N_8520,N_8411);
or U9032 (N_9032,N_8405,N_8367);
nor U9033 (N_9033,N_8506,N_8462);
nor U9034 (N_9034,N_8125,N_7914);
xor U9035 (N_9035,N_7668,N_7736);
nor U9036 (N_9036,N_8186,N_8212);
nand U9037 (N_9037,N_8013,N_8084);
nand U9038 (N_9038,N_8202,N_7503);
or U9039 (N_9039,N_8696,N_8595);
xnor U9040 (N_9040,N_8427,N_8498);
nand U9041 (N_9041,N_8155,N_7702);
and U9042 (N_9042,N_7853,N_7572);
and U9043 (N_9043,N_8145,N_7858);
and U9044 (N_9044,N_8016,N_8081);
nor U9045 (N_9045,N_7862,N_7750);
nand U9046 (N_9046,N_7894,N_8741);
nand U9047 (N_9047,N_8109,N_8283);
or U9048 (N_9048,N_8655,N_8613);
xor U9049 (N_9049,N_8459,N_7623);
xor U9050 (N_9050,N_8356,N_8584);
nor U9051 (N_9051,N_7887,N_7731);
and U9052 (N_9052,N_8386,N_7751);
nand U9053 (N_9053,N_7592,N_8264);
and U9054 (N_9054,N_7539,N_7545);
nand U9055 (N_9055,N_8015,N_8318);
nand U9056 (N_9056,N_7534,N_7690);
or U9057 (N_9057,N_8438,N_7840);
xor U9058 (N_9058,N_7856,N_8476);
nand U9059 (N_9059,N_8701,N_8596);
or U9060 (N_9060,N_7812,N_8419);
nand U9061 (N_9061,N_8138,N_7665);
and U9062 (N_9062,N_7748,N_8087);
nor U9063 (N_9063,N_8543,N_7588);
or U9064 (N_9064,N_8653,N_8445);
and U9065 (N_9065,N_8612,N_8552);
or U9066 (N_9066,N_8492,N_8489);
and U9067 (N_9067,N_7854,N_7817);
and U9068 (N_9068,N_8416,N_8639);
and U9069 (N_9069,N_7867,N_8395);
nand U9070 (N_9070,N_8102,N_8574);
xnor U9071 (N_9071,N_8521,N_8147);
xnor U9072 (N_9072,N_7728,N_7594);
nand U9073 (N_9073,N_8251,N_8700);
nand U9074 (N_9074,N_8528,N_8398);
nand U9075 (N_9075,N_8660,N_7569);
or U9076 (N_9076,N_8188,N_8749);
nor U9077 (N_9077,N_7574,N_7884);
nand U9078 (N_9078,N_8110,N_8354);
nand U9079 (N_9079,N_7971,N_7776);
nand U9080 (N_9080,N_8114,N_7939);
and U9081 (N_9081,N_7747,N_8096);
or U9082 (N_9082,N_8123,N_8676);
and U9083 (N_9083,N_8633,N_8630);
or U9084 (N_9084,N_8339,N_8142);
nand U9085 (N_9085,N_8407,N_7710);
nand U9086 (N_9086,N_8611,N_7641);
nor U9087 (N_9087,N_7610,N_8434);
and U9088 (N_9088,N_8345,N_8053);
and U9089 (N_9089,N_8042,N_7657);
xnor U9090 (N_9090,N_7777,N_7829);
nor U9091 (N_9091,N_8553,N_8632);
nor U9092 (N_9092,N_7717,N_7602);
nand U9093 (N_9093,N_8184,N_8547);
nor U9094 (N_9094,N_8241,N_8629);
and U9095 (N_9095,N_8267,N_8695);
xnor U9096 (N_9096,N_7861,N_7553);
and U9097 (N_9097,N_7739,N_8285);
and U9098 (N_9098,N_7550,N_8176);
nor U9099 (N_9099,N_8185,N_7720);
xor U9100 (N_9100,N_8456,N_8035);
nand U9101 (N_9101,N_8466,N_8286);
xor U9102 (N_9102,N_7988,N_8593);
nor U9103 (N_9103,N_8276,N_7558);
nand U9104 (N_9104,N_8250,N_8392);
and U9105 (N_9105,N_8618,N_8171);
nor U9106 (N_9106,N_7771,N_7842);
nor U9107 (N_9107,N_7631,N_7960);
or U9108 (N_9108,N_7625,N_7634);
or U9109 (N_9109,N_7648,N_8495);
and U9110 (N_9110,N_7729,N_7689);
or U9111 (N_9111,N_8448,N_8621);
or U9112 (N_9112,N_7787,N_8108);
xor U9113 (N_9113,N_7638,N_8361);
xor U9114 (N_9114,N_7836,N_7766);
nor U9115 (N_9115,N_8510,N_8204);
nor U9116 (N_9116,N_8422,N_7589);
nor U9117 (N_9117,N_7925,N_7513);
and U9118 (N_9118,N_7727,N_7943);
xor U9119 (N_9119,N_7783,N_7686);
nand U9120 (N_9120,N_7519,N_7599);
and U9121 (N_9121,N_7563,N_8073);
nand U9122 (N_9122,N_8450,N_8733);
xnor U9123 (N_9123,N_7597,N_8663);
nand U9124 (N_9124,N_8402,N_8308);
and U9125 (N_9125,N_7913,N_7627);
or U9126 (N_9126,N_8141,N_7950);
xnor U9127 (N_9127,N_7618,N_7643);
or U9128 (N_9128,N_8369,N_7514);
nor U9129 (N_9129,N_8297,N_7886);
or U9130 (N_9130,N_8735,N_8681);
xnor U9131 (N_9131,N_7980,N_8239);
nand U9132 (N_9132,N_7834,N_7561);
nor U9133 (N_9133,N_8646,N_8381);
or U9134 (N_9134,N_8368,N_8376);
and U9135 (N_9135,N_8351,N_7926);
nor U9136 (N_9136,N_8182,N_8739);
or U9137 (N_9137,N_8519,N_8662);
or U9138 (N_9138,N_8127,N_7612);
nand U9139 (N_9139,N_7660,N_7909);
nand U9140 (N_9140,N_7521,N_8451);
nor U9141 (N_9141,N_8270,N_8275);
and U9142 (N_9142,N_7835,N_8732);
nand U9143 (N_9143,N_8400,N_7724);
xor U9144 (N_9144,N_7547,N_8085);
or U9145 (N_9145,N_8022,N_8296);
nor U9146 (N_9146,N_7566,N_8304);
and U9147 (N_9147,N_8470,N_8689);
nand U9148 (N_9148,N_8314,N_8399);
nand U9149 (N_9149,N_7581,N_7890);
nand U9150 (N_9150,N_8716,N_7865);
nand U9151 (N_9151,N_7595,N_8403);
xnor U9152 (N_9152,N_8014,N_8316);
nor U9153 (N_9153,N_7786,N_7680);
xor U9154 (N_9154,N_8116,N_7556);
nor U9155 (N_9155,N_8271,N_8332);
xnor U9156 (N_9156,N_7679,N_8065);
or U9157 (N_9157,N_8209,N_7557);
xor U9158 (N_9158,N_8502,N_7935);
and U9159 (N_9159,N_8707,N_7929);
or U9160 (N_9160,N_8215,N_7818);
and U9161 (N_9161,N_8457,N_7742);
nand U9162 (N_9162,N_7828,N_7528);
and U9163 (N_9163,N_8467,N_8169);
or U9164 (N_9164,N_8664,N_7723);
and U9165 (N_9165,N_8217,N_8068);
xnor U9166 (N_9166,N_7855,N_8500);
nand U9167 (N_9167,N_7523,N_7620);
or U9168 (N_9168,N_7934,N_7694);
and U9169 (N_9169,N_8651,N_7809);
nor U9170 (N_9170,N_7949,N_7788);
nor U9171 (N_9171,N_8281,N_8740);
and U9172 (N_9172,N_7808,N_8069);
xor U9173 (N_9173,N_8530,N_8527);
and U9174 (N_9174,N_8683,N_7763);
or U9175 (N_9175,N_7764,N_8525);
xnor U9176 (N_9176,N_7758,N_7883);
or U9177 (N_9177,N_7898,N_8203);
xor U9178 (N_9178,N_8418,N_7873);
or U9179 (N_9179,N_7502,N_8247);
and U9180 (N_9180,N_7956,N_8210);
and U9181 (N_9181,N_8341,N_8688);
or U9182 (N_9182,N_8055,N_8570);
xnor U9183 (N_9183,N_8298,N_8153);
xnor U9184 (N_9184,N_8321,N_7922);
nand U9185 (N_9185,N_8317,N_8248);
nand U9186 (N_9186,N_8719,N_8693);
and U9187 (N_9187,N_7616,N_8736);
and U9188 (N_9188,N_7876,N_7779);
and U9189 (N_9189,N_8037,N_8483);
or U9190 (N_9190,N_7624,N_8628);
nor U9191 (N_9191,N_8556,N_7967);
and U9192 (N_9192,N_8643,N_8706);
nand U9193 (N_9193,N_8666,N_7559);
xnor U9194 (N_9194,N_8559,N_8261);
nand U9195 (N_9195,N_7650,N_8323);
or U9196 (N_9196,N_8344,N_8228);
and U9197 (N_9197,N_7942,N_7506);
or U9198 (N_9198,N_8365,N_8609);
nand U9199 (N_9199,N_7591,N_8272);
nor U9200 (N_9200,N_7684,N_8737);
nand U9201 (N_9201,N_8097,N_8353);
nor U9202 (N_9202,N_8563,N_8526);
and U9203 (N_9203,N_8117,N_7930);
or U9204 (N_9204,N_8047,N_8718);
nor U9205 (N_9205,N_7517,N_8292);
xor U9206 (N_9206,N_8441,N_7527);
or U9207 (N_9207,N_8307,N_7637);
nand U9208 (N_9208,N_7645,N_7654);
xnor U9209 (N_9209,N_7985,N_7770);
or U9210 (N_9210,N_7500,N_8019);
and U9211 (N_9211,N_7646,N_7981);
nor U9212 (N_9212,N_8415,N_8436);
or U9213 (N_9213,N_7961,N_7986);
nand U9214 (N_9214,N_7683,N_8335);
or U9215 (N_9215,N_7979,N_8118);
and U9216 (N_9216,N_7851,N_7596);
and U9217 (N_9217,N_8698,N_8469);
and U9218 (N_9218,N_8254,N_7580);
xor U9219 (N_9219,N_8558,N_8011);
and U9220 (N_9220,N_8277,N_7565);
nand U9221 (N_9221,N_8179,N_7587);
and U9222 (N_9222,N_7614,N_8352);
and U9223 (N_9223,N_8576,N_8113);
or U9224 (N_9224,N_8192,N_8610);
or U9225 (N_9225,N_8299,N_8095);
xor U9226 (N_9226,N_7632,N_8207);
nor U9227 (N_9227,N_7870,N_8151);
nand U9228 (N_9228,N_7605,N_7761);
and U9229 (N_9229,N_7518,N_8690);
nor U9230 (N_9230,N_7991,N_7501);
nor U9231 (N_9231,N_8379,N_7791);
xor U9232 (N_9232,N_8624,N_7780);
nand U9233 (N_9233,N_7891,N_7948);
and U9234 (N_9234,N_7541,N_8033);
nor U9235 (N_9235,N_8534,N_8359);
xor U9236 (N_9236,N_8614,N_7999);
nor U9237 (N_9237,N_8566,N_7936);
and U9238 (N_9238,N_8714,N_8126);
and U9239 (N_9239,N_7613,N_8330);
or U9240 (N_9240,N_8668,N_7918);
xnor U9241 (N_9241,N_8106,N_8748);
nand U9242 (N_9242,N_7687,N_8742);
and U9243 (N_9243,N_7921,N_8501);
nor U9244 (N_9244,N_8604,N_8046);
xor U9245 (N_9245,N_8156,N_7701);
or U9246 (N_9246,N_8417,N_8350);
or U9247 (N_9247,N_7601,N_8389);
or U9248 (N_9248,N_8190,N_8052);
and U9249 (N_9249,N_8699,N_7642);
or U9250 (N_9250,N_8018,N_7585);
nand U9251 (N_9251,N_8729,N_8200);
or U9252 (N_9252,N_8375,N_8377);
xnor U9253 (N_9253,N_8030,N_7792);
or U9254 (N_9254,N_7789,N_8522);
and U9255 (N_9255,N_8551,N_8636);
nand U9256 (N_9256,N_8133,N_8002);
nor U9257 (N_9257,N_8464,N_7911);
nor U9258 (N_9258,N_8708,N_7782);
nor U9259 (N_9259,N_7721,N_8545);
xor U9260 (N_9260,N_8183,N_8245);
and U9261 (N_9261,N_8583,N_8230);
and U9262 (N_9262,N_7895,N_7830);
nand U9263 (N_9263,N_8573,N_8723);
or U9264 (N_9264,N_7677,N_8649);
and U9265 (N_9265,N_7705,N_7905);
nand U9266 (N_9266,N_7726,N_8004);
and U9267 (N_9267,N_7978,N_7806);
xor U9268 (N_9268,N_8461,N_8447);
nor U9269 (N_9269,N_7966,N_7744);
or U9270 (N_9270,N_8020,N_7711);
or U9271 (N_9271,N_7946,N_7544);
or U9272 (N_9272,N_8591,N_7639);
or U9273 (N_9273,N_8220,N_7997);
xnor U9274 (N_9274,N_8565,N_8507);
xor U9275 (N_9275,N_8320,N_8579);
xnor U9276 (N_9276,N_7713,N_8051);
nor U9277 (N_9277,N_7972,N_7857);
and U9278 (N_9278,N_7907,N_8623);
nand U9279 (N_9279,N_7590,N_7807);
or U9280 (N_9280,N_7917,N_8694);
nor U9281 (N_9281,N_8588,N_8174);
nor U9282 (N_9282,N_7871,N_8571);
nor U9283 (N_9283,N_8064,N_8430);
and U9284 (N_9284,N_8432,N_7804);
or U9285 (N_9285,N_8066,N_8164);
nor U9286 (N_9286,N_7756,N_7504);
xor U9287 (N_9287,N_7671,N_8244);
nand U9288 (N_9288,N_8007,N_8026);
xor U9289 (N_9289,N_7915,N_8092);
and U9290 (N_9290,N_8561,N_8711);
nor U9291 (N_9291,N_7709,N_7965);
nor U9292 (N_9292,N_8225,N_7802);
nand U9293 (N_9293,N_7560,N_8374);
and U9294 (N_9294,N_8687,N_7832);
nand U9295 (N_9295,N_8535,N_8269);
nand U9296 (N_9296,N_8326,N_7682);
or U9297 (N_9297,N_7611,N_8468);
or U9298 (N_9298,N_8421,N_8414);
nor U9299 (N_9299,N_7993,N_8119);
nand U9300 (N_9300,N_8490,N_7707);
xnor U9301 (N_9301,N_7838,N_8435);
nand U9302 (N_9302,N_7515,N_8088);
nor U9303 (N_9303,N_8665,N_8677);
nand U9304 (N_9304,N_8197,N_8008);
xnor U9305 (N_9305,N_8306,N_8463);
nor U9306 (N_9306,N_8157,N_8582);
and U9307 (N_9307,N_8067,N_7904);
xnor U9308 (N_9308,N_8036,N_7582);
nand U9309 (N_9309,N_8581,N_7951);
nand U9310 (N_9310,N_8263,N_8334);
and U9311 (N_9311,N_8722,N_8257);
or U9312 (N_9312,N_8045,N_7507);
xnor U9313 (N_9313,N_8218,N_8074);
nor U9314 (N_9314,N_7968,N_8238);
nand U9315 (N_9315,N_7765,N_8337);
xnor U9316 (N_9316,N_8122,N_7703);
xnor U9317 (N_9317,N_8642,N_8482);
or U9318 (N_9318,N_7888,N_8311);
nor U9319 (N_9319,N_7604,N_7652);
nand U9320 (N_9320,N_8252,N_7510);
nand U9321 (N_9321,N_8536,N_7688);
nor U9322 (N_9322,N_8143,N_8167);
nand U9323 (N_9323,N_8031,N_8236);
nor U9324 (N_9324,N_8533,N_8442);
or U9325 (N_9325,N_8680,N_8532);
xnor U9326 (N_9326,N_7945,N_7897);
nor U9327 (N_9327,N_7511,N_8303);
nand U9328 (N_9328,N_8494,N_7655);
nor U9329 (N_9329,N_8038,N_8211);
nor U9330 (N_9330,N_8322,N_7669);
and U9331 (N_9331,N_8154,N_8006);
xnor U9332 (N_9332,N_8331,N_8216);
and U9333 (N_9333,N_8541,N_8743);
xor U9334 (N_9334,N_7880,N_8150);
nor U9335 (N_9335,N_8647,N_8268);
and U9336 (N_9336,N_7901,N_7629);
xnor U9337 (N_9337,N_8262,N_7827);
xnor U9338 (N_9338,N_7622,N_7760);
or U9339 (N_9339,N_7735,N_8100);
nand U9340 (N_9340,N_8166,N_8288);
xnor U9341 (N_9341,N_8715,N_7636);
xnor U9342 (N_9342,N_8539,N_8315);
nor U9343 (N_9343,N_8062,N_8028);
or U9344 (N_9344,N_8473,N_8479);
or U9345 (N_9345,N_7902,N_7977);
or U9346 (N_9346,N_8509,N_7959);
xnor U9347 (N_9347,N_8139,N_7795);
or U9348 (N_9348,N_8305,N_8348);
nor U9349 (N_9349,N_7543,N_7524);
nor U9350 (N_9350,N_7869,N_8458);
and U9351 (N_9351,N_7989,N_7796);
nor U9352 (N_9352,N_7676,N_8024);
nand U9353 (N_9353,N_7754,N_7598);
nor U9354 (N_9354,N_8396,N_8487);
or U9355 (N_9355,N_8181,N_8734);
xor U9356 (N_9356,N_8309,N_8023);
nand U9357 (N_9357,N_7874,N_8384);
or U9358 (N_9358,N_7878,N_7797);
or U9359 (N_9359,N_8504,N_8302);
nand U9360 (N_9360,N_8364,N_7530);
nand U9361 (N_9361,N_8355,N_8371);
or U9362 (N_9362,N_8137,N_7615);
nand U9363 (N_9363,N_8219,N_7617);
or U9364 (N_9364,N_8728,N_8333);
or U9365 (N_9365,N_8423,N_8437);
or U9366 (N_9366,N_8709,N_8342);
nor U9367 (N_9367,N_7609,N_8234);
or U9368 (N_9368,N_7697,N_7778);
or U9369 (N_9369,N_8503,N_8208);
or U9370 (N_9370,N_7576,N_8738);
and U9371 (N_9371,N_7593,N_8703);
or U9372 (N_9372,N_8717,N_7546);
nand U9373 (N_9373,N_8602,N_8372);
xnor U9374 (N_9374,N_8380,N_7877);
xnor U9375 (N_9375,N_7624,N_8458);
xnor U9376 (N_9376,N_8474,N_8440);
or U9377 (N_9377,N_7715,N_8091);
nand U9378 (N_9378,N_7974,N_7780);
nor U9379 (N_9379,N_7602,N_8573);
and U9380 (N_9380,N_8130,N_8673);
or U9381 (N_9381,N_8080,N_8076);
nand U9382 (N_9382,N_8394,N_8688);
xor U9383 (N_9383,N_8418,N_7962);
nor U9384 (N_9384,N_7605,N_8460);
and U9385 (N_9385,N_7598,N_8108);
and U9386 (N_9386,N_8338,N_7595);
and U9387 (N_9387,N_8267,N_8710);
or U9388 (N_9388,N_8119,N_7771);
nand U9389 (N_9389,N_8187,N_7932);
or U9390 (N_9390,N_7895,N_8627);
nand U9391 (N_9391,N_8223,N_7886);
and U9392 (N_9392,N_8100,N_8596);
or U9393 (N_9393,N_7974,N_7883);
xor U9394 (N_9394,N_7814,N_8207);
xor U9395 (N_9395,N_7537,N_8543);
and U9396 (N_9396,N_8375,N_8210);
or U9397 (N_9397,N_8419,N_8523);
xnor U9398 (N_9398,N_8472,N_7673);
nor U9399 (N_9399,N_8701,N_7582);
or U9400 (N_9400,N_7881,N_8171);
or U9401 (N_9401,N_7506,N_8112);
nand U9402 (N_9402,N_8548,N_8565);
xor U9403 (N_9403,N_7913,N_7823);
nand U9404 (N_9404,N_8121,N_7602);
nand U9405 (N_9405,N_7929,N_8003);
or U9406 (N_9406,N_8548,N_8035);
xnor U9407 (N_9407,N_8447,N_8357);
xor U9408 (N_9408,N_8015,N_8478);
xor U9409 (N_9409,N_8153,N_7717);
or U9410 (N_9410,N_7518,N_7936);
or U9411 (N_9411,N_8653,N_7581);
nor U9412 (N_9412,N_7792,N_7580);
nand U9413 (N_9413,N_7965,N_8269);
xor U9414 (N_9414,N_7579,N_7500);
nor U9415 (N_9415,N_7821,N_8579);
or U9416 (N_9416,N_7657,N_8396);
nor U9417 (N_9417,N_7718,N_7815);
or U9418 (N_9418,N_8304,N_7996);
or U9419 (N_9419,N_7788,N_7827);
xnor U9420 (N_9420,N_8403,N_8034);
nor U9421 (N_9421,N_8099,N_8166);
nand U9422 (N_9422,N_7811,N_8388);
nor U9423 (N_9423,N_7521,N_8394);
or U9424 (N_9424,N_7944,N_8105);
nor U9425 (N_9425,N_8685,N_7816);
nand U9426 (N_9426,N_8599,N_8406);
and U9427 (N_9427,N_8489,N_7721);
xnor U9428 (N_9428,N_7931,N_8592);
nand U9429 (N_9429,N_8362,N_8115);
nand U9430 (N_9430,N_8401,N_8491);
or U9431 (N_9431,N_7517,N_7706);
xnor U9432 (N_9432,N_8065,N_8429);
and U9433 (N_9433,N_7844,N_8664);
nor U9434 (N_9434,N_7535,N_8120);
and U9435 (N_9435,N_7764,N_8322);
and U9436 (N_9436,N_7630,N_8243);
xnor U9437 (N_9437,N_7548,N_8236);
nor U9438 (N_9438,N_7810,N_8028);
or U9439 (N_9439,N_8264,N_8081);
and U9440 (N_9440,N_7583,N_8051);
xnor U9441 (N_9441,N_8296,N_8671);
or U9442 (N_9442,N_8463,N_7694);
nand U9443 (N_9443,N_8279,N_7987);
xnor U9444 (N_9444,N_8417,N_8147);
nor U9445 (N_9445,N_8180,N_8605);
nand U9446 (N_9446,N_8540,N_7626);
nor U9447 (N_9447,N_8568,N_7640);
nor U9448 (N_9448,N_7581,N_8664);
and U9449 (N_9449,N_8350,N_8493);
and U9450 (N_9450,N_8133,N_7675);
and U9451 (N_9451,N_7542,N_8028);
and U9452 (N_9452,N_8249,N_8214);
xor U9453 (N_9453,N_7778,N_7501);
nand U9454 (N_9454,N_7710,N_8741);
and U9455 (N_9455,N_8456,N_8222);
nand U9456 (N_9456,N_8479,N_8239);
xor U9457 (N_9457,N_7872,N_8206);
nor U9458 (N_9458,N_8376,N_8221);
or U9459 (N_9459,N_8214,N_7923);
nor U9460 (N_9460,N_8530,N_8208);
or U9461 (N_9461,N_7629,N_8485);
nor U9462 (N_9462,N_8309,N_8282);
nor U9463 (N_9463,N_7662,N_8437);
and U9464 (N_9464,N_8684,N_8231);
nand U9465 (N_9465,N_8172,N_8748);
xor U9466 (N_9466,N_7618,N_8687);
nand U9467 (N_9467,N_8413,N_8281);
nor U9468 (N_9468,N_8204,N_8749);
xor U9469 (N_9469,N_8299,N_7731);
xor U9470 (N_9470,N_7686,N_8117);
nor U9471 (N_9471,N_7840,N_8079);
xor U9472 (N_9472,N_8288,N_7516);
or U9473 (N_9473,N_7672,N_8191);
xor U9474 (N_9474,N_8644,N_7867);
xnor U9475 (N_9475,N_8582,N_7891);
and U9476 (N_9476,N_8744,N_8292);
and U9477 (N_9477,N_8105,N_8171);
or U9478 (N_9478,N_7640,N_8252);
nor U9479 (N_9479,N_7641,N_8535);
xor U9480 (N_9480,N_7546,N_7614);
and U9481 (N_9481,N_7864,N_8725);
nand U9482 (N_9482,N_8299,N_8028);
or U9483 (N_9483,N_8043,N_8520);
nor U9484 (N_9484,N_8063,N_7694);
or U9485 (N_9485,N_7525,N_7945);
nand U9486 (N_9486,N_7892,N_8478);
and U9487 (N_9487,N_8293,N_7724);
xor U9488 (N_9488,N_8530,N_7653);
or U9489 (N_9489,N_7678,N_8033);
nor U9490 (N_9490,N_8353,N_8016);
and U9491 (N_9491,N_7934,N_7740);
nand U9492 (N_9492,N_8114,N_8470);
or U9493 (N_9493,N_8555,N_8747);
or U9494 (N_9494,N_8562,N_8421);
and U9495 (N_9495,N_7952,N_7568);
or U9496 (N_9496,N_8542,N_8366);
xor U9497 (N_9497,N_7920,N_8173);
xnor U9498 (N_9498,N_8514,N_8535);
and U9499 (N_9499,N_8097,N_7754);
and U9500 (N_9500,N_8435,N_8054);
or U9501 (N_9501,N_8334,N_8364);
or U9502 (N_9502,N_7756,N_8591);
nand U9503 (N_9503,N_7830,N_8694);
nand U9504 (N_9504,N_8077,N_7612);
nor U9505 (N_9505,N_8408,N_7925);
nand U9506 (N_9506,N_7973,N_8350);
xnor U9507 (N_9507,N_8071,N_8175);
nor U9508 (N_9508,N_8168,N_7908);
nor U9509 (N_9509,N_8425,N_7521);
and U9510 (N_9510,N_7922,N_8355);
nand U9511 (N_9511,N_8679,N_8646);
and U9512 (N_9512,N_7519,N_8202);
nor U9513 (N_9513,N_8484,N_7689);
nand U9514 (N_9514,N_7775,N_8558);
or U9515 (N_9515,N_8353,N_8049);
and U9516 (N_9516,N_7580,N_8634);
and U9517 (N_9517,N_7572,N_8103);
or U9518 (N_9518,N_8260,N_7695);
and U9519 (N_9519,N_8584,N_7508);
nand U9520 (N_9520,N_7580,N_8079);
nand U9521 (N_9521,N_7991,N_7734);
or U9522 (N_9522,N_7890,N_8341);
nand U9523 (N_9523,N_8458,N_8068);
xor U9524 (N_9524,N_8272,N_8385);
and U9525 (N_9525,N_7866,N_8608);
xnor U9526 (N_9526,N_7560,N_7825);
xor U9527 (N_9527,N_8056,N_7505);
or U9528 (N_9528,N_7750,N_7937);
xor U9529 (N_9529,N_7556,N_8376);
xor U9530 (N_9530,N_8329,N_8157);
xor U9531 (N_9531,N_7703,N_7514);
xnor U9532 (N_9532,N_7625,N_8705);
nand U9533 (N_9533,N_8640,N_8080);
xor U9534 (N_9534,N_8349,N_7868);
nor U9535 (N_9535,N_8097,N_7576);
xor U9536 (N_9536,N_8690,N_7993);
xor U9537 (N_9537,N_8411,N_8328);
nand U9538 (N_9538,N_7870,N_8527);
nand U9539 (N_9539,N_8361,N_8337);
nand U9540 (N_9540,N_7557,N_8476);
nand U9541 (N_9541,N_7884,N_7630);
and U9542 (N_9542,N_8224,N_8569);
nor U9543 (N_9543,N_8008,N_8176);
and U9544 (N_9544,N_7788,N_8514);
xnor U9545 (N_9545,N_8473,N_8356);
xor U9546 (N_9546,N_7926,N_8678);
nor U9547 (N_9547,N_7586,N_8193);
and U9548 (N_9548,N_8149,N_7583);
nor U9549 (N_9549,N_8166,N_7856);
or U9550 (N_9550,N_7588,N_8518);
nand U9551 (N_9551,N_7932,N_8324);
or U9552 (N_9552,N_7826,N_8027);
xnor U9553 (N_9553,N_8064,N_8168);
xnor U9554 (N_9554,N_7900,N_8597);
nor U9555 (N_9555,N_8264,N_7841);
and U9556 (N_9556,N_7592,N_8460);
and U9557 (N_9557,N_8616,N_7772);
and U9558 (N_9558,N_7809,N_8674);
nor U9559 (N_9559,N_8492,N_8532);
and U9560 (N_9560,N_8390,N_7547);
nand U9561 (N_9561,N_8366,N_7926);
and U9562 (N_9562,N_8026,N_8323);
nand U9563 (N_9563,N_8141,N_8169);
or U9564 (N_9564,N_8222,N_7927);
nor U9565 (N_9565,N_7635,N_8512);
nand U9566 (N_9566,N_8681,N_7672);
xor U9567 (N_9567,N_7527,N_8004);
nand U9568 (N_9568,N_7829,N_8564);
xor U9569 (N_9569,N_8198,N_8121);
nor U9570 (N_9570,N_8028,N_7632);
xor U9571 (N_9571,N_8518,N_8458);
xor U9572 (N_9572,N_8174,N_8525);
or U9573 (N_9573,N_7821,N_7800);
nor U9574 (N_9574,N_8389,N_8193);
nand U9575 (N_9575,N_8625,N_8421);
and U9576 (N_9576,N_8495,N_7791);
xnor U9577 (N_9577,N_7525,N_7811);
and U9578 (N_9578,N_7974,N_7674);
xnor U9579 (N_9579,N_7601,N_8395);
nand U9580 (N_9580,N_8240,N_7535);
and U9581 (N_9581,N_8428,N_7563);
xor U9582 (N_9582,N_8443,N_8140);
or U9583 (N_9583,N_8533,N_7500);
or U9584 (N_9584,N_8399,N_7963);
xnor U9585 (N_9585,N_8015,N_7820);
nand U9586 (N_9586,N_8516,N_8040);
nor U9587 (N_9587,N_7772,N_7759);
or U9588 (N_9588,N_8674,N_8523);
and U9589 (N_9589,N_8309,N_8598);
and U9590 (N_9590,N_8679,N_8642);
xor U9591 (N_9591,N_8711,N_7681);
nor U9592 (N_9592,N_7822,N_8517);
and U9593 (N_9593,N_8376,N_8452);
and U9594 (N_9594,N_8263,N_8099);
xnor U9595 (N_9595,N_8672,N_7606);
nand U9596 (N_9596,N_7854,N_7997);
nor U9597 (N_9597,N_8271,N_8214);
and U9598 (N_9598,N_8296,N_8535);
and U9599 (N_9599,N_8035,N_7559);
xor U9600 (N_9600,N_7560,N_8062);
and U9601 (N_9601,N_7904,N_8268);
nor U9602 (N_9602,N_8250,N_7837);
xnor U9603 (N_9603,N_7925,N_7667);
and U9604 (N_9604,N_8303,N_7813);
nand U9605 (N_9605,N_8522,N_8662);
xnor U9606 (N_9606,N_7981,N_8280);
nor U9607 (N_9607,N_7913,N_8279);
xnor U9608 (N_9608,N_8708,N_8475);
and U9609 (N_9609,N_7647,N_7700);
and U9610 (N_9610,N_8570,N_8698);
nand U9611 (N_9611,N_8218,N_8379);
and U9612 (N_9612,N_8277,N_8428);
and U9613 (N_9613,N_7591,N_8538);
nor U9614 (N_9614,N_7522,N_8370);
nor U9615 (N_9615,N_7880,N_8179);
and U9616 (N_9616,N_7647,N_7698);
nor U9617 (N_9617,N_8671,N_8599);
and U9618 (N_9618,N_8633,N_8020);
nor U9619 (N_9619,N_7714,N_7509);
or U9620 (N_9620,N_7788,N_8584);
nor U9621 (N_9621,N_8148,N_8406);
or U9622 (N_9622,N_8269,N_7635);
nand U9623 (N_9623,N_7878,N_8147);
nand U9624 (N_9624,N_7606,N_7897);
or U9625 (N_9625,N_7923,N_8743);
nand U9626 (N_9626,N_7861,N_7739);
nand U9627 (N_9627,N_8534,N_7907);
nor U9628 (N_9628,N_8415,N_8510);
or U9629 (N_9629,N_8577,N_8730);
nand U9630 (N_9630,N_7789,N_7604);
and U9631 (N_9631,N_8039,N_8251);
and U9632 (N_9632,N_8652,N_7579);
or U9633 (N_9633,N_7887,N_8730);
xnor U9634 (N_9634,N_8564,N_7788);
or U9635 (N_9635,N_8152,N_8616);
xnor U9636 (N_9636,N_7723,N_7610);
nand U9637 (N_9637,N_8370,N_7906);
xor U9638 (N_9638,N_7666,N_8396);
nor U9639 (N_9639,N_8067,N_8103);
xnor U9640 (N_9640,N_7731,N_8443);
nand U9641 (N_9641,N_8721,N_7977);
nor U9642 (N_9642,N_8069,N_7997);
xnor U9643 (N_9643,N_8656,N_7928);
or U9644 (N_9644,N_8682,N_7663);
and U9645 (N_9645,N_8557,N_8362);
xor U9646 (N_9646,N_7829,N_7736);
nor U9647 (N_9647,N_8214,N_7742);
and U9648 (N_9648,N_8484,N_7818);
and U9649 (N_9649,N_8629,N_7814);
nor U9650 (N_9650,N_7867,N_8176);
and U9651 (N_9651,N_7639,N_7643);
nor U9652 (N_9652,N_8090,N_8560);
or U9653 (N_9653,N_7877,N_8349);
or U9654 (N_9654,N_8640,N_7889);
nand U9655 (N_9655,N_8196,N_8208);
nor U9656 (N_9656,N_7530,N_7937);
and U9657 (N_9657,N_7931,N_8348);
and U9658 (N_9658,N_8583,N_8075);
xnor U9659 (N_9659,N_8169,N_8550);
xnor U9660 (N_9660,N_7854,N_7781);
or U9661 (N_9661,N_8217,N_7811);
and U9662 (N_9662,N_7551,N_7877);
or U9663 (N_9663,N_7635,N_7977);
xnor U9664 (N_9664,N_8614,N_7515);
and U9665 (N_9665,N_8592,N_8732);
and U9666 (N_9666,N_8603,N_8258);
and U9667 (N_9667,N_8140,N_8444);
nand U9668 (N_9668,N_7904,N_8525);
nor U9669 (N_9669,N_8216,N_8603);
xor U9670 (N_9670,N_7798,N_8348);
nand U9671 (N_9671,N_7648,N_7547);
and U9672 (N_9672,N_8223,N_7547);
nor U9673 (N_9673,N_8242,N_8271);
nor U9674 (N_9674,N_8017,N_8292);
and U9675 (N_9675,N_8206,N_8545);
xnor U9676 (N_9676,N_8030,N_7655);
nand U9677 (N_9677,N_8256,N_8218);
nand U9678 (N_9678,N_8608,N_7775);
xnor U9679 (N_9679,N_7558,N_8076);
nand U9680 (N_9680,N_8410,N_7829);
or U9681 (N_9681,N_7950,N_8429);
nor U9682 (N_9682,N_8464,N_8546);
nand U9683 (N_9683,N_7564,N_7936);
xnor U9684 (N_9684,N_7972,N_8235);
nand U9685 (N_9685,N_8054,N_8470);
xor U9686 (N_9686,N_8587,N_7794);
nor U9687 (N_9687,N_7654,N_7855);
and U9688 (N_9688,N_7856,N_7945);
nand U9689 (N_9689,N_8631,N_8404);
or U9690 (N_9690,N_7903,N_7798);
and U9691 (N_9691,N_7658,N_7566);
nand U9692 (N_9692,N_7652,N_8065);
or U9693 (N_9693,N_7698,N_8526);
and U9694 (N_9694,N_7941,N_8636);
nand U9695 (N_9695,N_7635,N_8681);
and U9696 (N_9696,N_8364,N_8077);
or U9697 (N_9697,N_8338,N_8255);
xor U9698 (N_9698,N_7859,N_7593);
xor U9699 (N_9699,N_8448,N_7627);
or U9700 (N_9700,N_7839,N_8045);
or U9701 (N_9701,N_8226,N_8353);
or U9702 (N_9702,N_7727,N_8718);
or U9703 (N_9703,N_7758,N_7709);
and U9704 (N_9704,N_7606,N_8588);
nand U9705 (N_9705,N_8412,N_8490);
xor U9706 (N_9706,N_8189,N_7650);
and U9707 (N_9707,N_8674,N_8130);
and U9708 (N_9708,N_8598,N_8583);
nor U9709 (N_9709,N_8397,N_7755);
and U9710 (N_9710,N_8096,N_7818);
nand U9711 (N_9711,N_7581,N_7590);
and U9712 (N_9712,N_7759,N_7577);
xor U9713 (N_9713,N_7750,N_8135);
nor U9714 (N_9714,N_8468,N_7957);
and U9715 (N_9715,N_8106,N_7818);
or U9716 (N_9716,N_8629,N_7955);
xnor U9717 (N_9717,N_7754,N_8624);
nor U9718 (N_9718,N_8670,N_7599);
and U9719 (N_9719,N_7928,N_7827);
xor U9720 (N_9720,N_7748,N_7557);
nand U9721 (N_9721,N_8198,N_8232);
and U9722 (N_9722,N_8319,N_8629);
nand U9723 (N_9723,N_7502,N_7879);
nor U9724 (N_9724,N_7532,N_8390);
xor U9725 (N_9725,N_8193,N_8692);
xor U9726 (N_9726,N_8346,N_7873);
nor U9727 (N_9727,N_7919,N_8357);
or U9728 (N_9728,N_8276,N_8202);
nand U9729 (N_9729,N_8468,N_8003);
and U9730 (N_9730,N_8745,N_7658);
xor U9731 (N_9731,N_8340,N_8370);
nor U9732 (N_9732,N_8661,N_8682);
nor U9733 (N_9733,N_7837,N_8447);
nor U9734 (N_9734,N_8398,N_7733);
xnor U9735 (N_9735,N_8484,N_8135);
nand U9736 (N_9736,N_8420,N_8727);
or U9737 (N_9737,N_7888,N_8177);
xnor U9738 (N_9738,N_8146,N_7779);
xnor U9739 (N_9739,N_7522,N_8658);
nand U9740 (N_9740,N_8252,N_8601);
nor U9741 (N_9741,N_7954,N_8120);
nand U9742 (N_9742,N_8058,N_7953);
or U9743 (N_9743,N_8650,N_7802);
nor U9744 (N_9744,N_8286,N_8665);
and U9745 (N_9745,N_8146,N_7571);
nand U9746 (N_9746,N_7943,N_8596);
nand U9747 (N_9747,N_8215,N_7925);
nor U9748 (N_9748,N_8592,N_8094);
nand U9749 (N_9749,N_8035,N_7703);
nor U9750 (N_9750,N_7514,N_8478);
nand U9751 (N_9751,N_8236,N_7621);
nand U9752 (N_9752,N_7923,N_8245);
and U9753 (N_9753,N_7739,N_8385);
or U9754 (N_9754,N_8017,N_7673);
xnor U9755 (N_9755,N_7724,N_7588);
and U9756 (N_9756,N_8180,N_8663);
nor U9757 (N_9757,N_8008,N_8672);
nand U9758 (N_9758,N_7910,N_8537);
xnor U9759 (N_9759,N_7617,N_7574);
nand U9760 (N_9760,N_8606,N_8469);
xnor U9761 (N_9761,N_7876,N_8730);
and U9762 (N_9762,N_8239,N_8147);
or U9763 (N_9763,N_8537,N_8412);
nand U9764 (N_9764,N_7777,N_7794);
xnor U9765 (N_9765,N_8148,N_7690);
xnor U9766 (N_9766,N_8132,N_8112);
or U9767 (N_9767,N_8076,N_7893);
nor U9768 (N_9768,N_7745,N_8204);
or U9769 (N_9769,N_8042,N_7893);
and U9770 (N_9770,N_8117,N_7513);
xnor U9771 (N_9771,N_8180,N_7911);
nand U9772 (N_9772,N_8141,N_8040);
xor U9773 (N_9773,N_8468,N_7616);
nand U9774 (N_9774,N_7849,N_7961);
or U9775 (N_9775,N_8705,N_8370);
xnor U9776 (N_9776,N_8680,N_8426);
nand U9777 (N_9777,N_8401,N_8037);
xor U9778 (N_9778,N_8241,N_8713);
nand U9779 (N_9779,N_8053,N_7862);
or U9780 (N_9780,N_8676,N_7798);
or U9781 (N_9781,N_8251,N_8552);
nor U9782 (N_9782,N_8742,N_7761);
nand U9783 (N_9783,N_7877,N_7752);
nor U9784 (N_9784,N_7660,N_8421);
or U9785 (N_9785,N_7840,N_8237);
nor U9786 (N_9786,N_7771,N_7745);
and U9787 (N_9787,N_7847,N_8332);
xor U9788 (N_9788,N_8104,N_8355);
nor U9789 (N_9789,N_7683,N_7720);
nor U9790 (N_9790,N_7724,N_8631);
xnor U9791 (N_9791,N_8717,N_7703);
and U9792 (N_9792,N_8496,N_8011);
xnor U9793 (N_9793,N_7748,N_7949);
nand U9794 (N_9794,N_8458,N_8425);
and U9795 (N_9795,N_7810,N_8042);
nor U9796 (N_9796,N_8489,N_7651);
and U9797 (N_9797,N_8289,N_8335);
nor U9798 (N_9798,N_8382,N_8254);
nor U9799 (N_9799,N_7649,N_8742);
nor U9800 (N_9800,N_8507,N_7507);
and U9801 (N_9801,N_8660,N_8566);
nor U9802 (N_9802,N_8556,N_8008);
and U9803 (N_9803,N_7832,N_7744);
nand U9804 (N_9804,N_8268,N_7515);
and U9805 (N_9805,N_8478,N_7707);
or U9806 (N_9806,N_8261,N_7866);
nand U9807 (N_9807,N_7512,N_8507);
nor U9808 (N_9808,N_7755,N_8518);
or U9809 (N_9809,N_8064,N_8404);
and U9810 (N_9810,N_8079,N_8347);
and U9811 (N_9811,N_7561,N_7837);
and U9812 (N_9812,N_7701,N_8258);
nor U9813 (N_9813,N_7512,N_7793);
nand U9814 (N_9814,N_7726,N_8022);
nand U9815 (N_9815,N_8044,N_8554);
xor U9816 (N_9816,N_7826,N_8227);
or U9817 (N_9817,N_7573,N_7541);
or U9818 (N_9818,N_8258,N_7622);
nor U9819 (N_9819,N_8144,N_8734);
or U9820 (N_9820,N_8258,N_8591);
xnor U9821 (N_9821,N_8568,N_8560);
nand U9822 (N_9822,N_8196,N_7629);
or U9823 (N_9823,N_8346,N_8746);
nand U9824 (N_9824,N_8461,N_7515);
or U9825 (N_9825,N_7696,N_7624);
and U9826 (N_9826,N_8561,N_7766);
nand U9827 (N_9827,N_8143,N_7668);
nand U9828 (N_9828,N_7859,N_8659);
nor U9829 (N_9829,N_8695,N_8288);
or U9830 (N_9830,N_7833,N_8511);
xor U9831 (N_9831,N_7533,N_7522);
xor U9832 (N_9832,N_7597,N_8681);
xnor U9833 (N_9833,N_8411,N_8073);
or U9834 (N_9834,N_8748,N_7525);
nand U9835 (N_9835,N_8200,N_7541);
and U9836 (N_9836,N_8309,N_8187);
nor U9837 (N_9837,N_8157,N_7856);
nor U9838 (N_9838,N_8516,N_7651);
or U9839 (N_9839,N_8721,N_7764);
or U9840 (N_9840,N_7557,N_8197);
and U9841 (N_9841,N_7720,N_7953);
or U9842 (N_9842,N_8627,N_8212);
nand U9843 (N_9843,N_7911,N_8071);
and U9844 (N_9844,N_8590,N_8401);
or U9845 (N_9845,N_8413,N_8337);
nand U9846 (N_9846,N_8661,N_7753);
and U9847 (N_9847,N_7823,N_8093);
nor U9848 (N_9848,N_7555,N_7732);
xnor U9849 (N_9849,N_7770,N_8309);
and U9850 (N_9850,N_8256,N_7854);
or U9851 (N_9851,N_7761,N_8399);
xor U9852 (N_9852,N_8573,N_8151);
nor U9853 (N_9853,N_7891,N_8558);
xnor U9854 (N_9854,N_8517,N_7899);
and U9855 (N_9855,N_8458,N_8405);
and U9856 (N_9856,N_8367,N_8369);
nor U9857 (N_9857,N_7846,N_8465);
xnor U9858 (N_9858,N_8276,N_7962);
xor U9859 (N_9859,N_7981,N_7760);
nor U9860 (N_9860,N_8460,N_7551);
and U9861 (N_9861,N_8522,N_8136);
and U9862 (N_9862,N_8321,N_8283);
nor U9863 (N_9863,N_8393,N_7552);
nor U9864 (N_9864,N_8172,N_7873);
xnor U9865 (N_9865,N_7971,N_8640);
and U9866 (N_9866,N_8610,N_7639);
xnor U9867 (N_9867,N_8168,N_8690);
nand U9868 (N_9868,N_7918,N_8611);
nor U9869 (N_9869,N_8140,N_8104);
xnor U9870 (N_9870,N_8344,N_8573);
xor U9871 (N_9871,N_8614,N_8587);
and U9872 (N_9872,N_7659,N_8689);
and U9873 (N_9873,N_7504,N_8466);
or U9874 (N_9874,N_8247,N_7616);
xnor U9875 (N_9875,N_8270,N_8301);
xnor U9876 (N_9876,N_8626,N_7636);
and U9877 (N_9877,N_8547,N_8041);
and U9878 (N_9878,N_7987,N_8264);
nor U9879 (N_9879,N_8373,N_7999);
nor U9880 (N_9880,N_8482,N_8582);
or U9881 (N_9881,N_7771,N_8085);
or U9882 (N_9882,N_8105,N_8013);
nor U9883 (N_9883,N_8717,N_8209);
nor U9884 (N_9884,N_8739,N_7961);
nor U9885 (N_9885,N_7940,N_8363);
nor U9886 (N_9886,N_8319,N_8548);
and U9887 (N_9887,N_8498,N_8670);
xor U9888 (N_9888,N_7539,N_8207);
nand U9889 (N_9889,N_8504,N_8231);
nor U9890 (N_9890,N_8095,N_7653);
nor U9891 (N_9891,N_8350,N_8021);
xor U9892 (N_9892,N_8254,N_7537);
nand U9893 (N_9893,N_8480,N_8549);
xnor U9894 (N_9894,N_8594,N_7906);
and U9895 (N_9895,N_8617,N_7919);
or U9896 (N_9896,N_7973,N_8102);
nor U9897 (N_9897,N_8081,N_8135);
nor U9898 (N_9898,N_7857,N_7991);
or U9899 (N_9899,N_8281,N_8213);
nor U9900 (N_9900,N_7606,N_8009);
and U9901 (N_9901,N_8517,N_7990);
nor U9902 (N_9902,N_7622,N_8074);
xor U9903 (N_9903,N_8712,N_8587);
nand U9904 (N_9904,N_7931,N_7707);
nor U9905 (N_9905,N_7692,N_8643);
and U9906 (N_9906,N_8194,N_8303);
or U9907 (N_9907,N_7984,N_7833);
nor U9908 (N_9908,N_8079,N_7645);
xnor U9909 (N_9909,N_8117,N_8628);
xnor U9910 (N_9910,N_7545,N_7988);
or U9911 (N_9911,N_8265,N_7905);
and U9912 (N_9912,N_7736,N_8105);
nand U9913 (N_9913,N_8681,N_8479);
nand U9914 (N_9914,N_7566,N_7851);
or U9915 (N_9915,N_8444,N_7563);
xor U9916 (N_9916,N_7557,N_7873);
or U9917 (N_9917,N_8612,N_7660);
xnor U9918 (N_9918,N_8735,N_7933);
nor U9919 (N_9919,N_8483,N_8269);
and U9920 (N_9920,N_7779,N_7987);
nand U9921 (N_9921,N_7755,N_7780);
or U9922 (N_9922,N_8367,N_8742);
nand U9923 (N_9923,N_7974,N_8677);
or U9924 (N_9924,N_8696,N_8706);
xnor U9925 (N_9925,N_8616,N_7726);
or U9926 (N_9926,N_7651,N_8671);
and U9927 (N_9927,N_8282,N_7750);
or U9928 (N_9928,N_8297,N_8121);
and U9929 (N_9929,N_7994,N_8190);
xnor U9930 (N_9930,N_8268,N_8164);
nor U9931 (N_9931,N_7564,N_8089);
nand U9932 (N_9932,N_8739,N_7877);
xnor U9933 (N_9933,N_8074,N_7902);
and U9934 (N_9934,N_8011,N_7506);
xnor U9935 (N_9935,N_8418,N_8375);
nor U9936 (N_9936,N_7850,N_7804);
xor U9937 (N_9937,N_8188,N_8485);
or U9938 (N_9938,N_7921,N_8353);
xor U9939 (N_9939,N_7657,N_7927);
and U9940 (N_9940,N_8075,N_8015);
nor U9941 (N_9941,N_7649,N_8523);
and U9942 (N_9942,N_8729,N_8068);
and U9943 (N_9943,N_8317,N_8065);
or U9944 (N_9944,N_7874,N_7827);
or U9945 (N_9945,N_7817,N_7850);
xnor U9946 (N_9946,N_8292,N_8443);
xnor U9947 (N_9947,N_7608,N_7605);
nand U9948 (N_9948,N_7866,N_7549);
xnor U9949 (N_9949,N_8242,N_7993);
nor U9950 (N_9950,N_7971,N_8589);
or U9951 (N_9951,N_7518,N_8110);
and U9952 (N_9952,N_8334,N_7969);
or U9953 (N_9953,N_8102,N_8359);
xor U9954 (N_9954,N_8434,N_8608);
nand U9955 (N_9955,N_8284,N_8298);
nor U9956 (N_9956,N_7915,N_8417);
nand U9957 (N_9957,N_7969,N_7817);
and U9958 (N_9958,N_8404,N_8395);
nand U9959 (N_9959,N_7707,N_8336);
xnor U9960 (N_9960,N_8281,N_7910);
and U9961 (N_9961,N_7832,N_8305);
xor U9962 (N_9962,N_8264,N_8705);
and U9963 (N_9963,N_8326,N_8616);
nand U9964 (N_9964,N_8739,N_7704);
and U9965 (N_9965,N_8003,N_8263);
nand U9966 (N_9966,N_7965,N_7881);
or U9967 (N_9967,N_7729,N_7795);
or U9968 (N_9968,N_7732,N_8596);
or U9969 (N_9969,N_7521,N_8159);
nand U9970 (N_9970,N_7848,N_8048);
nand U9971 (N_9971,N_7857,N_8211);
or U9972 (N_9972,N_8677,N_8651);
nor U9973 (N_9973,N_8047,N_8123);
nand U9974 (N_9974,N_8707,N_7825);
xnor U9975 (N_9975,N_7926,N_8208);
nand U9976 (N_9976,N_8341,N_7986);
nand U9977 (N_9977,N_8707,N_8185);
nand U9978 (N_9978,N_7665,N_7772);
nor U9979 (N_9979,N_7650,N_8311);
nand U9980 (N_9980,N_8701,N_8246);
or U9981 (N_9981,N_7721,N_7529);
nor U9982 (N_9982,N_8408,N_7664);
nor U9983 (N_9983,N_7764,N_7725);
nand U9984 (N_9984,N_8710,N_7782);
and U9985 (N_9985,N_8089,N_8387);
or U9986 (N_9986,N_7803,N_7643);
nor U9987 (N_9987,N_7549,N_8587);
and U9988 (N_9988,N_7600,N_8261);
and U9989 (N_9989,N_8525,N_7594);
and U9990 (N_9990,N_8398,N_7763);
xor U9991 (N_9991,N_7775,N_8682);
and U9992 (N_9992,N_7899,N_7847);
nand U9993 (N_9993,N_7865,N_8337);
or U9994 (N_9994,N_8084,N_8261);
nor U9995 (N_9995,N_7711,N_7710);
xnor U9996 (N_9996,N_8178,N_8484);
or U9997 (N_9997,N_7806,N_7817);
or U9998 (N_9998,N_8014,N_8001);
or U9999 (N_9999,N_8736,N_7656);
nand U10000 (N_10000,N_9377,N_9600);
nor U10001 (N_10001,N_9538,N_9098);
xor U10002 (N_10002,N_9728,N_9283);
and U10003 (N_10003,N_9925,N_9213);
xor U10004 (N_10004,N_9083,N_9466);
nor U10005 (N_10005,N_9504,N_8753);
and U10006 (N_10006,N_8860,N_9240);
and U10007 (N_10007,N_9481,N_9618);
or U10008 (N_10008,N_9069,N_9609);
xor U10009 (N_10009,N_9947,N_9631);
nand U10010 (N_10010,N_9917,N_9766);
or U10011 (N_10011,N_8849,N_9977);
xnor U10012 (N_10012,N_9445,N_9454);
nor U10013 (N_10013,N_8985,N_9603);
nand U10014 (N_10014,N_9404,N_9782);
nand U10015 (N_10015,N_9997,N_9918);
nand U10016 (N_10016,N_9934,N_9847);
nor U10017 (N_10017,N_8905,N_9510);
nand U10018 (N_10018,N_9543,N_9251);
and U10019 (N_10019,N_9806,N_9294);
xnor U10020 (N_10020,N_9812,N_8879);
or U10021 (N_10021,N_9329,N_9598);
xnor U10022 (N_10022,N_8940,N_9551);
nand U10023 (N_10023,N_9559,N_9172);
or U10024 (N_10024,N_9372,N_9010);
and U10025 (N_10025,N_8809,N_9170);
or U10026 (N_10026,N_9828,N_9760);
xor U10027 (N_10027,N_9422,N_9493);
xnor U10028 (N_10028,N_8930,N_9699);
nor U10029 (N_10029,N_9721,N_9672);
xor U10030 (N_10030,N_9502,N_9696);
or U10031 (N_10031,N_9425,N_9656);
and U10032 (N_10032,N_9430,N_9688);
or U10033 (N_10033,N_9558,N_9000);
nor U10034 (N_10034,N_9421,N_9714);
xnor U10035 (N_10035,N_9756,N_9767);
or U10036 (N_10036,N_9755,N_9439);
nor U10037 (N_10037,N_9307,N_9028);
and U10038 (N_10038,N_9886,N_8955);
xnor U10039 (N_10039,N_8865,N_9608);
or U10040 (N_10040,N_9096,N_9063);
xor U10041 (N_10041,N_9991,N_9239);
or U10042 (N_10042,N_9770,N_9254);
nor U10043 (N_10043,N_9219,N_9505);
xor U10044 (N_10044,N_8855,N_8901);
xnor U10045 (N_10045,N_9520,N_8772);
and U10046 (N_10046,N_9476,N_9854);
or U10047 (N_10047,N_9852,N_9084);
nor U10048 (N_10048,N_9380,N_9450);
nand U10049 (N_10049,N_8911,N_9326);
nand U10050 (N_10050,N_9796,N_9956);
and U10051 (N_10051,N_8981,N_9513);
and U10052 (N_10052,N_9318,N_9964);
or U10053 (N_10053,N_9826,N_9047);
nor U10054 (N_10054,N_9230,N_9507);
xnor U10055 (N_10055,N_8818,N_9641);
nand U10056 (N_10056,N_8993,N_9491);
nor U10057 (N_10057,N_8792,N_8874);
and U10058 (N_10058,N_9786,N_9601);
nor U10059 (N_10059,N_8757,N_9483);
nor U10060 (N_10060,N_8899,N_9410);
and U10061 (N_10061,N_8800,N_9521);
or U10062 (N_10062,N_8776,N_9857);
or U10063 (N_10063,N_9301,N_9071);
or U10064 (N_10064,N_9980,N_9815);
nor U10065 (N_10065,N_9398,N_9655);
xor U10066 (N_10066,N_9257,N_9075);
nor U10067 (N_10067,N_8934,N_9133);
or U10068 (N_10068,N_9942,N_9720);
nand U10069 (N_10069,N_9193,N_9937);
nand U10070 (N_10070,N_9892,N_8821);
nor U10071 (N_10071,N_9807,N_9820);
and U10072 (N_10072,N_9628,N_9617);
nor U10073 (N_10073,N_9958,N_9021);
nor U10074 (N_10074,N_9652,N_9646);
nor U10075 (N_10075,N_9431,N_9757);
nor U10076 (N_10076,N_9785,N_9031);
xnor U10077 (N_10077,N_9516,N_9356);
nor U10078 (N_10078,N_9435,N_9580);
xor U10079 (N_10079,N_8906,N_9588);
and U10080 (N_10080,N_8867,N_9223);
nand U10081 (N_10081,N_9933,N_9064);
nor U10082 (N_10082,N_9341,N_9006);
nor U10083 (N_10083,N_9761,N_8803);
nand U10084 (N_10084,N_9969,N_9582);
xor U10085 (N_10085,N_9461,N_8890);
xnor U10086 (N_10086,N_9371,N_8963);
or U10087 (N_10087,N_9141,N_9186);
nand U10088 (N_10088,N_8972,N_9633);
nor U10089 (N_10089,N_9774,N_9823);
xor U10090 (N_10090,N_9025,N_9358);
xor U10091 (N_10091,N_9040,N_9190);
nor U10092 (N_10092,N_9152,N_9490);
or U10093 (N_10093,N_9988,N_8882);
and U10094 (N_10094,N_9469,N_9634);
xor U10095 (N_10095,N_8765,N_9577);
nand U10096 (N_10096,N_9710,N_9973);
xor U10097 (N_10097,N_9198,N_8789);
nor U10098 (N_10098,N_8912,N_8777);
xnor U10099 (N_10099,N_8796,N_8898);
xnor U10100 (N_10100,N_8840,N_9093);
or U10101 (N_10101,N_9386,N_8866);
xnor U10102 (N_10102,N_9226,N_9471);
and U10103 (N_10103,N_8968,N_9196);
or U10104 (N_10104,N_9579,N_9821);
or U10105 (N_10105,N_8794,N_9347);
or U10106 (N_10106,N_8791,N_9967);
or U10107 (N_10107,N_9158,N_9395);
nor U10108 (N_10108,N_8990,N_9482);
and U10109 (N_10109,N_9142,N_8848);
nand U10110 (N_10110,N_9310,N_9676);
xor U10111 (N_10111,N_9108,N_8763);
or U10112 (N_10112,N_9492,N_9266);
nand U10113 (N_10113,N_9649,N_9290);
and U10114 (N_10114,N_9087,N_9355);
xor U10115 (N_10115,N_9692,N_9191);
nor U10116 (N_10116,N_8774,N_9352);
xnor U10117 (N_10117,N_9938,N_9565);
and U10118 (N_10118,N_9673,N_9053);
nor U10119 (N_10119,N_9700,N_8939);
nand U10120 (N_10120,N_9065,N_9263);
and U10121 (N_10121,N_9138,N_8945);
or U10122 (N_10122,N_9740,N_9512);
or U10123 (N_10123,N_9880,N_9725);
xnor U10124 (N_10124,N_9960,N_8769);
xor U10125 (N_10125,N_8980,N_8937);
nand U10126 (N_10126,N_8838,N_9405);
and U10127 (N_10127,N_9818,N_9667);
xnor U10128 (N_10128,N_9935,N_9836);
or U10129 (N_10129,N_9848,N_9636);
xor U10130 (N_10130,N_8870,N_9246);
xor U10131 (N_10131,N_9085,N_9549);
and U10132 (N_10132,N_9067,N_9293);
xor U10133 (N_10133,N_8761,N_9308);
xor U10134 (N_10134,N_9705,N_9914);
nand U10135 (N_10135,N_9130,N_9907);
xor U10136 (N_10136,N_8843,N_9206);
nand U10137 (N_10137,N_9550,N_8778);
nand U10138 (N_10138,N_9248,N_9055);
nor U10139 (N_10139,N_8862,N_9903);
and U10140 (N_10140,N_8891,N_9765);
nand U10141 (N_10141,N_9016,N_9954);
xnor U10142 (N_10142,N_8915,N_9204);
nand U10143 (N_10143,N_9680,N_9732);
nand U10144 (N_10144,N_9176,N_8759);
xor U10145 (N_10145,N_9607,N_8825);
or U10146 (N_10146,N_9234,N_9175);
nor U10147 (N_10147,N_9131,N_8982);
xnor U10148 (N_10148,N_9034,N_8752);
nor U10149 (N_10149,N_9181,N_8983);
and U10150 (N_10150,N_8973,N_8988);
and U10151 (N_10151,N_8847,N_9535);
nor U10152 (N_10152,N_9097,N_8986);
nand U10153 (N_10153,N_9218,N_9889);
nor U10154 (N_10154,N_9261,N_9870);
and U10155 (N_10155,N_8984,N_9153);
nor U10156 (N_10156,N_8839,N_9682);
xor U10157 (N_10157,N_9416,N_8768);
nand U10158 (N_10158,N_8815,N_9474);
xnor U10159 (N_10159,N_9208,N_9321);
xor U10160 (N_10160,N_9272,N_9477);
nand U10161 (N_10161,N_9072,N_9390);
or U10162 (N_10162,N_9173,N_8971);
xnor U10163 (N_10163,N_9136,N_9428);
xnor U10164 (N_10164,N_9424,N_9233);
and U10165 (N_10165,N_8970,N_9408);
nand U10166 (N_10166,N_9898,N_9018);
nor U10167 (N_10167,N_9165,N_8907);
nor U10168 (N_10168,N_9916,N_8767);
nand U10169 (N_10169,N_9091,N_9825);
nand U10170 (N_10170,N_9140,N_9397);
nor U10171 (N_10171,N_9999,N_9624);
or U10172 (N_10172,N_8947,N_9282);
and U10173 (N_10173,N_8927,N_8852);
nor U10174 (N_10174,N_9709,N_9645);
nand U10175 (N_10175,N_9773,N_9745);
xnor U10176 (N_10176,N_9707,N_9961);
and U10177 (N_10177,N_9941,N_9070);
or U10178 (N_10178,N_9361,N_9296);
nor U10179 (N_10179,N_8858,N_8903);
or U10180 (N_10180,N_9896,N_9210);
or U10181 (N_10181,N_9955,N_9831);
or U10182 (N_10182,N_9370,N_9434);
nor U10183 (N_10183,N_9269,N_8977);
and U10184 (N_10184,N_9503,N_9561);
xnor U10185 (N_10185,N_9320,N_9560);
or U10186 (N_10186,N_9702,N_8805);
xor U10187 (N_10187,N_9833,N_9401);
or U10188 (N_10188,N_9414,N_8959);
xor U10189 (N_10189,N_9730,N_9871);
and U10190 (N_10190,N_8808,N_9894);
nor U10191 (N_10191,N_9727,N_9129);
nand U10192 (N_10192,N_9494,N_9574);
or U10193 (N_10193,N_9719,N_9237);
xor U10194 (N_10194,N_8826,N_9703);
and U10195 (N_10195,N_8967,N_8935);
and U10196 (N_10196,N_9780,N_9027);
nor U10197 (N_10197,N_9841,N_9429);
nor U10198 (N_10198,N_9778,N_9723);
xor U10199 (N_10199,N_9548,N_9104);
nor U10200 (N_10200,N_9019,N_9332);
nor U10201 (N_10201,N_9791,N_9915);
nor U10202 (N_10202,N_9236,N_9923);
xnor U10203 (N_10203,N_9524,N_9242);
nor U10204 (N_10204,N_9529,N_9276);
xor U10205 (N_10205,N_9808,N_9241);
xnor U10206 (N_10206,N_9456,N_8975);
or U10207 (N_10207,N_9267,N_9930);
nor U10208 (N_10208,N_9333,N_9385);
xor U10209 (N_10209,N_8783,N_9351);
nand U10210 (N_10210,N_8762,N_8873);
and U10211 (N_10211,N_9389,N_8920);
and U10212 (N_10212,N_9953,N_9273);
nand U10213 (N_10213,N_9619,N_9217);
xnor U10214 (N_10214,N_8966,N_9073);
xnor U10215 (N_10215,N_9350,N_8878);
or U10216 (N_10216,N_8948,N_9575);
or U10217 (N_10217,N_8932,N_8928);
nor U10218 (N_10218,N_8964,N_9872);
xnor U10219 (N_10219,N_9748,N_9317);
and U10220 (N_10220,N_8869,N_9118);
nand U10221 (N_10221,N_9581,N_9771);
xnor U10222 (N_10222,N_9643,N_9909);
nor U10223 (N_10223,N_9527,N_8942);
or U10224 (N_10224,N_8962,N_9722);
and U10225 (N_10225,N_9620,N_9974);
and U10226 (N_10226,N_9144,N_9887);
or U10227 (N_10227,N_9354,N_9867);
or U10228 (N_10228,N_9994,N_9245);
nand U10229 (N_10229,N_8889,N_9962);
nor U10230 (N_10230,N_9982,N_9926);
and U10231 (N_10231,N_9418,N_9486);
and U10232 (N_10232,N_9384,N_8938);
and U10233 (N_10233,N_9260,N_8875);
or U10234 (N_10234,N_9216,N_9900);
or U10235 (N_10235,N_9866,N_9827);
nand U10236 (N_10236,N_9986,N_9837);
and U10237 (N_10237,N_8773,N_9675);
nand U10238 (N_10238,N_9274,N_9623);
xor U10239 (N_10239,N_9013,N_9314);
and U10240 (N_10240,N_9162,N_9455);
nor U10241 (N_10241,N_9048,N_9876);
xnor U10242 (N_10242,N_8900,N_9095);
nand U10243 (N_10243,N_8854,N_9076);
nor U10244 (N_10244,N_9570,N_9022);
xor U10245 (N_10245,N_9362,N_9465);
xnor U10246 (N_10246,N_9284,N_9920);
nand U10247 (N_10247,N_8979,N_9012);
and U10248 (N_10248,N_9768,N_9932);
and U10249 (N_10249,N_9004,N_9911);
nor U10250 (N_10250,N_9105,N_9519);
xnor U10251 (N_10251,N_9128,N_8976);
nand U10252 (N_10252,N_9840,N_9883);
nand U10253 (N_10253,N_9222,N_9984);
or U10254 (N_10254,N_8820,N_9100);
nor U10255 (N_10255,N_9050,N_9612);
or U10256 (N_10256,N_9146,N_9192);
xnor U10257 (N_10257,N_8782,N_9079);
xnor U10258 (N_10258,N_9211,N_9297);
xor U10259 (N_10259,N_9302,N_8965);
nor U10260 (N_10260,N_9739,N_9102);
or U10261 (N_10261,N_8958,N_9717);
or U10262 (N_10262,N_9875,N_9487);
and U10263 (N_10263,N_9992,N_8892);
nand U10264 (N_10264,N_9289,N_8833);
and U10265 (N_10265,N_9346,N_9790);
xor U10266 (N_10266,N_9082,N_9987);
xor U10267 (N_10267,N_9971,N_9413);
nand U10268 (N_10268,N_9342,N_9891);
xnor U10269 (N_10269,N_9605,N_8813);
nor U10270 (N_10270,N_9794,N_9194);
and U10271 (N_10271,N_8797,N_9674);
and U10272 (N_10272,N_8841,N_9859);
nand U10273 (N_10273,N_9446,N_9023);
and U10274 (N_10274,N_9906,N_8861);
and U10275 (N_10275,N_9749,N_9850);
nor U10276 (N_10276,N_9295,N_9968);
xor U10277 (N_10277,N_8863,N_8908);
xor U10278 (N_10278,N_9375,N_8832);
or U10279 (N_10279,N_9694,N_9929);
or U10280 (N_10280,N_8775,N_9275);
xnor U10281 (N_10281,N_8851,N_9981);
nand U10282 (N_10282,N_9174,N_9473);
xnor U10283 (N_10283,N_9374,N_9978);
nand U10284 (N_10284,N_9051,N_9331);
xor U10285 (N_10285,N_9737,N_8836);
and U10286 (N_10286,N_9957,N_8888);
nor U10287 (N_10287,N_9697,N_8902);
xnor U10288 (N_10288,N_9156,N_9411);
or U10289 (N_10289,N_9406,N_8956);
nor U10290 (N_10290,N_8853,N_9830);
nor U10291 (N_10291,N_9555,N_9863);
and U10292 (N_10292,N_9684,N_8929);
xnor U10293 (N_10293,N_9017,N_9689);
nand U10294 (N_10294,N_9713,N_9014);
xor U10295 (N_10295,N_9400,N_8894);
and U10296 (N_10296,N_9637,N_9563);
nor U10297 (N_10297,N_9243,N_9526);
and U10298 (N_10298,N_9249,N_9642);
nand U10299 (N_10299,N_9160,N_9062);
and U10300 (N_10300,N_9244,N_9921);
or U10301 (N_10301,N_9393,N_9412);
nor U10302 (N_10302,N_8916,N_9734);
nor U10303 (N_10303,N_9387,N_9793);
nor U10304 (N_10304,N_9166,N_9449);
and U10305 (N_10305,N_9338,N_8999);
xnor U10306 (N_10306,N_8790,N_9811);
nor U10307 (N_10307,N_9495,N_9865);
and U10308 (N_10308,N_9795,N_8857);
nor U10309 (N_10309,N_9458,N_9799);
nand U10310 (N_10310,N_8949,N_9077);
nor U10311 (N_10311,N_9797,N_9029);
nor U10312 (N_10312,N_9678,N_9666);
xnor U10313 (N_10313,N_9661,N_9724);
nor U10314 (N_10314,N_8953,N_9901);
nor U10315 (N_10315,N_9685,N_8770);
xnor U10316 (N_10316,N_9690,N_8917);
nand U10317 (N_10317,N_9154,N_8807);
nand U10318 (N_10318,N_9126,N_9665);
nand U10319 (N_10319,N_9200,N_9357);
xor U10320 (N_10320,N_8994,N_9189);
nor U10321 (N_10321,N_9202,N_8859);
xnor U10322 (N_10322,N_9718,N_9846);
nor U10323 (N_10323,N_9501,N_9037);
and U10324 (N_10324,N_9784,N_9810);
nor U10325 (N_10325,N_9115,N_9537);
nor U10326 (N_10326,N_9205,N_9147);
xor U10327 (N_10327,N_9285,N_9706);
and U10328 (N_10328,N_9985,N_9625);
and U10329 (N_10329,N_9670,N_9856);
nand U10330 (N_10330,N_9359,N_8779);
or U10331 (N_10331,N_9489,N_9541);
nor U10332 (N_10332,N_9530,N_9640);
xnor U10333 (N_10333,N_9658,N_9562);
and U10334 (N_10334,N_9168,N_8913);
nor U10335 (N_10335,N_9298,N_9292);
nor U10336 (N_10336,N_9256,N_9340);
and U10337 (N_10337,N_8845,N_8787);
nor U10338 (N_10338,N_9591,N_9125);
and U10339 (N_10339,N_9122,N_9769);
or U10340 (N_10340,N_9842,N_9878);
xnor U10341 (N_10341,N_9711,N_9998);
xnor U10342 (N_10342,N_9159,N_9695);
xor U10343 (N_10343,N_9905,N_9195);
and U10344 (N_10344,N_9804,N_9940);
nor U10345 (N_10345,N_9364,N_9809);
and U10346 (N_10346,N_9287,N_8886);
xor U10347 (N_10347,N_9975,N_9045);
xor U10348 (N_10348,N_8918,N_9895);
and U10349 (N_10349,N_8842,N_9776);
or U10350 (N_10350,N_8864,N_9451);
or U10351 (N_10351,N_9800,N_9902);
nand U10352 (N_10352,N_9651,N_9365);
nand U10353 (N_10353,N_9203,N_8780);
nor U10354 (N_10354,N_9970,N_9817);
xnor U10355 (N_10355,N_9533,N_9783);
nand U10356 (N_10356,N_9585,N_9819);
nand U10357 (N_10357,N_9966,N_8868);
nand U10358 (N_10358,N_9514,N_9394);
nor U10359 (N_10359,N_9539,N_9813);
and U10360 (N_10360,N_9103,N_8771);
nor U10361 (N_10361,N_9278,N_9151);
and U10362 (N_10362,N_8784,N_8996);
nand U10363 (N_10363,N_9030,N_9816);
and U10364 (N_10364,N_9214,N_8946);
nor U10365 (N_10365,N_9899,N_9518);
xor U10366 (N_10366,N_9306,N_9924);
nor U10367 (N_10367,N_9253,N_8895);
and U10368 (N_10368,N_9378,N_9508);
and U10369 (N_10369,N_9215,N_9113);
and U10370 (N_10370,N_9534,N_9838);
and U10371 (N_10371,N_9379,N_9388);
nand U10372 (N_10372,N_9345,N_9881);
nor U10373 (N_10373,N_9668,N_9648);
or U10374 (N_10374,N_9247,N_9092);
and U10375 (N_10375,N_9750,N_9046);
xnor U10376 (N_10376,N_9772,N_9726);
nor U10377 (N_10377,N_9177,N_8987);
or U10378 (N_10378,N_9110,N_9396);
nand U10379 (N_10379,N_8844,N_9528);
nor U10380 (N_10380,N_9252,N_9322);
nand U10381 (N_10381,N_9485,N_9270);
or U10382 (N_10382,N_9066,N_9369);
nand U10383 (N_10383,N_9259,N_9939);
nor U10384 (N_10384,N_9325,N_9313);
or U10385 (N_10385,N_9525,N_9928);
xor U10386 (N_10386,N_9207,N_9324);
xor U10387 (N_10387,N_9614,N_8764);
or U10388 (N_10388,N_8812,N_8837);
nand U10389 (N_10389,N_9931,N_9664);
or U10390 (N_10390,N_9758,N_9323);
nor U10391 (N_10391,N_9630,N_9989);
nor U10392 (N_10392,N_9462,N_9499);
and U10393 (N_10393,N_9546,N_9448);
and U10394 (N_10394,N_9179,N_9009);
nor U10395 (N_10395,N_9802,N_9644);
nor U10396 (N_10396,N_9033,N_9032);
xnor U10397 (N_10397,N_9877,N_9657);
nor U10398 (N_10398,N_9762,N_8933);
xnor U10399 (N_10399,N_9843,N_9348);
nand U10400 (N_10400,N_8756,N_9288);
nor U10401 (N_10401,N_9627,N_9209);
or U10402 (N_10402,N_9121,N_9080);
and U10403 (N_10403,N_9114,N_9669);
xor U10404 (N_10404,N_8883,N_9829);
and U10405 (N_10405,N_9036,N_8798);
xor U10406 (N_10406,N_9303,N_9407);
nand U10407 (N_10407,N_9123,N_9101);
xnor U10408 (N_10408,N_8755,N_9976);
nor U10409 (N_10409,N_9691,N_9650);
and U10410 (N_10410,N_9199,N_8991);
or U10411 (N_10411,N_8880,N_9155);
and U10412 (N_10412,N_9038,N_9759);
nand U10413 (N_10413,N_9751,N_9564);
and U10414 (N_10414,N_9291,N_9908);
nor U10415 (N_10415,N_8850,N_9169);
xnor U10416 (N_10416,N_8781,N_9059);
xor U10417 (N_10417,N_9343,N_9912);
and U10418 (N_10418,N_8969,N_9729);
xor U10419 (N_10419,N_8885,N_8926);
and U10420 (N_10420,N_9500,N_9498);
nor U10421 (N_10421,N_9316,N_9315);
nand U10422 (N_10422,N_8804,N_9629);
nand U10423 (N_10423,N_9792,N_9081);
xor U10424 (N_10424,N_9747,N_9573);
xor U10425 (N_10425,N_9480,N_9328);
xor U10426 (N_10426,N_9983,N_9304);
and U10427 (N_10427,N_8816,N_9221);
nand U10428 (N_10428,N_9467,N_9441);
nor U10429 (N_10429,N_9927,N_8814);
and U10430 (N_10430,N_9112,N_9044);
nand U10431 (N_10431,N_9090,N_9423);
nor U10432 (N_10432,N_9963,N_9787);
xor U10433 (N_10433,N_9002,N_9553);
or U10434 (N_10434,N_9610,N_9436);
nor U10435 (N_10435,N_9959,N_9148);
or U10436 (N_10436,N_9003,N_8827);
xnor U10437 (N_10437,N_9281,N_9229);
or U10438 (N_10438,N_9088,N_9693);
or U10439 (N_10439,N_9187,N_9074);
nor U10440 (N_10440,N_9861,N_9459);
nand U10441 (N_10441,N_8943,N_9381);
nand U10442 (N_10442,N_9382,N_8876);
nor U10443 (N_10443,N_9220,N_9227);
and U10444 (N_10444,N_9647,N_9803);
and U10445 (N_10445,N_9704,N_9754);
and U10446 (N_10446,N_9845,N_9137);
or U10447 (N_10447,N_8830,N_8824);
or U10448 (N_10448,N_9086,N_9255);
or U10449 (N_10449,N_9132,N_9035);
or U10450 (N_10450,N_9741,N_9515);
xor U10451 (N_10451,N_9157,N_8941);
xnor U10452 (N_10452,N_9595,N_8998);
nand U10453 (N_10453,N_8887,N_9862);
nand U10454 (N_10454,N_9544,N_9452);
and U10455 (N_10455,N_9265,N_9686);
nand U10456 (N_10456,N_9426,N_9327);
nor U10457 (N_10457,N_9788,N_9592);
and U10458 (N_10458,N_9586,N_9834);
nor U10459 (N_10459,N_9621,N_9662);
and U10460 (N_10460,N_9119,N_9238);
nor U10461 (N_10461,N_9008,N_9280);
nor U10462 (N_10462,N_8788,N_9433);
or U10463 (N_10463,N_8750,N_9532);
xor U10464 (N_10464,N_9910,N_9611);
or U10465 (N_10465,N_9116,N_9576);
nor U10466 (N_10466,N_9944,N_8914);
and U10467 (N_10467,N_9587,N_8978);
nor U10468 (N_10468,N_9736,N_9360);
or U10469 (N_10469,N_9007,N_8846);
or U10470 (N_10470,N_9305,N_9885);
nor U10471 (N_10471,N_9054,N_9279);
and U10472 (N_10472,N_8997,N_9654);
xor U10473 (N_10473,N_9569,N_9583);
nor U10474 (N_10474,N_9363,N_9590);
nor U10475 (N_10475,N_9596,N_9882);
and U10476 (N_10476,N_9475,N_9945);
or U10477 (N_10477,N_9599,N_9383);
or U10478 (N_10478,N_9185,N_9171);
xnor U10479 (N_10479,N_9026,N_9567);
and U10480 (N_10480,N_9965,N_9058);
or U10481 (N_10481,N_9443,N_9801);
nor U10482 (N_10482,N_9632,N_8904);
and U10483 (N_10483,N_9488,N_9687);
nor U10484 (N_10484,N_9742,N_8909);
nand U10485 (N_10485,N_9764,N_8922);
and U10486 (N_10486,N_8954,N_9188);
nor U10487 (N_10487,N_9716,N_9763);
or U10488 (N_10488,N_9890,N_9733);
nand U10489 (N_10489,N_9319,N_9164);
nor U10490 (N_10490,N_8828,N_9061);
nor U10491 (N_10491,N_9068,N_9120);
nand U10492 (N_10492,N_9869,N_8924);
nand U10493 (N_10493,N_9712,N_9224);
and U10494 (N_10494,N_8810,N_9698);
and U10495 (N_10495,N_9057,N_9904);
nor U10496 (N_10496,N_9552,N_8799);
xnor U10497 (N_10497,N_9484,N_9832);
or U10498 (N_10498,N_9453,N_9438);
nor U10499 (N_10499,N_9868,N_9679);
or U10500 (N_10500,N_9554,N_9309);
and U10501 (N_10501,N_8793,N_9178);
and U10502 (N_10502,N_9277,N_9183);
nand U10503 (N_10503,N_8856,N_9547);
or U10504 (N_10504,N_9184,N_9540);
and U10505 (N_10505,N_9020,N_9851);
nor U10506 (N_10506,N_9024,N_8893);
or U10507 (N_10507,N_8795,N_8871);
or U10508 (N_10508,N_9622,N_9855);
and U10509 (N_10509,N_9367,N_9677);
nand U10510 (N_10510,N_9052,N_9604);
xnor U10511 (N_10511,N_9948,N_9858);
xnor U10512 (N_10512,N_9212,N_9753);
and U10513 (N_10513,N_9258,N_8896);
and U10514 (N_10514,N_8952,N_9311);
and U10515 (N_10515,N_8995,N_9078);
nand U10516 (N_10516,N_9232,N_9545);
and U10517 (N_10517,N_8786,N_8823);
or U10518 (N_10518,N_9444,N_9135);
and U10519 (N_10519,N_9897,N_8957);
and U10520 (N_10520,N_9417,N_9336);
xor U10521 (N_10521,N_9995,N_9864);
or U10522 (N_10522,N_9874,N_9805);
nand U10523 (N_10523,N_9470,N_8835);
nor U10524 (N_10524,N_9015,N_9835);
and U10525 (N_10525,N_8802,N_8989);
nor U10526 (N_10526,N_9163,N_9368);
nor U10527 (N_10527,N_9578,N_9099);
nor U10528 (N_10528,N_8960,N_8760);
nor U10529 (N_10529,N_9506,N_9250);
xor U10530 (N_10530,N_9919,N_9523);
nor U10531 (N_10531,N_9432,N_9337);
nor U10532 (N_10532,N_8950,N_9615);
or U10533 (N_10533,N_9124,N_9653);
nor U10534 (N_10534,N_9638,N_9127);
and U10535 (N_10535,N_9913,N_9335);
nand U10536 (N_10536,N_9299,N_8961);
nor U10537 (N_10537,N_9049,N_9589);
and U10538 (N_10538,N_9979,N_8831);
nand U10539 (N_10539,N_9671,N_9635);
nor U10540 (N_10540,N_9043,N_8884);
nor U10541 (N_10541,N_9366,N_9743);
xor U10542 (N_10542,N_9522,N_9735);
nor U10543 (N_10543,N_9391,N_9660);
or U10544 (N_10544,N_9531,N_9197);
nand U10545 (N_10545,N_9117,N_9107);
and U10546 (N_10546,N_9264,N_9468);
nand U10547 (N_10547,N_9479,N_8801);
or U10548 (N_10548,N_8910,N_8751);
or U10549 (N_10549,N_9708,N_9775);
or U10550 (N_10550,N_9180,N_9089);
nor U10551 (N_10551,N_9572,N_9511);
nand U10552 (N_10552,N_9731,N_9789);
or U10553 (N_10553,N_9399,N_9951);
and U10554 (N_10554,N_9701,N_9557);
and U10555 (N_10555,N_9893,N_9225);
xor U10556 (N_10556,N_9150,N_9415);
or U10557 (N_10557,N_9464,N_9231);
nand U10558 (N_10558,N_9478,N_9779);
xor U10559 (N_10559,N_8817,N_9376);
nor U10560 (N_10560,N_9844,N_9134);
xnor U10561 (N_10561,N_9922,N_9349);
nand U10562 (N_10562,N_8822,N_9613);
or U10563 (N_10563,N_9271,N_8936);
and U10564 (N_10564,N_9509,N_9420);
and U10565 (N_10565,N_9946,N_9235);
and U10566 (N_10566,N_8785,N_9873);
nand U10567 (N_10567,N_8829,N_8925);
xor U10568 (N_10568,N_9286,N_9606);
nor U10569 (N_10569,N_9094,N_8766);
nor U10570 (N_10570,N_9566,N_9442);
and U10571 (N_10571,N_9106,N_9427);
nor U10572 (N_10572,N_9330,N_9597);
nor U10573 (N_10573,N_9143,N_9888);
or U10574 (N_10574,N_9145,N_8877);
and U10575 (N_10575,N_9402,N_9798);
nor U10576 (N_10576,N_8758,N_9571);
nor U10577 (N_10577,N_9042,N_9990);
xor U10578 (N_10578,N_8754,N_8923);
nand U10579 (N_10579,N_9952,N_9403);
xor U10580 (N_10580,N_9041,N_8944);
nor U10581 (N_10581,N_9594,N_9109);
nor U10582 (N_10582,N_9149,N_9616);
nor U10583 (N_10583,N_9011,N_8819);
or U10584 (N_10584,N_9496,N_8834);
or U10585 (N_10585,N_9860,N_9584);
xnor U10586 (N_10586,N_9344,N_9373);
and U10587 (N_10587,N_9659,N_8881);
nor U10588 (N_10588,N_9949,N_9853);
nor U10589 (N_10589,N_8921,N_8811);
nand U10590 (N_10590,N_9556,N_9626);
xnor U10591 (N_10591,N_9738,N_9312);
xnor U10592 (N_10592,N_9334,N_9392);
nand U10593 (N_10593,N_9936,N_9639);
nand U10594 (N_10594,N_9943,N_9752);
nand U10595 (N_10595,N_9593,N_9849);
or U10596 (N_10596,N_9228,N_9268);
nand U10597 (N_10597,N_9447,N_9005);
or U10598 (N_10598,N_9001,N_8919);
nor U10599 (N_10599,N_9822,N_9781);
nor U10600 (N_10600,N_8974,N_9182);
nand U10601 (N_10601,N_9457,N_9950);
xnor U10602 (N_10602,N_9300,N_9884);
or U10603 (N_10603,N_9681,N_9993);
and U10604 (N_10604,N_9463,N_9744);
nor U10605 (N_10605,N_9542,N_9111);
and U10606 (N_10606,N_8806,N_9996);
and U10607 (N_10607,N_9201,N_9139);
nor U10608 (N_10608,N_9353,N_8931);
nor U10609 (N_10609,N_9824,N_9262);
xnor U10610 (N_10610,N_9683,N_9472);
nor U10611 (N_10611,N_9056,N_9814);
nor U10612 (N_10612,N_9746,N_9602);
nor U10613 (N_10613,N_9715,N_9568);
and U10614 (N_10614,N_8951,N_9536);
nor U10615 (N_10615,N_9167,N_9339);
and U10616 (N_10616,N_9419,N_9440);
and U10617 (N_10617,N_8897,N_9972);
or U10618 (N_10618,N_9161,N_9437);
or U10619 (N_10619,N_9517,N_9409);
xor U10620 (N_10620,N_8872,N_9497);
xor U10621 (N_10621,N_9039,N_9460);
and U10622 (N_10622,N_9879,N_9839);
xor U10623 (N_10623,N_9663,N_9060);
or U10624 (N_10624,N_9777,N_8992);
nor U10625 (N_10625,N_8751,N_9132);
or U10626 (N_10626,N_9239,N_9303);
xnor U10627 (N_10627,N_9899,N_9925);
xnor U10628 (N_10628,N_9184,N_9390);
nor U10629 (N_10629,N_9537,N_9403);
and U10630 (N_10630,N_9475,N_8792);
nand U10631 (N_10631,N_9240,N_8828);
xnor U10632 (N_10632,N_9126,N_8786);
or U10633 (N_10633,N_9227,N_9798);
and U10634 (N_10634,N_8981,N_9161);
xnor U10635 (N_10635,N_9257,N_9516);
or U10636 (N_10636,N_8855,N_9976);
xnor U10637 (N_10637,N_9287,N_9402);
and U10638 (N_10638,N_8965,N_9862);
nand U10639 (N_10639,N_9728,N_9346);
and U10640 (N_10640,N_9677,N_9082);
xor U10641 (N_10641,N_8960,N_9677);
nor U10642 (N_10642,N_9227,N_9898);
xor U10643 (N_10643,N_9905,N_9324);
nand U10644 (N_10644,N_9801,N_8986);
or U10645 (N_10645,N_9308,N_8834);
xnor U10646 (N_10646,N_9030,N_8970);
or U10647 (N_10647,N_9521,N_9921);
and U10648 (N_10648,N_9248,N_8875);
xnor U10649 (N_10649,N_8893,N_9535);
nor U10650 (N_10650,N_9465,N_9813);
nor U10651 (N_10651,N_9982,N_9383);
xnor U10652 (N_10652,N_9273,N_9099);
and U10653 (N_10653,N_9502,N_9307);
nand U10654 (N_10654,N_8894,N_8850);
xor U10655 (N_10655,N_9791,N_9528);
or U10656 (N_10656,N_9153,N_9967);
and U10657 (N_10657,N_9595,N_9400);
xnor U10658 (N_10658,N_9717,N_9180);
xnor U10659 (N_10659,N_9047,N_9797);
nand U10660 (N_10660,N_9613,N_9800);
xnor U10661 (N_10661,N_9896,N_9025);
and U10662 (N_10662,N_9993,N_9600);
or U10663 (N_10663,N_9438,N_9956);
and U10664 (N_10664,N_9227,N_9033);
and U10665 (N_10665,N_9543,N_9507);
and U10666 (N_10666,N_9587,N_9332);
or U10667 (N_10667,N_9718,N_9965);
nand U10668 (N_10668,N_8914,N_9872);
xor U10669 (N_10669,N_9556,N_9615);
and U10670 (N_10670,N_9268,N_8903);
nor U10671 (N_10671,N_8893,N_9485);
nand U10672 (N_10672,N_8888,N_9608);
and U10673 (N_10673,N_9506,N_9004);
nor U10674 (N_10674,N_9213,N_8764);
xnor U10675 (N_10675,N_9916,N_9034);
nand U10676 (N_10676,N_9921,N_9258);
or U10677 (N_10677,N_8903,N_8956);
xnor U10678 (N_10678,N_9637,N_9735);
or U10679 (N_10679,N_9150,N_9420);
nor U10680 (N_10680,N_8771,N_8914);
nand U10681 (N_10681,N_9716,N_9810);
or U10682 (N_10682,N_9883,N_9578);
or U10683 (N_10683,N_9397,N_9513);
or U10684 (N_10684,N_9005,N_9721);
xor U10685 (N_10685,N_8786,N_9887);
or U10686 (N_10686,N_9136,N_9750);
or U10687 (N_10687,N_9200,N_9141);
xnor U10688 (N_10688,N_9120,N_8842);
nand U10689 (N_10689,N_9323,N_9126);
or U10690 (N_10690,N_9035,N_9408);
xor U10691 (N_10691,N_9286,N_9116);
xnor U10692 (N_10692,N_9614,N_9706);
nand U10693 (N_10693,N_9497,N_9859);
nor U10694 (N_10694,N_8929,N_8827);
nor U10695 (N_10695,N_9146,N_9599);
and U10696 (N_10696,N_9801,N_9678);
nand U10697 (N_10697,N_8842,N_8976);
nor U10698 (N_10698,N_9821,N_9259);
nand U10699 (N_10699,N_8890,N_9777);
nand U10700 (N_10700,N_8802,N_8996);
or U10701 (N_10701,N_9372,N_9832);
xor U10702 (N_10702,N_9385,N_8839);
nor U10703 (N_10703,N_9727,N_8823);
and U10704 (N_10704,N_9473,N_9111);
nor U10705 (N_10705,N_9677,N_9772);
nor U10706 (N_10706,N_9216,N_9407);
and U10707 (N_10707,N_9758,N_9568);
xnor U10708 (N_10708,N_9955,N_9897);
nand U10709 (N_10709,N_9829,N_9290);
nor U10710 (N_10710,N_9672,N_9572);
nor U10711 (N_10711,N_9650,N_9128);
nand U10712 (N_10712,N_9561,N_9078);
xnor U10713 (N_10713,N_9253,N_9619);
xor U10714 (N_10714,N_9451,N_9904);
xor U10715 (N_10715,N_9699,N_9088);
and U10716 (N_10716,N_9811,N_9493);
nand U10717 (N_10717,N_8775,N_9601);
xnor U10718 (N_10718,N_9209,N_9483);
nor U10719 (N_10719,N_9009,N_9256);
nand U10720 (N_10720,N_9911,N_9317);
nand U10721 (N_10721,N_9800,N_9003);
or U10722 (N_10722,N_9650,N_8857);
nand U10723 (N_10723,N_9579,N_9597);
xnor U10724 (N_10724,N_8916,N_8786);
nand U10725 (N_10725,N_9060,N_9552);
nor U10726 (N_10726,N_9793,N_9183);
or U10727 (N_10727,N_9033,N_9379);
or U10728 (N_10728,N_8817,N_9144);
or U10729 (N_10729,N_9186,N_9823);
nor U10730 (N_10730,N_9828,N_9717);
or U10731 (N_10731,N_9431,N_9086);
and U10732 (N_10732,N_8814,N_9776);
and U10733 (N_10733,N_9136,N_9032);
or U10734 (N_10734,N_9725,N_9619);
and U10735 (N_10735,N_9114,N_8800);
xnor U10736 (N_10736,N_9270,N_9638);
or U10737 (N_10737,N_9154,N_9927);
nand U10738 (N_10738,N_9871,N_8759);
nor U10739 (N_10739,N_8906,N_9101);
and U10740 (N_10740,N_9659,N_9289);
xnor U10741 (N_10741,N_9260,N_9291);
xnor U10742 (N_10742,N_9814,N_9182);
and U10743 (N_10743,N_9226,N_8949);
or U10744 (N_10744,N_8794,N_8828);
or U10745 (N_10745,N_9713,N_9910);
nor U10746 (N_10746,N_9173,N_8948);
nand U10747 (N_10747,N_9663,N_9588);
xnor U10748 (N_10748,N_9854,N_9498);
and U10749 (N_10749,N_9578,N_9490);
or U10750 (N_10750,N_9477,N_9936);
or U10751 (N_10751,N_9078,N_8880);
or U10752 (N_10752,N_9501,N_9725);
or U10753 (N_10753,N_8917,N_9130);
and U10754 (N_10754,N_8938,N_9428);
or U10755 (N_10755,N_9874,N_9646);
or U10756 (N_10756,N_9581,N_9616);
or U10757 (N_10757,N_8828,N_9478);
nand U10758 (N_10758,N_9243,N_9943);
and U10759 (N_10759,N_9068,N_9355);
or U10760 (N_10760,N_9405,N_9776);
nand U10761 (N_10761,N_9006,N_8868);
xor U10762 (N_10762,N_9267,N_9512);
nand U10763 (N_10763,N_8954,N_9608);
nand U10764 (N_10764,N_8782,N_9946);
or U10765 (N_10765,N_9135,N_9951);
and U10766 (N_10766,N_9793,N_9918);
xor U10767 (N_10767,N_9650,N_9988);
xnor U10768 (N_10768,N_8755,N_9984);
nor U10769 (N_10769,N_9528,N_9681);
xor U10770 (N_10770,N_9916,N_9215);
nand U10771 (N_10771,N_9640,N_9184);
and U10772 (N_10772,N_9443,N_9413);
or U10773 (N_10773,N_9430,N_9891);
nor U10774 (N_10774,N_9859,N_9485);
nand U10775 (N_10775,N_9300,N_9771);
or U10776 (N_10776,N_8807,N_9652);
nand U10777 (N_10777,N_8942,N_8761);
nor U10778 (N_10778,N_9801,N_9605);
nor U10779 (N_10779,N_8973,N_9659);
and U10780 (N_10780,N_8864,N_9870);
or U10781 (N_10781,N_9923,N_9056);
or U10782 (N_10782,N_8976,N_9863);
or U10783 (N_10783,N_9736,N_9407);
or U10784 (N_10784,N_9221,N_9085);
xor U10785 (N_10785,N_9601,N_9376);
nand U10786 (N_10786,N_9706,N_9423);
nor U10787 (N_10787,N_8956,N_9987);
and U10788 (N_10788,N_9777,N_9922);
and U10789 (N_10789,N_8965,N_9763);
and U10790 (N_10790,N_9428,N_9420);
xnor U10791 (N_10791,N_9131,N_9817);
nand U10792 (N_10792,N_9802,N_9076);
xnor U10793 (N_10793,N_9876,N_8890);
nand U10794 (N_10794,N_9542,N_9572);
nor U10795 (N_10795,N_8859,N_9676);
nand U10796 (N_10796,N_9424,N_8756);
and U10797 (N_10797,N_8987,N_9589);
nor U10798 (N_10798,N_9242,N_8810);
xnor U10799 (N_10799,N_9305,N_9696);
nor U10800 (N_10800,N_9504,N_9568);
xor U10801 (N_10801,N_9952,N_8769);
xnor U10802 (N_10802,N_9610,N_9110);
nand U10803 (N_10803,N_9265,N_9628);
nand U10804 (N_10804,N_9146,N_9898);
xor U10805 (N_10805,N_9491,N_9582);
or U10806 (N_10806,N_9692,N_9183);
nand U10807 (N_10807,N_9648,N_9545);
xnor U10808 (N_10808,N_9565,N_8875);
or U10809 (N_10809,N_9060,N_9499);
and U10810 (N_10810,N_9821,N_9128);
xor U10811 (N_10811,N_9580,N_9013);
or U10812 (N_10812,N_9198,N_9789);
nor U10813 (N_10813,N_9278,N_9619);
xor U10814 (N_10814,N_9029,N_9373);
and U10815 (N_10815,N_8810,N_9853);
nand U10816 (N_10816,N_9141,N_9494);
nand U10817 (N_10817,N_9191,N_9835);
xnor U10818 (N_10818,N_9770,N_9241);
xor U10819 (N_10819,N_9745,N_8876);
and U10820 (N_10820,N_9749,N_9470);
and U10821 (N_10821,N_9122,N_8766);
or U10822 (N_10822,N_9993,N_9521);
nor U10823 (N_10823,N_9172,N_9859);
nor U10824 (N_10824,N_9663,N_9642);
nand U10825 (N_10825,N_9925,N_9163);
and U10826 (N_10826,N_8927,N_9894);
xnor U10827 (N_10827,N_9250,N_9118);
xnor U10828 (N_10828,N_9954,N_9980);
xor U10829 (N_10829,N_8893,N_9808);
or U10830 (N_10830,N_9804,N_8938);
nand U10831 (N_10831,N_9523,N_9385);
and U10832 (N_10832,N_9719,N_8780);
nand U10833 (N_10833,N_9157,N_9749);
nor U10834 (N_10834,N_9485,N_8938);
nor U10835 (N_10835,N_9502,N_9379);
nor U10836 (N_10836,N_8823,N_8813);
or U10837 (N_10837,N_9210,N_9212);
nand U10838 (N_10838,N_9221,N_9458);
nand U10839 (N_10839,N_8835,N_9347);
nand U10840 (N_10840,N_9519,N_8939);
and U10841 (N_10841,N_9108,N_8964);
nor U10842 (N_10842,N_9856,N_9842);
or U10843 (N_10843,N_8788,N_9555);
nand U10844 (N_10844,N_9927,N_9950);
xor U10845 (N_10845,N_9544,N_9104);
and U10846 (N_10846,N_9164,N_8993);
nand U10847 (N_10847,N_9044,N_9457);
xnor U10848 (N_10848,N_9321,N_8890);
xnor U10849 (N_10849,N_9606,N_9993);
or U10850 (N_10850,N_9282,N_9078);
nor U10851 (N_10851,N_9490,N_9980);
nand U10852 (N_10852,N_9558,N_9058);
nand U10853 (N_10853,N_9849,N_9433);
xor U10854 (N_10854,N_9414,N_8996);
nand U10855 (N_10855,N_9193,N_9521);
xnor U10856 (N_10856,N_8884,N_9680);
nor U10857 (N_10857,N_9348,N_8881);
nor U10858 (N_10858,N_9976,N_9523);
nand U10859 (N_10859,N_9676,N_9677);
nand U10860 (N_10860,N_9887,N_9109);
and U10861 (N_10861,N_9863,N_9376);
xnor U10862 (N_10862,N_9433,N_9783);
xor U10863 (N_10863,N_9171,N_8778);
or U10864 (N_10864,N_9903,N_9720);
or U10865 (N_10865,N_9612,N_9818);
or U10866 (N_10866,N_9715,N_9463);
or U10867 (N_10867,N_9636,N_8993);
xor U10868 (N_10868,N_9052,N_9033);
nand U10869 (N_10869,N_9824,N_9730);
or U10870 (N_10870,N_9405,N_8972);
or U10871 (N_10871,N_9167,N_9768);
nand U10872 (N_10872,N_8834,N_8929);
or U10873 (N_10873,N_9878,N_9900);
or U10874 (N_10874,N_9694,N_8869);
nand U10875 (N_10875,N_9688,N_9842);
nor U10876 (N_10876,N_9770,N_9978);
and U10877 (N_10877,N_9568,N_9795);
and U10878 (N_10878,N_9826,N_9535);
nand U10879 (N_10879,N_9499,N_9604);
nor U10880 (N_10880,N_8906,N_9098);
nor U10881 (N_10881,N_8826,N_9727);
or U10882 (N_10882,N_9250,N_8957);
or U10883 (N_10883,N_9596,N_9723);
or U10884 (N_10884,N_9678,N_9737);
xor U10885 (N_10885,N_9482,N_9608);
xor U10886 (N_10886,N_9602,N_9555);
nor U10887 (N_10887,N_9628,N_9712);
and U10888 (N_10888,N_8873,N_9004);
nor U10889 (N_10889,N_9940,N_9326);
nor U10890 (N_10890,N_9457,N_9636);
nor U10891 (N_10891,N_9466,N_9612);
nor U10892 (N_10892,N_9349,N_9693);
and U10893 (N_10893,N_9679,N_9233);
nor U10894 (N_10894,N_9090,N_9293);
nand U10895 (N_10895,N_9651,N_9025);
nand U10896 (N_10896,N_9992,N_9561);
nor U10897 (N_10897,N_8952,N_9943);
nor U10898 (N_10898,N_9881,N_8876);
xor U10899 (N_10899,N_9270,N_9935);
and U10900 (N_10900,N_9293,N_9144);
nand U10901 (N_10901,N_9109,N_9309);
or U10902 (N_10902,N_9454,N_9593);
nand U10903 (N_10903,N_9240,N_9651);
and U10904 (N_10904,N_9838,N_9643);
nand U10905 (N_10905,N_8985,N_9301);
nor U10906 (N_10906,N_8874,N_9316);
and U10907 (N_10907,N_9570,N_9179);
nor U10908 (N_10908,N_9812,N_9855);
and U10909 (N_10909,N_8924,N_8814);
xnor U10910 (N_10910,N_9432,N_9305);
nand U10911 (N_10911,N_9476,N_9899);
nand U10912 (N_10912,N_9196,N_9881);
nand U10913 (N_10913,N_9758,N_9019);
nor U10914 (N_10914,N_9854,N_8942);
nand U10915 (N_10915,N_9288,N_9071);
and U10916 (N_10916,N_8900,N_9707);
nand U10917 (N_10917,N_9081,N_9501);
and U10918 (N_10918,N_8768,N_9594);
or U10919 (N_10919,N_8812,N_9561);
nor U10920 (N_10920,N_9911,N_9262);
or U10921 (N_10921,N_9834,N_9100);
xor U10922 (N_10922,N_9171,N_9188);
nor U10923 (N_10923,N_9548,N_9289);
xor U10924 (N_10924,N_9550,N_9576);
or U10925 (N_10925,N_9117,N_9609);
nand U10926 (N_10926,N_9001,N_9355);
and U10927 (N_10927,N_9507,N_9681);
nor U10928 (N_10928,N_9877,N_8932);
or U10929 (N_10929,N_8834,N_8910);
xnor U10930 (N_10930,N_8817,N_9530);
nand U10931 (N_10931,N_9293,N_8768);
nor U10932 (N_10932,N_8975,N_9346);
or U10933 (N_10933,N_9943,N_9967);
nor U10934 (N_10934,N_9418,N_9451);
or U10935 (N_10935,N_9756,N_9474);
nand U10936 (N_10936,N_9157,N_9093);
nand U10937 (N_10937,N_9241,N_8776);
and U10938 (N_10938,N_9559,N_9245);
xor U10939 (N_10939,N_9712,N_9591);
nor U10940 (N_10940,N_8801,N_8769);
nand U10941 (N_10941,N_9306,N_9161);
xor U10942 (N_10942,N_9172,N_9339);
nor U10943 (N_10943,N_9154,N_9308);
and U10944 (N_10944,N_9614,N_9607);
nand U10945 (N_10945,N_8908,N_8958);
and U10946 (N_10946,N_9592,N_9161);
or U10947 (N_10947,N_9567,N_9445);
or U10948 (N_10948,N_9089,N_9316);
xor U10949 (N_10949,N_9104,N_9965);
or U10950 (N_10950,N_9204,N_8853);
nor U10951 (N_10951,N_8884,N_9529);
nor U10952 (N_10952,N_8932,N_9293);
nand U10953 (N_10953,N_8917,N_9497);
and U10954 (N_10954,N_9172,N_9389);
nand U10955 (N_10955,N_9543,N_9985);
or U10956 (N_10956,N_9651,N_8996);
nor U10957 (N_10957,N_9215,N_9132);
and U10958 (N_10958,N_9450,N_9820);
or U10959 (N_10959,N_8897,N_9812);
xnor U10960 (N_10960,N_9272,N_8940);
nand U10961 (N_10961,N_9683,N_9474);
nand U10962 (N_10962,N_9102,N_9608);
or U10963 (N_10963,N_9529,N_9789);
xor U10964 (N_10964,N_9362,N_8782);
nand U10965 (N_10965,N_9246,N_9719);
or U10966 (N_10966,N_9848,N_9756);
xor U10967 (N_10967,N_9323,N_9182);
xnor U10968 (N_10968,N_9447,N_8961);
nand U10969 (N_10969,N_9098,N_8936);
nand U10970 (N_10970,N_9506,N_9397);
nand U10971 (N_10971,N_9927,N_9850);
nor U10972 (N_10972,N_9713,N_8956);
and U10973 (N_10973,N_9746,N_9025);
and U10974 (N_10974,N_9674,N_9797);
nand U10975 (N_10975,N_9812,N_8823);
nor U10976 (N_10976,N_9190,N_8929);
and U10977 (N_10977,N_9416,N_9033);
xnor U10978 (N_10978,N_8752,N_9023);
nor U10979 (N_10979,N_9354,N_8905);
nand U10980 (N_10980,N_9146,N_9894);
nor U10981 (N_10981,N_9609,N_9759);
nand U10982 (N_10982,N_9899,N_8770);
nor U10983 (N_10983,N_9296,N_9995);
xnor U10984 (N_10984,N_9523,N_9931);
and U10985 (N_10985,N_8999,N_9811);
nand U10986 (N_10986,N_8829,N_9544);
nand U10987 (N_10987,N_9443,N_9458);
and U10988 (N_10988,N_9893,N_8978);
xor U10989 (N_10989,N_9685,N_9261);
or U10990 (N_10990,N_9102,N_9636);
xnor U10991 (N_10991,N_9903,N_9695);
or U10992 (N_10992,N_8804,N_8955);
nor U10993 (N_10993,N_9691,N_9209);
or U10994 (N_10994,N_9833,N_8929);
xnor U10995 (N_10995,N_9763,N_9227);
nand U10996 (N_10996,N_9360,N_9551);
nor U10997 (N_10997,N_8967,N_9537);
xnor U10998 (N_10998,N_9864,N_9898);
and U10999 (N_10999,N_9051,N_8918);
xnor U11000 (N_11000,N_8894,N_8766);
nor U11001 (N_11001,N_9026,N_9028);
nand U11002 (N_11002,N_8901,N_9072);
xnor U11003 (N_11003,N_9489,N_9014);
or U11004 (N_11004,N_9697,N_8752);
nand U11005 (N_11005,N_9827,N_9783);
or U11006 (N_11006,N_9079,N_9544);
xnor U11007 (N_11007,N_9332,N_9865);
or U11008 (N_11008,N_9316,N_9564);
nor U11009 (N_11009,N_9007,N_9738);
nand U11010 (N_11010,N_9793,N_9541);
or U11011 (N_11011,N_9875,N_8795);
nand U11012 (N_11012,N_9466,N_9358);
nand U11013 (N_11013,N_9090,N_9601);
xor U11014 (N_11014,N_9063,N_9177);
and U11015 (N_11015,N_8828,N_9824);
nand U11016 (N_11016,N_9267,N_9177);
or U11017 (N_11017,N_9700,N_8896);
or U11018 (N_11018,N_9544,N_9100);
nor U11019 (N_11019,N_9065,N_9973);
and U11020 (N_11020,N_9824,N_9495);
and U11021 (N_11021,N_9575,N_9522);
xnor U11022 (N_11022,N_9227,N_9562);
nor U11023 (N_11023,N_8828,N_9379);
nor U11024 (N_11024,N_9346,N_8797);
xnor U11025 (N_11025,N_9741,N_9270);
nor U11026 (N_11026,N_9625,N_9555);
nand U11027 (N_11027,N_9342,N_8758);
and U11028 (N_11028,N_9213,N_8890);
nand U11029 (N_11029,N_8856,N_9961);
and U11030 (N_11030,N_9089,N_8925);
and U11031 (N_11031,N_9929,N_9901);
nor U11032 (N_11032,N_9342,N_9370);
xnor U11033 (N_11033,N_9908,N_9602);
and U11034 (N_11034,N_9184,N_9457);
nor U11035 (N_11035,N_9645,N_9970);
and U11036 (N_11036,N_8865,N_8907);
nor U11037 (N_11037,N_8804,N_9433);
or U11038 (N_11038,N_9345,N_9839);
xnor U11039 (N_11039,N_9991,N_9063);
nand U11040 (N_11040,N_9310,N_9904);
and U11041 (N_11041,N_9279,N_9370);
or U11042 (N_11042,N_8850,N_9647);
nand U11043 (N_11043,N_9482,N_9389);
or U11044 (N_11044,N_9219,N_9471);
and U11045 (N_11045,N_8805,N_9083);
nor U11046 (N_11046,N_9412,N_9831);
or U11047 (N_11047,N_9758,N_8874);
or U11048 (N_11048,N_9640,N_8992);
and U11049 (N_11049,N_9460,N_9152);
or U11050 (N_11050,N_9266,N_9329);
and U11051 (N_11051,N_9240,N_8858);
or U11052 (N_11052,N_9126,N_9868);
or U11053 (N_11053,N_8866,N_9374);
xor U11054 (N_11054,N_9306,N_8839);
nand U11055 (N_11055,N_9186,N_8758);
and U11056 (N_11056,N_8912,N_9796);
xnor U11057 (N_11057,N_9565,N_9613);
xnor U11058 (N_11058,N_8898,N_9378);
nor U11059 (N_11059,N_8897,N_9457);
nand U11060 (N_11060,N_9623,N_9320);
nand U11061 (N_11061,N_9022,N_9872);
or U11062 (N_11062,N_9878,N_9606);
nor U11063 (N_11063,N_8913,N_9337);
nor U11064 (N_11064,N_9375,N_9406);
xor U11065 (N_11065,N_8902,N_9940);
nand U11066 (N_11066,N_9447,N_9033);
or U11067 (N_11067,N_9504,N_9354);
and U11068 (N_11068,N_8936,N_9766);
nand U11069 (N_11069,N_9244,N_8922);
xor U11070 (N_11070,N_9105,N_9229);
nor U11071 (N_11071,N_9601,N_9754);
and U11072 (N_11072,N_8799,N_9640);
or U11073 (N_11073,N_8992,N_9080);
and U11074 (N_11074,N_9906,N_9157);
and U11075 (N_11075,N_9892,N_9896);
nand U11076 (N_11076,N_9369,N_9312);
and U11077 (N_11077,N_9253,N_9097);
and U11078 (N_11078,N_9613,N_8922);
and U11079 (N_11079,N_9722,N_9090);
nand U11080 (N_11080,N_9606,N_9117);
nor U11081 (N_11081,N_9182,N_9292);
nand U11082 (N_11082,N_9687,N_9737);
and U11083 (N_11083,N_9374,N_9156);
or U11084 (N_11084,N_9486,N_9238);
nor U11085 (N_11085,N_8804,N_9547);
xnor U11086 (N_11086,N_9615,N_9359);
and U11087 (N_11087,N_8858,N_9625);
and U11088 (N_11088,N_9868,N_9912);
or U11089 (N_11089,N_8918,N_9785);
xnor U11090 (N_11090,N_9577,N_9302);
nor U11091 (N_11091,N_9841,N_8920);
nand U11092 (N_11092,N_9036,N_9895);
and U11093 (N_11093,N_9774,N_9686);
or U11094 (N_11094,N_9857,N_9512);
and U11095 (N_11095,N_9001,N_8903);
and U11096 (N_11096,N_9307,N_9467);
or U11097 (N_11097,N_9333,N_8856);
nand U11098 (N_11098,N_8881,N_8898);
and U11099 (N_11099,N_9035,N_9856);
nand U11100 (N_11100,N_9311,N_9168);
or U11101 (N_11101,N_9777,N_9249);
xor U11102 (N_11102,N_8751,N_9851);
and U11103 (N_11103,N_9255,N_9117);
and U11104 (N_11104,N_8858,N_9056);
nor U11105 (N_11105,N_9305,N_8794);
and U11106 (N_11106,N_9654,N_8939);
and U11107 (N_11107,N_9500,N_9237);
nand U11108 (N_11108,N_9527,N_9488);
or U11109 (N_11109,N_9167,N_9988);
and U11110 (N_11110,N_9040,N_9333);
xor U11111 (N_11111,N_9392,N_9512);
or U11112 (N_11112,N_9084,N_9487);
nor U11113 (N_11113,N_8837,N_8826);
and U11114 (N_11114,N_8851,N_9951);
or U11115 (N_11115,N_9835,N_9109);
and U11116 (N_11116,N_9976,N_9080);
or U11117 (N_11117,N_8762,N_9400);
xor U11118 (N_11118,N_9810,N_9465);
and U11119 (N_11119,N_9192,N_8853);
and U11120 (N_11120,N_9339,N_9037);
and U11121 (N_11121,N_9718,N_9112);
or U11122 (N_11122,N_9603,N_8938);
or U11123 (N_11123,N_9565,N_9423);
or U11124 (N_11124,N_9006,N_9822);
or U11125 (N_11125,N_9501,N_9815);
xnor U11126 (N_11126,N_8979,N_9299);
xnor U11127 (N_11127,N_9588,N_9492);
or U11128 (N_11128,N_9474,N_9912);
nor U11129 (N_11129,N_9548,N_9476);
or U11130 (N_11130,N_8994,N_9764);
nor U11131 (N_11131,N_9911,N_9101);
nor U11132 (N_11132,N_9693,N_8912);
or U11133 (N_11133,N_8985,N_9560);
nand U11134 (N_11134,N_9589,N_9360);
nor U11135 (N_11135,N_9354,N_9164);
xnor U11136 (N_11136,N_9884,N_9234);
or U11137 (N_11137,N_9430,N_9150);
and U11138 (N_11138,N_9028,N_9125);
and U11139 (N_11139,N_9461,N_8986);
nand U11140 (N_11140,N_9554,N_8758);
or U11141 (N_11141,N_9836,N_9498);
xnor U11142 (N_11142,N_9600,N_8786);
nor U11143 (N_11143,N_9679,N_8772);
xnor U11144 (N_11144,N_8803,N_9165);
and U11145 (N_11145,N_9742,N_9111);
and U11146 (N_11146,N_9497,N_9352);
xnor U11147 (N_11147,N_9439,N_8806);
or U11148 (N_11148,N_8901,N_9167);
nor U11149 (N_11149,N_9124,N_8992);
nand U11150 (N_11150,N_8951,N_8996);
nand U11151 (N_11151,N_9815,N_9435);
or U11152 (N_11152,N_9198,N_9159);
nor U11153 (N_11153,N_9277,N_9197);
xnor U11154 (N_11154,N_9760,N_9946);
or U11155 (N_11155,N_9828,N_9340);
xor U11156 (N_11156,N_9681,N_9369);
or U11157 (N_11157,N_8858,N_9051);
xor U11158 (N_11158,N_9987,N_9193);
xnor U11159 (N_11159,N_8854,N_9280);
or U11160 (N_11160,N_9935,N_9563);
and U11161 (N_11161,N_9871,N_8804);
or U11162 (N_11162,N_9765,N_9517);
or U11163 (N_11163,N_9923,N_8832);
nand U11164 (N_11164,N_9554,N_9534);
or U11165 (N_11165,N_9368,N_9895);
xor U11166 (N_11166,N_9321,N_9961);
nor U11167 (N_11167,N_9902,N_9080);
nor U11168 (N_11168,N_9721,N_9685);
nor U11169 (N_11169,N_9806,N_9038);
nand U11170 (N_11170,N_9372,N_9804);
or U11171 (N_11171,N_9914,N_8995);
xnor U11172 (N_11172,N_9855,N_9061);
nand U11173 (N_11173,N_9298,N_9851);
xnor U11174 (N_11174,N_9495,N_8902);
nor U11175 (N_11175,N_8991,N_9974);
or U11176 (N_11176,N_9565,N_9438);
nor U11177 (N_11177,N_8755,N_9272);
nand U11178 (N_11178,N_9773,N_9336);
and U11179 (N_11179,N_9271,N_9558);
nor U11180 (N_11180,N_9542,N_9262);
nand U11181 (N_11181,N_8967,N_9734);
and U11182 (N_11182,N_9523,N_9015);
xnor U11183 (N_11183,N_9412,N_9887);
and U11184 (N_11184,N_9338,N_9355);
or U11185 (N_11185,N_9408,N_9341);
xnor U11186 (N_11186,N_9269,N_8793);
and U11187 (N_11187,N_9463,N_9394);
and U11188 (N_11188,N_9021,N_9120);
nor U11189 (N_11189,N_8767,N_9336);
nand U11190 (N_11190,N_9450,N_8905);
or U11191 (N_11191,N_8929,N_9594);
or U11192 (N_11192,N_9808,N_9457);
and U11193 (N_11193,N_9912,N_9228);
nand U11194 (N_11194,N_9825,N_8915);
nor U11195 (N_11195,N_9112,N_9288);
and U11196 (N_11196,N_8990,N_8901);
xor U11197 (N_11197,N_9218,N_8956);
or U11198 (N_11198,N_9054,N_8753);
nand U11199 (N_11199,N_9564,N_9623);
nand U11200 (N_11200,N_9729,N_9201);
and U11201 (N_11201,N_8774,N_9936);
xor U11202 (N_11202,N_9174,N_9975);
nand U11203 (N_11203,N_9123,N_9351);
nand U11204 (N_11204,N_9135,N_8877);
and U11205 (N_11205,N_9948,N_8786);
nor U11206 (N_11206,N_9648,N_9877);
xnor U11207 (N_11207,N_8902,N_8953);
and U11208 (N_11208,N_9645,N_9796);
nor U11209 (N_11209,N_9417,N_9387);
or U11210 (N_11210,N_9125,N_9827);
nor U11211 (N_11211,N_9886,N_9670);
and U11212 (N_11212,N_9685,N_9457);
and U11213 (N_11213,N_9627,N_9647);
nor U11214 (N_11214,N_9742,N_8903);
xnor U11215 (N_11215,N_9747,N_9731);
nand U11216 (N_11216,N_8806,N_9326);
nor U11217 (N_11217,N_8874,N_9464);
nand U11218 (N_11218,N_9551,N_9389);
and U11219 (N_11219,N_9997,N_9527);
or U11220 (N_11220,N_9352,N_8905);
xnor U11221 (N_11221,N_9353,N_9055);
nand U11222 (N_11222,N_8881,N_9641);
or U11223 (N_11223,N_9681,N_9510);
and U11224 (N_11224,N_9881,N_9880);
xnor U11225 (N_11225,N_9555,N_9535);
or U11226 (N_11226,N_8814,N_9407);
and U11227 (N_11227,N_8996,N_9242);
nand U11228 (N_11228,N_9934,N_9093);
nand U11229 (N_11229,N_9011,N_8824);
xnor U11230 (N_11230,N_9704,N_8905);
nor U11231 (N_11231,N_9142,N_9071);
and U11232 (N_11232,N_9916,N_9095);
nand U11233 (N_11233,N_9623,N_8762);
nand U11234 (N_11234,N_9910,N_9479);
nor U11235 (N_11235,N_9903,N_9828);
nand U11236 (N_11236,N_9930,N_9310);
nor U11237 (N_11237,N_8872,N_8908);
xor U11238 (N_11238,N_9404,N_8973);
and U11239 (N_11239,N_9418,N_9619);
xor U11240 (N_11240,N_8793,N_9157);
or U11241 (N_11241,N_9199,N_9761);
or U11242 (N_11242,N_9559,N_9782);
and U11243 (N_11243,N_9690,N_9341);
and U11244 (N_11244,N_9980,N_9459);
nor U11245 (N_11245,N_9189,N_9284);
and U11246 (N_11246,N_9440,N_9883);
xor U11247 (N_11247,N_9608,N_9176);
nor U11248 (N_11248,N_8969,N_8898);
nor U11249 (N_11249,N_9753,N_9818);
or U11250 (N_11250,N_10742,N_10984);
and U11251 (N_11251,N_10830,N_10212);
nor U11252 (N_11252,N_10911,N_10128);
or U11253 (N_11253,N_11089,N_11153);
nand U11254 (N_11254,N_11021,N_10546);
nand U11255 (N_11255,N_11129,N_10088);
nor U11256 (N_11256,N_10424,N_10447);
and U11257 (N_11257,N_10065,N_11006);
and U11258 (N_11258,N_10127,N_10502);
and U11259 (N_11259,N_10946,N_11057);
xnor U11260 (N_11260,N_11144,N_10098);
nor U11261 (N_11261,N_10862,N_10720);
nand U11262 (N_11262,N_10311,N_10285);
nor U11263 (N_11263,N_10225,N_10522);
or U11264 (N_11264,N_10988,N_10373);
and U11265 (N_11265,N_10171,N_10589);
nand U11266 (N_11266,N_10387,N_10467);
xnor U11267 (N_11267,N_10487,N_10086);
and U11268 (N_11268,N_10395,N_10158);
and U11269 (N_11269,N_11123,N_10622);
and U11270 (N_11270,N_10433,N_10140);
or U11271 (N_11271,N_11192,N_10631);
nand U11272 (N_11272,N_10020,N_10030);
or U11273 (N_11273,N_10340,N_10381);
nor U11274 (N_11274,N_10841,N_10796);
xor U11275 (N_11275,N_10904,N_10397);
and U11276 (N_11276,N_10644,N_11062);
and U11277 (N_11277,N_10723,N_10084);
nand U11278 (N_11278,N_11172,N_10312);
and U11279 (N_11279,N_10174,N_11186);
and U11280 (N_11280,N_10139,N_10001);
nor U11281 (N_11281,N_10492,N_11064);
and U11282 (N_11282,N_10846,N_10951);
nor U11283 (N_11283,N_10221,N_11048);
or U11284 (N_11284,N_11245,N_10439);
or U11285 (N_11285,N_10822,N_10563);
nor U11286 (N_11286,N_10787,N_10462);
and U11287 (N_11287,N_11247,N_10364);
nor U11288 (N_11288,N_10125,N_10935);
nand U11289 (N_11289,N_11105,N_10168);
or U11290 (N_11290,N_10993,N_10342);
and U11291 (N_11291,N_10069,N_11157);
and U11292 (N_11292,N_10678,N_10251);
and U11293 (N_11293,N_10129,N_10294);
nor U11294 (N_11294,N_11097,N_10777);
nand U11295 (N_11295,N_10775,N_10421);
or U11296 (N_11296,N_10934,N_10949);
nand U11297 (N_11297,N_10277,N_10301);
xnor U11298 (N_11298,N_10386,N_10704);
nor U11299 (N_11299,N_10580,N_10976);
or U11300 (N_11300,N_11221,N_10436);
nand U11301 (N_11301,N_10363,N_11060);
or U11302 (N_11302,N_10121,N_10407);
and U11303 (N_11303,N_10246,N_11036);
and U11304 (N_11304,N_10416,N_11027);
and U11305 (N_11305,N_10939,N_11068);
or U11306 (N_11306,N_10728,N_11082);
or U11307 (N_11307,N_10006,N_10960);
nor U11308 (N_11308,N_10553,N_10926);
or U11309 (N_11309,N_10019,N_10990);
or U11310 (N_11310,N_11205,N_11076);
nand U11311 (N_11311,N_10972,N_10017);
nand U11312 (N_11312,N_10942,N_10235);
nor U11313 (N_11313,N_10901,N_10895);
or U11314 (N_11314,N_10769,N_11067);
and U11315 (N_11315,N_10076,N_11026);
and U11316 (N_11316,N_10996,N_10481);
and U11317 (N_11317,N_10583,N_10443);
or U11318 (N_11318,N_10919,N_11243);
or U11319 (N_11319,N_10037,N_10776);
xnor U11320 (N_11320,N_10913,N_11104);
xnor U11321 (N_11321,N_11019,N_10666);
nor U11322 (N_11322,N_10551,N_10152);
or U11323 (N_11323,N_11053,N_10864);
nand U11324 (N_11324,N_10741,N_10422);
nand U11325 (N_11325,N_10555,N_11229);
and U11326 (N_11326,N_10708,N_10624);
and U11327 (N_11327,N_10727,N_10784);
nor U11328 (N_11328,N_10890,N_11035);
and U11329 (N_11329,N_10718,N_11179);
xnor U11330 (N_11330,N_10535,N_10073);
or U11331 (N_11331,N_10119,N_11195);
and U11332 (N_11332,N_10560,N_10157);
xnor U11333 (N_11333,N_10928,N_10593);
or U11334 (N_11334,N_11014,N_10868);
nor U11335 (N_11335,N_10420,N_11239);
xor U11336 (N_11336,N_10645,N_10962);
and U11337 (N_11337,N_10595,N_10449);
nor U11338 (N_11338,N_10191,N_11156);
nor U11339 (N_11339,N_10562,N_10520);
nor U11340 (N_11340,N_10791,N_10240);
or U11341 (N_11341,N_10968,N_10599);
and U11342 (N_11342,N_11093,N_10078);
and U11343 (N_11343,N_10346,N_10237);
nor U11344 (N_11344,N_10423,N_10401);
xor U11345 (N_11345,N_10063,N_10557);
and U11346 (N_11346,N_10686,N_10501);
and U11347 (N_11347,N_10307,N_10893);
nor U11348 (N_11348,N_10305,N_10513);
nor U11349 (N_11349,N_10500,N_10012);
and U11350 (N_11350,N_10573,N_10412);
or U11351 (N_11351,N_10596,N_10924);
nand U11352 (N_11352,N_10350,N_11161);
nand U11353 (N_11353,N_10998,N_11016);
xnor U11354 (N_11354,N_10007,N_10041);
or U11355 (N_11355,N_10915,N_11199);
and U11356 (N_11356,N_11244,N_10751);
and U11357 (N_11357,N_10837,N_10612);
and U11358 (N_11358,N_10633,N_10630);
nand U11359 (N_11359,N_10605,N_10179);
xnor U11360 (N_11360,N_10690,N_10441);
nand U11361 (N_11361,N_11023,N_10014);
or U11362 (N_11362,N_10679,N_10745);
nor U11363 (N_11363,N_10571,N_10877);
and U11364 (N_11364,N_10002,N_10556);
xor U11365 (N_11365,N_11041,N_10315);
xnor U11366 (N_11366,N_10023,N_10714);
nand U11367 (N_11367,N_11081,N_10493);
and U11368 (N_11368,N_10117,N_11102);
nand U11369 (N_11369,N_11071,N_10232);
xnor U11370 (N_11370,N_10146,N_11055);
or U11371 (N_11371,N_10840,N_11003);
xor U11372 (N_11372,N_10101,N_10133);
xor U11373 (N_11373,N_10731,N_10115);
and U11374 (N_11374,N_11122,N_10565);
nor U11375 (N_11375,N_11086,N_10411);
and U11376 (N_11376,N_10740,N_10602);
or U11377 (N_11377,N_11240,N_10124);
nand U11378 (N_11378,N_10961,N_11131);
and U11379 (N_11379,N_11002,N_10244);
or U11380 (N_11380,N_10061,N_10752);
or U11381 (N_11381,N_11040,N_10626);
nor U11382 (N_11382,N_11018,N_10808);
nand U11383 (N_11383,N_10943,N_10722);
nor U11384 (N_11384,N_10349,N_10313);
xor U11385 (N_11385,N_10814,N_10999);
xor U11386 (N_11386,N_10217,N_10187);
nor U11387 (N_11387,N_10706,N_10032);
nand U11388 (N_11388,N_11181,N_11098);
and U11389 (N_11389,N_11127,N_10149);
xnor U11390 (N_11390,N_10974,N_11012);
or U11391 (N_11391,N_10995,N_11106);
nand U11392 (N_11392,N_11201,N_10569);
or U11393 (N_11393,N_10445,N_10184);
and U11394 (N_11394,N_11237,N_10647);
and U11395 (N_11395,N_10668,N_11162);
xnor U11396 (N_11396,N_11078,N_10483);
or U11397 (N_11397,N_10224,N_10248);
or U11398 (N_11398,N_10850,N_10883);
nor U11399 (N_11399,N_10338,N_10711);
or U11400 (N_11400,N_10189,N_10074);
nor U11401 (N_11401,N_10444,N_10105);
nor U11402 (N_11402,N_10749,N_11169);
xor U11403 (N_11403,N_10255,N_10729);
nor U11404 (N_11404,N_11167,N_10800);
nand U11405 (N_11405,N_10495,N_10818);
or U11406 (N_11406,N_10476,N_10035);
or U11407 (N_11407,N_10498,N_10308);
nor U11408 (N_11408,N_10427,N_10732);
nand U11409 (N_11409,N_10337,N_10709);
nand U11410 (N_11410,N_10151,N_10587);
nand U11411 (N_11411,N_10440,N_10458);
and U11412 (N_11412,N_10572,N_10684);
and U11413 (N_11413,N_11015,N_10652);
or U11414 (N_11414,N_10180,N_10537);
or U11415 (N_11415,N_10639,N_10812);
nor U11416 (N_11416,N_10548,N_10888);
nand U11417 (N_11417,N_10543,N_11143);
nor U11418 (N_11418,N_10003,N_10432);
nand U11419 (N_11419,N_11159,N_10102);
xor U11420 (N_11420,N_10403,N_10056);
nor U11421 (N_11421,N_10024,N_11005);
xor U11422 (N_11422,N_11045,N_10053);
and U11423 (N_11423,N_10369,N_10468);
and U11424 (N_11424,N_10733,N_10821);
nor U11425 (N_11425,N_11059,N_10504);
xnor U11426 (N_11426,N_10638,N_11158);
nor U11427 (N_11427,N_10717,N_11100);
nor U11428 (N_11428,N_11011,N_10849);
nand U11429 (N_11429,N_11017,N_10848);
and U11430 (N_11430,N_11185,N_10524);
or U11431 (N_11431,N_10887,N_10367);
nand U11432 (N_11432,N_10092,N_10667);
xnor U11433 (N_11433,N_11032,N_10320);
xnor U11434 (N_11434,N_10527,N_11038);
and U11435 (N_11435,N_10044,N_10496);
or U11436 (N_11436,N_10170,N_10173);
xnor U11437 (N_11437,N_10585,N_10229);
nand U11438 (N_11438,N_11217,N_11149);
or U11439 (N_11439,N_10798,N_10021);
xor U11440 (N_11440,N_10721,N_10907);
and U11441 (N_11441,N_10809,N_11058);
and U11442 (N_11442,N_10159,N_10860);
nand U11443 (N_11443,N_10402,N_10955);
and U11444 (N_11444,N_11160,N_10760);
xor U11445 (N_11445,N_10870,N_10788);
and U11446 (N_11446,N_10190,N_11213);
xor U11447 (N_11447,N_10687,N_10245);
nor U11448 (N_11448,N_10658,N_10163);
xor U11449 (N_11449,N_10810,N_10359);
nor U11450 (N_11450,N_11171,N_10997);
nor U11451 (N_11451,N_11147,N_10811);
nor U11452 (N_11452,N_11218,N_10641);
xnor U11453 (N_11453,N_10634,N_10176);
nor U11454 (N_11454,N_10361,N_10792);
xor U11455 (N_11455,N_10561,N_10451);
or U11456 (N_11456,N_10750,N_10748);
nand U11457 (N_11457,N_11065,N_10842);
nor U11458 (N_11458,N_10754,N_10653);
and U11459 (N_11459,N_11096,N_10396);
nand U11460 (N_11460,N_10620,N_10828);
nor U11461 (N_11461,N_10122,N_11173);
nand U11462 (N_11462,N_10735,N_11091);
or U11463 (N_11463,N_11142,N_10430);
nand U11464 (N_11464,N_10558,N_10651);
nor U11465 (N_11465,N_11043,N_10486);
nor U11466 (N_11466,N_11232,N_10867);
xnor U11467 (N_11467,N_10912,N_10210);
xnor U11468 (N_11468,N_10592,N_11025);
nand U11469 (N_11469,N_10082,N_10511);
nand U11470 (N_11470,N_10043,N_10103);
nand U11471 (N_11471,N_10414,N_10448);
nand U11472 (N_11472,N_11154,N_10167);
nand U11473 (N_11473,N_11226,N_10576);
nand U11474 (N_11474,N_10485,N_10050);
or U11475 (N_11475,N_10616,N_10113);
nand U11476 (N_11476,N_10966,N_11155);
nor U11477 (N_11477,N_10204,N_11128);
nor U11478 (N_11478,N_11108,N_11052);
nand U11479 (N_11479,N_10869,N_10259);
and U11480 (N_11480,N_10781,N_10896);
nand U11481 (N_11481,N_10534,N_10286);
nand U11482 (N_11482,N_10034,N_10797);
xnor U11483 (N_11483,N_10953,N_11180);
and U11484 (N_11484,N_10209,N_10695);
or U11485 (N_11485,N_10820,N_10093);
xor U11486 (N_11486,N_11175,N_10405);
xnor U11487 (N_11487,N_11223,N_10713);
xnor U11488 (N_11488,N_10354,N_10083);
xnor U11489 (N_11489,N_10670,N_10692);
xor U11490 (N_11490,N_10264,N_10959);
and U11491 (N_11491,N_10197,N_10952);
or U11492 (N_11492,N_10525,N_10282);
nor U11493 (N_11493,N_10637,N_11116);
nor U11494 (N_11494,N_10300,N_10835);
or U11495 (N_11495,N_10676,N_10270);
nand U11496 (N_11496,N_10833,N_10619);
and U11497 (N_11497,N_10819,N_10280);
and U11498 (N_11498,N_10150,N_10391);
xor U11499 (N_11499,N_10856,N_10623);
or U11500 (N_11500,N_10091,N_10400);
and U11501 (N_11501,N_10202,N_10823);
and U11502 (N_11502,N_10118,N_10393);
nor U11503 (N_11503,N_10505,N_10028);
or U11504 (N_11504,N_10080,N_10773);
nor U11505 (N_11505,N_10591,N_10298);
xor U11506 (N_11506,N_10989,N_10594);
xor U11507 (N_11507,N_10372,N_10060);
and U11508 (N_11508,N_10330,N_10097);
xnor U11509 (N_11509,N_10610,N_11024);
and U11510 (N_11510,N_10747,N_10764);
or U11511 (N_11511,N_10816,N_10243);
nand U11512 (N_11512,N_10757,N_11050);
nand U11513 (N_11513,N_11196,N_10902);
or U11514 (N_11514,N_10077,N_10921);
nor U11515 (N_11515,N_10135,N_10710);
nor U11516 (N_11516,N_10892,N_10323);
nor U11517 (N_11517,N_10662,N_10213);
or U11518 (N_11518,N_10654,N_10183);
nor U11519 (N_11519,N_10681,N_10130);
nand U11520 (N_11520,N_10107,N_10618);
xnor U11521 (N_11521,N_10753,N_10287);
xnor U11522 (N_11522,N_11051,N_10343);
xor U11523 (N_11523,N_11073,N_10697);
xor U11524 (N_11524,N_10854,N_10490);
or U11525 (N_11525,N_10656,N_10109);
or U11526 (N_11526,N_10971,N_10419);
nand U11527 (N_11527,N_10375,N_11039);
nand U11528 (N_11528,N_11085,N_10166);
and U11529 (N_11529,N_10872,N_10873);
nor U11530 (N_11530,N_10774,N_10807);
or U11531 (N_11531,N_10977,N_10459);
and U11532 (N_11532,N_10607,N_10409);
or U11533 (N_11533,N_10712,N_10611);
and U11534 (N_11534,N_10138,N_11044);
xnor U11535 (N_11535,N_10328,N_10033);
or U11536 (N_11536,N_11029,N_10322);
and U11537 (N_11537,N_10013,N_10965);
and U11538 (N_11538,N_11033,N_10529);
or U11539 (N_11539,N_10929,N_10805);
and U11540 (N_11540,N_11111,N_10577);
xnor U11541 (N_11541,N_10378,N_10040);
nand U11542 (N_11542,N_11008,N_10702);
nand U11543 (N_11543,N_10917,N_10694);
nand U11544 (N_11544,N_10208,N_11120);
xor U11545 (N_11545,N_10200,N_10910);
or U11546 (N_11546,N_11214,N_10446);
nand U11547 (N_11547,N_10269,N_10779);
xor U11548 (N_11548,N_10426,N_10164);
nor U11549 (N_11549,N_10780,N_10068);
nor U11550 (N_11550,N_10859,N_10880);
or U11551 (N_11551,N_10582,N_10234);
nand U11552 (N_11552,N_10242,N_10940);
or U11553 (N_11553,N_11238,N_10699);
and U11554 (N_11554,N_11004,N_10782);
and U11555 (N_11555,N_11207,N_10148);
nand U11556 (N_11556,N_10029,N_10096);
or U11557 (N_11557,N_10601,N_10434);
or U11558 (N_11558,N_10855,N_10256);
nand U11559 (N_11559,N_10112,N_10539);
nor U11560 (N_11560,N_10108,N_10356);
or U11561 (N_11561,N_10010,N_10042);
xnor U11562 (N_11562,N_10052,N_10332);
and U11563 (N_11563,N_10273,N_11231);
nor U11564 (N_11564,N_10743,N_10431);
xor U11565 (N_11565,N_10199,N_10665);
or U11566 (N_11566,N_10005,N_10734);
or U11567 (N_11567,N_10874,N_11031);
and U11568 (N_11568,N_10716,N_10516);
and U11569 (N_11569,N_10278,N_11136);
and U11570 (N_11570,N_10351,N_10969);
xnor U11571 (N_11571,N_10636,N_10648);
xor U11572 (N_11572,N_10978,N_10055);
and U11573 (N_11573,N_10628,N_10933);
and U11574 (N_11574,N_10066,N_10321);
and U11575 (N_11575,N_10228,N_11049);
nor U11576 (N_11576,N_10983,N_11152);
or U11577 (N_11577,N_10374,N_10507);
or U11578 (N_11578,N_11203,N_10172);
nor U11579 (N_11579,N_10613,N_10087);
nor U11580 (N_11580,N_10206,N_10215);
and U11581 (N_11581,N_10897,N_11204);
or U11582 (N_11582,N_11188,N_10008);
xor U11583 (N_11583,N_10932,N_10655);
nand U11584 (N_11584,N_10975,N_10844);
or U11585 (N_11585,N_10203,N_10494);
nand U11586 (N_11586,N_10478,N_10759);
or U11587 (N_11587,N_11099,N_10145);
nor U11588 (N_11588,N_10991,N_10009);
or U11589 (N_11589,N_10049,N_11084);
xnor U11590 (N_11590,N_10579,N_11125);
xnor U11591 (N_11591,N_10196,N_11242);
nor U11592 (N_11592,N_10182,N_11109);
or U11593 (N_11593,N_11061,N_10746);
or U11594 (N_11594,N_11148,N_10967);
xor U11595 (N_11595,N_11110,N_10266);
nand U11596 (N_11596,N_10536,N_10394);
nand U11597 (N_11597,N_10909,N_10480);
and U11598 (N_11598,N_11227,N_11168);
xor U11599 (N_11599,N_10786,N_10847);
nor U11600 (N_11600,N_10464,N_11133);
or U11601 (N_11601,N_10889,N_10362);
and U11602 (N_11602,N_11080,N_10227);
and U11603 (N_11603,N_10241,N_11087);
xnor U11604 (N_11604,N_10506,N_10861);
and U11605 (N_11605,N_11177,N_10011);
or U11606 (N_11606,N_10914,N_10884);
xor U11607 (N_11607,N_10303,N_10114);
nand U11608 (N_11608,N_10894,N_10958);
or U11609 (N_11609,N_10169,N_10326);
nor U11610 (N_11610,N_10472,N_10039);
nand U11611 (N_11611,N_10154,N_10540);
and U11612 (N_11612,N_10437,N_10194);
or U11613 (N_11613,N_11113,N_11077);
or U11614 (N_11614,N_10726,N_10992);
nand U11615 (N_11615,N_10964,N_10768);
nor U11616 (N_11616,N_10371,N_10070);
and U11617 (N_11617,N_11241,N_10790);
xnor U11618 (N_11618,N_11206,N_11178);
nor U11619 (N_11619,N_11197,N_10143);
xnor U11620 (N_11620,N_10886,N_10382);
nand U11621 (N_11621,N_10508,N_10260);
nor U11622 (N_11622,N_10094,N_10185);
xor U11623 (N_11623,N_10578,N_10239);
or U11624 (N_11624,N_10765,N_10477);
xor U11625 (N_11625,N_10650,N_11103);
nor U11626 (N_11626,N_10415,N_10250);
nand U11627 (N_11627,N_10568,N_10205);
and U11628 (N_11628,N_10570,N_10761);
or U11629 (N_11629,N_10045,N_10484);
and U11630 (N_11630,N_10025,N_10575);
or U11631 (N_11631,N_10198,N_11212);
xnor U11632 (N_11632,N_10353,N_10131);
nor U11633 (N_11633,N_10542,N_10418);
or U11634 (N_11634,N_10925,N_10789);
or U11635 (N_11635,N_11165,N_10193);
xor U11636 (N_11636,N_10763,N_10365);
xnor U11637 (N_11637,N_10425,N_10675);
nand U11638 (N_11638,N_11164,N_10899);
xnor U11639 (N_11639,N_10519,N_10987);
nor U11640 (N_11640,N_11117,N_10022);
or U11641 (N_11641,N_10274,N_10288);
nor U11642 (N_11642,N_10120,N_11037);
xor U11643 (N_11643,N_10755,N_11174);
or U11644 (N_11644,N_10606,N_10089);
nand U11645 (N_11645,N_10701,N_10026);
nand U11646 (N_11646,N_10707,N_10559);
or U11647 (N_11647,N_10465,N_10175);
or U11648 (N_11648,N_10360,N_10106);
nor U11649 (N_11649,N_10253,N_10302);
xor U11650 (N_11650,N_10642,N_11001);
nand U11651 (N_11651,N_10839,N_10267);
or U11652 (N_11652,N_10314,N_10640);
xnor U11653 (N_11653,N_10461,N_10071);
nor U11654 (N_11654,N_10454,N_10165);
and U11655 (N_11655,N_10345,N_10898);
xnor U11656 (N_11656,N_10178,N_10455);
nor U11657 (N_11657,N_10900,N_10016);
nand U11658 (N_11658,N_10689,N_11184);
nand U11659 (N_11659,N_10671,N_10804);
xor U11660 (N_11660,N_11225,N_10715);
xnor U11661 (N_11661,N_10906,N_10292);
and U11662 (N_11662,N_10147,N_11092);
nor U11663 (N_11663,N_10388,N_10329);
nand U11664 (N_11664,N_10905,N_10018);
and U11665 (N_11665,N_10470,N_10584);
nor U11666 (N_11666,N_10903,N_10272);
and U11667 (N_11667,N_10801,N_10738);
xor U11668 (N_11668,N_10730,N_11190);
xor U11669 (N_11669,N_10230,N_10218);
xor U11670 (N_11670,N_10110,N_10155);
xnor U11671 (N_11671,N_11182,N_10499);
nand U11672 (N_11672,N_10116,N_10317);
xnor U11673 (N_11673,N_10247,N_10857);
or U11674 (N_11674,N_11230,N_10104);
nor U11675 (N_11675,N_10072,N_10564);
or U11676 (N_11676,N_11009,N_11194);
and U11677 (N_11677,N_11215,N_10980);
nor U11678 (N_11678,N_10973,N_10680);
nor U11679 (N_11679,N_10799,N_11047);
xnor U11680 (N_11680,N_10211,N_10567);
xor U11681 (N_11681,N_11094,N_10673);
and U11682 (N_11682,N_10986,N_10325);
or U11683 (N_11683,N_10471,N_10383);
nor U11684 (N_11684,N_10258,N_10876);
nor U11685 (N_11685,N_10324,N_10979);
nand U11686 (N_11686,N_10336,N_11137);
or U11687 (N_11687,N_10297,N_10309);
nand U11688 (N_11688,N_10566,N_10806);
and U11689 (N_11689,N_10825,N_10696);
or U11690 (N_11690,N_10136,N_10355);
nor U11691 (N_11691,N_10834,N_10836);
nor U11692 (N_11692,N_11189,N_10144);
nand U11693 (N_11693,N_11090,N_10523);
nor U11694 (N_11694,N_10526,N_10703);
nor U11695 (N_11695,N_11236,N_10532);
nor U11696 (N_11696,N_10685,N_11072);
and U11697 (N_11697,N_10879,N_11145);
xnor U11698 (N_11698,N_10460,N_10469);
or U11699 (N_11699,N_10719,N_11166);
nand U11700 (N_11700,N_10134,N_10463);
and U11701 (N_11701,N_10456,N_11208);
nor U11702 (N_11702,N_10453,N_10829);
and U11703 (N_11703,N_10123,N_10099);
xnor U11704 (N_11704,N_10263,N_10793);
xor U11705 (N_11705,N_10268,N_10442);
or U11706 (N_11706,N_10223,N_11191);
xor U11707 (N_11707,N_11030,N_10015);
nand U11708 (N_11708,N_10963,N_11235);
xnor U11709 (N_11709,N_10950,N_10762);
or U11710 (N_11710,N_10588,N_11070);
or U11711 (N_11711,N_10054,N_10881);
nor U11712 (N_11712,N_10408,N_11146);
xor U11713 (N_11713,N_10380,N_10661);
nor U11714 (N_11714,N_10766,N_10186);
xor U11715 (N_11715,N_10698,N_10772);
nor U11716 (N_11716,N_10331,N_10352);
nor U11717 (N_11717,N_10908,N_10852);
xor U11718 (N_11718,N_10058,N_10682);
or U11719 (N_11719,N_10882,N_10756);
nor U11720 (N_11720,N_11209,N_10137);
nor U11721 (N_11721,N_10257,N_10428);
xor U11722 (N_11722,N_10177,N_10473);
and U11723 (N_11723,N_10236,N_10489);
and U11724 (N_11724,N_10509,N_10528);
and U11725 (N_11725,N_10095,N_10188);
nor U11726 (N_11726,N_10544,N_10586);
and U11727 (N_11727,N_11119,N_11132);
xor U11728 (N_11728,N_10803,N_10057);
or U11729 (N_11729,N_10550,N_10944);
or U11730 (N_11730,N_10770,N_10614);
nor U11731 (N_11731,N_11220,N_11124);
xnor U11732 (N_11732,N_10417,N_10920);
nor U11733 (N_11733,N_10366,N_11150);
and U11734 (N_11734,N_10275,N_10664);
xor U11735 (N_11735,N_10347,N_10126);
nand U11736 (N_11736,N_10067,N_10276);
xor U11737 (N_11737,N_11000,N_10252);
nor U11738 (N_11738,N_11042,N_11056);
xnor U11739 (N_11739,N_10609,N_10141);
xnor U11740 (N_11740,N_11249,N_10831);
nor U11741 (N_11741,N_10435,N_10438);
nand U11742 (N_11742,N_10254,N_10370);
xor U11743 (N_11743,N_11075,N_11101);
or U11744 (N_11744,N_10413,N_10310);
xnor U11745 (N_11745,N_11007,N_10161);
and U11746 (N_11746,N_10758,N_10000);
or U11747 (N_11747,N_11246,N_11046);
xnor U11748 (N_11748,N_10604,N_10938);
nand U11749 (N_11749,N_10948,N_10406);
nand U11750 (N_11750,N_10344,N_10838);
and U11751 (N_11751,N_11112,N_11183);
nand U11752 (N_11752,N_11202,N_10918);
and U11753 (N_11753,N_10339,N_10085);
nor U11754 (N_11754,N_10956,N_10457);
and U11755 (N_11755,N_10357,N_10142);
and U11756 (N_11756,N_10865,N_10216);
nand U11757 (N_11757,N_11107,N_11234);
nand U11758 (N_11758,N_11079,N_11224);
nand U11759 (N_11759,N_10482,N_10794);
nand U11760 (N_11760,N_10475,N_10004);
or U11761 (N_11761,N_10318,N_10214);
nand U11762 (N_11762,N_10517,N_10474);
and U11763 (N_11763,N_10657,N_10027);
and U11764 (N_11764,N_10295,N_10659);
and U11765 (N_11765,N_10885,N_10545);
or U11766 (N_11766,N_11233,N_10289);
xnor U11767 (N_11767,N_10736,N_10574);
xor U11768 (N_11768,N_11140,N_10541);
and U11769 (N_11769,N_10866,N_10632);
nor U11770 (N_11770,N_10878,N_10334);
nand U11771 (N_11771,N_10261,N_10552);
and U11772 (N_11772,N_10220,N_11219);
nand U11773 (N_11773,N_10497,N_10389);
and U11774 (N_11774,N_10488,N_10479);
nand U11775 (N_11775,N_10047,N_10700);
and U11776 (N_11776,N_10672,N_11248);
nor U11777 (N_11777,N_10802,N_11126);
and U11778 (N_11778,N_10875,N_10724);
xnor U11779 (N_11779,N_10646,N_10547);
nor U11780 (N_11780,N_10265,N_10510);
or U11781 (N_11781,N_11022,N_10038);
and U11782 (N_11782,N_10090,N_10100);
or U11783 (N_11783,N_10737,N_10615);
nand U11784 (N_11784,N_11121,N_10299);
nor U11785 (N_11785,N_10663,N_10674);
xnor U11786 (N_11786,N_10348,N_10693);
and U11787 (N_11787,N_10195,N_10392);
nand U11788 (N_11788,N_10581,N_10281);
xor U11789 (N_11789,N_10219,N_10597);
or U11790 (N_11790,N_10333,N_10238);
xnor U11791 (N_11791,N_10064,N_10994);
nand U11792 (N_11792,N_10785,N_10081);
nor U11793 (N_11793,N_11170,N_11187);
and U11794 (N_11794,N_10132,N_11141);
or U11795 (N_11795,N_10304,N_10384);
or U11796 (N_11796,N_10767,N_10669);
nand U11797 (N_11797,N_10845,N_11216);
nor U11798 (N_11798,N_11088,N_11010);
nor U11799 (N_11799,N_11228,N_10284);
nor U11800 (N_11800,N_10410,N_10923);
nand U11801 (N_11801,N_10390,N_10739);
nand U11802 (N_11802,N_10533,N_11222);
xor U11803 (N_11803,N_11066,N_10404);
nor U11804 (N_11804,N_10429,N_10853);
nand U11805 (N_11805,N_10783,N_10036);
or U11806 (N_11806,N_10937,N_10600);
or U11807 (N_11807,N_10945,N_11063);
or U11808 (N_11808,N_10271,N_10503);
nor U11809 (N_11809,N_10279,N_10771);
or U11810 (N_11810,N_10922,N_10377);
or U11811 (N_11811,N_10262,N_10341);
xnor U11812 (N_11812,N_10832,N_11083);
nor U11813 (N_11813,N_10319,N_10931);
and U11814 (N_11814,N_10629,N_10970);
nor U11815 (N_11815,N_10518,N_10627);
or U11816 (N_11816,N_10621,N_11034);
nor U11817 (N_11817,N_10936,N_10851);
or U11818 (N_11818,N_11069,N_10514);
and U11819 (N_11819,N_10891,N_10683);
xor U11820 (N_11820,N_10233,N_10059);
or U11821 (N_11821,N_10691,N_10725);
or U11822 (N_11822,N_10062,N_10981);
and U11823 (N_11823,N_10515,N_10826);
and U11824 (N_11824,N_10531,N_10954);
and U11825 (N_11825,N_10744,N_11028);
nor U11826 (N_11826,N_10466,N_11135);
and U11827 (N_11827,N_10927,N_10231);
nor U11828 (N_11828,N_10530,N_10947);
or U11829 (N_11829,N_11118,N_10385);
xnor U11830 (N_11830,N_10290,N_10598);
and U11831 (N_11831,N_11198,N_11176);
xor U11832 (N_11832,N_10379,N_10450);
xor U11833 (N_11833,N_10824,N_10296);
xor U11834 (N_11834,N_10813,N_10871);
or U11835 (N_11835,N_10222,N_10643);
nand U11836 (N_11836,N_11138,N_10635);
xor U11837 (N_11837,N_10982,N_10590);
nor U11838 (N_11838,N_10554,N_10778);
xor U11839 (N_11839,N_10031,N_10293);
or U11840 (N_11840,N_10625,N_10399);
nand U11841 (N_11841,N_10603,N_10863);
nand U11842 (N_11842,N_10815,N_10452);
xnor U11843 (N_11843,N_10291,N_10985);
or U11844 (N_11844,N_10358,N_10538);
nor U11845 (N_11845,N_11130,N_10051);
xor U11846 (N_11846,N_10705,N_10111);
nand U11847 (N_11847,N_11020,N_10649);
nor U11848 (N_11848,N_11074,N_11193);
nand U11849 (N_11849,N_10941,N_10249);
or U11850 (N_11850,N_10181,N_11163);
nand U11851 (N_11851,N_11054,N_10207);
nand U11852 (N_11852,N_10376,N_10226);
or U11853 (N_11853,N_10283,N_10688);
xnor U11854 (N_11854,N_10160,N_11114);
nor U11855 (N_11855,N_10827,N_10957);
nor U11856 (N_11856,N_11013,N_10075);
and U11857 (N_11857,N_10048,N_11200);
nor U11858 (N_11858,N_10549,N_10046);
nor U11859 (N_11859,N_10192,N_10162);
and U11860 (N_11860,N_10491,N_10512);
xnor U11861 (N_11861,N_10201,N_10677);
nor U11862 (N_11862,N_10608,N_10795);
nor U11863 (N_11863,N_10156,N_10327);
nor U11864 (N_11864,N_10368,N_10335);
and U11865 (N_11865,N_11211,N_10617);
xor U11866 (N_11866,N_10521,N_11139);
xor U11867 (N_11867,N_10398,N_10930);
xnor U11868 (N_11868,N_10306,N_10660);
nand U11869 (N_11869,N_10079,N_11095);
xnor U11870 (N_11870,N_10153,N_10817);
xnor U11871 (N_11871,N_11210,N_10316);
nand U11872 (N_11872,N_10858,N_11151);
nand U11873 (N_11873,N_10916,N_10843);
nor U11874 (N_11874,N_11134,N_11115);
nor U11875 (N_11875,N_10607,N_11106);
or U11876 (N_11876,N_10649,N_10900);
and U11877 (N_11877,N_10440,N_11158);
or U11878 (N_11878,N_10237,N_10051);
nand U11879 (N_11879,N_10447,N_11134);
nand U11880 (N_11880,N_10485,N_10331);
or U11881 (N_11881,N_10314,N_10634);
or U11882 (N_11882,N_10926,N_10110);
nand U11883 (N_11883,N_11065,N_10610);
and U11884 (N_11884,N_10467,N_10514);
or U11885 (N_11885,N_10411,N_10712);
xor U11886 (N_11886,N_10756,N_10527);
and U11887 (N_11887,N_10644,N_10518);
xor U11888 (N_11888,N_10722,N_10094);
xor U11889 (N_11889,N_10382,N_11190);
xor U11890 (N_11890,N_10896,N_10454);
or U11891 (N_11891,N_10374,N_10752);
and U11892 (N_11892,N_10206,N_10027);
and U11893 (N_11893,N_10694,N_10771);
nand U11894 (N_11894,N_10469,N_10203);
xor U11895 (N_11895,N_10380,N_10852);
and U11896 (N_11896,N_10756,N_10472);
nand U11897 (N_11897,N_10775,N_10310);
and U11898 (N_11898,N_10785,N_10915);
nor U11899 (N_11899,N_10106,N_10556);
nor U11900 (N_11900,N_10879,N_11001);
xnor U11901 (N_11901,N_10659,N_10463);
xnor U11902 (N_11902,N_10110,N_10868);
nor U11903 (N_11903,N_10711,N_10938);
and U11904 (N_11904,N_10062,N_10571);
xor U11905 (N_11905,N_10352,N_10573);
nand U11906 (N_11906,N_10341,N_10233);
nor U11907 (N_11907,N_10812,N_10073);
nor U11908 (N_11908,N_10282,N_10210);
nand U11909 (N_11909,N_10831,N_10941);
and U11910 (N_11910,N_10726,N_11079);
and U11911 (N_11911,N_10967,N_11140);
nor U11912 (N_11912,N_11235,N_10980);
nand U11913 (N_11913,N_10798,N_10409);
and U11914 (N_11914,N_10906,N_10497);
nand U11915 (N_11915,N_10236,N_11234);
or U11916 (N_11916,N_10914,N_10963);
nor U11917 (N_11917,N_10189,N_11096);
nor U11918 (N_11918,N_10317,N_10440);
and U11919 (N_11919,N_11151,N_11184);
xor U11920 (N_11920,N_10544,N_10995);
nand U11921 (N_11921,N_10448,N_10214);
and U11922 (N_11922,N_10722,N_11210);
and U11923 (N_11923,N_10460,N_11187);
or U11924 (N_11924,N_10141,N_10336);
nand U11925 (N_11925,N_10094,N_10926);
nand U11926 (N_11926,N_10819,N_11136);
or U11927 (N_11927,N_10436,N_11172);
or U11928 (N_11928,N_11172,N_10528);
xnor U11929 (N_11929,N_10328,N_10362);
nand U11930 (N_11930,N_10251,N_10793);
nor U11931 (N_11931,N_10563,N_11158);
and U11932 (N_11932,N_11195,N_10922);
nand U11933 (N_11933,N_10591,N_10819);
xor U11934 (N_11934,N_10508,N_11043);
and U11935 (N_11935,N_10289,N_10161);
or U11936 (N_11936,N_11131,N_10191);
or U11937 (N_11937,N_10275,N_10193);
xnor U11938 (N_11938,N_10910,N_10613);
xor U11939 (N_11939,N_11060,N_10197);
nor U11940 (N_11940,N_10651,N_10435);
xor U11941 (N_11941,N_10765,N_10270);
and U11942 (N_11942,N_10873,N_10136);
xnor U11943 (N_11943,N_10933,N_11118);
nor U11944 (N_11944,N_10148,N_10699);
and U11945 (N_11945,N_10186,N_10791);
and U11946 (N_11946,N_10114,N_10622);
xnor U11947 (N_11947,N_10394,N_10325);
and U11948 (N_11948,N_10933,N_10518);
and U11949 (N_11949,N_10840,N_10507);
nor U11950 (N_11950,N_10074,N_10606);
xor U11951 (N_11951,N_10733,N_11131);
nor U11952 (N_11952,N_10995,N_10892);
nand U11953 (N_11953,N_10674,N_10798);
nand U11954 (N_11954,N_10400,N_10431);
nand U11955 (N_11955,N_10973,N_10247);
nor U11956 (N_11956,N_10016,N_10102);
nand U11957 (N_11957,N_10822,N_10359);
or U11958 (N_11958,N_10346,N_11010);
nor U11959 (N_11959,N_10844,N_10225);
nand U11960 (N_11960,N_11126,N_10192);
nor U11961 (N_11961,N_10892,N_11183);
and U11962 (N_11962,N_10748,N_10342);
nand U11963 (N_11963,N_10463,N_11103);
or U11964 (N_11964,N_11222,N_10625);
or U11965 (N_11965,N_10502,N_10659);
nor U11966 (N_11966,N_11027,N_10021);
xnor U11967 (N_11967,N_10831,N_10004);
and U11968 (N_11968,N_10183,N_10850);
nand U11969 (N_11969,N_10855,N_10898);
nand U11970 (N_11970,N_11222,N_11143);
nand U11971 (N_11971,N_10205,N_10636);
and U11972 (N_11972,N_11132,N_10904);
or U11973 (N_11973,N_10437,N_11231);
and U11974 (N_11974,N_10175,N_10289);
nor U11975 (N_11975,N_10002,N_11183);
xor U11976 (N_11976,N_10459,N_10912);
or U11977 (N_11977,N_10761,N_11238);
xnor U11978 (N_11978,N_10943,N_10511);
or U11979 (N_11979,N_10556,N_10530);
xor U11980 (N_11980,N_10698,N_10373);
or U11981 (N_11981,N_11019,N_10174);
xnor U11982 (N_11982,N_10828,N_10123);
and U11983 (N_11983,N_10643,N_11221);
nor U11984 (N_11984,N_11087,N_10530);
and U11985 (N_11985,N_10136,N_10439);
xnor U11986 (N_11986,N_11182,N_10743);
and U11987 (N_11987,N_10816,N_10754);
nand U11988 (N_11988,N_10274,N_11113);
nand U11989 (N_11989,N_10145,N_10592);
and U11990 (N_11990,N_11192,N_10115);
nand U11991 (N_11991,N_11139,N_10351);
xor U11992 (N_11992,N_11079,N_10385);
or U11993 (N_11993,N_10591,N_10939);
nand U11994 (N_11994,N_10068,N_10943);
nand U11995 (N_11995,N_10817,N_10845);
xor U11996 (N_11996,N_10277,N_10454);
xnor U11997 (N_11997,N_11220,N_10084);
nand U11998 (N_11998,N_10149,N_10223);
nand U11999 (N_11999,N_10987,N_10646);
and U12000 (N_12000,N_10672,N_10557);
or U12001 (N_12001,N_10305,N_10848);
xnor U12002 (N_12002,N_10443,N_10638);
and U12003 (N_12003,N_10457,N_10040);
xor U12004 (N_12004,N_10121,N_10172);
or U12005 (N_12005,N_10606,N_10923);
nor U12006 (N_12006,N_10629,N_10384);
nand U12007 (N_12007,N_11209,N_10894);
nand U12008 (N_12008,N_10108,N_10935);
nor U12009 (N_12009,N_10521,N_10442);
nand U12010 (N_12010,N_10838,N_10357);
and U12011 (N_12011,N_10616,N_10293);
nand U12012 (N_12012,N_10325,N_10565);
and U12013 (N_12013,N_10698,N_10129);
nand U12014 (N_12014,N_10732,N_10175);
and U12015 (N_12015,N_10248,N_10908);
nor U12016 (N_12016,N_10706,N_10735);
and U12017 (N_12017,N_10508,N_10535);
or U12018 (N_12018,N_10855,N_10148);
xor U12019 (N_12019,N_10693,N_10768);
nor U12020 (N_12020,N_10758,N_10495);
and U12021 (N_12021,N_10693,N_10971);
nand U12022 (N_12022,N_10189,N_10252);
nand U12023 (N_12023,N_10273,N_11212);
or U12024 (N_12024,N_10460,N_10531);
nand U12025 (N_12025,N_11219,N_10219);
nand U12026 (N_12026,N_10057,N_10570);
and U12027 (N_12027,N_10657,N_10391);
nor U12028 (N_12028,N_11029,N_10495);
nand U12029 (N_12029,N_10473,N_10933);
or U12030 (N_12030,N_10456,N_11223);
or U12031 (N_12031,N_10033,N_10508);
xor U12032 (N_12032,N_10518,N_11014);
xor U12033 (N_12033,N_10888,N_10206);
and U12034 (N_12034,N_10215,N_10285);
xnor U12035 (N_12035,N_10753,N_10126);
nor U12036 (N_12036,N_10187,N_10889);
or U12037 (N_12037,N_10599,N_11200);
xnor U12038 (N_12038,N_10850,N_10191);
and U12039 (N_12039,N_10290,N_11071);
nand U12040 (N_12040,N_10259,N_10358);
nand U12041 (N_12041,N_10551,N_10436);
xnor U12042 (N_12042,N_11110,N_10901);
or U12043 (N_12043,N_10641,N_10629);
xor U12044 (N_12044,N_10990,N_11149);
nor U12045 (N_12045,N_11175,N_11036);
nand U12046 (N_12046,N_11052,N_10537);
nor U12047 (N_12047,N_10586,N_11185);
or U12048 (N_12048,N_10352,N_10054);
nand U12049 (N_12049,N_10976,N_10728);
nand U12050 (N_12050,N_11185,N_10050);
or U12051 (N_12051,N_10589,N_10193);
nand U12052 (N_12052,N_10536,N_11122);
nand U12053 (N_12053,N_11167,N_10878);
or U12054 (N_12054,N_10001,N_11132);
nor U12055 (N_12055,N_10210,N_11173);
xnor U12056 (N_12056,N_10202,N_10201);
xor U12057 (N_12057,N_11043,N_10296);
and U12058 (N_12058,N_11096,N_10900);
xnor U12059 (N_12059,N_10204,N_11220);
xnor U12060 (N_12060,N_10094,N_10223);
nor U12061 (N_12061,N_11079,N_10347);
nand U12062 (N_12062,N_10019,N_10789);
nand U12063 (N_12063,N_10202,N_10118);
and U12064 (N_12064,N_10092,N_10475);
and U12065 (N_12065,N_10816,N_10643);
xnor U12066 (N_12066,N_10866,N_11118);
xnor U12067 (N_12067,N_10632,N_10560);
xnor U12068 (N_12068,N_10085,N_10720);
xor U12069 (N_12069,N_10383,N_10311);
xor U12070 (N_12070,N_10938,N_10165);
nand U12071 (N_12071,N_10645,N_11082);
nor U12072 (N_12072,N_10704,N_11175);
and U12073 (N_12073,N_10192,N_10508);
or U12074 (N_12074,N_10124,N_11187);
xor U12075 (N_12075,N_10505,N_10534);
nor U12076 (N_12076,N_10405,N_10104);
nand U12077 (N_12077,N_11235,N_10404);
or U12078 (N_12078,N_10082,N_10991);
xor U12079 (N_12079,N_10058,N_10444);
or U12080 (N_12080,N_11167,N_10989);
and U12081 (N_12081,N_10499,N_10343);
and U12082 (N_12082,N_10474,N_11040);
or U12083 (N_12083,N_10092,N_10151);
nor U12084 (N_12084,N_10871,N_10475);
nand U12085 (N_12085,N_10013,N_10992);
nand U12086 (N_12086,N_10666,N_10912);
nand U12087 (N_12087,N_10338,N_10639);
or U12088 (N_12088,N_10337,N_10884);
nand U12089 (N_12089,N_10263,N_10302);
nand U12090 (N_12090,N_10538,N_10565);
xor U12091 (N_12091,N_11005,N_10215);
nand U12092 (N_12092,N_10397,N_10658);
or U12093 (N_12093,N_10042,N_10631);
nand U12094 (N_12094,N_10145,N_10482);
nor U12095 (N_12095,N_10571,N_10245);
or U12096 (N_12096,N_10969,N_10032);
and U12097 (N_12097,N_10410,N_10091);
xor U12098 (N_12098,N_10285,N_10279);
or U12099 (N_12099,N_10238,N_10407);
nand U12100 (N_12100,N_10483,N_10981);
or U12101 (N_12101,N_10963,N_10449);
and U12102 (N_12102,N_10737,N_10261);
nor U12103 (N_12103,N_10623,N_10039);
or U12104 (N_12104,N_10434,N_10767);
nand U12105 (N_12105,N_10174,N_10030);
or U12106 (N_12106,N_10781,N_10569);
or U12107 (N_12107,N_10764,N_11000);
nand U12108 (N_12108,N_10140,N_10096);
nand U12109 (N_12109,N_10866,N_10107);
nand U12110 (N_12110,N_10101,N_10301);
xor U12111 (N_12111,N_11103,N_11116);
or U12112 (N_12112,N_11042,N_10554);
nor U12113 (N_12113,N_10694,N_11022);
nor U12114 (N_12114,N_11014,N_10605);
xnor U12115 (N_12115,N_11067,N_10694);
nor U12116 (N_12116,N_11161,N_10449);
and U12117 (N_12117,N_10259,N_10346);
nor U12118 (N_12118,N_10901,N_11212);
and U12119 (N_12119,N_10182,N_10861);
nor U12120 (N_12120,N_10570,N_11040);
or U12121 (N_12121,N_10919,N_10925);
or U12122 (N_12122,N_11229,N_10591);
and U12123 (N_12123,N_10757,N_10472);
nor U12124 (N_12124,N_10023,N_11063);
xor U12125 (N_12125,N_10155,N_10575);
or U12126 (N_12126,N_10339,N_10203);
nand U12127 (N_12127,N_10758,N_11187);
xor U12128 (N_12128,N_10458,N_10954);
xor U12129 (N_12129,N_10493,N_10320);
or U12130 (N_12130,N_10741,N_11215);
xor U12131 (N_12131,N_10249,N_10736);
xnor U12132 (N_12132,N_10465,N_10384);
or U12133 (N_12133,N_11065,N_10299);
nand U12134 (N_12134,N_10450,N_10902);
or U12135 (N_12135,N_11021,N_11227);
or U12136 (N_12136,N_10240,N_10019);
nand U12137 (N_12137,N_10398,N_10406);
nor U12138 (N_12138,N_10697,N_10295);
xor U12139 (N_12139,N_10930,N_10633);
and U12140 (N_12140,N_10707,N_10633);
nand U12141 (N_12141,N_10117,N_10717);
xnor U12142 (N_12142,N_10861,N_11013);
xor U12143 (N_12143,N_11045,N_11053);
and U12144 (N_12144,N_10218,N_10581);
or U12145 (N_12145,N_10438,N_10038);
nand U12146 (N_12146,N_10992,N_10818);
nand U12147 (N_12147,N_10265,N_10744);
nor U12148 (N_12148,N_10555,N_10617);
nand U12149 (N_12149,N_10951,N_10363);
xor U12150 (N_12150,N_10540,N_10496);
nor U12151 (N_12151,N_11210,N_10098);
nor U12152 (N_12152,N_10448,N_10502);
or U12153 (N_12153,N_10430,N_11113);
xor U12154 (N_12154,N_10435,N_11088);
xnor U12155 (N_12155,N_10420,N_10484);
nand U12156 (N_12156,N_10748,N_10559);
and U12157 (N_12157,N_10986,N_11058);
nor U12158 (N_12158,N_10483,N_10546);
or U12159 (N_12159,N_10976,N_11007);
nand U12160 (N_12160,N_11028,N_10108);
or U12161 (N_12161,N_10111,N_11146);
and U12162 (N_12162,N_10973,N_10443);
nor U12163 (N_12163,N_10876,N_10536);
nand U12164 (N_12164,N_10121,N_10342);
nand U12165 (N_12165,N_10814,N_11155);
and U12166 (N_12166,N_10977,N_10401);
nor U12167 (N_12167,N_10420,N_10510);
xor U12168 (N_12168,N_10967,N_10682);
nor U12169 (N_12169,N_10640,N_10822);
nand U12170 (N_12170,N_10348,N_10088);
and U12171 (N_12171,N_10953,N_10937);
nand U12172 (N_12172,N_10738,N_10441);
or U12173 (N_12173,N_10813,N_11140);
and U12174 (N_12174,N_10393,N_10340);
nand U12175 (N_12175,N_10508,N_10308);
nor U12176 (N_12176,N_11177,N_10641);
or U12177 (N_12177,N_10233,N_11109);
and U12178 (N_12178,N_10716,N_10900);
or U12179 (N_12179,N_10374,N_10334);
and U12180 (N_12180,N_10372,N_10862);
nor U12181 (N_12181,N_10799,N_10206);
nor U12182 (N_12182,N_10606,N_10912);
nand U12183 (N_12183,N_10699,N_10475);
xnor U12184 (N_12184,N_10285,N_10305);
or U12185 (N_12185,N_10620,N_10816);
or U12186 (N_12186,N_11232,N_11066);
xnor U12187 (N_12187,N_10611,N_10553);
or U12188 (N_12188,N_10030,N_10345);
xor U12189 (N_12189,N_11035,N_10248);
nand U12190 (N_12190,N_10864,N_10602);
or U12191 (N_12191,N_10305,N_10423);
nand U12192 (N_12192,N_10748,N_10842);
xor U12193 (N_12193,N_10413,N_11012);
nand U12194 (N_12194,N_11133,N_10658);
nand U12195 (N_12195,N_11246,N_10607);
nand U12196 (N_12196,N_10872,N_10959);
xor U12197 (N_12197,N_10913,N_10004);
xnor U12198 (N_12198,N_10616,N_10829);
xor U12199 (N_12199,N_10570,N_11045);
nand U12200 (N_12200,N_10802,N_11085);
xor U12201 (N_12201,N_10586,N_10841);
xor U12202 (N_12202,N_10760,N_10475);
and U12203 (N_12203,N_10315,N_10710);
nor U12204 (N_12204,N_10687,N_10817);
nand U12205 (N_12205,N_10676,N_10410);
xnor U12206 (N_12206,N_10030,N_10144);
xnor U12207 (N_12207,N_10473,N_10304);
nand U12208 (N_12208,N_10078,N_10497);
or U12209 (N_12209,N_10435,N_11105);
and U12210 (N_12210,N_10692,N_10351);
nand U12211 (N_12211,N_10656,N_11049);
nand U12212 (N_12212,N_10739,N_11003);
and U12213 (N_12213,N_10997,N_11125);
nand U12214 (N_12214,N_10892,N_10260);
xor U12215 (N_12215,N_10185,N_10630);
nor U12216 (N_12216,N_10215,N_10090);
xor U12217 (N_12217,N_10264,N_10756);
or U12218 (N_12218,N_10399,N_10428);
nor U12219 (N_12219,N_10097,N_10266);
and U12220 (N_12220,N_11021,N_10753);
or U12221 (N_12221,N_11233,N_11248);
nor U12222 (N_12222,N_10097,N_11128);
and U12223 (N_12223,N_10035,N_11179);
or U12224 (N_12224,N_10937,N_10408);
or U12225 (N_12225,N_10369,N_10190);
xnor U12226 (N_12226,N_10225,N_10192);
xor U12227 (N_12227,N_10178,N_10725);
or U12228 (N_12228,N_10643,N_11220);
nand U12229 (N_12229,N_10539,N_10602);
and U12230 (N_12230,N_10358,N_10775);
xor U12231 (N_12231,N_10574,N_10382);
and U12232 (N_12232,N_10400,N_10255);
and U12233 (N_12233,N_10731,N_10979);
nand U12234 (N_12234,N_11081,N_10516);
xor U12235 (N_12235,N_10593,N_10170);
xor U12236 (N_12236,N_10450,N_11151);
or U12237 (N_12237,N_10575,N_10773);
and U12238 (N_12238,N_10855,N_10004);
nor U12239 (N_12239,N_10335,N_10747);
and U12240 (N_12240,N_11123,N_10408);
xnor U12241 (N_12241,N_10267,N_10756);
and U12242 (N_12242,N_10271,N_10775);
xnor U12243 (N_12243,N_10399,N_11055);
nand U12244 (N_12244,N_10310,N_10277);
xnor U12245 (N_12245,N_10874,N_10274);
or U12246 (N_12246,N_11026,N_10825);
and U12247 (N_12247,N_10038,N_10817);
or U12248 (N_12248,N_10336,N_10007);
or U12249 (N_12249,N_11112,N_10951);
nor U12250 (N_12250,N_11110,N_10918);
nor U12251 (N_12251,N_11129,N_10369);
nand U12252 (N_12252,N_10158,N_11187);
and U12253 (N_12253,N_10528,N_10810);
or U12254 (N_12254,N_11127,N_10659);
xor U12255 (N_12255,N_10893,N_10635);
and U12256 (N_12256,N_10019,N_10456);
nor U12257 (N_12257,N_10172,N_10682);
xor U12258 (N_12258,N_10276,N_10230);
nor U12259 (N_12259,N_10341,N_11179);
nand U12260 (N_12260,N_10086,N_10326);
and U12261 (N_12261,N_10663,N_11055);
xor U12262 (N_12262,N_10551,N_10608);
or U12263 (N_12263,N_10997,N_10794);
xnor U12264 (N_12264,N_10621,N_10145);
and U12265 (N_12265,N_10783,N_10778);
xor U12266 (N_12266,N_10805,N_11136);
xor U12267 (N_12267,N_10260,N_10533);
or U12268 (N_12268,N_10543,N_10120);
nand U12269 (N_12269,N_10236,N_10086);
xnor U12270 (N_12270,N_10224,N_10700);
and U12271 (N_12271,N_10269,N_11137);
and U12272 (N_12272,N_10065,N_11232);
and U12273 (N_12273,N_10194,N_10244);
nor U12274 (N_12274,N_10684,N_10354);
nor U12275 (N_12275,N_10006,N_10895);
nor U12276 (N_12276,N_10766,N_10944);
xor U12277 (N_12277,N_10044,N_10494);
xnor U12278 (N_12278,N_10004,N_11182);
xnor U12279 (N_12279,N_10142,N_10653);
and U12280 (N_12280,N_10257,N_10986);
and U12281 (N_12281,N_11163,N_10394);
nand U12282 (N_12282,N_10495,N_11169);
or U12283 (N_12283,N_11167,N_11031);
nand U12284 (N_12284,N_10528,N_11069);
and U12285 (N_12285,N_10021,N_11064);
nand U12286 (N_12286,N_11012,N_10500);
nor U12287 (N_12287,N_10276,N_10028);
or U12288 (N_12288,N_11114,N_10499);
nor U12289 (N_12289,N_10471,N_11169);
nor U12290 (N_12290,N_10430,N_11006);
xnor U12291 (N_12291,N_10198,N_11184);
xor U12292 (N_12292,N_10322,N_10806);
nand U12293 (N_12293,N_11175,N_10178);
nand U12294 (N_12294,N_10097,N_10400);
or U12295 (N_12295,N_10020,N_11186);
and U12296 (N_12296,N_10022,N_11226);
or U12297 (N_12297,N_10049,N_10489);
nand U12298 (N_12298,N_10241,N_11223);
and U12299 (N_12299,N_10735,N_10531);
and U12300 (N_12300,N_10314,N_10786);
nor U12301 (N_12301,N_11024,N_10805);
nor U12302 (N_12302,N_11028,N_10900);
nor U12303 (N_12303,N_10148,N_11200);
nand U12304 (N_12304,N_10623,N_10841);
nand U12305 (N_12305,N_10072,N_11064);
xnor U12306 (N_12306,N_11145,N_10481);
nor U12307 (N_12307,N_10123,N_10307);
xnor U12308 (N_12308,N_10825,N_10662);
nand U12309 (N_12309,N_10766,N_10416);
and U12310 (N_12310,N_10675,N_11225);
nor U12311 (N_12311,N_10008,N_10182);
nor U12312 (N_12312,N_10548,N_11198);
nor U12313 (N_12313,N_10101,N_10926);
xnor U12314 (N_12314,N_10039,N_11232);
nand U12315 (N_12315,N_10758,N_10560);
nand U12316 (N_12316,N_10640,N_10392);
or U12317 (N_12317,N_10275,N_10959);
nor U12318 (N_12318,N_10848,N_11010);
nor U12319 (N_12319,N_10464,N_11245);
or U12320 (N_12320,N_10783,N_10123);
and U12321 (N_12321,N_10599,N_11163);
xnor U12322 (N_12322,N_10247,N_10727);
xor U12323 (N_12323,N_10154,N_10956);
and U12324 (N_12324,N_11136,N_10594);
nand U12325 (N_12325,N_11078,N_11143);
or U12326 (N_12326,N_10047,N_10399);
or U12327 (N_12327,N_10149,N_10992);
nor U12328 (N_12328,N_11181,N_10990);
nor U12329 (N_12329,N_10817,N_10321);
nand U12330 (N_12330,N_10915,N_10251);
xnor U12331 (N_12331,N_10268,N_10685);
and U12332 (N_12332,N_11150,N_10477);
or U12333 (N_12333,N_10729,N_10634);
xnor U12334 (N_12334,N_10918,N_10065);
and U12335 (N_12335,N_10136,N_11235);
and U12336 (N_12336,N_10979,N_11036);
xor U12337 (N_12337,N_10587,N_10410);
or U12338 (N_12338,N_10437,N_10261);
and U12339 (N_12339,N_10124,N_11175);
nor U12340 (N_12340,N_11191,N_11204);
xnor U12341 (N_12341,N_10602,N_11005);
nor U12342 (N_12342,N_11155,N_11181);
xnor U12343 (N_12343,N_10552,N_10276);
nand U12344 (N_12344,N_11017,N_10348);
and U12345 (N_12345,N_10559,N_10957);
nor U12346 (N_12346,N_10124,N_10027);
or U12347 (N_12347,N_10580,N_10179);
nand U12348 (N_12348,N_10557,N_10520);
nand U12349 (N_12349,N_10329,N_10495);
nor U12350 (N_12350,N_10496,N_10216);
or U12351 (N_12351,N_10353,N_11016);
nor U12352 (N_12352,N_11185,N_10322);
or U12353 (N_12353,N_11199,N_10995);
and U12354 (N_12354,N_10568,N_10900);
or U12355 (N_12355,N_10160,N_10673);
or U12356 (N_12356,N_10515,N_11228);
or U12357 (N_12357,N_10982,N_11164);
xor U12358 (N_12358,N_11056,N_10042);
and U12359 (N_12359,N_10874,N_10035);
nor U12360 (N_12360,N_10109,N_11034);
nor U12361 (N_12361,N_10706,N_10093);
nor U12362 (N_12362,N_10295,N_11202);
nor U12363 (N_12363,N_10322,N_11061);
or U12364 (N_12364,N_11038,N_10255);
nand U12365 (N_12365,N_10043,N_10144);
or U12366 (N_12366,N_11037,N_11186);
nand U12367 (N_12367,N_10352,N_10659);
xnor U12368 (N_12368,N_10107,N_10277);
nor U12369 (N_12369,N_10425,N_10814);
nand U12370 (N_12370,N_10824,N_11033);
or U12371 (N_12371,N_11180,N_10192);
xor U12372 (N_12372,N_10117,N_10723);
xor U12373 (N_12373,N_10174,N_10120);
or U12374 (N_12374,N_10622,N_10860);
xor U12375 (N_12375,N_11142,N_11247);
and U12376 (N_12376,N_10502,N_10813);
and U12377 (N_12377,N_11224,N_10197);
and U12378 (N_12378,N_10398,N_11075);
xor U12379 (N_12379,N_10262,N_10301);
nand U12380 (N_12380,N_10688,N_10798);
xnor U12381 (N_12381,N_11080,N_10350);
and U12382 (N_12382,N_10961,N_10398);
xor U12383 (N_12383,N_10765,N_10543);
nor U12384 (N_12384,N_11185,N_10581);
or U12385 (N_12385,N_10089,N_10323);
and U12386 (N_12386,N_11049,N_10304);
and U12387 (N_12387,N_10577,N_11036);
xor U12388 (N_12388,N_10233,N_10004);
and U12389 (N_12389,N_10512,N_10532);
nor U12390 (N_12390,N_10741,N_10560);
nor U12391 (N_12391,N_11185,N_10099);
nor U12392 (N_12392,N_10629,N_10595);
xor U12393 (N_12393,N_10839,N_10578);
and U12394 (N_12394,N_11041,N_10924);
xnor U12395 (N_12395,N_10774,N_11103);
or U12396 (N_12396,N_10511,N_10199);
and U12397 (N_12397,N_10739,N_10617);
nand U12398 (N_12398,N_10299,N_11048);
nor U12399 (N_12399,N_11099,N_10194);
xnor U12400 (N_12400,N_10787,N_10201);
nor U12401 (N_12401,N_11018,N_10755);
and U12402 (N_12402,N_10739,N_10447);
nor U12403 (N_12403,N_10107,N_10656);
nand U12404 (N_12404,N_10681,N_10450);
nand U12405 (N_12405,N_10038,N_10260);
nor U12406 (N_12406,N_10731,N_11239);
and U12407 (N_12407,N_10977,N_10452);
and U12408 (N_12408,N_10436,N_11121);
nand U12409 (N_12409,N_10520,N_10037);
nand U12410 (N_12410,N_10987,N_10718);
nor U12411 (N_12411,N_10040,N_11142);
nand U12412 (N_12412,N_10231,N_11227);
and U12413 (N_12413,N_11199,N_10808);
nand U12414 (N_12414,N_10872,N_10059);
xnor U12415 (N_12415,N_11095,N_10584);
and U12416 (N_12416,N_10316,N_10930);
xor U12417 (N_12417,N_11001,N_10826);
and U12418 (N_12418,N_10612,N_10879);
or U12419 (N_12419,N_11001,N_11071);
xnor U12420 (N_12420,N_11036,N_10619);
nor U12421 (N_12421,N_10319,N_10603);
xnor U12422 (N_12422,N_10392,N_10050);
and U12423 (N_12423,N_11015,N_10483);
and U12424 (N_12424,N_10030,N_10092);
or U12425 (N_12425,N_10348,N_10514);
nand U12426 (N_12426,N_11180,N_11243);
or U12427 (N_12427,N_10082,N_11156);
and U12428 (N_12428,N_10774,N_11040);
nand U12429 (N_12429,N_11122,N_10121);
and U12430 (N_12430,N_10970,N_10829);
or U12431 (N_12431,N_10658,N_10327);
nand U12432 (N_12432,N_10229,N_10679);
and U12433 (N_12433,N_10048,N_10462);
xor U12434 (N_12434,N_11129,N_10064);
and U12435 (N_12435,N_11208,N_10888);
or U12436 (N_12436,N_10656,N_10801);
nor U12437 (N_12437,N_10308,N_10458);
or U12438 (N_12438,N_10332,N_10489);
nand U12439 (N_12439,N_10264,N_10367);
and U12440 (N_12440,N_10080,N_10738);
or U12441 (N_12441,N_10112,N_11155);
and U12442 (N_12442,N_10980,N_11209);
nor U12443 (N_12443,N_11198,N_10002);
nor U12444 (N_12444,N_11025,N_10103);
nand U12445 (N_12445,N_10622,N_10898);
nor U12446 (N_12446,N_10203,N_10409);
or U12447 (N_12447,N_10659,N_10984);
or U12448 (N_12448,N_11201,N_11006);
nor U12449 (N_12449,N_10376,N_10045);
and U12450 (N_12450,N_11248,N_11174);
nor U12451 (N_12451,N_10967,N_10427);
nor U12452 (N_12452,N_10625,N_10423);
and U12453 (N_12453,N_10508,N_10913);
and U12454 (N_12454,N_10961,N_10878);
nor U12455 (N_12455,N_10824,N_11227);
or U12456 (N_12456,N_10164,N_11004);
nand U12457 (N_12457,N_10307,N_11232);
and U12458 (N_12458,N_10813,N_11132);
xor U12459 (N_12459,N_10760,N_10721);
or U12460 (N_12460,N_11026,N_10872);
or U12461 (N_12461,N_10528,N_10061);
xor U12462 (N_12462,N_10718,N_10307);
nand U12463 (N_12463,N_11039,N_10007);
xnor U12464 (N_12464,N_10089,N_10794);
nor U12465 (N_12465,N_10551,N_10458);
nor U12466 (N_12466,N_10696,N_11077);
nand U12467 (N_12467,N_10192,N_10041);
and U12468 (N_12468,N_10095,N_10294);
and U12469 (N_12469,N_10427,N_10925);
and U12470 (N_12470,N_11059,N_10476);
nand U12471 (N_12471,N_11214,N_11227);
nand U12472 (N_12472,N_10321,N_10525);
nand U12473 (N_12473,N_10766,N_10899);
or U12474 (N_12474,N_10842,N_10329);
nor U12475 (N_12475,N_10673,N_10425);
nand U12476 (N_12476,N_10024,N_10475);
or U12477 (N_12477,N_10322,N_10011);
nand U12478 (N_12478,N_10375,N_10316);
or U12479 (N_12479,N_10176,N_11086);
nand U12480 (N_12480,N_11195,N_10804);
nand U12481 (N_12481,N_10598,N_10300);
or U12482 (N_12482,N_10434,N_11006);
nor U12483 (N_12483,N_10042,N_10694);
nand U12484 (N_12484,N_10892,N_11137);
and U12485 (N_12485,N_10489,N_10906);
xnor U12486 (N_12486,N_11197,N_10317);
xor U12487 (N_12487,N_10851,N_11159);
nand U12488 (N_12488,N_10034,N_10075);
nand U12489 (N_12489,N_11228,N_11001);
nor U12490 (N_12490,N_11160,N_10075);
or U12491 (N_12491,N_11145,N_10531);
xor U12492 (N_12492,N_10716,N_10959);
nand U12493 (N_12493,N_10733,N_10220);
nand U12494 (N_12494,N_10101,N_10454);
xor U12495 (N_12495,N_11139,N_10185);
nor U12496 (N_12496,N_10095,N_10351);
nand U12497 (N_12497,N_10668,N_11170);
or U12498 (N_12498,N_10702,N_10617);
or U12499 (N_12499,N_10571,N_10821);
or U12500 (N_12500,N_12062,N_12316);
xor U12501 (N_12501,N_12145,N_12467);
nand U12502 (N_12502,N_11757,N_11777);
nand U12503 (N_12503,N_12143,N_12172);
or U12504 (N_12504,N_11369,N_11420);
and U12505 (N_12505,N_11254,N_11590);
nand U12506 (N_12506,N_11610,N_12404);
or U12507 (N_12507,N_11354,N_11300);
xnor U12508 (N_12508,N_12155,N_11325);
or U12509 (N_12509,N_11648,N_12478);
or U12510 (N_12510,N_11412,N_11501);
xnor U12511 (N_12511,N_12068,N_11982);
xnor U12512 (N_12512,N_11364,N_11406);
or U12513 (N_12513,N_11569,N_12270);
and U12514 (N_12514,N_11820,N_11441);
nor U12515 (N_12515,N_11802,N_11552);
or U12516 (N_12516,N_11658,N_12452);
and U12517 (N_12517,N_11267,N_12198);
or U12518 (N_12518,N_11398,N_11755);
or U12519 (N_12519,N_12051,N_12135);
and U12520 (N_12520,N_11459,N_11840);
xor U12521 (N_12521,N_12326,N_12146);
nor U12522 (N_12522,N_12387,N_11293);
and U12523 (N_12523,N_12071,N_11960);
xor U12524 (N_12524,N_11916,N_11438);
nand U12525 (N_12525,N_12016,N_12355);
xnor U12526 (N_12526,N_11323,N_12003);
nand U12527 (N_12527,N_11490,N_11404);
nor U12528 (N_12528,N_11463,N_12108);
xor U12529 (N_12529,N_12253,N_12086);
nand U12530 (N_12530,N_11460,N_11301);
xor U12531 (N_12531,N_11432,N_11657);
nand U12532 (N_12532,N_12047,N_12219);
nor U12533 (N_12533,N_12396,N_11667);
nor U12534 (N_12534,N_11938,N_11389);
xnor U12535 (N_12535,N_11799,N_12353);
and U12536 (N_12536,N_12189,N_12288);
and U12537 (N_12537,N_11918,N_11319);
xor U12538 (N_12538,N_12491,N_11679);
or U12539 (N_12539,N_11291,N_11603);
nand U12540 (N_12540,N_11548,N_11942);
xor U12541 (N_12541,N_11280,N_11791);
xnor U12542 (N_12542,N_12426,N_11595);
nor U12543 (N_12543,N_11661,N_12165);
or U12544 (N_12544,N_11919,N_11915);
nand U12545 (N_12545,N_11401,N_12224);
or U12546 (N_12546,N_11593,N_12241);
or U12547 (N_12547,N_11456,N_11874);
nor U12548 (N_12548,N_12262,N_11591);
and U12549 (N_12549,N_11341,N_11475);
nor U12550 (N_12550,N_11542,N_12366);
nand U12551 (N_12551,N_11746,N_11442);
and U12552 (N_12552,N_11886,N_12249);
nand U12553 (N_12553,N_12328,N_12177);
xor U12554 (N_12554,N_12179,N_11952);
and U12555 (N_12555,N_11798,N_12390);
xor U12556 (N_12556,N_11640,N_12096);
nand U12557 (N_12557,N_11635,N_12461);
and U12558 (N_12558,N_12321,N_11786);
nand U12559 (N_12559,N_12411,N_12073);
xnor U12560 (N_12560,N_12476,N_11421);
xnor U12561 (N_12561,N_11643,N_11846);
or U12562 (N_12562,N_11864,N_11829);
and U12563 (N_12563,N_12379,N_12124);
nand U12564 (N_12564,N_11264,N_11959);
or U12565 (N_12565,N_11894,N_12091);
and U12566 (N_12566,N_11517,N_12239);
or U12567 (N_12567,N_11743,N_11531);
nand U12568 (N_12568,N_12414,N_12251);
nor U12569 (N_12569,N_11447,N_12268);
xor U12570 (N_12570,N_12254,N_11434);
or U12571 (N_12571,N_12325,N_11549);
or U12572 (N_12572,N_12159,N_11493);
or U12573 (N_12573,N_11586,N_11858);
xor U12574 (N_12574,N_12066,N_12103);
nor U12575 (N_12575,N_12056,N_12152);
or U12576 (N_12576,N_11998,N_11662);
xnor U12577 (N_12577,N_12136,N_12450);
and U12578 (N_12578,N_11578,N_12458);
nor U12579 (N_12579,N_11939,N_11741);
xnor U12580 (N_12580,N_11892,N_12474);
xnor U12581 (N_12581,N_11540,N_11350);
nor U12582 (N_12582,N_11399,N_11298);
and U12583 (N_12583,N_12279,N_12349);
nor U12584 (N_12584,N_11677,N_11813);
nand U12585 (N_12585,N_11303,N_12197);
or U12586 (N_12586,N_11506,N_12186);
nand U12587 (N_12587,N_12225,N_11943);
and U12588 (N_12588,N_11855,N_11415);
and U12589 (N_12589,N_11682,N_12149);
and U12590 (N_12590,N_12115,N_12246);
or U12591 (N_12591,N_12256,N_11397);
xor U12592 (N_12592,N_11674,N_11538);
nand U12593 (N_12593,N_11931,N_11841);
and U12594 (N_12594,N_12214,N_11464);
nor U12595 (N_12595,N_12290,N_12301);
nand U12596 (N_12596,N_11435,N_12295);
xor U12597 (N_12597,N_11678,N_12208);
or U12598 (N_12598,N_12076,N_11411);
or U12599 (N_12599,N_12111,N_12485);
and U12600 (N_12600,N_11532,N_11896);
nor U12601 (N_12601,N_12050,N_11822);
nand U12602 (N_12602,N_11659,N_11419);
and U12603 (N_12603,N_12240,N_12057);
nor U12604 (N_12604,N_11413,N_12154);
or U12605 (N_12605,N_11262,N_11486);
and U12606 (N_12606,N_11541,N_12082);
nand U12607 (N_12607,N_12020,N_11946);
nand U12608 (N_12608,N_12403,N_11685);
nand U12609 (N_12609,N_12369,N_12244);
nand U12610 (N_12610,N_11545,N_11808);
and U12611 (N_12611,N_11990,N_11366);
xnor U12612 (N_12612,N_12131,N_11269);
nand U12613 (N_12613,N_11525,N_11634);
nand U12614 (N_12614,N_11676,N_11870);
xor U12615 (N_12615,N_11535,N_11430);
xnor U12616 (N_12616,N_11418,N_11736);
and U12617 (N_12617,N_12227,N_12188);
or U12618 (N_12618,N_11407,N_11365);
nand U12619 (N_12619,N_11543,N_11878);
nand U12620 (N_12620,N_11932,N_11480);
or U12621 (N_12621,N_12490,N_12294);
nand U12622 (N_12622,N_12049,N_12106);
nand U12623 (N_12623,N_12032,N_12213);
xnor U12624 (N_12624,N_11934,N_11324);
xor U12625 (N_12625,N_12178,N_11315);
or U12626 (N_12626,N_11471,N_11580);
or U12627 (N_12627,N_11513,N_11284);
xnor U12628 (N_12628,N_12303,N_11842);
nor U12629 (N_12629,N_12202,N_11704);
xnor U12630 (N_12630,N_12024,N_11868);
and U12631 (N_12631,N_11276,N_12389);
and U12632 (N_12632,N_11694,N_12342);
and U12633 (N_12633,N_12412,N_11974);
and U12634 (N_12634,N_11347,N_11554);
xor U12635 (N_12635,N_11993,N_12228);
nand U12636 (N_12636,N_12237,N_12109);
xnor U12637 (N_12637,N_11718,N_11912);
and U12638 (N_12638,N_11391,N_11779);
nor U12639 (N_12639,N_11848,N_11646);
nand U12640 (N_12640,N_12304,N_11817);
nor U12641 (N_12641,N_11948,N_12469);
nand U12642 (N_12642,N_12015,N_11830);
and U12643 (N_12643,N_11362,N_11902);
or U12644 (N_12644,N_12243,N_12218);
nor U12645 (N_12645,N_11452,N_12431);
xor U12646 (N_12646,N_11865,N_11964);
nand U12647 (N_12647,N_11334,N_12477);
and U12648 (N_12648,N_12454,N_11614);
and U12649 (N_12649,N_11929,N_11805);
nand U12650 (N_12650,N_11526,N_11423);
or U12651 (N_12651,N_11877,N_12498);
xor U12652 (N_12652,N_11984,N_11905);
nand U12653 (N_12653,N_12421,N_11722);
nor U12654 (N_12654,N_12409,N_12022);
or U12655 (N_12655,N_11283,N_11336);
or U12656 (N_12656,N_11408,N_11875);
and U12657 (N_12657,N_11955,N_11266);
nand U12658 (N_12658,N_11473,N_11520);
and U12659 (N_12659,N_12487,N_11606);
nor U12660 (N_12660,N_11379,N_12479);
and U12661 (N_12661,N_11876,N_11827);
or U12662 (N_12662,N_11986,N_11706);
nand U12663 (N_12663,N_11385,N_11331);
nor U12664 (N_12664,N_11563,N_11689);
nand U12665 (N_12665,N_12418,N_11771);
nor U12666 (N_12666,N_11668,N_12433);
and U12667 (N_12667,N_11812,N_11485);
and U12668 (N_12668,N_11286,N_12181);
or U12669 (N_12669,N_11832,N_12245);
xor U12670 (N_12670,N_12141,N_12074);
or U12671 (N_12671,N_11624,N_11346);
nor U12672 (N_12672,N_12098,N_11901);
nor U12673 (N_12673,N_11458,N_11833);
xnor U12674 (N_12674,N_12345,N_11680);
nor U12675 (N_12675,N_12392,N_11382);
xnor U12676 (N_12676,N_11496,N_12119);
and U12677 (N_12677,N_11601,N_11428);
and U12678 (N_12678,N_11655,N_11255);
or U12679 (N_12679,N_11781,N_12105);
nor U12680 (N_12680,N_11395,N_11922);
nand U12681 (N_12681,N_11321,N_11512);
xor U12682 (N_12682,N_11288,N_12144);
or U12683 (N_12683,N_11550,N_11568);
xnor U12684 (N_12684,N_12424,N_12116);
nand U12685 (N_12685,N_12417,N_11769);
nand U12686 (N_12686,N_12045,N_11815);
nor U12687 (N_12687,N_11356,N_12297);
nand U12688 (N_12688,N_12460,N_11363);
nand U12689 (N_12689,N_12038,N_11523);
nor U12690 (N_12690,N_12435,N_12238);
nor U12691 (N_12691,N_11733,N_12367);
nor U12692 (N_12692,N_11978,N_12267);
nand U12693 (N_12693,N_11673,N_12457);
and U12694 (N_12694,N_12271,N_12191);
and U12695 (N_12695,N_12089,N_11927);
nand U12696 (N_12696,N_11565,N_11866);
nor U12697 (N_12697,N_11417,N_11429);
and U12698 (N_12698,N_11756,N_11695);
xnor U12699 (N_12699,N_12161,N_11923);
and U12700 (N_12700,N_12215,N_12110);
or U12701 (N_12701,N_12069,N_12204);
nand U12702 (N_12702,N_11744,N_11951);
nor U12703 (N_12703,N_11339,N_12012);
nor U12704 (N_12704,N_11845,N_12026);
nand U12705 (N_12705,N_12455,N_11883);
or U12706 (N_12706,N_12329,N_11814);
or U12707 (N_12707,N_11304,N_11602);
nand U12708 (N_12708,N_11509,N_11328);
xnor U12709 (N_12709,N_11597,N_12453);
nand U12710 (N_12710,N_11904,N_12230);
xor U12711 (N_12711,N_12148,N_12185);
nand U12712 (N_12712,N_11312,N_11309);
nor U12713 (N_12713,N_11313,N_12083);
xor U12714 (N_12714,N_11282,N_12407);
and U12715 (N_12715,N_12255,N_11329);
nor U12716 (N_12716,N_12233,N_11281);
xnor U12717 (N_12717,N_11553,N_11575);
or U12718 (N_12718,N_11446,N_11774);
nor U12719 (N_12719,N_11966,N_12497);
xor U12720 (N_12720,N_11612,N_12440);
nor U12721 (N_12721,N_11594,N_12350);
nand U12722 (N_12722,N_12093,N_12284);
nand U12723 (N_12723,N_11271,N_11872);
and U12724 (N_12724,N_11748,N_12129);
nand U12725 (N_12725,N_11310,N_11305);
and U12726 (N_12726,N_12216,N_11763);
or U12727 (N_12727,N_12483,N_11386);
nor U12728 (N_12728,N_12019,N_11294);
and U12729 (N_12729,N_12397,N_12158);
xor U12730 (N_12730,N_11273,N_12042);
and U12731 (N_12731,N_12285,N_12030);
xor U12732 (N_12732,N_12322,N_11863);
nor U12733 (N_12733,N_12346,N_11387);
and U12734 (N_12734,N_11476,N_12176);
xnor U12735 (N_12735,N_11852,N_11592);
xnor U12736 (N_12736,N_11383,N_11732);
nand U12737 (N_12737,N_11274,N_11436);
and U12738 (N_12738,N_12383,N_11857);
nand U12739 (N_12739,N_11616,N_11712);
xor U12740 (N_12740,N_12337,N_11360);
xnor U12741 (N_12741,N_11585,N_12283);
and U12742 (N_12742,N_11720,N_11937);
nor U12743 (N_12743,N_11311,N_12359);
and U12744 (N_12744,N_12365,N_11344);
or U12745 (N_12745,N_11700,N_11307);
or U12746 (N_12746,N_11469,N_11751);
or U12747 (N_12747,N_11261,N_11353);
nor U12748 (N_12748,N_12211,N_12087);
and U12749 (N_12749,N_11348,N_11994);
xor U12750 (N_12750,N_12332,N_12247);
and U12751 (N_12751,N_11800,N_12391);
or U12752 (N_12752,N_12043,N_11772);
nand U12753 (N_12753,N_11913,N_11619);
or U12754 (N_12754,N_11596,N_12427);
or U12755 (N_12755,N_11598,N_11738);
or U12756 (N_12756,N_12223,N_11851);
and U12757 (N_12757,N_11831,N_11579);
and U12758 (N_12758,N_11270,N_12482);
and U12759 (N_12759,N_11317,N_11296);
nand U12760 (N_12760,N_11839,N_11729);
and U12761 (N_12761,N_12384,N_11767);
xor U12762 (N_12762,N_12331,N_11971);
xor U12763 (N_12763,N_12085,N_12099);
xor U12764 (N_12764,N_11450,N_11470);
nand U12765 (N_12765,N_11881,N_11416);
and U12766 (N_12766,N_11519,N_12272);
nand U12767 (N_12767,N_12462,N_12001);
or U12768 (N_12768,N_12274,N_12192);
and U12769 (N_12769,N_11775,N_11691);
or U12770 (N_12770,N_11654,N_11547);
xnor U12771 (N_12771,N_11696,N_11534);
nor U12772 (N_12772,N_12336,N_11836);
xor U12773 (N_12773,N_11454,N_12092);
nor U12774 (N_12774,N_11873,N_12348);
and U12775 (N_12775,N_11882,N_11638);
nor U12776 (N_12776,N_11715,N_12286);
nor U12777 (N_12777,N_12395,N_11749);
nor U12778 (N_12778,N_11675,N_12101);
nand U12779 (N_12779,N_11975,N_12293);
nand U12780 (N_12780,N_11316,N_11518);
nand U12781 (N_12781,N_11489,N_12125);
nand U12782 (N_12782,N_12037,N_11394);
or U12783 (N_12783,N_11745,N_11641);
or U12784 (N_12784,N_11465,N_12318);
and U12785 (N_12785,N_11622,N_11561);
nand U12786 (N_12786,N_12021,N_11926);
nand U12787 (N_12787,N_11494,N_11488);
nand U12788 (N_12788,N_11268,N_11265);
nor U12789 (N_12789,N_12370,N_11925);
or U12790 (N_12790,N_11589,N_11508);
nor U12791 (N_12791,N_12220,N_11789);
nand U12792 (N_12792,N_11965,N_11295);
nor U12793 (N_12793,N_11425,N_12430);
xnor U12794 (N_12794,N_12190,N_12472);
xnor U12795 (N_12795,N_12343,N_11500);
and U12796 (N_12796,N_11867,N_11482);
xnor U12797 (N_12797,N_11507,N_11697);
xor U12798 (N_12798,N_11910,N_12394);
nor U12799 (N_12799,N_11289,N_11390);
and U12800 (N_12800,N_12040,N_11530);
nor U12801 (N_12801,N_11686,N_11726);
or U12802 (N_12802,N_11803,N_12356);
and U12803 (N_12803,N_11987,N_12234);
nand U12804 (N_12804,N_12481,N_12182);
nor U12805 (N_12805,N_12084,N_12088);
and U12806 (N_12806,N_11967,N_12195);
nand U12807 (N_12807,N_11451,N_11914);
nand U12808 (N_12808,N_12364,N_12381);
nor U12809 (N_12809,N_11809,N_11725);
xor U12810 (N_12810,N_11721,N_12072);
or U12811 (N_12811,N_11539,N_12444);
nor U12812 (N_12812,N_12232,N_12296);
nand U12813 (N_12813,N_11613,N_11357);
nor U12814 (N_12814,N_11380,N_12419);
and U12815 (N_12815,N_11976,N_12480);
or U12816 (N_12816,N_11853,N_11797);
and U12817 (N_12817,N_12107,N_11544);
or U12818 (N_12818,N_12277,N_11327);
and U12819 (N_12819,N_11514,N_11997);
or U12820 (N_12820,N_11524,N_12063);
xor U12821 (N_12821,N_11761,N_12323);
and U12822 (N_12822,N_11834,N_12058);
and U12823 (N_12823,N_11377,N_12064);
xnor U12824 (N_12824,N_11367,N_11630);
or U12825 (N_12825,N_12416,N_11587);
nor U12826 (N_12826,N_12017,N_11707);
xnor U12827 (N_12827,N_12206,N_11818);
nand U12828 (N_12828,N_11933,N_12493);
and U12829 (N_12829,N_11605,N_11502);
nand U12830 (N_12830,N_12305,N_11448);
and U12831 (N_12831,N_12126,N_11555);
or U12832 (N_12832,N_11989,N_11566);
nand U12833 (N_12833,N_11690,N_12121);
xnor U12834 (N_12834,N_11302,N_12281);
nand U12835 (N_12835,N_11628,N_12079);
nand U12836 (N_12836,N_11664,N_11497);
or U12837 (N_12837,N_12077,N_11437);
nor U12838 (N_12838,N_11393,N_12432);
or U12839 (N_12839,N_12464,N_12425);
xnor U12840 (N_12840,N_12446,N_12250);
or U12841 (N_12841,N_12229,N_12180);
nand U12842 (N_12842,N_12330,N_12385);
or U12843 (N_12843,N_12499,N_11887);
nand U12844 (N_12844,N_11862,N_11449);
and U12845 (N_12845,N_12226,N_11995);
xor U12846 (N_12846,N_11625,N_12489);
and U12847 (N_12847,N_11631,N_12210);
and U12848 (N_12848,N_12036,N_11468);
nand U12849 (N_12849,N_11361,N_11272);
or U12850 (N_12850,N_11467,N_11637);
or U12851 (N_12851,N_11376,N_11670);
nand U12852 (N_12852,N_11889,N_11278);
nand U12853 (N_12853,N_11533,N_11623);
nand U12854 (N_12854,N_12203,N_11576);
and U12855 (N_12855,N_11402,N_12171);
or U12856 (N_12856,N_11935,N_12339);
nand U12857 (N_12857,N_11433,N_12142);
and U12858 (N_12858,N_11895,N_12127);
or U12859 (N_12859,N_11957,N_11478);
or U12860 (N_12860,N_12122,N_11522);
nor U12861 (N_12861,N_11856,N_11521);
or U12862 (N_12862,N_11285,N_12368);
and U12863 (N_12863,N_12495,N_11396);
or U12864 (N_12864,N_12002,N_11252);
nand U12865 (N_12865,N_12200,N_12023);
and U12866 (N_12866,N_12441,N_12352);
or U12867 (N_12867,N_12357,N_11322);
and U12868 (N_12868,N_11351,N_11621);
or U12869 (N_12869,N_12187,N_11735);
xnor U12870 (N_12870,N_12335,N_12486);
xor U12871 (N_12871,N_11516,N_11861);
and U12872 (N_12872,N_11880,N_11961);
nor U12873 (N_12873,N_11983,N_11871);
or U12874 (N_12874,N_12298,N_11709);
nor U12875 (N_12875,N_11843,N_11571);
nor U12876 (N_12876,N_11705,N_11345);
and U12877 (N_12877,N_12222,N_11826);
nor U12878 (N_12878,N_11992,N_11343);
nor U12879 (N_12879,N_12013,N_12398);
nand U12880 (N_12880,N_12118,N_11949);
nor U12881 (N_12881,N_11936,N_12340);
xnor U12882 (N_12882,N_11649,N_12338);
xor U12883 (N_12883,N_11823,N_11588);
or U12884 (N_12884,N_11849,N_11556);
xnor U12885 (N_12885,N_12217,N_11794);
nor U12886 (N_12886,N_12371,N_12428);
or U12887 (N_12887,N_11979,N_12437);
nor U12888 (N_12888,N_12196,N_12278);
or U12889 (N_12889,N_12362,N_11666);
nor U12890 (N_12890,N_11374,N_12488);
and U12891 (N_12891,N_11573,N_12170);
or U12892 (N_12892,N_11899,N_11713);
nor U12893 (N_12893,N_12408,N_12302);
and U12894 (N_12894,N_12194,N_11251);
and U12895 (N_12895,N_11584,N_11711);
xor U12896 (N_12896,N_12166,N_11338);
or U12897 (N_12897,N_12263,N_11629);
nand U12898 (N_12898,N_11708,N_11981);
and U12899 (N_12899,N_12175,N_11609);
and U12900 (N_12900,N_12094,N_11962);
nor U12901 (N_12901,N_12150,N_12162);
and U12902 (N_12902,N_12313,N_11956);
xnor U12903 (N_12903,N_11947,N_11941);
nand U12904 (N_12904,N_12117,N_11632);
xor U12905 (N_12905,N_12014,N_12434);
nor U12906 (N_12906,N_12028,N_12377);
or U12907 (N_12907,N_11444,N_11615);
nor U12908 (N_12908,N_11945,N_12132);
or U12909 (N_12909,N_11639,N_11930);
nand U12910 (N_12910,N_11299,N_11297);
or U12911 (N_12911,N_12386,N_11859);
or U12912 (N_12912,N_11600,N_11422);
nand U12913 (N_12913,N_12496,N_11734);
nor U12914 (N_12914,N_11907,N_11292);
nor U12915 (N_12915,N_11636,N_11810);
and U12916 (N_12916,N_11985,N_11504);
or U12917 (N_12917,N_12445,N_12358);
and U12918 (N_12918,N_12265,N_11320);
nand U12919 (N_12919,N_11776,N_12231);
nor U12920 (N_12920,N_11647,N_11567);
nand U12921 (N_12921,N_11620,N_12120);
xor U12922 (N_12922,N_12374,N_11250);
nand U12923 (N_12923,N_12341,N_12449);
or U12924 (N_12924,N_11788,N_12059);
nor U12925 (N_12925,N_11515,N_11760);
or U12926 (N_12926,N_11660,N_12311);
or U12927 (N_12927,N_11906,N_11766);
nand U12928 (N_12928,N_11352,N_11801);
or U12929 (N_12929,N_11572,N_11381);
nand U12930 (N_12930,N_11972,N_12209);
nor U12931 (N_12931,N_11717,N_11409);
or U12932 (N_12932,N_11375,N_11977);
and U12933 (N_12933,N_12029,N_12090);
or U12934 (N_12934,N_11893,N_11577);
or U12935 (N_12935,N_12307,N_11884);
and U12936 (N_12936,N_11642,N_11258);
nor U12937 (N_12937,N_12112,N_11693);
or U12938 (N_12938,N_11821,N_11644);
xnor U12939 (N_12939,N_11944,N_12004);
nand U12940 (N_12940,N_12317,N_12102);
nand U12941 (N_12941,N_12448,N_11495);
nor U12942 (N_12942,N_11728,N_11570);
nor U12943 (N_12943,N_11400,N_12309);
nand U12944 (N_12944,N_11607,N_11558);
or U12945 (N_12945,N_11479,N_11672);
xnor U12946 (N_12946,N_12123,N_11969);
nor U12947 (N_12947,N_11770,N_12252);
or U12948 (N_12948,N_11681,N_11703);
and U12949 (N_12949,N_11332,N_11671);
or U12950 (N_12950,N_11890,N_12306);
or U12951 (N_12951,N_11740,N_12269);
nand U12952 (N_12952,N_11928,N_11727);
nor U12953 (N_12953,N_11359,N_12054);
and U12954 (N_12954,N_12423,N_11804);
nand U12955 (N_12955,N_12048,N_11940);
and U12956 (N_12956,N_12199,N_12291);
nand U12957 (N_12957,N_11529,N_11318);
nand U12958 (N_12958,N_12468,N_12308);
and U12959 (N_12959,N_12041,N_12201);
or U12960 (N_12960,N_12010,N_11773);
nand U12961 (N_12961,N_12360,N_11279);
nor U12962 (N_12962,N_12055,N_11466);
or U12963 (N_12963,N_11692,N_11780);
or U12964 (N_12964,N_12018,N_11378);
nand U12965 (N_12965,N_12459,N_11795);
nand U12966 (N_12966,N_11574,N_11807);
xnor U12967 (N_12967,N_12128,N_11909);
or U12968 (N_12968,N_12168,N_11753);
nor U12969 (N_12969,N_11701,N_12157);
nand U12970 (N_12970,N_12280,N_11499);
and U12971 (N_12971,N_12070,N_12053);
nor U12972 (N_12972,N_11869,N_11954);
or U12973 (N_12973,N_11988,N_11492);
and U12974 (N_12974,N_12212,N_12034);
nor U12975 (N_12975,N_11793,N_12205);
and U12976 (N_12976,N_12393,N_12315);
and U12977 (N_12977,N_11527,N_12324);
xnor U12978 (N_12978,N_12465,N_11443);
xnor U12979 (N_12979,N_12439,N_11627);
and U12980 (N_12980,N_12033,N_12410);
or U12981 (N_12981,N_11716,N_11669);
nor U12982 (N_12982,N_12282,N_12429);
nor U12983 (N_12983,N_12372,N_12422);
and U12984 (N_12984,N_11903,N_12382);
nand U12985 (N_12985,N_12031,N_11950);
xnor U12986 (N_12986,N_11958,N_11474);
xor U12987 (N_12987,N_11739,N_11604);
nand U12988 (N_12988,N_12327,N_11684);
nand U12989 (N_12989,N_11330,N_12139);
xnor U12990 (N_12990,N_11487,N_11503);
or U12991 (N_12991,N_12320,N_12137);
or U12992 (N_12992,N_11340,N_11306);
nand U12993 (N_12993,N_12471,N_12438);
and U12994 (N_12994,N_11663,N_11439);
and U12995 (N_12995,N_12451,N_11483);
nor U12996 (N_12996,N_11431,N_11996);
nand U12997 (N_12997,N_12242,N_11440);
and U12998 (N_12998,N_12035,N_11888);
nor U12999 (N_12999,N_12275,N_12163);
nand U13000 (N_13000,N_11263,N_11645);
and U13001 (N_13001,N_11838,N_12261);
or U13002 (N_13002,N_12314,N_11759);
nand U13003 (N_13003,N_11308,N_11275);
nand U13004 (N_13004,N_11453,N_12011);
nand U13005 (N_13005,N_11472,N_11498);
and U13006 (N_13006,N_12046,N_11844);
nand U13007 (N_13007,N_11260,N_11891);
and U13008 (N_13008,N_12065,N_11665);
xnor U13009 (N_13009,N_12130,N_11368);
xor U13010 (N_13010,N_11783,N_12344);
or U13011 (N_13011,N_11358,N_11618);
nor U13012 (N_13012,N_11557,N_11999);
xor U13013 (N_13013,N_11414,N_11650);
xor U13014 (N_13014,N_11920,N_11683);
nor U13015 (N_13015,N_11427,N_12008);
or U13016 (N_13016,N_11617,N_11764);
xnor U13017 (N_13017,N_12378,N_12273);
and U13018 (N_13018,N_11714,N_12260);
or U13019 (N_13019,N_11461,N_12147);
nand U13020 (N_13020,N_11900,N_11737);
nor U13021 (N_13021,N_12221,N_11564);
nor U13022 (N_13022,N_12380,N_11626);
xnor U13023 (N_13023,N_11384,N_12114);
or U13024 (N_13024,N_11599,N_12044);
nor U13025 (N_13025,N_11698,N_11765);
nand U13026 (N_13026,N_12061,N_11898);
and U13027 (N_13027,N_12151,N_11333);
nand U13028 (N_13028,N_11611,N_11491);
or U13029 (N_13029,N_11560,N_12363);
nor U13030 (N_13030,N_12492,N_12494);
xor U13031 (N_13031,N_12375,N_11816);
and U13032 (N_13032,N_12399,N_11392);
nand U13033 (N_13033,N_11811,N_11651);
and U13034 (N_13034,N_11768,N_11253);
or U13035 (N_13035,N_11924,N_12388);
xor U13036 (N_13036,N_11652,N_12401);
nor U13037 (N_13037,N_11562,N_12443);
and U13038 (N_13038,N_12039,N_12095);
or U13039 (N_13039,N_12400,N_11687);
and U13040 (N_13040,N_12405,N_12470);
or U13041 (N_13041,N_12183,N_12299);
or U13042 (N_13042,N_11723,N_11835);
or U13043 (N_13043,N_12264,N_11410);
xor U13044 (N_13044,N_12276,N_11256);
and U13045 (N_13045,N_11973,N_11583);
and U13046 (N_13046,N_11980,N_11455);
nor U13047 (N_13047,N_12361,N_11911);
nor U13048 (N_13048,N_11477,N_12447);
nor U13049 (N_13049,N_11370,N_12140);
xor U13050 (N_13050,N_12258,N_11806);
and U13051 (N_13051,N_12259,N_12484);
nand U13052 (N_13052,N_11917,N_11426);
nand U13053 (N_13053,N_11719,N_11373);
xor U13054 (N_13054,N_12456,N_11963);
nand U13055 (N_13055,N_11752,N_11656);
or U13056 (N_13056,N_11785,N_11837);
nor U13057 (N_13057,N_12138,N_11824);
xor U13058 (N_13058,N_12266,N_11762);
xnor U13059 (N_13059,N_11314,N_11921);
or U13060 (N_13060,N_11758,N_11287);
and U13061 (N_13061,N_12153,N_11259);
or U13062 (N_13062,N_11326,N_11699);
and U13063 (N_13063,N_12248,N_12000);
and U13064 (N_13064,N_12333,N_11854);
xor U13065 (N_13065,N_11608,N_11349);
xor U13066 (N_13066,N_11742,N_11991);
nand U13067 (N_13067,N_11825,N_11730);
or U13068 (N_13068,N_11850,N_11510);
xor U13069 (N_13069,N_12027,N_11582);
nor U13070 (N_13070,N_11782,N_12067);
or U13071 (N_13071,N_11970,N_11953);
nand U13072 (N_13072,N_11403,N_12257);
nand U13073 (N_13073,N_11968,N_12236);
nand U13074 (N_13074,N_11787,N_12402);
nor U13075 (N_13075,N_11388,N_11537);
nor U13076 (N_13076,N_11342,N_11828);
xor U13077 (N_13077,N_11702,N_12006);
or U13078 (N_13078,N_12292,N_11747);
xnor U13079 (N_13079,N_12160,N_12052);
and U13080 (N_13080,N_12475,N_11546);
and U13081 (N_13081,N_12354,N_12312);
or U13082 (N_13082,N_12347,N_12463);
or U13083 (N_13083,N_12406,N_11633);
xnor U13084 (N_13084,N_11445,N_12174);
or U13085 (N_13085,N_11796,N_12100);
nor U13086 (N_13086,N_11457,N_11790);
and U13087 (N_13087,N_11462,N_11528);
and U13088 (N_13088,N_12081,N_11257);
nand U13089 (N_13089,N_11536,N_11290);
xor U13090 (N_13090,N_11337,N_12097);
or U13091 (N_13091,N_12442,N_11897);
nand U13092 (N_13092,N_11710,N_12413);
or U13093 (N_13093,N_11754,N_11505);
nand U13094 (N_13094,N_12436,N_12080);
and U13095 (N_13095,N_12376,N_11885);
xnor U13096 (N_13096,N_12169,N_12164);
nor U13097 (N_13097,N_12319,N_11481);
or U13098 (N_13098,N_12007,N_11511);
and U13099 (N_13099,N_11484,N_11372);
nor U13100 (N_13100,N_12334,N_12173);
and U13101 (N_13101,N_12415,N_11551);
and U13102 (N_13102,N_11879,N_11355);
nor U13103 (N_13103,N_12420,N_12287);
xnor U13104 (N_13104,N_11750,N_11792);
or U13105 (N_13105,N_11653,N_11778);
nor U13106 (N_13106,N_12113,N_11847);
and U13107 (N_13107,N_12473,N_12104);
or U13108 (N_13108,N_11724,N_12351);
or U13109 (N_13109,N_12373,N_12466);
and U13110 (N_13110,N_11860,N_12009);
nand U13111 (N_13111,N_11371,N_11908);
nor U13112 (N_13112,N_11277,N_12075);
xor U13113 (N_13113,N_12060,N_11581);
or U13114 (N_13114,N_12133,N_11731);
xor U13115 (N_13115,N_11559,N_11405);
nand U13116 (N_13116,N_12300,N_12167);
nor U13117 (N_13117,N_11424,N_12184);
xnor U13118 (N_13118,N_11819,N_12235);
nor U13119 (N_13119,N_12134,N_12025);
nor U13120 (N_13120,N_12078,N_12310);
nand U13121 (N_13121,N_12193,N_12156);
xnor U13122 (N_13122,N_11335,N_11688);
nor U13123 (N_13123,N_12207,N_12005);
or U13124 (N_13124,N_12289,N_11784);
nand U13125 (N_13125,N_11252,N_12463);
and U13126 (N_13126,N_11317,N_11353);
nand U13127 (N_13127,N_12392,N_11388);
or U13128 (N_13128,N_11755,N_11939);
and U13129 (N_13129,N_11553,N_11418);
and U13130 (N_13130,N_12118,N_11921);
or U13131 (N_13131,N_11863,N_12071);
xnor U13132 (N_13132,N_12466,N_12267);
nor U13133 (N_13133,N_12125,N_11736);
nor U13134 (N_13134,N_11541,N_12061);
and U13135 (N_13135,N_11796,N_11771);
nand U13136 (N_13136,N_12473,N_11714);
xor U13137 (N_13137,N_12287,N_12201);
nand U13138 (N_13138,N_11259,N_12058);
and U13139 (N_13139,N_11977,N_11483);
or U13140 (N_13140,N_11911,N_11503);
xor U13141 (N_13141,N_11773,N_11964);
nor U13142 (N_13142,N_11737,N_12306);
xnor U13143 (N_13143,N_11901,N_11470);
xor U13144 (N_13144,N_12269,N_11640);
nand U13145 (N_13145,N_11409,N_11354);
or U13146 (N_13146,N_11435,N_11324);
xor U13147 (N_13147,N_11993,N_11256);
nor U13148 (N_13148,N_12465,N_11935);
nor U13149 (N_13149,N_12005,N_11647);
nand U13150 (N_13150,N_12425,N_11509);
xnor U13151 (N_13151,N_11311,N_12329);
nor U13152 (N_13152,N_11590,N_11486);
nor U13153 (N_13153,N_11333,N_11739);
xor U13154 (N_13154,N_11918,N_12376);
nand U13155 (N_13155,N_12492,N_11627);
xnor U13156 (N_13156,N_12156,N_11437);
xor U13157 (N_13157,N_11390,N_12428);
nor U13158 (N_13158,N_11481,N_12110);
or U13159 (N_13159,N_12414,N_11395);
and U13160 (N_13160,N_12004,N_11786);
or U13161 (N_13161,N_11281,N_12110);
and U13162 (N_13162,N_12449,N_11905);
xnor U13163 (N_13163,N_11401,N_11967);
xor U13164 (N_13164,N_12011,N_12463);
and U13165 (N_13165,N_12218,N_11354);
or U13166 (N_13166,N_11783,N_11651);
and U13167 (N_13167,N_11393,N_11848);
and U13168 (N_13168,N_12371,N_11891);
xor U13169 (N_13169,N_11490,N_11823);
nand U13170 (N_13170,N_12116,N_11790);
nor U13171 (N_13171,N_12192,N_12216);
nand U13172 (N_13172,N_11983,N_12318);
and U13173 (N_13173,N_11613,N_11315);
nor U13174 (N_13174,N_11488,N_11699);
or U13175 (N_13175,N_11670,N_11560);
or U13176 (N_13176,N_12208,N_12006);
and U13177 (N_13177,N_11793,N_11344);
xor U13178 (N_13178,N_12056,N_11555);
nor U13179 (N_13179,N_11415,N_11889);
and U13180 (N_13180,N_11801,N_11288);
and U13181 (N_13181,N_12007,N_12217);
or U13182 (N_13182,N_12003,N_11479);
nor U13183 (N_13183,N_11414,N_12460);
or U13184 (N_13184,N_11785,N_11485);
and U13185 (N_13185,N_12316,N_11610);
nor U13186 (N_13186,N_11754,N_11333);
or U13187 (N_13187,N_12001,N_11285);
xnor U13188 (N_13188,N_11575,N_11579);
xor U13189 (N_13189,N_11549,N_11805);
and U13190 (N_13190,N_11661,N_12407);
and U13191 (N_13191,N_11513,N_12290);
nor U13192 (N_13192,N_12233,N_12251);
nand U13193 (N_13193,N_11540,N_12132);
and U13194 (N_13194,N_12277,N_12200);
nand U13195 (N_13195,N_12406,N_12218);
xnor U13196 (N_13196,N_12011,N_11470);
nand U13197 (N_13197,N_11362,N_11270);
nand U13198 (N_13198,N_11609,N_12062);
nand U13199 (N_13199,N_12435,N_12443);
nor U13200 (N_13200,N_12275,N_12114);
xor U13201 (N_13201,N_11392,N_11506);
nor U13202 (N_13202,N_12415,N_12344);
nand U13203 (N_13203,N_11600,N_11546);
nor U13204 (N_13204,N_11922,N_12209);
nor U13205 (N_13205,N_11902,N_11342);
xor U13206 (N_13206,N_11956,N_11291);
or U13207 (N_13207,N_12050,N_12302);
nor U13208 (N_13208,N_12205,N_11501);
or U13209 (N_13209,N_12037,N_11632);
nand U13210 (N_13210,N_12172,N_12399);
and U13211 (N_13211,N_11366,N_11369);
nand U13212 (N_13212,N_11405,N_11776);
and U13213 (N_13213,N_11932,N_11974);
and U13214 (N_13214,N_11871,N_12310);
and U13215 (N_13215,N_12028,N_11678);
nor U13216 (N_13216,N_11256,N_12324);
and U13217 (N_13217,N_12114,N_11655);
and U13218 (N_13218,N_12170,N_12274);
nand U13219 (N_13219,N_11417,N_11955);
xnor U13220 (N_13220,N_12376,N_11411);
nand U13221 (N_13221,N_12345,N_11957);
nand U13222 (N_13222,N_11578,N_11993);
xor U13223 (N_13223,N_11595,N_11468);
nand U13224 (N_13224,N_11260,N_11967);
xor U13225 (N_13225,N_11825,N_11572);
xor U13226 (N_13226,N_11380,N_12488);
or U13227 (N_13227,N_12205,N_11900);
nor U13228 (N_13228,N_12485,N_11874);
and U13229 (N_13229,N_11948,N_11300);
xor U13230 (N_13230,N_12370,N_12038);
nand U13231 (N_13231,N_11445,N_11376);
nand U13232 (N_13232,N_11554,N_11405);
and U13233 (N_13233,N_12399,N_11316);
or U13234 (N_13234,N_12367,N_12262);
and U13235 (N_13235,N_12109,N_11704);
and U13236 (N_13236,N_12030,N_12182);
or U13237 (N_13237,N_11807,N_11337);
and U13238 (N_13238,N_11946,N_11891);
or U13239 (N_13239,N_12288,N_11944);
nor U13240 (N_13240,N_12206,N_11431);
and U13241 (N_13241,N_11421,N_12169);
and U13242 (N_13242,N_11480,N_11698);
xor U13243 (N_13243,N_11603,N_11866);
nor U13244 (N_13244,N_11942,N_11517);
nor U13245 (N_13245,N_12140,N_12058);
nor U13246 (N_13246,N_11447,N_11288);
nor U13247 (N_13247,N_11360,N_12028);
nor U13248 (N_13248,N_12087,N_11335);
nor U13249 (N_13249,N_12452,N_12060);
and U13250 (N_13250,N_12492,N_11904);
or U13251 (N_13251,N_11291,N_12223);
or U13252 (N_13252,N_11889,N_11990);
or U13253 (N_13253,N_12444,N_12419);
or U13254 (N_13254,N_11928,N_11293);
and U13255 (N_13255,N_11420,N_11429);
nand U13256 (N_13256,N_11720,N_12416);
nand U13257 (N_13257,N_12044,N_11773);
xnor U13258 (N_13258,N_11933,N_11992);
and U13259 (N_13259,N_11345,N_11270);
and U13260 (N_13260,N_11671,N_12186);
or U13261 (N_13261,N_11576,N_11747);
and U13262 (N_13262,N_12248,N_11258);
or U13263 (N_13263,N_11777,N_11772);
or U13264 (N_13264,N_11667,N_11320);
nand U13265 (N_13265,N_11692,N_11923);
or U13266 (N_13266,N_11302,N_12222);
xnor U13267 (N_13267,N_12245,N_11642);
nand U13268 (N_13268,N_11991,N_11431);
nand U13269 (N_13269,N_11848,N_11853);
xnor U13270 (N_13270,N_11632,N_11375);
or U13271 (N_13271,N_11980,N_11966);
or U13272 (N_13272,N_11623,N_11348);
xor U13273 (N_13273,N_11804,N_11936);
nand U13274 (N_13274,N_12326,N_11462);
xnor U13275 (N_13275,N_12028,N_12127);
nor U13276 (N_13276,N_11526,N_11394);
nand U13277 (N_13277,N_11595,N_11348);
or U13278 (N_13278,N_12350,N_12426);
and U13279 (N_13279,N_11707,N_11259);
and U13280 (N_13280,N_12353,N_12100);
nor U13281 (N_13281,N_12391,N_11921);
and U13282 (N_13282,N_12421,N_11506);
nand U13283 (N_13283,N_12453,N_11550);
or U13284 (N_13284,N_12096,N_11483);
or U13285 (N_13285,N_12013,N_11601);
or U13286 (N_13286,N_12263,N_12240);
nor U13287 (N_13287,N_11677,N_11257);
nor U13288 (N_13288,N_11808,N_12322);
nor U13289 (N_13289,N_11317,N_12026);
xnor U13290 (N_13290,N_11773,N_11958);
and U13291 (N_13291,N_11374,N_12161);
nor U13292 (N_13292,N_12096,N_11428);
nand U13293 (N_13293,N_12025,N_12304);
and U13294 (N_13294,N_12010,N_11390);
nand U13295 (N_13295,N_12309,N_11637);
nand U13296 (N_13296,N_11562,N_11356);
nor U13297 (N_13297,N_12240,N_12148);
or U13298 (N_13298,N_12483,N_12227);
xnor U13299 (N_13299,N_11625,N_11814);
xnor U13300 (N_13300,N_11357,N_12128);
nor U13301 (N_13301,N_11855,N_12186);
and U13302 (N_13302,N_12360,N_11812);
xnor U13303 (N_13303,N_11883,N_11757);
or U13304 (N_13304,N_11257,N_12393);
and U13305 (N_13305,N_12187,N_11282);
nand U13306 (N_13306,N_12471,N_12429);
nand U13307 (N_13307,N_11544,N_12234);
or U13308 (N_13308,N_11945,N_12489);
nand U13309 (N_13309,N_12418,N_12066);
nand U13310 (N_13310,N_12335,N_11892);
nor U13311 (N_13311,N_12296,N_11923);
nor U13312 (N_13312,N_12266,N_11726);
or U13313 (N_13313,N_11439,N_11674);
or U13314 (N_13314,N_11257,N_12479);
and U13315 (N_13315,N_11621,N_12059);
or U13316 (N_13316,N_12446,N_11418);
nor U13317 (N_13317,N_12107,N_12164);
nor U13318 (N_13318,N_12441,N_11882);
nand U13319 (N_13319,N_11554,N_12373);
and U13320 (N_13320,N_11865,N_11689);
or U13321 (N_13321,N_12120,N_11695);
or U13322 (N_13322,N_12324,N_12205);
nor U13323 (N_13323,N_12085,N_11666);
nor U13324 (N_13324,N_12276,N_12038);
or U13325 (N_13325,N_11625,N_11788);
xor U13326 (N_13326,N_12028,N_12393);
and U13327 (N_13327,N_12390,N_11593);
and U13328 (N_13328,N_12119,N_11357);
nand U13329 (N_13329,N_11658,N_11319);
nand U13330 (N_13330,N_11904,N_12448);
xor U13331 (N_13331,N_11925,N_12162);
nand U13332 (N_13332,N_12240,N_11709);
or U13333 (N_13333,N_11915,N_12207);
and U13334 (N_13334,N_12463,N_12121);
xor U13335 (N_13335,N_12386,N_12078);
nor U13336 (N_13336,N_11833,N_11775);
nor U13337 (N_13337,N_12014,N_11979);
and U13338 (N_13338,N_11666,N_11326);
xor U13339 (N_13339,N_12162,N_11453);
or U13340 (N_13340,N_12375,N_12074);
nand U13341 (N_13341,N_11677,N_12380);
and U13342 (N_13342,N_12278,N_11345);
or U13343 (N_13343,N_12484,N_12396);
xnor U13344 (N_13344,N_11656,N_11505);
or U13345 (N_13345,N_12043,N_11718);
xor U13346 (N_13346,N_11735,N_12468);
nor U13347 (N_13347,N_12083,N_11478);
or U13348 (N_13348,N_12091,N_12010);
or U13349 (N_13349,N_11377,N_11762);
and U13350 (N_13350,N_11542,N_12440);
nor U13351 (N_13351,N_11685,N_11990);
xor U13352 (N_13352,N_11693,N_11796);
nand U13353 (N_13353,N_12400,N_12142);
and U13354 (N_13354,N_11515,N_11926);
nor U13355 (N_13355,N_12241,N_12072);
xnor U13356 (N_13356,N_11889,N_12298);
nand U13357 (N_13357,N_12313,N_11623);
nand U13358 (N_13358,N_11646,N_11946);
nor U13359 (N_13359,N_12495,N_12060);
nand U13360 (N_13360,N_12263,N_11304);
and U13361 (N_13361,N_12348,N_12201);
nand U13362 (N_13362,N_11588,N_11988);
xor U13363 (N_13363,N_11704,N_11253);
and U13364 (N_13364,N_11418,N_11352);
nand U13365 (N_13365,N_11378,N_11844);
or U13366 (N_13366,N_12203,N_12309);
and U13367 (N_13367,N_12097,N_11259);
nand U13368 (N_13368,N_12136,N_11842);
and U13369 (N_13369,N_12267,N_12197);
xor U13370 (N_13370,N_11864,N_11746);
xor U13371 (N_13371,N_12249,N_12226);
nand U13372 (N_13372,N_11821,N_11469);
nand U13373 (N_13373,N_12228,N_12384);
or U13374 (N_13374,N_12406,N_12161);
nor U13375 (N_13375,N_12417,N_12416);
xnor U13376 (N_13376,N_11867,N_12439);
xnor U13377 (N_13377,N_11604,N_11945);
nand U13378 (N_13378,N_11259,N_11400);
nor U13379 (N_13379,N_11996,N_12199);
and U13380 (N_13380,N_11838,N_12264);
and U13381 (N_13381,N_11489,N_11538);
xor U13382 (N_13382,N_11507,N_11610);
and U13383 (N_13383,N_12452,N_12031);
nand U13384 (N_13384,N_12423,N_11557);
or U13385 (N_13385,N_11614,N_12282);
xor U13386 (N_13386,N_12231,N_11564);
nand U13387 (N_13387,N_11261,N_11687);
nand U13388 (N_13388,N_12298,N_11851);
and U13389 (N_13389,N_11919,N_12059);
or U13390 (N_13390,N_12130,N_11447);
and U13391 (N_13391,N_12422,N_11928);
nand U13392 (N_13392,N_11536,N_11744);
xnor U13393 (N_13393,N_12005,N_11409);
xor U13394 (N_13394,N_12181,N_11882);
and U13395 (N_13395,N_12408,N_11414);
nand U13396 (N_13396,N_12028,N_11418);
nor U13397 (N_13397,N_11785,N_12295);
nor U13398 (N_13398,N_11551,N_12379);
xor U13399 (N_13399,N_11995,N_11464);
xor U13400 (N_13400,N_11919,N_11808);
or U13401 (N_13401,N_11616,N_12296);
xnor U13402 (N_13402,N_11605,N_11369);
nand U13403 (N_13403,N_11650,N_11280);
nor U13404 (N_13404,N_11528,N_11968);
or U13405 (N_13405,N_12004,N_12018);
and U13406 (N_13406,N_11492,N_12023);
or U13407 (N_13407,N_11411,N_12358);
xor U13408 (N_13408,N_12377,N_11427);
nand U13409 (N_13409,N_11271,N_11335);
xor U13410 (N_13410,N_12247,N_11355);
nor U13411 (N_13411,N_11730,N_12109);
nor U13412 (N_13412,N_12007,N_11575);
nor U13413 (N_13413,N_12206,N_11827);
or U13414 (N_13414,N_11360,N_11999);
and U13415 (N_13415,N_12407,N_11856);
or U13416 (N_13416,N_11565,N_12316);
or U13417 (N_13417,N_12236,N_11355);
or U13418 (N_13418,N_11413,N_12284);
and U13419 (N_13419,N_11321,N_11413);
xor U13420 (N_13420,N_11658,N_11503);
and U13421 (N_13421,N_12419,N_12412);
or U13422 (N_13422,N_12251,N_12115);
and U13423 (N_13423,N_11308,N_11254);
xor U13424 (N_13424,N_11840,N_11827);
and U13425 (N_13425,N_11618,N_12352);
nor U13426 (N_13426,N_12181,N_12028);
and U13427 (N_13427,N_11286,N_12319);
nor U13428 (N_13428,N_11669,N_11546);
and U13429 (N_13429,N_11474,N_11813);
or U13430 (N_13430,N_11851,N_12109);
nand U13431 (N_13431,N_11483,N_11367);
xnor U13432 (N_13432,N_11642,N_11627);
xor U13433 (N_13433,N_11328,N_11978);
or U13434 (N_13434,N_11287,N_12057);
xnor U13435 (N_13435,N_12101,N_11784);
nand U13436 (N_13436,N_12072,N_12251);
nand U13437 (N_13437,N_12140,N_12237);
and U13438 (N_13438,N_11848,N_11402);
xnor U13439 (N_13439,N_11290,N_11433);
or U13440 (N_13440,N_11625,N_11630);
and U13441 (N_13441,N_11886,N_11939);
xor U13442 (N_13442,N_12294,N_11754);
nor U13443 (N_13443,N_12269,N_11458);
nand U13444 (N_13444,N_11763,N_12474);
and U13445 (N_13445,N_12321,N_12307);
nand U13446 (N_13446,N_11502,N_11342);
xor U13447 (N_13447,N_12317,N_12353);
nor U13448 (N_13448,N_12181,N_11415);
nand U13449 (N_13449,N_12196,N_12271);
nand U13450 (N_13450,N_12202,N_11358);
or U13451 (N_13451,N_11321,N_12431);
nand U13452 (N_13452,N_12275,N_12234);
and U13453 (N_13453,N_12150,N_11394);
xnor U13454 (N_13454,N_11842,N_11308);
nand U13455 (N_13455,N_11685,N_11421);
xnor U13456 (N_13456,N_12391,N_11688);
or U13457 (N_13457,N_12467,N_12067);
xnor U13458 (N_13458,N_12392,N_12379);
or U13459 (N_13459,N_12301,N_11604);
or U13460 (N_13460,N_12135,N_11606);
nor U13461 (N_13461,N_11370,N_12094);
xnor U13462 (N_13462,N_12492,N_11841);
and U13463 (N_13463,N_11430,N_11633);
nand U13464 (N_13464,N_11842,N_12472);
xnor U13465 (N_13465,N_11684,N_11418);
xnor U13466 (N_13466,N_11455,N_11407);
xor U13467 (N_13467,N_11627,N_11768);
xor U13468 (N_13468,N_11997,N_11272);
xor U13469 (N_13469,N_11819,N_12482);
or U13470 (N_13470,N_11423,N_12278);
or U13471 (N_13471,N_12029,N_12010);
xor U13472 (N_13472,N_12272,N_11407);
nor U13473 (N_13473,N_11991,N_11351);
nand U13474 (N_13474,N_12207,N_11909);
or U13475 (N_13475,N_12310,N_12017);
and U13476 (N_13476,N_11975,N_12328);
xor U13477 (N_13477,N_11444,N_11788);
nand U13478 (N_13478,N_11288,N_12103);
xor U13479 (N_13479,N_11313,N_11662);
xnor U13480 (N_13480,N_11985,N_11928);
nor U13481 (N_13481,N_12380,N_11278);
nand U13482 (N_13482,N_11566,N_11545);
xnor U13483 (N_13483,N_12238,N_11251);
and U13484 (N_13484,N_12415,N_11661);
nor U13485 (N_13485,N_11936,N_12258);
and U13486 (N_13486,N_12348,N_11765);
xnor U13487 (N_13487,N_11943,N_11379);
nor U13488 (N_13488,N_11838,N_11395);
nor U13489 (N_13489,N_11383,N_11425);
nor U13490 (N_13490,N_12038,N_11608);
xnor U13491 (N_13491,N_11607,N_12223);
nand U13492 (N_13492,N_11934,N_11551);
xor U13493 (N_13493,N_12053,N_12304);
or U13494 (N_13494,N_12340,N_12079);
nand U13495 (N_13495,N_12126,N_11734);
or U13496 (N_13496,N_12213,N_12184);
or U13497 (N_13497,N_12153,N_12428);
nand U13498 (N_13498,N_12467,N_11649);
nor U13499 (N_13499,N_11632,N_11864);
xor U13500 (N_13500,N_12478,N_12179);
xnor U13501 (N_13501,N_12317,N_12302);
xor U13502 (N_13502,N_11608,N_11335);
nand U13503 (N_13503,N_11287,N_12352);
nand U13504 (N_13504,N_11491,N_12249);
xnor U13505 (N_13505,N_12448,N_12042);
and U13506 (N_13506,N_12127,N_11311);
nor U13507 (N_13507,N_11446,N_11518);
nand U13508 (N_13508,N_11802,N_12073);
nor U13509 (N_13509,N_12447,N_12115);
xnor U13510 (N_13510,N_12106,N_12073);
nor U13511 (N_13511,N_12034,N_12440);
and U13512 (N_13512,N_12390,N_11465);
nor U13513 (N_13513,N_11596,N_12396);
nand U13514 (N_13514,N_11479,N_12473);
and U13515 (N_13515,N_11393,N_11720);
nand U13516 (N_13516,N_11749,N_11426);
xor U13517 (N_13517,N_11702,N_11511);
nand U13518 (N_13518,N_11519,N_11970);
nand U13519 (N_13519,N_11498,N_11425);
or U13520 (N_13520,N_11489,N_12471);
nor U13521 (N_13521,N_12426,N_11314);
xor U13522 (N_13522,N_11724,N_11501);
nand U13523 (N_13523,N_11599,N_12073);
nand U13524 (N_13524,N_12432,N_11688);
or U13525 (N_13525,N_11951,N_11270);
or U13526 (N_13526,N_11485,N_11733);
nor U13527 (N_13527,N_11383,N_12115);
xnor U13528 (N_13528,N_11389,N_11724);
and U13529 (N_13529,N_12193,N_12310);
and U13530 (N_13530,N_11550,N_11600);
or U13531 (N_13531,N_11487,N_12083);
xor U13532 (N_13532,N_11529,N_12395);
and U13533 (N_13533,N_11806,N_11630);
nor U13534 (N_13534,N_11923,N_12095);
nand U13535 (N_13535,N_11744,N_12331);
nand U13536 (N_13536,N_11585,N_12144);
or U13537 (N_13537,N_11571,N_12029);
or U13538 (N_13538,N_12418,N_12298);
and U13539 (N_13539,N_11288,N_12457);
nor U13540 (N_13540,N_11832,N_11494);
and U13541 (N_13541,N_12046,N_11525);
nor U13542 (N_13542,N_12385,N_12055);
or U13543 (N_13543,N_11345,N_12287);
and U13544 (N_13544,N_12116,N_12126);
or U13545 (N_13545,N_11604,N_11795);
nor U13546 (N_13546,N_11408,N_12186);
nand U13547 (N_13547,N_11426,N_11283);
xor U13548 (N_13548,N_12127,N_11313);
or U13549 (N_13549,N_12400,N_12095);
xnor U13550 (N_13550,N_12152,N_12332);
nand U13551 (N_13551,N_12463,N_11759);
and U13552 (N_13552,N_12176,N_11641);
and U13553 (N_13553,N_11350,N_12029);
xnor U13554 (N_13554,N_11423,N_12328);
or U13555 (N_13555,N_11253,N_11817);
nor U13556 (N_13556,N_11793,N_12247);
and U13557 (N_13557,N_12382,N_11398);
and U13558 (N_13558,N_12349,N_11900);
nand U13559 (N_13559,N_12028,N_12386);
or U13560 (N_13560,N_11595,N_12131);
nor U13561 (N_13561,N_11437,N_12458);
and U13562 (N_13562,N_11458,N_12413);
xor U13563 (N_13563,N_11787,N_12367);
and U13564 (N_13564,N_11757,N_11687);
nand U13565 (N_13565,N_11359,N_11265);
and U13566 (N_13566,N_12316,N_11865);
and U13567 (N_13567,N_12189,N_11764);
nor U13568 (N_13568,N_11437,N_12320);
and U13569 (N_13569,N_12412,N_11667);
nor U13570 (N_13570,N_12398,N_12040);
xnor U13571 (N_13571,N_11441,N_11956);
nor U13572 (N_13572,N_11525,N_11603);
and U13573 (N_13573,N_11634,N_11377);
nand U13574 (N_13574,N_11727,N_11448);
xnor U13575 (N_13575,N_11356,N_12277);
nor U13576 (N_13576,N_11642,N_11382);
or U13577 (N_13577,N_11780,N_12206);
nand U13578 (N_13578,N_12471,N_11831);
nand U13579 (N_13579,N_11294,N_11943);
xor U13580 (N_13580,N_11917,N_12454);
and U13581 (N_13581,N_12217,N_12329);
nor U13582 (N_13582,N_12066,N_11828);
and U13583 (N_13583,N_11384,N_11393);
xor U13584 (N_13584,N_12385,N_12442);
xnor U13585 (N_13585,N_11347,N_11581);
xor U13586 (N_13586,N_11970,N_12425);
xnor U13587 (N_13587,N_11903,N_12018);
nand U13588 (N_13588,N_12094,N_11935);
nand U13589 (N_13589,N_11620,N_11673);
or U13590 (N_13590,N_11689,N_11980);
and U13591 (N_13591,N_11561,N_11921);
nand U13592 (N_13592,N_12020,N_12156);
or U13593 (N_13593,N_12055,N_12293);
nand U13594 (N_13594,N_11962,N_11296);
and U13595 (N_13595,N_12453,N_12168);
nand U13596 (N_13596,N_11323,N_11339);
nor U13597 (N_13597,N_11836,N_11434);
nor U13598 (N_13598,N_11413,N_11879);
or U13599 (N_13599,N_12316,N_12484);
and U13600 (N_13600,N_11690,N_11440);
nand U13601 (N_13601,N_11356,N_12320);
xnor U13602 (N_13602,N_11346,N_11890);
or U13603 (N_13603,N_11936,N_11791);
xor U13604 (N_13604,N_11341,N_11692);
nor U13605 (N_13605,N_12408,N_12010);
and U13606 (N_13606,N_12349,N_12479);
and U13607 (N_13607,N_11254,N_11733);
nand U13608 (N_13608,N_11726,N_12274);
and U13609 (N_13609,N_12009,N_11278);
nand U13610 (N_13610,N_11273,N_12470);
xor U13611 (N_13611,N_11524,N_12043);
xor U13612 (N_13612,N_11333,N_11321);
nand U13613 (N_13613,N_12486,N_11393);
nor U13614 (N_13614,N_12292,N_12249);
xor U13615 (N_13615,N_11958,N_11692);
nand U13616 (N_13616,N_12133,N_12384);
and U13617 (N_13617,N_12288,N_11669);
xor U13618 (N_13618,N_12163,N_11328);
or U13619 (N_13619,N_11907,N_11958);
or U13620 (N_13620,N_12200,N_11833);
and U13621 (N_13621,N_12051,N_12366);
nand U13622 (N_13622,N_11575,N_12146);
and U13623 (N_13623,N_11330,N_11907);
nor U13624 (N_13624,N_11714,N_12241);
and U13625 (N_13625,N_11693,N_12492);
or U13626 (N_13626,N_11516,N_11771);
or U13627 (N_13627,N_11920,N_12300);
and U13628 (N_13628,N_11977,N_12498);
xnor U13629 (N_13629,N_11681,N_11637);
or U13630 (N_13630,N_11565,N_11518);
xor U13631 (N_13631,N_11259,N_12322);
and U13632 (N_13632,N_11784,N_12262);
and U13633 (N_13633,N_11376,N_11963);
or U13634 (N_13634,N_12340,N_11324);
xor U13635 (N_13635,N_11364,N_11322);
and U13636 (N_13636,N_11480,N_11934);
xnor U13637 (N_13637,N_12001,N_11286);
xor U13638 (N_13638,N_11854,N_11280);
nor U13639 (N_13639,N_12401,N_11842);
or U13640 (N_13640,N_11300,N_11998);
nor U13641 (N_13641,N_11884,N_11879);
and U13642 (N_13642,N_12068,N_12349);
nand U13643 (N_13643,N_11825,N_11391);
xnor U13644 (N_13644,N_11884,N_12305);
xnor U13645 (N_13645,N_12196,N_11333);
nor U13646 (N_13646,N_11536,N_12069);
or U13647 (N_13647,N_12372,N_12344);
nor U13648 (N_13648,N_12273,N_11971);
and U13649 (N_13649,N_11805,N_11480);
xnor U13650 (N_13650,N_11652,N_11656);
or U13651 (N_13651,N_11510,N_12090);
nand U13652 (N_13652,N_11631,N_11679);
nand U13653 (N_13653,N_11430,N_12466);
xor U13654 (N_13654,N_11957,N_12448);
nor U13655 (N_13655,N_12389,N_11509);
nor U13656 (N_13656,N_11756,N_11950);
nor U13657 (N_13657,N_11979,N_11924);
xnor U13658 (N_13658,N_12107,N_12352);
nor U13659 (N_13659,N_11436,N_11746);
and U13660 (N_13660,N_11615,N_12295);
or U13661 (N_13661,N_12018,N_11915);
nor U13662 (N_13662,N_12213,N_12327);
or U13663 (N_13663,N_11945,N_11420);
and U13664 (N_13664,N_11869,N_11498);
or U13665 (N_13665,N_12301,N_11666);
or U13666 (N_13666,N_11916,N_11743);
and U13667 (N_13667,N_11964,N_12284);
nand U13668 (N_13668,N_11495,N_11914);
or U13669 (N_13669,N_11825,N_12443);
xor U13670 (N_13670,N_11335,N_11480);
and U13671 (N_13671,N_11455,N_12027);
nand U13672 (N_13672,N_12178,N_11427);
nand U13673 (N_13673,N_11578,N_11890);
and U13674 (N_13674,N_12470,N_12130);
xor U13675 (N_13675,N_11338,N_11923);
xnor U13676 (N_13676,N_12332,N_12104);
or U13677 (N_13677,N_11759,N_11543);
xnor U13678 (N_13678,N_11856,N_11317);
and U13679 (N_13679,N_11486,N_11549);
nand U13680 (N_13680,N_11848,N_12226);
and U13681 (N_13681,N_12099,N_12210);
xnor U13682 (N_13682,N_12088,N_11865);
nor U13683 (N_13683,N_11349,N_11523);
nor U13684 (N_13684,N_12368,N_11297);
nand U13685 (N_13685,N_11773,N_12375);
nor U13686 (N_13686,N_12075,N_11521);
nand U13687 (N_13687,N_11852,N_11483);
nor U13688 (N_13688,N_12139,N_12488);
nor U13689 (N_13689,N_11721,N_11646);
or U13690 (N_13690,N_11349,N_11935);
nand U13691 (N_13691,N_11753,N_11638);
xor U13692 (N_13692,N_12381,N_12372);
or U13693 (N_13693,N_11830,N_12254);
xor U13694 (N_13694,N_12364,N_12239);
nor U13695 (N_13695,N_11577,N_12152);
nand U13696 (N_13696,N_11391,N_12377);
xor U13697 (N_13697,N_12372,N_12414);
nand U13698 (N_13698,N_12338,N_11870);
nand U13699 (N_13699,N_12478,N_11622);
xor U13700 (N_13700,N_11943,N_11951);
and U13701 (N_13701,N_12316,N_12438);
and U13702 (N_13702,N_11519,N_12152);
nand U13703 (N_13703,N_11792,N_11625);
nand U13704 (N_13704,N_11873,N_11949);
or U13705 (N_13705,N_11542,N_12312);
or U13706 (N_13706,N_11853,N_12479);
xor U13707 (N_13707,N_11764,N_12437);
or U13708 (N_13708,N_12429,N_11281);
xnor U13709 (N_13709,N_11497,N_11256);
xnor U13710 (N_13710,N_12047,N_12194);
and U13711 (N_13711,N_12119,N_11865);
xor U13712 (N_13712,N_11492,N_11630);
and U13713 (N_13713,N_12209,N_11285);
nor U13714 (N_13714,N_11272,N_11943);
nor U13715 (N_13715,N_11976,N_11333);
xor U13716 (N_13716,N_11981,N_11308);
or U13717 (N_13717,N_11621,N_11599);
nand U13718 (N_13718,N_11263,N_11800);
xor U13719 (N_13719,N_12036,N_12333);
nand U13720 (N_13720,N_12166,N_12152);
xor U13721 (N_13721,N_12121,N_11851);
or U13722 (N_13722,N_11996,N_12084);
nand U13723 (N_13723,N_12355,N_12352);
nor U13724 (N_13724,N_11607,N_12279);
xor U13725 (N_13725,N_11462,N_12221);
nand U13726 (N_13726,N_11457,N_12306);
and U13727 (N_13727,N_11848,N_11556);
nor U13728 (N_13728,N_12319,N_11449);
nand U13729 (N_13729,N_11602,N_12250);
xnor U13730 (N_13730,N_11377,N_11437);
and U13731 (N_13731,N_12213,N_11257);
and U13732 (N_13732,N_11880,N_12497);
and U13733 (N_13733,N_12347,N_11333);
and U13734 (N_13734,N_12023,N_12048);
nand U13735 (N_13735,N_12186,N_11952);
nand U13736 (N_13736,N_11611,N_11461);
nor U13737 (N_13737,N_11856,N_11417);
xor U13738 (N_13738,N_12113,N_12327);
nor U13739 (N_13739,N_12122,N_11338);
or U13740 (N_13740,N_12108,N_11653);
and U13741 (N_13741,N_12083,N_12324);
nand U13742 (N_13742,N_11953,N_12480);
or U13743 (N_13743,N_11904,N_12368);
or U13744 (N_13744,N_12266,N_12110);
and U13745 (N_13745,N_12206,N_12055);
xnor U13746 (N_13746,N_11452,N_12375);
and U13747 (N_13747,N_11349,N_11872);
xor U13748 (N_13748,N_11519,N_12301);
nand U13749 (N_13749,N_11546,N_11297);
nor U13750 (N_13750,N_13007,N_13433);
xor U13751 (N_13751,N_12845,N_12571);
xor U13752 (N_13752,N_13147,N_13135);
and U13753 (N_13753,N_12713,N_13096);
and U13754 (N_13754,N_13390,N_13425);
and U13755 (N_13755,N_12536,N_12873);
nor U13756 (N_13756,N_13735,N_13294);
and U13757 (N_13757,N_13391,N_12519);
xor U13758 (N_13758,N_13153,N_12911);
nor U13759 (N_13759,N_12527,N_13132);
nor U13760 (N_13760,N_13671,N_12586);
nor U13761 (N_13761,N_12743,N_13033);
nor U13762 (N_13762,N_13497,N_12952);
xor U13763 (N_13763,N_12630,N_13495);
nand U13764 (N_13764,N_13193,N_12990);
or U13765 (N_13765,N_13436,N_12682);
xnor U13766 (N_13766,N_13550,N_12782);
and U13767 (N_13767,N_12705,N_12644);
or U13768 (N_13768,N_12720,N_13219);
and U13769 (N_13769,N_12589,N_13378);
nor U13770 (N_13770,N_12746,N_13694);
nor U13771 (N_13771,N_12617,N_13571);
and U13772 (N_13772,N_13612,N_13696);
nand U13773 (N_13773,N_13240,N_13343);
nor U13774 (N_13774,N_13558,N_12701);
and U13775 (N_13775,N_13261,N_13077);
xor U13776 (N_13776,N_13573,N_12723);
nor U13777 (N_13777,N_12725,N_12554);
nor U13778 (N_13778,N_12729,N_13095);
xnor U13779 (N_13779,N_12798,N_12836);
and U13780 (N_13780,N_12735,N_12807);
xnor U13781 (N_13781,N_12766,N_12711);
nand U13782 (N_13782,N_13318,N_13600);
or U13783 (N_13783,N_13282,N_12904);
nand U13784 (N_13784,N_13144,N_13145);
or U13785 (N_13785,N_13129,N_12759);
xor U13786 (N_13786,N_12956,N_12815);
nand U13787 (N_13787,N_13496,N_13723);
xnor U13788 (N_13788,N_13593,N_12728);
nor U13789 (N_13789,N_13202,N_12737);
or U13790 (N_13790,N_12906,N_13368);
xnor U13791 (N_13791,N_12754,N_12504);
and U13792 (N_13792,N_13189,N_13321);
xnor U13793 (N_13793,N_13664,N_12605);
or U13794 (N_13794,N_13310,N_13625);
nand U13795 (N_13795,N_13383,N_12539);
nor U13796 (N_13796,N_12982,N_13471);
or U13797 (N_13797,N_12581,N_13716);
nand U13798 (N_13798,N_13233,N_12667);
or U13799 (N_13799,N_12645,N_13686);
nor U13800 (N_13800,N_13708,N_13340);
xnor U13801 (N_13801,N_13181,N_13553);
nor U13802 (N_13802,N_13229,N_12913);
nor U13803 (N_13803,N_13355,N_12719);
nor U13804 (N_13804,N_13161,N_13413);
nand U13805 (N_13805,N_13268,N_12893);
nand U13806 (N_13806,N_13725,N_12840);
xor U13807 (N_13807,N_12526,N_12665);
xnor U13808 (N_13808,N_12817,N_12934);
nand U13809 (N_13809,N_12602,N_13342);
and U13810 (N_13810,N_13747,N_13247);
and U13811 (N_13811,N_13592,N_13088);
and U13812 (N_13812,N_13207,N_13498);
and U13813 (N_13813,N_12769,N_13464);
and U13814 (N_13814,N_12640,N_13692);
xor U13815 (N_13815,N_13020,N_13273);
xor U13816 (N_13816,N_12681,N_13641);
nor U13817 (N_13817,N_13512,N_13490);
nor U13818 (N_13818,N_13289,N_13002);
nand U13819 (N_13819,N_12613,N_13094);
nor U13820 (N_13820,N_12578,N_13572);
nand U13821 (N_13821,N_13414,N_13394);
nor U13822 (N_13822,N_13638,N_13618);
xor U13823 (N_13823,N_13109,N_13103);
nor U13824 (N_13824,N_13659,N_13112);
or U13825 (N_13825,N_12827,N_13595);
and U13826 (N_13826,N_12570,N_13503);
nor U13827 (N_13827,N_12594,N_12981);
nand U13828 (N_13828,N_13663,N_13691);
or U13829 (N_13829,N_13209,N_13395);
nand U13830 (N_13830,N_12622,N_12610);
xor U13831 (N_13831,N_13004,N_13203);
xor U13832 (N_13832,N_12727,N_12888);
and U13833 (N_13833,N_12706,N_13622);
nand U13834 (N_13834,N_13645,N_12755);
nand U13835 (N_13835,N_13393,N_13700);
and U13836 (N_13836,N_13005,N_13561);
or U13837 (N_13837,N_12661,N_13734);
nand U13838 (N_13838,N_12511,N_13339);
nor U13839 (N_13839,N_13200,N_13257);
or U13840 (N_13840,N_12968,N_13741);
nor U13841 (N_13841,N_12524,N_13110);
nor U13842 (N_13842,N_12812,N_12659);
nor U13843 (N_13843,N_12700,N_12903);
xor U13844 (N_13844,N_12690,N_13420);
xor U13845 (N_13845,N_12677,N_13398);
and U13846 (N_13846,N_13465,N_13720);
nand U13847 (N_13847,N_13055,N_13548);
or U13848 (N_13848,N_13250,N_13400);
xor U13849 (N_13849,N_12621,N_13479);
nand U13850 (N_13850,N_13246,N_13149);
xnor U13851 (N_13851,N_12916,N_13107);
nand U13852 (N_13852,N_12804,N_12612);
xnor U13853 (N_13853,N_12859,N_13260);
and U13854 (N_13854,N_13669,N_13124);
nor U13855 (N_13855,N_13026,N_12865);
nor U13856 (N_13856,N_13565,N_13141);
nand U13857 (N_13857,N_12939,N_12533);
and U13858 (N_13858,N_13048,N_12799);
xnor U13859 (N_13859,N_13163,N_13045);
nor U13860 (N_13860,N_12598,N_13627);
nand U13861 (N_13861,N_13348,N_13482);
nor U13862 (N_13862,N_12978,N_13080);
nor U13863 (N_13863,N_12858,N_13346);
and U13864 (N_13864,N_12707,N_13293);
nand U13865 (N_13865,N_12693,N_12940);
nand U13866 (N_13866,N_12717,N_13316);
and U13867 (N_13867,N_13381,N_12509);
nor U13868 (N_13868,N_13644,N_13427);
xnor U13869 (N_13869,N_12877,N_13486);
nor U13870 (N_13870,N_13173,N_13411);
nand U13871 (N_13871,N_13320,N_13577);
xnor U13872 (N_13872,N_12558,N_13643);
xnor U13873 (N_13873,N_13126,N_13673);
nand U13874 (N_13874,N_12672,N_13234);
nand U13875 (N_13875,N_13035,N_13705);
xnor U13876 (N_13876,N_12999,N_12662);
nand U13877 (N_13877,N_12569,N_12651);
nand U13878 (N_13878,N_13501,N_13102);
and U13879 (N_13879,N_13249,N_12547);
xor U13880 (N_13880,N_13265,N_13041);
and U13881 (N_13881,N_12931,N_12738);
nand U13882 (N_13882,N_13211,N_13204);
nor U13883 (N_13883,N_13443,N_13067);
or U13884 (N_13884,N_13043,N_13419);
and U13885 (N_13885,N_13054,N_12748);
xor U13886 (N_13886,N_13730,N_13307);
nor U13887 (N_13887,N_12574,N_12673);
and U13888 (N_13888,N_13380,N_13605);
xor U13889 (N_13889,N_13507,N_12830);
xor U13890 (N_13890,N_12878,N_12823);
or U13891 (N_13891,N_13567,N_13746);
nor U13892 (N_13892,N_12587,N_13323);
xnor U13893 (N_13893,N_12715,N_12795);
nand U13894 (N_13894,N_13025,N_12953);
nand U13895 (N_13895,N_13668,N_13210);
nand U13896 (N_13896,N_13376,N_13500);
or U13897 (N_13897,N_12943,N_13629);
nor U13898 (N_13898,N_12584,N_12801);
or U13899 (N_13899,N_12508,N_12559);
nand U13900 (N_13900,N_12819,N_13016);
xor U13901 (N_13901,N_13604,N_13442);
or U13902 (N_13902,N_12638,N_12593);
xnor U13903 (N_13903,N_13559,N_13712);
nand U13904 (N_13904,N_12868,N_13703);
or U13905 (N_13905,N_12550,N_13542);
or U13906 (N_13906,N_12698,N_13356);
nand U13907 (N_13907,N_13366,N_13676);
xor U13908 (N_13908,N_13201,N_13177);
and U13909 (N_13909,N_12994,N_13475);
xnor U13910 (N_13910,N_13682,N_13529);
and U13911 (N_13911,N_12803,N_13483);
or U13912 (N_13912,N_12595,N_13502);
nand U13913 (N_13913,N_13586,N_12641);
xor U13914 (N_13914,N_12933,N_13369);
xnor U13915 (N_13915,N_13259,N_12542);
nor U13916 (N_13916,N_13737,N_13707);
xor U13917 (N_13917,N_13563,N_13402);
xor U13918 (N_13918,N_12575,N_13008);
xnor U13919 (N_13919,N_13373,N_12747);
nor U13920 (N_13920,N_12518,N_12902);
and U13921 (N_13921,N_12632,N_13727);
xnor U13922 (N_13922,N_13587,N_13040);
and U13923 (N_13923,N_13736,N_13424);
and U13924 (N_13924,N_13162,N_13679);
nand U13925 (N_13925,N_13560,N_12709);
xnor U13926 (N_13926,N_13030,N_12631);
nand U13927 (N_13927,N_13151,N_13171);
nand U13928 (N_13928,N_12629,N_13416);
xor U13929 (N_13929,N_13185,N_13142);
xor U13930 (N_13930,N_12771,N_12660);
nand U13931 (N_13931,N_12826,N_12973);
and U13932 (N_13932,N_13687,N_12699);
or U13933 (N_13933,N_12988,N_13570);
nand U13934 (N_13934,N_13311,N_12505);
or U13935 (N_13935,N_12867,N_13387);
nor U13936 (N_13936,N_13731,N_13599);
and U13937 (N_13937,N_13389,N_13699);
and U13938 (N_13938,N_13410,N_12643);
xor U13939 (N_13939,N_12576,N_12653);
nand U13940 (N_13940,N_13444,N_13613);
xnor U13941 (N_13941,N_12758,N_13401);
nor U13942 (N_13942,N_12680,N_12927);
xnor U13943 (N_13943,N_13066,N_13574);
xnor U13944 (N_13944,N_13062,N_13590);
and U13945 (N_13945,N_13295,N_13286);
and U13946 (N_13946,N_13452,N_13421);
nand U13947 (N_13947,N_12566,N_13336);
and U13948 (N_13948,N_13217,N_12765);
xnor U13949 (N_13949,N_12831,N_12742);
and U13950 (N_13950,N_12712,N_13639);
xor U13951 (N_13951,N_13205,N_13218);
nand U13952 (N_13952,N_12532,N_13438);
xor U13953 (N_13953,N_12863,N_13078);
nor U13954 (N_13954,N_13722,N_13683);
and U13955 (N_13955,N_12838,N_13404);
nor U13956 (N_13956,N_12548,N_13271);
xor U13957 (N_13957,N_13059,N_13596);
and U13958 (N_13958,N_12549,N_12676);
or U13959 (N_13959,N_13417,N_12557);
nor U13960 (N_13960,N_13408,N_13199);
or U13961 (N_13961,N_13693,N_13430);
nor U13962 (N_13962,N_13509,N_13674);
and U13963 (N_13963,N_13034,N_13037);
and U13964 (N_13964,N_13540,N_13685);
xnor U13965 (N_13965,N_12851,N_13051);
or U13966 (N_13966,N_12962,N_12787);
xnor U13967 (N_13967,N_13384,N_13583);
nor U13968 (N_13968,N_12828,N_13224);
xnor U13969 (N_13969,N_13702,N_13511);
xnor U13970 (N_13970,N_12960,N_13350);
nand U13971 (N_13971,N_13491,N_13481);
nor U13972 (N_13972,N_12683,N_13531);
xor U13973 (N_13973,N_13654,N_13517);
nand U13974 (N_13974,N_13704,N_13695);
nand U13975 (N_13975,N_12618,N_13620);
nand U13976 (N_13976,N_12503,N_13575);
nand U13977 (N_13977,N_12739,N_12507);
nand U13978 (N_13978,N_13049,N_13183);
and U13979 (N_13979,N_13354,N_13283);
nor U13980 (N_13980,N_12937,N_13023);
and U13981 (N_13981,N_12780,N_12615);
and U13982 (N_13982,N_13182,N_13729);
nor U13983 (N_13983,N_13225,N_13473);
and U13984 (N_13984,N_13235,N_13073);
and U13985 (N_13985,N_13174,N_12976);
xnor U13986 (N_13986,N_13603,N_13415);
xnor U13987 (N_13987,N_12567,N_13140);
or U13988 (N_13988,N_12875,N_13630);
xor U13989 (N_13989,N_13285,N_13435);
nand U13990 (N_13990,N_13422,N_12984);
xor U13991 (N_13991,N_12991,N_13352);
nor U13992 (N_13992,N_13423,N_12761);
and U13993 (N_13993,N_13290,N_12871);
xnor U13994 (N_13994,N_13636,N_12963);
nand U13995 (N_13995,N_13278,N_13231);
xor U13996 (N_13996,N_12920,N_12521);
nand U13997 (N_13997,N_12704,N_12750);
nand U13998 (N_13998,N_13510,N_13439);
xnor U13999 (N_13999,N_12540,N_12797);
or U14000 (N_14000,N_13370,N_13098);
and U14001 (N_14001,N_13585,N_12919);
and U14002 (N_14002,N_12995,N_13166);
or U14003 (N_14003,N_13714,N_12535);
or U14004 (N_14004,N_13546,N_12773);
nand U14005 (N_14005,N_13226,N_13221);
or U14006 (N_14006,N_12918,N_12620);
or U14007 (N_14007,N_13099,N_12987);
nor U14008 (N_14008,N_12914,N_13480);
and U14009 (N_14009,N_13215,N_12512);
xnor U14010 (N_14010,N_12796,N_13656);
nand U14011 (N_14011,N_12652,N_13313);
nor U14012 (N_14012,N_13065,N_13287);
nand U14013 (N_14013,N_12718,N_12627);
nor U14014 (N_14014,N_13309,N_12528);
and U14015 (N_14015,N_12910,N_12543);
xnor U14016 (N_14016,N_13003,N_13168);
xnor U14017 (N_14017,N_13184,N_12948);
or U14018 (N_14018,N_13544,N_13169);
and U14019 (N_14019,N_13076,N_13709);
nand U14020 (N_14020,N_13523,N_13634);
xnor U14021 (N_14021,N_12970,N_12545);
and U14022 (N_14022,N_12697,N_13114);
nand U14023 (N_14023,N_13091,N_12730);
nor U14024 (N_14024,N_13052,N_13602);
or U14025 (N_14025,N_12912,N_13374);
or U14026 (N_14026,N_12614,N_13305);
or U14027 (N_14027,N_13158,N_12998);
nor U14028 (N_14028,N_12696,N_13324);
xnor U14029 (N_14029,N_13506,N_13533);
xor U14030 (N_14030,N_13057,N_12997);
nor U14031 (N_14031,N_13392,N_13299);
nand U14032 (N_14032,N_12928,N_13665);
or U14033 (N_14033,N_12800,N_13453);
and U14034 (N_14034,N_13155,N_12552);
or U14035 (N_14035,N_13713,N_13063);
and U14036 (N_14036,N_13056,N_12789);
nand U14037 (N_14037,N_13176,N_13172);
nor U14038 (N_14038,N_12992,N_13397);
nor U14039 (N_14039,N_12942,N_13266);
or U14040 (N_14040,N_13554,N_12885);
nor U14041 (N_14041,N_12702,N_13027);
and U14042 (N_14042,N_12961,N_13079);
and U14043 (N_14043,N_13578,N_13270);
and U14044 (N_14044,N_13363,N_13661);
or U14045 (N_14045,N_13418,N_13469);
nor U14046 (N_14046,N_13127,N_12657);
and U14047 (N_14047,N_13576,N_12608);
nor U14048 (N_14048,N_13032,N_12733);
nand U14049 (N_14049,N_12861,N_12710);
or U14050 (N_14050,N_13726,N_12517);
nand U14051 (N_14051,N_13082,N_12779);
nand U14052 (N_14052,N_12772,N_12784);
and U14053 (N_14053,N_13749,N_12989);
or U14054 (N_14054,N_12929,N_13101);
xnor U14055 (N_14055,N_12694,N_13616);
nand U14056 (N_14056,N_12749,N_12882);
nand U14057 (N_14057,N_12901,N_13262);
nor U14058 (N_14058,N_12597,N_13120);
or U14059 (N_14059,N_13549,N_13615);
or U14060 (N_14060,N_12808,N_13635);
nand U14061 (N_14061,N_12624,N_13123);
or U14062 (N_14062,N_12930,N_13297);
or U14063 (N_14063,N_13388,N_12506);
xnor U14064 (N_14064,N_13637,N_13308);
nor U14065 (N_14065,N_13006,N_13118);
nand U14066 (N_14066,N_13489,N_13721);
nand U14067 (N_14067,N_13300,N_13432);
nand U14068 (N_14068,N_12588,N_12553);
and U14069 (N_14069,N_12513,N_13198);
xor U14070 (N_14070,N_12932,N_13197);
and U14071 (N_14071,N_13655,N_13684);
nor U14072 (N_14072,N_13000,N_13125);
and U14073 (N_14073,N_12607,N_13180);
nand U14074 (N_14074,N_12609,N_12825);
or U14075 (N_14075,N_13680,N_13108);
xor U14076 (N_14076,N_13191,N_12726);
or U14077 (N_14077,N_13719,N_12670);
and U14078 (N_14078,N_12894,N_12688);
or U14079 (N_14079,N_12977,N_12949);
nand U14080 (N_14080,N_13322,N_13351);
or U14081 (N_14081,N_13557,N_12896);
nand U14082 (N_14082,N_12854,N_12834);
xnor U14083 (N_14083,N_13396,N_13681);
nor U14084 (N_14084,N_13284,N_12767);
or U14085 (N_14085,N_13449,N_13254);
or U14086 (N_14086,N_13434,N_13164);
nor U14087 (N_14087,N_13357,N_13196);
nor U14088 (N_14088,N_13068,N_12568);
and U14089 (N_14089,N_12551,N_13190);
or U14090 (N_14090,N_13640,N_13532);
nor U14091 (N_14091,N_12900,N_13441);
xnor U14092 (N_14092,N_13539,N_13446);
and U14093 (N_14093,N_13188,N_13258);
or U14094 (N_14094,N_13632,N_13515);
or U14095 (N_14095,N_13711,N_12611);
or U14096 (N_14096,N_13238,N_12664);
or U14097 (N_14097,N_12541,N_13521);
nand U14098 (N_14098,N_13334,N_12768);
xor U14099 (N_14099,N_13678,N_12975);
nand U14100 (N_14100,N_13535,N_12646);
nor U14101 (N_14101,N_12908,N_13304);
nor U14102 (N_14102,N_13150,N_12879);
and U14103 (N_14103,N_12841,N_13508);
nor U14104 (N_14104,N_13677,N_13071);
and U14105 (N_14105,N_13484,N_12855);
nor U14106 (N_14106,N_12634,N_13360);
nor U14107 (N_14107,N_13089,N_13454);
and U14108 (N_14108,N_12510,N_13298);
nor U14109 (N_14109,N_12866,N_13044);
nor U14110 (N_14110,N_12616,N_12502);
or U14111 (N_14111,N_13038,N_13156);
nor U14112 (N_14112,N_13302,N_13347);
and U14113 (N_14113,N_12674,N_12721);
nand U14114 (N_14114,N_13013,N_13328);
xor U14115 (N_14115,N_12781,N_13488);
nor U14116 (N_14116,N_13545,N_13117);
nor U14117 (N_14117,N_13021,N_13522);
nand U14118 (N_14118,N_13628,N_13462);
xor U14119 (N_14119,N_12955,N_13236);
and U14120 (N_14120,N_13241,N_13146);
and U14121 (N_14121,N_12760,N_12647);
and U14122 (N_14122,N_13216,N_13519);
and U14123 (N_14123,N_13303,N_12501);
xnor U14124 (N_14124,N_13649,N_13213);
or U14125 (N_14125,N_12816,N_12560);
xor U14126 (N_14126,N_13743,N_12935);
and U14127 (N_14127,N_13251,N_13119);
nand U14128 (N_14128,N_13459,N_13256);
nand U14129 (N_14129,N_12666,N_13195);
xor U14130 (N_14130,N_12687,N_13551);
nand U14131 (N_14131,N_13223,N_13105);
xor U14132 (N_14132,N_12778,N_13745);
nand U14133 (N_14133,N_12898,N_13252);
or U14134 (N_14134,N_13122,N_12764);
xnor U14135 (N_14135,N_13154,N_12907);
nor U14136 (N_14136,N_13648,N_13279);
xnor U14137 (N_14137,N_13019,N_12870);
nand U14138 (N_14138,N_12599,N_12722);
and U14139 (N_14139,N_12658,N_12923);
nand U14140 (N_14140,N_13242,N_13706);
nor U14141 (N_14141,N_12774,N_12947);
nor U14142 (N_14142,N_13428,N_13740);
nand U14143 (N_14143,N_12964,N_12529);
xnor U14144 (N_14144,N_13513,N_13160);
nor U14145 (N_14145,N_12969,N_12600);
xor U14146 (N_14146,N_13106,N_12635);
xor U14147 (N_14147,N_12966,N_13072);
xnor U14148 (N_14148,N_13010,N_12892);
and U14149 (N_14149,N_13333,N_13710);
nand U14150 (N_14150,N_12573,N_13569);
nor U14151 (N_14151,N_12785,N_12751);
xnor U14152 (N_14152,N_12736,N_13461);
nand U14153 (N_14153,N_12835,N_13028);
nand U14154 (N_14154,N_13385,N_13371);
nor U14155 (N_14155,N_12983,N_13058);
xnor U14156 (N_14156,N_12520,N_12703);
nand U14157 (N_14157,N_13597,N_13212);
nor U14158 (N_14158,N_13619,N_12788);
nand U14159 (N_14159,N_12818,N_12564);
or U14160 (N_14160,N_13437,N_12957);
nor U14161 (N_14161,N_13598,N_13525);
nor U14162 (N_14162,N_13301,N_12996);
and U14163 (N_14163,N_13275,N_13601);
nand U14164 (N_14164,N_13192,N_12864);
nor U14165 (N_14165,N_13607,N_13591);
or U14166 (N_14166,N_13412,N_12663);
and U14167 (N_14167,N_13253,N_13450);
and U14168 (N_14168,N_13042,N_13291);
nand U14169 (N_14169,N_13315,N_13748);
or U14170 (N_14170,N_13296,N_13097);
or U14171 (N_14171,N_13335,N_13022);
nand U14172 (N_14172,N_13670,N_12905);
nand U14173 (N_14173,N_13232,N_13012);
or U14174 (N_14174,N_13060,N_13326);
or U14175 (N_14175,N_12656,N_12824);
nand U14176 (N_14176,N_12791,N_13594);
or U14177 (N_14177,N_13227,N_13514);
and U14178 (N_14178,N_13739,N_13175);
xnor U14179 (N_14179,N_13222,N_12856);
and U14180 (N_14180,N_13157,N_13248);
nand U14181 (N_14181,N_13582,N_13306);
xor U14182 (N_14182,N_13092,N_13447);
and U14183 (N_14183,N_13194,N_12924);
nand U14184 (N_14184,N_12886,N_13332);
or U14185 (N_14185,N_13552,N_12887);
nand U14186 (N_14186,N_13470,N_12980);
nand U14187 (N_14187,N_13505,N_12654);
or U14188 (N_14188,N_13431,N_13588);
xor U14189 (N_14189,N_13319,N_12649);
xor U14190 (N_14190,N_12809,N_12740);
or U14191 (N_14191,N_12692,N_12897);
xor U14192 (N_14192,N_12745,N_12850);
or U14193 (N_14193,N_13472,N_13667);
or U14194 (N_14194,N_13646,N_12921);
and U14195 (N_14195,N_13379,N_13349);
or U14196 (N_14196,N_13492,N_13093);
xnor U14197 (N_14197,N_13264,N_13086);
and U14198 (N_14198,N_12691,N_13167);
and U14199 (N_14199,N_12708,N_13139);
nor U14200 (N_14200,N_13015,N_13104);
nand U14201 (N_14201,N_12849,N_13128);
or U14202 (N_14202,N_13527,N_12744);
and U14203 (N_14203,N_13621,N_13317);
xor U14204 (N_14204,N_12585,N_13466);
nand U14205 (N_14205,N_13014,N_12872);
nand U14206 (N_14206,N_12793,N_13455);
and U14207 (N_14207,N_12986,N_12639);
nand U14208 (N_14208,N_13715,N_13467);
nor U14209 (N_14209,N_12514,N_12731);
nor U14210 (N_14210,N_13130,N_13244);
and U14211 (N_14211,N_12689,N_13362);
xnor U14212 (N_14212,N_13624,N_13672);
and U14213 (N_14213,N_12794,N_13243);
or U14214 (N_14214,N_12899,N_12805);
nor U14215 (N_14215,N_12917,N_12876);
nand U14216 (N_14216,N_13485,N_12786);
nand U14217 (N_14217,N_12626,N_12813);
xor U14218 (N_14218,N_13372,N_13272);
nand U14219 (N_14219,N_13345,N_12883);
xor U14220 (N_14220,N_12844,N_12579);
or U14221 (N_14221,N_13353,N_13732);
xor U14222 (N_14222,N_12926,N_12842);
xnor U14223 (N_14223,N_12770,N_13170);
nand U14224 (N_14224,N_12974,N_13090);
or U14225 (N_14225,N_13724,N_12783);
nor U14226 (N_14226,N_13288,N_12633);
xor U14227 (N_14227,N_12941,N_12814);
nor U14228 (N_14228,N_13083,N_13543);
nor U14229 (N_14229,N_13115,N_12846);
nand U14230 (N_14230,N_13657,N_13516);
and U14231 (N_14231,N_13133,N_12822);
xnor U14232 (N_14232,N_13245,N_13658);
nand U14233 (N_14233,N_13113,N_13136);
and U14234 (N_14234,N_12839,N_12909);
xor U14235 (N_14235,N_12732,N_13220);
xnor U14236 (N_14236,N_13487,N_13579);
nand U14237 (N_14237,N_12648,N_13566);
xnor U14238 (N_14238,N_12577,N_13738);
xnor U14239 (N_14239,N_13581,N_13623);
and U14240 (N_14240,N_12555,N_13409);
xnor U14241 (N_14241,N_12678,N_13642);
or U14242 (N_14242,N_13292,N_12592);
xnor U14243 (N_14243,N_13239,N_12837);
or U14244 (N_14244,N_12946,N_13688);
nand U14245 (N_14245,N_13405,N_12958);
xnor U14246 (N_14246,N_13580,N_13001);
or U14247 (N_14247,N_13518,N_13460);
nor U14248 (N_14248,N_12762,N_12884);
nand U14249 (N_14249,N_12852,N_13276);
and U14250 (N_14250,N_13018,N_13137);
or U14251 (N_14251,N_12843,N_12874);
or U14252 (N_14252,N_13403,N_13609);
xnor U14253 (N_14253,N_12860,N_12675);
xnor U14254 (N_14254,N_13267,N_13152);
or U14255 (N_14255,N_13457,N_12583);
and U14256 (N_14256,N_12582,N_13650);
nand U14257 (N_14257,N_12596,N_13331);
or U14258 (N_14258,N_12833,N_13131);
and U14259 (N_14259,N_12716,N_13478);
nor U14260 (N_14260,N_12679,N_12776);
xnor U14261 (N_14261,N_13338,N_12763);
or U14262 (N_14262,N_13399,N_12938);
or U14263 (N_14263,N_12636,N_12810);
nor U14264 (N_14264,N_13186,N_12625);
nor U14265 (N_14265,N_12891,N_12811);
nor U14266 (N_14266,N_13728,N_12869);
nor U14267 (N_14267,N_12538,N_13382);
nor U14268 (N_14268,N_13476,N_13230);
and U14269 (N_14269,N_13365,N_13662);
nand U14270 (N_14270,N_12847,N_13237);
and U14271 (N_14271,N_12628,N_13329);
and U14272 (N_14272,N_13214,N_12790);
nand U14273 (N_14273,N_12853,N_12525);
nor U14274 (N_14274,N_13359,N_13036);
and U14275 (N_14275,N_12944,N_12848);
or U14276 (N_14276,N_13589,N_13024);
or U14277 (N_14277,N_13451,N_13074);
or U14278 (N_14278,N_13228,N_13556);
nand U14279 (N_14279,N_12590,N_13718);
and U14280 (N_14280,N_13187,N_12637);
nand U14281 (N_14281,N_12734,N_13653);
or U14282 (N_14282,N_13584,N_12523);
nand U14283 (N_14283,N_13358,N_13406);
nand U14284 (N_14284,N_12515,N_13504);
nand U14285 (N_14285,N_12563,N_13468);
nand U14286 (N_14286,N_12655,N_13337);
or U14287 (N_14287,N_13555,N_13047);
and U14288 (N_14288,N_12603,N_13263);
xor U14289 (N_14289,N_13697,N_13341);
nor U14290 (N_14290,N_13081,N_12959);
nor U14291 (N_14291,N_13690,N_13327);
and U14292 (N_14292,N_13009,N_13330);
nand U14293 (N_14293,N_12880,N_12752);
or U14294 (N_14294,N_13562,N_13536);
and U14295 (N_14295,N_12642,N_13280);
xnor U14296 (N_14296,N_13547,N_12945);
or U14297 (N_14297,N_12829,N_13717);
nor U14298 (N_14298,N_13617,N_13138);
nand U14299 (N_14299,N_13344,N_12965);
and U14300 (N_14300,N_13477,N_13029);
nand U14301 (N_14301,N_12686,N_13742);
or U14302 (N_14302,N_13698,N_13143);
or U14303 (N_14303,N_12922,N_13528);
nor U14304 (N_14304,N_12516,N_13524);
nor U14305 (N_14305,N_12685,N_13701);
xnor U14306 (N_14306,N_13116,N_13568);
or U14307 (N_14307,N_12562,N_13429);
nand U14308 (N_14308,N_12695,N_13312);
xor U14309 (N_14309,N_13611,N_12669);
nor U14310 (N_14310,N_12775,N_12522);
xnor U14311 (N_14311,N_13085,N_12757);
or U14312 (N_14312,N_13651,N_13610);
nor U14313 (N_14313,N_13314,N_12950);
xnor U14314 (N_14314,N_12993,N_13325);
xnor U14315 (N_14315,N_12580,N_13064);
or U14316 (N_14316,N_12971,N_13277);
xor U14317 (N_14317,N_13631,N_12756);
or U14318 (N_14318,N_12936,N_13608);
or U14319 (N_14319,N_13255,N_12967);
nor U14320 (N_14320,N_13011,N_12604);
and U14321 (N_14321,N_13606,N_12561);
xor U14322 (N_14322,N_13053,N_13538);
nand U14323 (N_14323,N_13017,N_13520);
or U14324 (N_14324,N_12544,N_12777);
nand U14325 (N_14325,N_12862,N_13534);
nor U14326 (N_14326,N_12530,N_12890);
nor U14327 (N_14327,N_13061,N_12714);
and U14328 (N_14328,N_13031,N_13208);
or U14329 (N_14329,N_13165,N_13386);
or U14330 (N_14330,N_13361,N_12951);
or U14331 (N_14331,N_12925,N_13274);
and U14332 (N_14332,N_13647,N_13046);
or U14333 (N_14333,N_13069,N_13526);
xnor U14334 (N_14334,N_13474,N_12623);
nand U14335 (N_14335,N_13499,N_13426);
or U14336 (N_14336,N_12537,N_13364);
and U14337 (N_14337,N_13458,N_12619);
or U14338 (N_14338,N_12591,N_12792);
nand U14339 (N_14339,N_13689,N_12972);
or U14340 (N_14340,N_12724,N_13463);
nor U14341 (N_14341,N_12979,N_13179);
xnor U14342 (N_14342,N_12820,N_13134);
and U14343 (N_14343,N_13070,N_13564);
or U14344 (N_14344,N_12546,N_13448);
and U14345 (N_14345,N_13541,N_13614);
or U14346 (N_14346,N_13075,N_12741);
and U14347 (N_14347,N_13744,N_12650);
xnor U14348 (N_14348,N_13626,N_12915);
nand U14349 (N_14349,N_12500,N_13407);
nand U14350 (N_14350,N_13159,N_13440);
and U14351 (N_14351,N_13100,N_13050);
xor U14352 (N_14352,N_12753,N_13675);
xor U14353 (N_14353,N_12556,N_13087);
or U14354 (N_14354,N_12565,N_12806);
and U14355 (N_14355,N_12601,N_13084);
and U14356 (N_14356,N_12534,N_13660);
nand U14357 (N_14357,N_13733,N_13375);
xor U14358 (N_14358,N_13666,N_13039);
or U14359 (N_14359,N_13494,N_13633);
and U14360 (N_14360,N_13445,N_13269);
xor U14361 (N_14361,N_12832,N_12802);
xor U14362 (N_14362,N_13121,N_13206);
xor U14363 (N_14363,N_13178,N_12985);
or U14364 (N_14364,N_12821,N_12572);
or U14365 (N_14365,N_13456,N_13111);
or U14366 (N_14366,N_12606,N_12954);
nand U14367 (N_14367,N_12881,N_13493);
xnor U14368 (N_14368,N_13377,N_12684);
nor U14369 (N_14369,N_13367,N_12531);
nand U14370 (N_14370,N_13281,N_13537);
nand U14371 (N_14371,N_13148,N_13652);
or U14372 (N_14372,N_13530,N_12857);
nand U14373 (N_14373,N_12895,N_12889);
or U14374 (N_14374,N_12668,N_12671);
xor U14375 (N_14375,N_12897,N_13698);
nand U14376 (N_14376,N_12583,N_13404);
xor U14377 (N_14377,N_12527,N_13099);
nor U14378 (N_14378,N_13734,N_13404);
nand U14379 (N_14379,N_13393,N_13376);
nand U14380 (N_14380,N_12755,N_12836);
nand U14381 (N_14381,N_13040,N_12735);
or U14382 (N_14382,N_12911,N_12525);
or U14383 (N_14383,N_13113,N_13000);
xnor U14384 (N_14384,N_12959,N_13171);
nand U14385 (N_14385,N_13315,N_13428);
xnor U14386 (N_14386,N_13612,N_13014);
or U14387 (N_14387,N_12757,N_12532);
nor U14388 (N_14388,N_13226,N_13020);
and U14389 (N_14389,N_12567,N_12598);
xnor U14390 (N_14390,N_12992,N_13509);
or U14391 (N_14391,N_13354,N_13306);
or U14392 (N_14392,N_13407,N_13538);
nand U14393 (N_14393,N_12872,N_13352);
xor U14394 (N_14394,N_13288,N_13606);
or U14395 (N_14395,N_13379,N_12637);
and U14396 (N_14396,N_13033,N_12784);
nor U14397 (N_14397,N_13254,N_13607);
nand U14398 (N_14398,N_12797,N_13502);
nor U14399 (N_14399,N_13440,N_13061);
xor U14400 (N_14400,N_13195,N_13031);
and U14401 (N_14401,N_13136,N_12595);
and U14402 (N_14402,N_12977,N_13183);
and U14403 (N_14403,N_12644,N_13008);
nand U14404 (N_14404,N_13082,N_12949);
xnor U14405 (N_14405,N_12900,N_13247);
xnor U14406 (N_14406,N_12508,N_13199);
xor U14407 (N_14407,N_13565,N_12562);
nor U14408 (N_14408,N_13232,N_13390);
nand U14409 (N_14409,N_13253,N_13601);
nor U14410 (N_14410,N_13061,N_12542);
or U14411 (N_14411,N_13651,N_12995);
xor U14412 (N_14412,N_12878,N_12985);
and U14413 (N_14413,N_13123,N_12939);
or U14414 (N_14414,N_13540,N_13015);
nand U14415 (N_14415,N_13477,N_13347);
nand U14416 (N_14416,N_13272,N_13416);
nand U14417 (N_14417,N_12692,N_12910);
and U14418 (N_14418,N_13371,N_12582);
nor U14419 (N_14419,N_12727,N_12968);
nand U14420 (N_14420,N_12588,N_12604);
and U14421 (N_14421,N_12604,N_13278);
and U14422 (N_14422,N_13274,N_12944);
xnor U14423 (N_14423,N_13564,N_13630);
nand U14424 (N_14424,N_12832,N_13064);
or U14425 (N_14425,N_12779,N_13302);
nor U14426 (N_14426,N_13337,N_12909);
or U14427 (N_14427,N_13553,N_13529);
or U14428 (N_14428,N_12778,N_13452);
xnor U14429 (N_14429,N_12897,N_13629);
nand U14430 (N_14430,N_13538,N_13482);
nand U14431 (N_14431,N_13166,N_13147);
nor U14432 (N_14432,N_13537,N_12738);
xnor U14433 (N_14433,N_12988,N_13538);
xor U14434 (N_14434,N_13637,N_12868);
nand U14435 (N_14435,N_12658,N_12666);
and U14436 (N_14436,N_13715,N_13738);
or U14437 (N_14437,N_13151,N_13080);
and U14438 (N_14438,N_13118,N_12990);
xnor U14439 (N_14439,N_12724,N_12909);
or U14440 (N_14440,N_12641,N_12983);
nor U14441 (N_14441,N_13124,N_13227);
nand U14442 (N_14442,N_13609,N_13728);
or U14443 (N_14443,N_12745,N_13475);
nor U14444 (N_14444,N_13726,N_12837);
xnor U14445 (N_14445,N_13289,N_13038);
or U14446 (N_14446,N_12821,N_12504);
and U14447 (N_14447,N_12837,N_13410);
nand U14448 (N_14448,N_13608,N_12848);
xor U14449 (N_14449,N_12517,N_13481);
and U14450 (N_14450,N_12598,N_13146);
nand U14451 (N_14451,N_12744,N_13030);
nor U14452 (N_14452,N_13638,N_12880);
and U14453 (N_14453,N_13046,N_12778);
nor U14454 (N_14454,N_13546,N_13180);
or U14455 (N_14455,N_12976,N_13238);
and U14456 (N_14456,N_13479,N_13396);
and U14457 (N_14457,N_13213,N_12983);
or U14458 (N_14458,N_13258,N_13210);
or U14459 (N_14459,N_13303,N_12600);
nor U14460 (N_14460,N_13004,N_13502);
xnor U14461 (N_14461,N_13330,N_13225);
nand U14462 (N_14462,N_13346,N_13232);
xnor U14463 (N_14463,N_13358,N_12930);
nand U14464 (N_14464,N_12931,N_13192);
nand U14465 (N_14465,N_13211,N_13151);
nor U14466 (N_14466,N_13546,N_13693);
or U14467 (N_14467,N_12696,N_13413);
xnor U14468 (N_14468,N_13497,N_12999);
or U14469 (N_14469,N_13567,N_13108);
nand U14470 (N_14470,N_12853,N_12828);
or U14471 (N_14471,N_13432,N_12540);
xor U14472 (N_14472,N_13306,N_12590);
nand U14473 (N_14473,N_13631,N_13669);
nand U14474 (N_14474,N_12617,N_12678);
nor U14475 (N_14475,N_12839,N_12798);
nor U14476 (N_14476,N_13433,N_12938);
and U14477 (N_14477,N_13400,N_13706);
nor U14478 (N_14478,N_13150,N_12909);
nand U14479 (N_14479,N_12789,N_13410);
nor U14480 (N_14480,N_12738,N_13313);
xor U14481 (N_14481,N_12870,N_13641);
or U14482 (N_14482,N_13003,N_13072);
xor U14483 (N_14483,N_12562,N_13591);
or U14484 (N_14484,N_13387,N_12983);
nand U14485 (N_14485,N_12639,N_13468);
or U14486 (N_14486,N_12945,N_13029);
xor U14487 (N_14487,N_12835,N_13442);
and U14488 (N_14488,N_13721,N_13127);
and U14489 (N_14489,N_13446,N_13707);
nand U14490 (N_14490,N_12578,N_13237);
and U14491 (N_14491,N_12752,N_13352);
xor U14492 (N_14492,N_13496,N_13318);
nand U14493 (N_14493,N_13248,N_12531);
nand U14494 (N_14494,N_13420,N_13440);
nand U14495 (N_14495,N_12912,N_12961);
nor U14496 (N_14496,N_13717,N_13676);
xnor U14497 (N_14497,N_12618,N_12531);
nor U14498 (N_14498,N_13081,N_13548);
and U14499 (N_14499,N_12672,N_13155);
nand U14500 (N_14500,N_13220,N_13630);
and U14501 (N_14501,N_13596,N_13408);
nor U14502 (N_14502,N_12860,N_13145);
xor U14503 (N_14503,N_13341,N_13674);
nor U14504 (N_14504,N_13455,N_13591);
nand U14505 (N_14505,N_13051,N_13045);
nand U14506 (N_14506,N_13430,N_13001);
xor U14507 (N_14507,N_12774,N_13264);
nand U14508 (N_14508,N_13437,N_12855);
xor U14509 (N_14509,N_12973,N_13544);
nand U14510 (N_14510,N_13619,N_12644);
nand U14511 (N_14511,N_13511,N_13122);
nand U14512 (N_14512,N_13534,N_13630);
and U14513 (N_14513,N_13148,N_12726);
and U14514 (N_14514,N_12720,N_13213);
xnor U14515 (N_14515,N_12890,N_12650);
xor U14516 (N_14516,N_13358,N_13577);
nand U14517 (N_14517,N_13193,N_12637);
and U14518 (N_14518,N_13042,N_13553);
xnor U14519 (N_14519,N_13355,N_13537);
or U14520 (N_14520,N_13512,N_13263);
xor U14521 (N_14521,N_13009,N_12888);
or U14522 (N_14522,N_13689,N_13231);
or U14523 (N_14523,N_12925,N_13381);
nand U14524 (N_14524,N_13300,N_12637);
nor U14525 (N_14525,N_12897,N_13366);
nand U14526 (N_14526,N_13581,N_13225);
or U14527 (N_14527,N_12781,N_13535);
and U14528 (N_14528,N_12772,N_13680);
nand U14529 (N_14529,N_12577,N_12840);
xnor U14530 (N_14530,N_13180,N_13143);
nand U14531 (N_14531,N_12501,N_13186);
nor U14532 (N_14532,N_13591,N_13576);
xnor U14533 (N_14533,N_13104,N_12574);
xor U14534 (N_14534,N_13404,N_12670);
or U14535 (N_14535,N_12843,N_12635);
and U14536 (N_14536,N_13683,N_12660);
nor U14537 (N_14537,N_13470,N_13171);
and U14538 (N_14538,N_12609,N_13449);
and U14539 (N_14539,N_13364,N_12750);
and U14540 (N_14540,N_12535,N_13285);
nand U14541 (N_14541,N_13221,N_13198);
nor U14542 (N_14542,N_13214,N_13102);
or U14543 (N_14543,N_13675,N_13149);
nand U14544 (N_14544,N_12725,N_13063);
or U14545 (N_14545,N_12570,N_12887);
xor U14546 (N_14546,N_13214,N_13317);
or U14547 (N_14547,N_13209,N_13509);
nand U14548 (N_14548,N_13022,N_12974);
xnor U14549 (N_14549,N_12585,N_13346);
xor U14550 (N_14550,N_12703,N_13577);
and U14551 (N_14551,N_13256,N_13282);
and U14552 (N_14552,N_12657,N_13148);
or U14553 (N_14553,N_13467,N_13676);
xor U14554 (N_14554,N_12889,N_12807);
or U14555 (N_14555,N_12628,N_12732);
nand U14556 (N_14556,N_13416,N_12813);
nand U14557 (N_14557,N_13158,N_12969);
nor U14558 (N_14558,N_12573,N_12961);
nand U14559 (N_14559,N_12523,N_13484);
nor U14560 (N_14560,N_13652,N_13112);
and U14561 (N_14561,N_12769,N_13594);
or U14562 (N_14562,N_12570,N_12843);
and U14563 (N_14563,N_13048,N_13691);
xor U14564 (N_14564,N_12693,N_13702);
xnor U14565 (N_14565,N_13687,N_13347);
and U14566 (N_14566,N_13599,N_13244);
or U14567 (N_14567,N_12853,N_13061);
and U14568 (N_14568,N_12635,N_13034);
xnor U14569 (N_14569,N_13102,N_13517);
or U14570 (N_14570,N_13043,N_12662);
nand U14571 (N_14571,N_12739,N_12719);
nand U14572 (N_14572,N_13279,N_13479);
nor U14573 (N_14573,N_13234,N_13345);
nand U14574 (N_14574,N_13406,N_13305);
and U14575 (N_14575,N_13387,N_13746);
nor U14576 (N_14576,N_13691,N_12541);
and U14577 (N_14577,N_13078,N_13270);
xnor U14578 (N_14578,N_13254,N_12647);
nor U14579 (N_14579,N_13645,N_13699);
nand U14580 (N_14580,N_13513,N_12796);
or U14581 (N_14581,N_12844,N_13373);
nor U14582 (N_14582,N_13724,N_13417);
and U14583 (N_14583,N_13730,N_13619);
nand U14584 (N_14584,N_12978,N_13289);
xnor U14585 (N_14585,N_12777,N_13193);
or U14586 (N_14586,N_13358,N_12521);
nor U14587 (N_14587,N_12553,N_12688);
nor U14588 (N_14588,N_12814,N_13046);
nor U14589 (N_14589,N_12966,N_12840);
nand U14590 (N_14590,N_13594,N_13715);
and U14591 (N_14591,N_13121,N_12612);
or U14592 (N_14592,N_13467,N_13357);
nand U14593 (N_14593,N_13572,N_12752);
xor U14594 (N_14594,N_13632,N_12560);
or U14595 (N_14595,N_12940,N_12500);
xnor U14596 (N_14596,N_12870,N_12582);
or U14597 (N_14597,N_13527,N_12897);
or U14598 (N_14598,N_13218,N_12877);
and U14599 (N_14599,N_12751,N_12652);
xnor U14600 (N_14600,N_13299,N_13522);
nor U14601 (N_14601,N_12954,N_13480);
and U14602 (N_14602,N_12613,N_13623);
and U14603 (N_14603,N_13092,N_13692);
nand U14604 (N_14604,N_13568,N_13263);
and U14605 (N_14605,N_13513,N_12525);
nand U14606 (N_14606,N_13536,N_12656);
and U14607 (N_14607,N_12575,N_13000);
or U14608 (N_14608,N_13597,N_13344);
nor U14609 (N_14609,N_13559,N_13360);
nand U14610 (N_14610,N_13518,N_12611);
nand U14611 (N_14611,N_12733,N_12759);
nand U14612 (N_14612,N_12761,N_13248);
nor U14613 (N_14613,N_12518,N_12712);
and U14614 (N_14614,N_12798,N_12919);
or U14615 (N_14615,N_13109,N_12873);
nor U14616 (N_14616,N_12831,N_12690);
or U14617 (N_14617,N_13551,N_13180);
xnor U14618 (N_14618,N_12974,N_12704);
and U14619 (N_14619,N_13567,N_13298);
nor U14620 (N_14620,N_12815,N_13717);
or U14621 (N_14621,N_12557,N_13327);
nand U14622 (N_14622,N_13461,N_13430);
nand U14623 (N_14623,N_13697,N_13456);
nand U14624 (N_14624,N_13319,N_13273);
xnor U14625 (N_14625,N_13653,N_12882);
nand U14626 (N_14626,N_13613,N_12636);
nor U14627 (N_14627,N_12965,N_13165);
nor U14628 (N_14628,N_13540,N_12963);
xnor U14629 (N_14629,N_13725,N_13690);
nand U14630 (N_14630,N_12657,N_13548);
nor U14631 (N_14631,N_12554,N_12569);
or U14632 (N_14632,N_13747,N_12835);
nor U14633 (N_14633,N_12649,N_13542);
or U14634 (N_14634,N_12501,N_13679);
or U14635 (N_14635,N_13447,N_12567);
xnor U14636 (N_14636,N_13169,N_13354);
and U14637 (N_14637,N_12726,N_13047);
and U14638 (N_14638,N_12720,N_13118);
xnor U14639 (N_14639,N_13701,N_12532);
nand U14640 (N_14640,N_12995,N_12928);
nor U14641 (N_14641,N_13278,N_12994);
nor U14642 (N_14642,N_13279,N_12670);
and U14643 (N_14643,N_12842,N_12828);
nor U14644 (N_14644,N_13430,N_12773);
xnor U14645 (N_14645,N_13339,N_12963);
and U14646 (N_14646,N_12811,N_13430);
xnor U14647 (N_14647,N_13541,N_12710);
and U14648 (N_14648,N_12908,N_13028);
nor U14649 (N_14649,N_12580,N_12868);
nor U14650 (N_14650,N_12576,N_13714);
nand U14651 (N_14651,N_12836,N_13045);
and U14652 (N_14652,N_12902,N_13382);
and U14653 (N_14653,N_12521,N_13524);
nand U14654 (N_14654,N_13428,N_13619);
xnor U14655 (N_14655,N_13054,N_12843);
and U14656 (N_14656,N_13001,N_13649);
nand U14657 (N_14657,N_13674,N_12660);
nand U14658 (N_14658,N_13126,N_12996);
nor U14659 (N_14659,N_12756,N_13590);
or U14660 (N_14660,N_13494,N_12552);
nand U14661 (N_14661,N_12945,N_13454);
xor U14662 (N_14662,N_12884,N_13457);
and U14663 (N_14663,N_13696,N_13263);
nand U14664 (N_14664,N_12600,N_13652);
nand U14665 (N_14665,N_12750,N_13550);
and U14666 (N_14666,N_13115,N_13515);
or U14667 (N_14667,N_12802,N_13650);
nor U14668 (N_14668,N_13513,N_13525);
or U14669 (N_14669,N_13503,N_13544);
or U14670 (N_14670,N_12933,N_13190);
nand U14671 (N_14671,N_12805,N_13241);
and U14672 (N_14672,N_13235,N_12642);
xnor U14673 (N_14673,N_13002,N_13530);
and U14674 (N_14674,N_12936,N_12519);
nand U14675 (N_14675,N_12518,N_13745);
nand U14676 (N_14676,N_12682,N_12920);
and U14677 (N_14677,N_12900,N_13035);
nand U14678 (N_14678,N_13149,N_13264);
or U14679 (N_14679,N_13516,N_13069);
nor U14680 (N_14680,N_12835,N_12722);
nor U14681 (N_14681,N_13223,N_13188);
xnor U14682 (N_14682,N_12583,N_13069);
and U14683 (N_14683,N_12976,N_13204);
xor U14684 (N_14684,N_12829,N_12905);
xor U14685 (N_14685,N_12562,N_13733);
nor U14686 (N_14686,N_13082,N_12978);
and U14687 (N_14687,N_13339,N_12599);
and U14688 (N_14688,N_13062,N_12683);
nand U14689 (N_14689,N_13406,N_13747);
nand U14690 (N_14690,N_12613,N_13599);
or U14691 (N_14691,N_13076,N_13646);
and U14692 (N_14692,N_13112,N_12737);
nor U14693 (N_14693,N_12824,N_12948);
xnor U14694 (N_14694,N_13077,N_13628);
xor U14695 (N_14695,N_12859,N_13729);
and U14696 (N_14696,N_12905,N_12599);
and U14697 (N_14697,N_12862,N_13356);
or U14698 (N_14698,N_12966,N_13087);
nand U14699 (N_14699,N_12852,N_12751);
xnor U14700 (N_14700,N_13479,N_13235);
nand U14701 (N_14701,N_12962,N_13247);
or U14702 (N_14702,N_13240,N_12836);
and U14703 (N_14703,N_12665,N_12898);
xnor U14704 (N_14704,N_13496,N_12591);
nor U14705 (N_14705,N_13527,N_13623);
nand U14706 (N_14706,N_13665,N_13466);
and U14707 (N_14707,N_13714,N_13492);
nor U14708 (N_14708,N_13409,N_12529);
or U14709 (N_14709,N_12783,N_13085);
xor U14710 (N_14710,N_13222,N_13307);
nor U14711 (N_14711,N_12515,N_13238);
nand U14712 (N_14712,N_13436,N_13555);
and U14713 (N_14713,N_12534,N_13038);
nor U14714 (N_14714,N_13309,N_12738);
xnor U14715 (N_14715,N_13205,N_13137);
xor U14716 (N_14716,N_13205,N_13399);
nand U14717 (N_14717,N_12745,N_12959);
xor U14718 (N_14718,N_12917,N_12512);
nor U14719 (N_14719,N_12988,N_13317);
or U14720 (N_14720,N_12757,N_12955);
nand U14721 (N_14721,N_13715,N_12685);
xnor U14722 (N_14722,N_13153,N_13658);
nor U14723 (N_14723,N_12954,N_13037);
or U14724 (N_14724,N_13537,N_13116);
and U14725 (N_14725,N_13661,N_12544);
nor U14726 (N_14726,N_13010,N_13208);
nand U14727 (N_14727,N_12715,N_13291);
and U14728 (N_14728,N_13674,N_13665);
and U14729 (N_14729,N_13340,N_13121);
or U14730 (N_14730,N_12524,N_13288);
nand U14731 (N_14731,N_13493,N_13237);
and U14732 (N_14732,N_12712,N_12546);
and U14733 (N_14733,N_12737,N_13530);
or U14734 (N_14734,N_13632,N_12821);
nand U14735 (N_14735,N_12747,N_13348);
xnor U14736 (N_14736,N_12797,N_13003);
nand U14737 (N_14737,N_12834,N_13098);
or U14738 (N_14738,N_12710,N_12538);
nor U14739 (N_14739,N_13439,N_12966);
nor U14740 (N_14740,N_12918,N_12665);
nor U14741 (N_14741,N_12919,N_13467);
or U14742 (N_14742,N_13444,N_12966);
or U14743 (N_14743,N_12578,N_13052);
nor U14744 (N_14744,N_13587,N_12578);
and U14745 (N_14745,N_13200,N_12543);
xnor U14746 (N_14746,N_12980,N_13577);
and U14747 (N_14747,N_13469,N_12866);
or U14748 (N_14748,N_13503,N_13158);
or U14749 (N_14749,N_13711,N_12547);
nor U14750 (N_14750,N_13145,N_13443);
nand U14751 (N_14751,N_13292,N_12792);
nor U14752 (N_14752,N_12863,N_13668);
or U14753 (N_14753,N_12825,N_13412);
nor U14754 (N_14754,N_12982,N_13027);
or U14755 (N_14755,N_12629,N_13686);
or U14756 (N_14756,N_13365,N_12940);
nor U14757 (N_14757,N_12854,N_12820);
and U14758 (N_14758,N_13698,N_13138);
or U14759 (N_14759,N_12534,N_13183);
and U14760 (N_14760,N_13008,N_12951);
nor U14761 (N_14761,N_13728,N_12769);
nand U14762 (N_14762,N_12635,N_13474);
or U14763 (N_14763,N_12694,N_12682);
nor U14764 (N_14764,N_13207,N_13576);
and U14765 (N_14765,N_13355,N_12733);
xor U14766 (N_14766,N_12896,N_13749);
xor U14767 (N_14767,N_13365,N_13544);
nand U14768 (N_14768,N_12801,N_12717);
and U14769 (N_14769,N_12857,N_13176);
and U14770 (N_14770,N_13649,N_13142);
and U14771 (N_14771,N_13659,N_13234);
and U14772 (N_14772,N_13149,N_12512);
and U14773 (N_14773,N_12876,N_13128);
nand U14774 (N_14774,N_13196,N_12722);
nand U14775 (N_14775,N_12944,N_13482);
xnor U14776 (N_14776,N_13311,N_12510);
or U14777 (N_14777,N_13268,N_12858);
xor U14778 (N_14778,N_13622,N_13707);
nor U14779 (N_14779,N_13303,N_12777);
nand U14780 (N_14780,N_13031,N_12505);
nor U14781 (N_14781,N_12505,N_13075);
and U14782 (N_14782,N_13384,N_12815);
nand U14783 (N_14783,N_13475,N_13094);
nor U14784 (N_14784,N_12829,N_13370);
and U14785 (N_14785,N_13312,N_12816);
xnor U14786 (N_14786,N_12599,N_13297);
nor U14787 (N_14787,N_12652,N_13088);
or U14788 (N_14788,N_12968,N_12774);
nand U14789 (N_14789,N_12562,N_13069);
and U14790 (N_14790,N_13192,N_13636);
or U14791 (N_14791,N_13122,N_12763);
nor U14792 (N_14792,N_13410,N_13581);
xor U14793 (N_14793,N_12913,N_13375);
nor U14794 (N_14794,N_13141,N_13663);
nor U14795 (N_14795,N_13088,N_12961);
and U14796 (N_14796,N_13396,N_13539);
or U14797 (N_14797,N_12916,N_13103);
nor U14798 (N_14798,N_12583,N_13490);
xnor U14799 (N_14799,N_12827,N_13353);
nor U14800 (N_14800,N_12872,N_13709);
nor U14801 (N_14801,N_13594,N_12666);
nor U14802 (N_14802,N_13598,N_13608);
or U14803 (N_14803,N_13251,N_13346);
nand U14804 (N_14804,N_13062,N_12761);
or U14805 (N_14805,N_13155,N_12782);
or U14806 (N_14806,N_12546,N_12854);
or U14807 (N_14807,N_13309,N_13194);
nor U14808 (N_14808,N_13692,N_12731);
nand U14809 (N_14809,N_13603,N_12606);
xnor U14810 (N_14810,N_13218,N_13121);
nand U14811 (N_14811,N_12614,N_13321);
nor U14812 (N_14812,N_12719,N_13138);
nand U14813 (N_14813,N_12869,N_13383);
and U14814 (N_14814,N_13729,N_12702);
and U14815 (N_14815,N_12954,N_12770);
nor U14816 (N_14816,N_13066,N_13184);
xor U14817 (N_14817,N_13397,N_13150);
xor U14818 (N_14818,N_13549,N_12975);
and U14819 (N_14819,N_13210,N_13358);
nand U14820 (N_14820,N_13229,N_13738);
and U14821 (N_14821,N_12824,N_12580);
and U14822 (N_14822,N_13274,N_12770);
and U14823 (N_14823,N_12513,N_13341);
nand U14824 (N_14824,N_13634,N_13436);
or U14825 (N_14825,N_12980,N_12746);
or U14826 (N_14826,N_13205,N_12980);
xor U14827 (N_14827,N_12905,N_12885);
nand U14828 (N_14828,N_13073,N_12639);
xor U14829 (N_14829,N_13542,N_12982);
xor U14830 (N_14830,N_12706,N_13533);
and U14831 (N_14831,N_13276,N_12541);
xor U14832 (N_14832,N_13560,N_12820);
nand U14833 (N_14833,N_13303,N_13379);
xnor U14834 (N_14834,N_12810,N_13389);
nor U14835 (N_14835,N_13272,N_12674);
nor U14836 (N_14836,N_12848,N_13411);
nor U14837 (N_14837,N_13401,N_12819);
xnor U14838 (N_14838,N_13052,N_13018);
nor U14839 (N_14839,N_12637,N_12972);
nand U14840 (N_14840,N_12941,N_13220);
xor U14841 (N_14841,N_13589,N_13126);
or U14842 (N_14842,N_12796,N_13403);
or U14843 (N_14843,N_13320,N_13125);
and U14844 (N_14844,N_13171,N_12883);
or U14845 (N_14845,N_13550,N_12574);
or U14846 (N_14846,N_13537,N_12728);
xor U14847 (N_14847,N_12704,N_13497);
and U14848 (N_14848,N_12989,N_13201);
nor U14849 (N_14849,N_13524,N_12837);
nand U14850 (N_14850,N_13459,N_13193);
nor U14851 (N_14851,N_13184,N_13467);
nand U14852 (N_14852,N_13606,N_12502);
nand U14853 (N_14853,N_13541,N_13236);
nand U14854 (N_14854,N_12808,N_12592);
xor U14855 (N_14855,N_13578,N_12631);
and U14856 (N_14856,N_12753,N_13661);
xor U14857 (N_14857,N_12642,N_12701);
nor U14858 (N_14858,N_13693,N_13155);
and U14859 (N_14859,N_13066,N_12679);
nor U14860 (N_14860,N_12870,N_13216);
xnor U14861 (N_14861,N_13600,N_13735);
and U14862 (N_14862,N_13236,N_12576);
nand U14863 (N_14863,N_12892,N_12974);
xor U14864 (N_14864,N_13413,N_12839);
xor U14865 (N_14865,N_13335,N_12951);
xnor U14866 (N_14866,N_13557,N_13034);
and U14867 (N_14867,N_13298,N_12818);
nor U14868 (N_14868,N_13403,N_13343);
nor U14869 (N_14869,N_13693,N_12949);
nor U14870 (N_14870,N_12713,N_12559);
nand U14871 (N_14871,N_12811,N_13528);
xnor U14872 (N_14872,N_13403,N_13732);
nand U14873 (N_14873,N_13086,N_12641);
xor U14874 (N_14874,N_13638,N_13663);
nor U14875 (N_14875,N_12891,N_13195);
xnor U14876 (N_14876,N_13336,N_12533);
nand U14877 (N_14877,N_13471,N_13678);
nor U14878 (N_14878,N_12683,N_13053);
or U14879 (N_14879,N_13001,N_13595);
and U14880 (N_14880,N_13415,N_13593);
and U14881 (N_14881,N_13443,N_12525);
nor U14882 (N_14882,N_13024,N_12844);
nor U14883 (N_14883,N_13606,N_12880);
nand U14884 (N_14884,N_12875,N_12876);
or U14885 (N_14885,N_13490,N_13145);
and U14886 (N_14886,N_13121,N_13196);
and U14887 (N_14887,N_13421,N_13114);
nor U14888 (N_14888,N_12926,N_13232);
or U14889 (N_14889,N_13321,N_12617);
nand U14890 (N_14890,N_12989,N_12735);
nand U14891 (N_14891,N_13064,N_13692);
xor U14892 (N_14892,N_13665,N_13670);
or U14893 (N_14893,N_12553,N_12574);
and U14894 (N_14894,N_13403,N_12772);
and U14895 (N_14895,N_12710,N_13491);
nand U14896 (N_14896,N_13667,N_13409);
xnor U14897 (N_14897,N_13720,N_12828);
and U14898 (N_14898,N_13048,N_13404);
nand U14899 (N_14899,N_13301,N_12999);
nand U14900 (N_14900,N_13303,N_12901);
and U14901 (N_14901,N_13316,N_12688);
xnor U14902 (N_14902,N_13620,N_13372);
nor U14903 (N_14903,N_12745,N_13606);
nand U14904 (N_14904,N_13335,N_12657);
nand U14905 (N_14905,N_13580,N_12828);
or U14906 (N_14906,N_13630,N_13358);
nand U14907 (N_14907,N_13279,N_13408);
or U14908 (N_14908,N_12522,N_12967);
and U14909 (N_14909,N_13507,N_13060);
and U14910 (N_14910,N_13647,N_12568);
nand U14911 (N_14911,N_13485,N_12642);
nand U14912 (N_14912,N_13654,N_12543);
nor U14913 (N_14913,N_12901,N_13385);
or U14914 (N_14914,N_13307,N_13346);
and U14915 (N_14915,N_12900,N_13180);
or U14916 (N_14916,N_13216,N_13394);
nand U14917 (N_14917,N_13322,N_12739);
and U14918 (N_14918,N_12895,N_13505);
xnor U14919 (N_14919,N_13338,N_13386);
and U14920 (N_14920,N_13122,N_12988);
xnor U14921 (N_14921,N_12736,N_12583);
and U14922 (N_14922,N_12591,N_12518);
nand U14923 (N_14923,N_13376,N_13725);
nand U14924 (N_14924,N_12937,N_13209);
and U14925 (N_14925,N_12992,N_13314);
nand U14926 (N_14926,N_12975,N_13503);
or U14927 (N_14927,N_13237,N_13007);
or U14928 (N_14928,N_12642,N_13608);
nor U14929 (N_14929,N_13091,N_13208);
nor U14930 (N_14930,N_13334,N_12978);
or U14931 (N_14931,N_13509,N_13198);
nand U14932 (N_14932,N_13090,N_13747);
nor U14933 (N_14933,N_13104,N_12911);
xor U14934 (N_14934,N_12733,N_13010);
xor U14935 (N_14935,N_13028,N_12973);
and U14936 (N_14936,N_13086,N_13107);
and U14937 (N_14937,N_12821,N_13371);
or U14938 (N_14938,N_13162,N_13465);
nor U14939 (N_14939,N_13316,N_13673);
and U14940 (N_14940,N_12974,N_12781);
nor U14941 (N_14941,N_13420,N_13319);
nand U14942 (N_14942,N_13193,N_12501);
nor U14943 (N_14943,N_13360,N_12523);
or U14944 (N_14944,N_12894,N_13490);
or U14945 (N_14945,N_13545,N_12573);
xnor U14946 (N_14946,N_12817,N_13681);
and U14947 (N_14947,N_12684,N_13304);
nor U14948 (N_14948,N_13568,N_12992);
and U14949 (N_14949,N_13176,N_13043);
nor U14950 (N_14950,N_12676,N_13108);
and U14951 (N_14951,N_13576,N_13629);
xnor U14952 (N_14952,N_13082,N_12672);
nor U14953 (N_14953,N_13306,N_13275);
and U14954 (N_14954,N_12702,N_13648);
and U14955 (N_14955,N_13492,N_13547);
nand U14956 (N_14956,N_13552,N_13449);
or U14957 (N_14957,N_12833,N_13423);
xor U14958 (N_14958,N_13492,N_12818);
and U14959 (N_14959,N_13402,N_13332);
or U14960 (N_14960,N_13078,N_13422);
nor U14961 (N_14961,N_12581,N_12640);
nor U14962 (N_14962,N_13250,N_12953);
or U14963 (N_14963,N_12970,N_13529);
or U14964 (N_14964,N_13710,N_13661);
nand U14965 (N_14965,N_13041,N_13297);
nor U14966 (N_14966,N_12894,N_13602);
or U14967 (N_14967,N_12610,N_13547);
and U14968 (N_14968,N_12850,N_13717);
nand U14969 (N_14969,N_12757,N_13514);
or U14970 (N_14970,N_13668,N_12574);
and U14971 (N_14971,N_12613,N_13050);
nor U14972 (N_14972,N_13092,N_13023);
nand U14973 (N_14973,N_12745,N_12780);
xor U14974 (N_14974,N_13744,N_12646);
nand U14975 (N_14975,N_13663,N_12821);
or U14976 (N_14976,N_13555,N_13544);
nor U14977 (N_14977,N_13392,N_12943);
xor U14978 (N_14978,N_13702,N_13327);
xnor U14979 (N_14979,N_13280,N_12776);
or U14980 (N_14980,N_12841,N_13436);
xnor U14981 (N_14981,N_13526,N_13631);
xnor U14982 (N_14982,N_12573,N_12684);
and U14983 (N_14983,N_13441,N_13207);
nand U14984 (N_14984,N_12880,N_12549);
or U14985 (N_14985,N_13410,N_13086);
nand U14986 (N_14986,N_12946,N_13616);
nand U14987 (N_14987,N_13547,N_13472);
nor U14988 (N_14988,N_12802,N_13619);
and U14989 (N_14989,N_13184,N_13373);
or U14990 (N_14990,N_12603,N_13720);
and U14991 (N_14991,N_12812,N_13139);
xnor U14992 (N_14992,N_13585,N_12725);
nand U14993 (N_14993,N_13461,N_13016);
or U14994 (N_14994,N_12682,N_12551);
xor U14995 (N_14995,N_12580,N_13733);
nor U14996 (N_14996,N_12601,N_12548);
and U14997 (N_14997,N_13110,N_13603);
xnor U14998 (N_14998,N_13100,N_12951);
nor U14999 (N_14999,N_12515,N_12839);
nor U15000 (N_15000,N_14762,N_14740);
and U15001 (N_15001,N_14590,N_14685);
and U15002 (N_15002,N_14222,N_14727);
or U15003 (N_15003,N_14441,N_14787);
and U15004 (N_15004,N_14113,N_14194);
nor U15005 (N_15005,N_13911,N_14996);
or U15006 (N_15006,N_14843,N_13868);
nor U15007 (N_15007,N_14298,N_14451);
xnor U15008 (N_15008,N_14535,N_14087);
xnor U15009 (N_15009,N_14306,N_14970);
nand U15010 (N_15010,N_14079,N_14892);
and U15011 (N_15011,N_14127,N_14687);
nor U15012 (N_15012,N_14405,N_14242);
and U15013 (N_15013,N_14159,N_14058);
or U15014 (N_15014,N_14689,N_13850);
nand U15015 (N_15015,N_14603,N_14784);
xor U15016 (N_15016,N_14406,N_14557);
or U15017 (N_15017,N_13859,N_13865);
and U15018 (N_15018,N_13781,N_14522);
or U15019 (N_15019,N_14790,N_14385);
or U15020 (N_15020,N_14882,N_13949);
or U15021 (N_15021,N_14846,N_13934);
or U15022 (N_15022,N_14981,N_14749);
nor U15023 (N_15023,N_13766,N_14481);
or U15024 (N_15024,N_14110,N_14682);
and U15025 (N_15025,N_14773,N_14263);
and U15026 (N_15026,N_14855,N_13957);
nor U15027 (N_15027,N_14177,N_14273);
nand U15028 (N_15028,N_14346,N_14761);
nand U15029 (N_15029,N_13816,N_14443);
or U15030 (N_15030,N_13935,N_14029);
nand U15031 (N_15031,N_14398,N_13822);
or U15032 (N_15032,N_14512,N_14941);
and U15033 (N_15033,N_14449,N_14847);
and U15034 (N_15034,N_14126,N_13847);
and U15035 (N_15035,N_14008,N_14577);
nand U15036 (N_15036,N_14561,N_13933);
and U15037 (N_15037,N_14477,N_14460);
xnor U15038 (N_15038,N_14560,N_14114);
or U15039 (N_15039,N_14310,N_14433);
and U15040 (N_15040,N_14951,N_14384);
nand U15041 (N_15041,N_14878,N_14276);
nand U15042 (N_15042,N_14658,N_14142);
nor U15043 (N_15043,N_14170,N_14818);
nor U15044 (N_15044,N_14622,N_14387);
xor U15045 (N_15045,N_14389,N_14529);
nand U15046 (N_15046,N_14038,N_14738);
and U15047 (N_15047,N_14821,N_13893);
and U15048 (N_15048,N_14674,N_13999);
or U15049 (N_15049,N_14399,N_14181);
and U15050 (N_15050,N_14753,N_14305);
nor U15051 (N_15051,N_14615,N_14457);
or U15052 (N_15052,N_13972,N_14012);
and U15053 (N_15053,N_14286,N_14144);
xor U15054 (N_15054,N_14748,N_13839);
xor U15055 (N_15055,N_14219,N_13925);
or U15056 (N_15056,N_14272,N_14108);
and U15057 (N_15057,N_14115,N_13846);
xnor U15058 (N_15058,N_14329,N_14018);
nor U15059 (N_15059,N_14936,N_14418);
or U15060 (N_15060,N_14665,N_13989);
nand U15061 (N_15061,N_14171,N_14388);
or U15062 (N_15062,N_14549,N_14509);
nand U15063 (N_15063,N_14432,N_13821);
or U15064 (N_15064,N_14120,N_13945);
xnor U15065 (N_15065,N_14214,N_14424);
or U15066 (N_15066,N_14813,N_14799);
or U15067 (N_15067,N_14505,N_14200);
nand U15068 (N_15068,N_13755,N_14641);
nor U15069 (N_15069,N_14092,N_14327);
nand U15070 (N_15070,N_14478,N_14401);
or U15071 (N_15071,N_14905,N_14606);
and U15072 (N_15072,N_14428,N_14750);
or U15073 (N_15073,N_14720,N_14123);
xor U15074 (N_15074,N_14921,N_14624);
or U15075 (N_15075,N_14902,N_14434);
nor U15076 (N_15076,N_14050,N_14035);
or U15077 (N_15077,N_14781,N_14332);
xor U15078 (N_15078,N_14836,N_14667);
nand U15079 (N_15079,N_13940,N_14514);
nand U15080 (N_15080,N_13825,N_14059);
and U15081 (N_15081,N_14380,N_14218);
xnor U15082 (N_15082,N_13771,N_14985);
nand U15083 (N_15083,N_14160,N_14786);
nor U15084 (N_15084,N_14645,N_14884);
nor U15085 (N_15085,N_14098,N_14107);
and U15086 (N_15086,N_14281,N_14541);
xor U15087 (N_15087,N_13956,N_14832);
nand U15088 (N_15088,N_13904,N_14677);
and U15089 (N_15089,N_13950,N_14162);
and U15090 (N_15090,N_13962,N_14005);
or U15091 (N_15091,N_14660,N_14206);
or U15092 (N_15092,N_14595,N_14109);
and U15093 (N_15093,N_13759,N_14986);
nor U15094 (N_15094,N_14835,N_14935);
nand U15095 (N_15095,N_14618,N_13762);
xnor U15096 (N_15096,N_14845,N_14354);
nand U15097 (N_15097,N_14780,N_14456);
and U15098 (N_15098,N_13835,N_14890);
xnor U15099 (N_15099,N_14006,N_13845);
and U15100 (N_15100,N_14349,N_14516);
and U15101 (N_15101,N_14152,N_14202);
nor U15102 (N_15102,N_14148,N_14971);
nor U15103 (N_15103,N_14554,N_14021);
and U15104 (N_15104,N_14984,N_14437);
nor U15105 (N_15105,N_14719,N_14414);
and U15106 (N_15106,N_14643,N_13866);
and U15107 (N_15107,N_14896,N_14596);
xor U15108 (N_15108,N_14779,N_14679);
nand U15109 (N_15109,N_14246,N_14716);
xnor U15110 (N_15110,N_14138,N_14724);
nor U15111 (N_15111,N_13778,N_14866);
nor U15112 (N_15112,N_14334,N_14331);
and U15113 (N_15113,N_13974,N_14807);
and U15114 (N_15114,N_14531,N_13967);
or U15115 (N_15115,N_14544,N_13902);
and U15116 (N_15116,N_13784,N_13907);
nor U15117 (N_15117,N_14849,N_13774);
or U15118 (N_15118,N_14711,N_13796);
nand U15119 (N_15119,N_14503,N_14867);
xor U15120 (N_15120,N_14469,N_14062);
or U15121 (N_15121,N_14788,N_14841);
nand U15122 (N_15122,N_13889,N_14237);
and U15123 (N_15123,N_13862,N_14684);
nor U15124 (N_15124,N_14511,N_14956);
xor U15125 (N_15125,N_14454,N_14259);
nand U15126 (N_15126,N_14484,N_13751);
and U15127 (N_15127,N_13946,N_14657);
xor U15128 (N_15128,N_14351,N_14187);
nand U15129 (N_15129,N_14423,N_14859);
nor U15130 (N_15130,N_13992,N_14267);
nand U15131 (N_15131,N_14186,N_13764);
nor U15132 (N_15132,N_14407,N_14492);
or U15133 (N_15133,N_14759,N_14736);
nor U15134 (N_15134,N_14096,N_14838);
xnor U15135 (N_15135,N_13963,N_14542);
nand U15136 (N_15136,N_13873,N_14774);
nor U15137 (N_15137,N_13838,N_14819);
xor U15138 (N_15138,N_14810,N_14284);
xor U15139 (N_15139,N_14722,N_13938);
xor U15140 (N_15140,N_14872,N_14105);
or U15141 (N_15141,N_14963,N_14967);
and U15142 (N_15142,N_14101,N_13970);
or U15143 (N_15143,N_13998,N_14532);
and U15144 (N_15144,N_14493,N_14545);
or U15145 (N_15145,N_14572,N_14704);
or U15146 (N_15146,N_14309,N_14323);
xnor U15147 (N_15147,N_14376,N_14906);
and U15148 (N_15148,N_14536,N_13895);
or U15149 (N_15149,N_14770,N_14369);
or U15150 (N_15150,N_14909,N_14559);
xnor U15151 (N_15151,N_14257,N_13906);
or U15152 (N_15152,N_14697,N_14692);
xor U15153 (N_15153,N_14778,N_14256);
or U15154 (N_15154,N_14969,N_14293);
xor U15155 (N_15155,N_14232,N_14065);
nand U15156 (N_15156,N_14605,N_14172);
and U15157 (N_15157,N_14041,N_14016);
or U15158 (N_15158,N_14515,N_14993);
nor U15159 (N_15159,N_13777,N_14390);
and U15160 (N_15160,N_13758,N_14347);
nor U15161 (N_15161,N_14919,N_14060);
or U15162 (N_15162,N_14483,N_14049);
and U15163 (N_15163,N_14285,N_14015);
xor U15164 (N_15164,N_14798,N_14772);
xor U15165 (N_15165,N_14485,N_14491);
xnor U15166 (N_15166,N_14494,N_14416);
xnor U15167 (N_15167,N_14883,N_14031);
nand U15168 (N_15168,N_13948,N_13763);
xnor U15169 (N_15169,N_14173,N_14464);
xnor U15170 (N_15170,N_14961,N_14634);
and U15171 (N_15171,N_14208,N_14973);
nand U15172 (N_15172,N_14592,N_14964);
and U15173 (N_15173,N_14023,N_13982);
nor U15174 (N_15174,N_13811,N_14497);
or U15175 (N_15175,N_14928,N_14600);
and U15176 (N_15176,N_14335,N_14254);
nor U15177 (N_15177,N_14757,N_14487);
xor U15178 (N_15178,N_14095,N_14420);
xnor U15179 (N_15179,N_14240,N_14694);
nor U15180 (N_15180,N_14977,N_14249);
and U15181 (N_15181,N_14308,N_14301);
nand U15182 (N_15182,N_14213,N_14816);
and U15183 (N_15183,N_14506,N_14582);
xnor U15184 (N_15184,N_14315,N_14988);
nand U15185 (N_15185,N_13915,N_14203);
nand U15186 (N_15186,N_14876,N_14279);
nor U15187 (N_15187,N_14467,N_14893);
nor U15188 (N_15188,N_14940,N_13750);
nand U15189 (N_15189,N_14910,N_14994);
nor U15190 (N_15190,N_14189,N_13802);
or U15191 (N_15191,N_14359,N_13908);
nor U15192 (N_15192,N_14507,N_14410);
and U15193 (N_15193,N_14562,N_14299);
or U15194 (N_15194,N_14375,N_14363);
xnor U15195 (N_15195,N_14201,N_14234);
nor U15196 (N_15196,N_14630,N_14934);
and U15197 (N_15197,N_14192,N_13857);
or U15198 (N_15198,N_14937,N_14621);
nand U15199 (N_15199,N_14198,N_14862);
and U15200 (N_15200,N_14633,N_14373);
or U15201 (N_15201,N_14135,N_13830);
nand U15202 (N_15202,N_13941,N_14378);
xnor U15203 (N_15203,N_14093,N_14668);
nor U15204 (N_15204,N_14944,N_14785);
and U15205 (N_15205,N_14009,N_14881);
and U15206 (N_15206,N_13772,N_14502);
and U15207 (N_15207,N_14631,N_14425);
nand U15208 (N_15208,N_14094,N_13884);
nor U15209 (N_15209,N_13837,N_14737);
xnor U15210 (N_15210,N_14607,N_14860);
nor U15211 (N_15211,N_14221,N_14104);
nand U15212 (N_15212,N_14955,N_14612);
or U15213 (N_15213,N_14320,N_14806);
and U15214 (N_15214,N_14337,N_13973);
xor U15215 (N_15215,N_14116,N_14394);
and U15216 (N_15216,N_14980,N_14132);
nor U15217 (N_15217,N_14765,N_13975);
nor U15218 (N_15218,N_14353,N_14472);
or U15219 (N_15219,N_14990,N_13798);
and U15220 (N_15220,N_14611,N_14576);
nor U15221 (N_15221,N_14854,N_13888);
or U15222 (N_15222,N_14945,N_13870);
nor U15223 (N_15223,N_14574,N_14251);
or U15224 (N_15224,N_14077,N_14666);
or U15225 (N_15225,N_14297,N_14448);
nor U15226 (N_15226,N_14158,N_14962);
and U15227 (N_15227,N_14828,N_13815);
or U15228 (N_15228,N_14649,N_13879);
nand U15229 (N_15229,N_14681,N_13819);
xor U15230 (N_15230,N_14508,N_14648);
nor U15231 (N_15231,N_13787,N_14047);
and U15232 (N_15232,N_14731,N_14356);
xor U15233 (N_15233,N_14371,N_14814);
nand U15234 (N_15234,N_14530,N_14243);
nor U15235 (N_15235,N_14693,N_14043);
and U15236 (N_15236,N_14030,N_14669);
nand U15237 (N_15237,N_13797,N_14037);
nand U15238 (N_15238,N_14654,N_14118);
xnor U15239 (N_15239,N_14475,N_13881);
xnor U15240 (N_15240,N_14024,N_14071);
and U15241 (N_15241,N_13969,N_14717);
and U15242 (N_15242,N_14145,N_14244);
nor U15243 (N_15243,N_13997,N_14217);
nand U15244 (N_15244,N_14436,N_14250);
nor U15245 (N_15245,N_13858,N_14129);
nor U15246 (N_15246,N_14408,N_14708);
or U15247 (N_15247,N_14580,N_14156);
or U15248 (N_15248,N_14879,N_14480);
nand U15249 (N_15249,N_14887,N_13978);
or U15250 (N_15250,N_14972,N_14803);
or U15251 (N_15251,N_14775,N_13990);
nor U15252 (N_15252,N_13814,N_14721);
nand U15253 (N_15253,N_13760,N_14943);
xnor U15254 (N_15254,N_13891,N_14207);
and U15255 (N_15255,N_13840,N_14199);
and U15256 (N_15256,N_14235,N_13932);
and U15257 (N_15257,N_13885,N_14820);
xor U15258 (N_15258,N_14161,N_13878);
and U15259 (N_15259,N_14230,N_13936);
or U15260 (N_15260,N_14482,N_14412);
xnor U15261 (N_15261,N_14918,N_14880);
or U15262 (N_15262,N_14524,N_14976);
xnor U15263 (N_15263,N_14520,N_13768);
and U15264 (N_15264,N_14625,N_14997);
and U15265 (N_15265,N_14652,N_14473);
xnor U15266 (N_15266,N_14080,N_14551);
xnor U15267 (N_15267,N_13991,N_13836);
nand U15268 (N_15268,N_14715,N_14122);
or U15269 (N_15269,N_14463,N_14730);
or U15270 (N_15270,N_14510,N_14318);
and U15271 (N_15271,N_14007,N_14446);
nand U15272 (N_15272,N_14155,N_13921);
nand U15273 (N_15273,N_13867,N_14383);
or U15274 (N_15274,N_14193,N_14195);
or U15275 (N_15275,N_14588,N_14056);
or U15276 (N_15276,N_14744,N_13916);
nor U15277 (N_15277,N_14034,N_14552);
nor U15278 (N_15278,N_14261,N_14771);
nand U15279 (N_15279,N_14061,N_14236);
xor U15280 (N_15280,N_14450,N_14646);
or U15281 (N_15281,N_14072,N_14823);
nor U15282 (N_15282,N_14324,N_14274);
nand U15283 (N_15283,N_14258,N_13898);
and U15284 (N_15284,N_14166,N_13789);
nand U15285 (N_15285,N_14864,N_14995);
and U15286 (N_15286,N_14670,N_14100);
and U15287 (N_15287,N_14989,N_14314);
or U15288 (N_15288,N_14302,N_14567);
nor U15289 (N_15289,N_14703,N_14002);
nand U15290 (N_15290,N_14713,N_14081);
and U15291 (N_15291,N_13849,N_14931);
nand U15292 (N_15292,N_14534,N_14139);
or U15293 (N_15293,N_14579,N_13880);
and U15294 (N_15294,N_14957,N_14225);
or U15295 (N_15295,N_13799,N_14556);
and U15296 (N_15296,N_14476,N_14468);
nor U15297 (N_15297,N_14069,N_14523);
nor U15298 (N_15298,N_14102,N_13791);
or U15299 (N_15299,N_14877,N_14404);
xnor U15300 (N_15300,N_14465,N_14678);
nand U15301 (N_15301,N_14231,N_13918);
nand U15302 (N_15302,N_14891,N_13788);
nand U15303 (N_15303,N_14794,N_13909);
or U15304 (N_15304,N_13954,N_14339);
xor U15305 (N_15305,N_14924,N_14733);
or U15306 (N_15306,N_13965,N_14117);
nand U15307 (N_15307,N_14010,N_14644);
nor U15308 (N_15308,N_13852,N_14136);
xor U15309 (N_15309,N_14526,N_14452);
nor U15310 (N_15310,N_14601,N_14718);
and U15311 (N_15311,N_14900,N_14812);
nand U15312 (N_15312,N_13813,N_13905);
nor U15313 (N_15313,N_14435,N_14429);
xnor U15314 (N_15314,N_14589,N_14564);
nand U15315 (N_15315,N_14063,N_13753);
or U15316 (N_15316,N_14265,N_14760);
nand U15317 (N_15317,N_14333,N_14789);
or U15318 (N_15318,N_14271,N_14929);
nand U15319 (N_15319,N_14856,N_13923);
nor U15320 (N_15320,N_14547,N_14741);
and U15321 (N_15321,N_13912,N_13988);
nand U15322 (N_15322,N_13993,N_14090);
and U15323 (N_15323,N_14952,N_14444);
and U15324 (N_15324,N_14826,N_14851);
xnor U15325 (N_15325,N_14125,N_14455);
or U15326 (N_15326,N_14958,N_14504);
nor U15327 (N_15327,N_14723,N_14525);
xnor U15328 (N_15328,N_14728,N_14459);
nand U15329 (N_15329,N_13810,N_13937);
or U15330 (N_15330,N_13900,N_14179);
or U15331 (N_15331,N_13994,N_14022);
and U15332 (N_15332,N_14974,N_14130);
nor U15333 (N_15333,N_14946,N_14647);
xor U15334 (N_15334,N_14197,N_14586);
and U15335 (N_15335,N_14707,N_14915);
and U15336 (N_15336,N_13977,N_13869);
and U15337 (N_15337,N_13757,N_14431);
nor U15338 (N_15338,N_14540,N_13775);
nand U15339 (N_15339,N_13812,N_14344);
or U15340 (N_15340,N_14539,N_13770);
nor U15341 (N_15341,N_14640,N_14747);
nor U15342 (N_15342,N_14280,N_14853);
xor U15343 (N_15343,N_14427,N_13872);
xnor U15344 (N_15344,N_14362,N_14488);
or U15345 (N_15345,N_14874,N_13981);
nor U15346 (N_15346,N_14563,N_14048);
nand U15347 (N_15347,N_14758,N_13984);
xnor U15348 (N_15348,N_13919,N_14099);
nor U15349 (N_15349,N_14157,N_14968);
nand U15350 (N_15350,N_14489,N_14312);
and U15351 (N_15351,N_14290,N_14714);
nor U15352 (N_15352,N_13928,N_13996);
xnor U15353 (N_15353,N_13790,N_14367);
or U15354 (N_15354,N_14863,N_14374);
or U15355 (N_15355,N_14147,N_14252);
nand U15356 (N_15356,N_14212,N_14495);
nor U15357 (N_15357,N_14073,N_14141);
nand U15358 (N_15358,N_14569,N_14777);
and U15359 (N_15359,N_14260,N_14501);
or U15360 (N_15360,N_14415,N_13808);
or U15361 (N_15361,N_14822,N_14690);
or U15362 (N_15362,N_14602,N_14154);
xor U15363 (N_15363,N_14040,N_14277);
nand U15364 (N_15364,N_14188,N_13961);
or U15365 (N_15365,N_13761,N_14519);
and U15366 (N_15366,N_14581,N_14184);
and U15367 (N_15367,N_14051,N_14833);
and U15368 (N_15368,N_14191,N_14637);
or U15369 (N_15369,N_13931,N_14289);
nand U15370 (N_15370,N_14017,N_14732);
nor U15371 (N_15371,N_14850,N_14421);
or U15372 (N_15372,N_14817,N_14671);
and U15373 (N_15373,N_13848,N_14764);
and U15374 (N_15374,N_14638,N_13875);
nor U15375 (N_15375,N_14597,N_14322);
nand U15376 (N_15376,N_14782,N_14165);
and U15377 (N_15377,N_14528,N_14325);
nand U15378 (N_15378,N_14223,N_14975);
xnor U15379 (N_15379,N_14829,N_14583);
xnor U15380 (N_15380,N_14870,N_14121);
or U15381 (N_15381,N_14471,N_14283);
xor U15382 (N_15382,N_14247,N_14411);
and U15383 (N_15383,N_13929,N_13843);
nor U15384 (N_15384,N_14185,N_14584);
and U15385 (N_15385,N_14869,N_14655);
and U15386 (N_15386,N_14861,N_14046);
or U15387 (N_15387,N_14783,N_14033);
or U15388 (N_15388,N_14889,N_13924);
or U15389 (N_15389,N_14635,N_13960);
xnor U15390 (N_15390,N_14167,N_14793);
nand U15391 (N_15391,N_13827,N_14548);
or U15392 (N_15392,N_14953,N_13947);
xor U15393 (N_15393,N_14922,N_14438);
nand U15394 (N_15394,N_14294,N_13824);
nor U15395 (N_15395,N_14233,N_14701);
xnor U15396 (N_15396,N_14000,N_14146);
xnor U15397 (N_15397,N_14313,N_14550);
nor U15398 (N_15398,N_13942,N_14453);
nand U15399 (N_15399,N_14983,N_14766);
xor U15400 (N_15400,N_14393,N_14183);
xnor U15401 (N_15401,N_14763,N_14656);
nor U15402 (N_15402,N_14124,N_14262);
nor U15403 (N_15403,N_14568,N_14565);
and U15404 (N_15404,N_14627,N_14133);
and U15405 (N_15405,N_14287,N_14176);
or U15406 (N_15406,N_14078,N_13886);
nand U15407 (N_15407,N_14119,N_13979);
nor U15408 (N_15408,N_14699,N_14517);
or U15409 (N_15409,N_14527,N_13754);
and U15410 (N_15410,N_14089,N_14917);
xor U15411 (N_15411,N_14227,N_14521);
nor U15412 (N_15412,N_14796,N_14791);
nor U15413 (N_15413,N_14672,N_13876);
and U15414 (N_15414,N_14011,N_14003);
and U15415 (N_15415,N_13800,N_14663);
xor U15416 (N_15416,N_14397,N_14026);
nor U15417 (N_15417,N_13951,N_14661);
nand U15418 (N_15418,N_14885,N_14614);
nand U15419 (N_15419,N_14609,N_14074);
xnor U15420 (N_15420,N_14848,N_14128);
nor U15421 (N_15421,N_13769,N_14111);
nand U15422 (N_15422,N_14868,N_14895);
nand U15423 (N_15423,N_14904,N_14311);
nor U15424 (N_15424,N_14462,N_13897);
and U15425 (N_15425,N_14844,N_13795);
nor U15426 (N_15426,N_14266,N_13958);
nor U15427 (N_15427,N_14134,N_14756);
nor U15428 (N_15428,N_14066,N_14623);
xnor U15429 (N_15429,N_14933,N_14028);
or U15430 (N_15430,N_14735,N_13776);
or U15431 (N_15431,N_14386,N_14920);
nor U15432 (N_15432,N_14422,N_14573);
nand U15433 (N_15433,N_14248,N_14149);
nor U15434 (N_15434,N_13959,N_14377);
nor U15435 (N_15435,N_13817,N_13855);
xnor U15436 (N_15436,N_14705,N_13971);
and U15437 (N_15437,N_14409,N_14898);
nand U15438 (N_15438,N_14365,N_14215);
or U15439 (N_15439,N_14675,N_14053);
and U15440 (N_15440,N_14224,N_13922);
nor U15441 (N_15441,N_13914,N_14330);
and U15442 (N_15442,N_14057,N_14537);
nor U15443 (N_15443,N_13890,N_14912);
or U15444 (N_15444,N_14417,N_13926);
and U15445 (N_15445,N_14131,N_14370);
xnor U15446 (N_15446,N_13851,N_13809);
and U15447 (N_15447,N_14831,N_14486);
and U15448 (N_15448,N_14593,N_14361);
xor U15449 (N_15449,N_14020,N_14769);
nand U15450 (N_15450,N_14350,N_13818);
nand U15451 (N_15451,N_14680,N_14558);
nor U15452 (N_15452,N_14960,N_14402);
nand U15453 (N_15453,N_14804,N_14808);
and U15454 (N_15454,N_14391,N_14470);
or U15455 (N_15455,N_14419,N_13831);
or U15456 (N_15456,N_14479,N_14364);
nor U15457 (N_15457,N_14288,N_14695);
xor U15458 (N_15458,N_14282,N_13844);
nand U15459 (N_15459,N_13986,N_14295);
nand U15460 (N_15460,N_13983,N_14499);
nor U15461 (N_15461,N_14070,N_14543);
or U15462 (N_15462,N_14691,N_14599);
xnor U15463 (N_15463,N_14927,N_14939);
and U15464 (N_15464,N_14982,N_14269);
xor U15465 (N_15465,N_14076,N_13860);
nor U15466 (N_15466,N_13783,N_14103);
nor U15467 (N_15467,N_14304,N_14916);
or U15468 (N_15468,N_14710,N_14268);
or U15469 (N_15469,N_13805,N_14241);
nand U15470 (N_15470,N_14317,N_14802);
and U15471 (N_15471,N_13968,N_14696);
and U15472 (N_15472,N_14538,N_14088);
or U15473 (N_15473,N_14992,N_14746);
xnor U15474 (N_15474,N_14987,N_14360);
nor U15475 (N_15475,N_14533,N_14342);
nand U15476 (N_15476,N_13871,N_13930);
xor U15477 (N_15477,N_14151,N_14068);
or U15478 (N_15478,N_14903,N_14204);
and U15479 (N_15479,N_13939,N_13917);
nor U15480 (N_15480,N_13792,N_14965);
or U15481 (N_15481,N_14358,N_14616);
and U15482 (N_15482,N_14575,N_14620);
nand U15483 (N_15483,N_13841,N_14182);
xnor U15484 (N_15484,N_14013,N_14923);
and U15485 (N_15485,N_14742,N_14343);
or U15486 (N_15486,N_14555,N_14932);
or U15487 (N_15487,N_14513,N_14570);
xor U15488 (N_15488,N_14888,N_13887);
nand U15489 (N_15489,N_14585,N_13807);
and U15490 (N_15490,N_14825,N_14998);
nor U15491 (N_15491,N_14871,N_14296);
or U15492 (N_15492,N_14164,N_14617);
and U15493 (N_15493,N_14837,N_14840);
xor U15494 (N_15494,N_14636,N_14852);
nand U15495 (N_15495,N_14834,N_14253);
xor U15496 (N_15496,N_14886,N_14925);
nand U15497 (N_15497,N_14726,N_13842);
xor U15498 (N_15498,N_14729,N_14067);
and U15499 (N_15499,N_14001,N_14083);
nand U15500 (N_15500,N_14842,N_14914);
xor U15501 (N_15501,N_13861,N_13803);
or U15502 (N_15502,N_14300,N_13806);
xor U15503 (N_15503,N_14651,N_13976);
nand U15504 (N_15504,N_14712,N_14084);
nor U15505 (N_15505,N_14153,N_14291);
nand U15506 (N_15506,N_14400,N_14571);
nor U15507 (N_15507,N_14163,N_14014);
nand U15508 (N_15508,N_14054,N_14150);
nand U15509 (N_15509,N_14591,N_14178);
or U15510 (N_15510,N_14379,N_13980);
xnor U15511 (N_15511,N_14395,N_14303);
nand U15512 (N_15512,N_14447,N_13874);
or U15513 (N_15513,N_14911,N_14174);
or U15514 (N_15514,N_14991,N_13793);
nor U15515 (N_15515,N_14245,N_14875);
nor U15516 (N_15516,N_13953,N_14815);
or U15517 (N_15517,N_14355,N_14440);
and U15518 (N_15518,N_13780,N_14938);
xnor U15519 (N_15519,N_13899,N_14426);
nand U15520 (N_15520,N_13952,N_13794);
and U15521 (N_15521,N_14019,N_14264);
nor U15522 (N_15522,N_13877,N_14025);
xnor U15523 (N_15523,N_14950,N_14055);
and U15524 (N_15524,N_14445,N_14216);
and U15525 (N_15525,N_14948,N_14664);
nor U15526 (N_15526,N_14328,N_13985);
and U15527 (N_15527,N_14036,N_13910);
xnor U15528 (N_15528,N_14345,N_13863);
and U15529 (N_15529,N_14897,N_14381);
and U15530 (N_15530,N_14220,N_14653);
and U15531 (N_15531,N_14097,N_14908);
nand U15532 (N_15532,N_14439,N_14619);
and U15533 (N_15533,N_13944,N_14776);
nand U15534 (N_15534,N_14700,N_14743);
nor U15535 (N_15535,N_14211,N_14755);
or U15536 (N_15536,N_14795,N_13964);
or U15537 (N_15537,N_14546,N_14926);
nor U15538 (N_15538,N_13756,N_14673);
and U15539 (N_15539,N_14734,N_14566);
and U15540 (N_15540,N_14316,N_14966);
xnor U15541 (N_15541,N_14598,N_14064);
xnor U15542 (N_15542,N_14827,N_13892);
and U15543 (N_15543,N_14413,N_13804);
nor U15544 (N_15544,N_14239,N_14461);
or U15545 (N_15545,N_14382,N_14085);
and U15546 (N_15546,N_14754,N_14209);
nand U15547 (N_15547,N_14137,N_13853);
or U15548 (N_15548,N_14702,N_14578);
xnor U15549 (N_15549,N_14858,N_14594);
nand U15550 (N_15550,N_14430,N_14352);
nand U15551 (N_15551,N_13801,N_14751);
nor U15552 (N_15552,N_14949,N_14045);
or U15553 (N_15553,N_13779,N_14608);
xnor U15554 (N_15554,N_14270,N_14901);
nand U15555 (N_15555,N_13913,N_14091);
xnor U15556 (N_15556,N_14086,N_14709);
nand U15557 (N_15557,N_14659,N_14238);
nand U15558 (N_15558,N_13833,N_14210);
or U15559 (N_15559,N_14112,N_13995);
xnor U15560 (N_15560,N_13765,N_14336);
nand U15561 (N_15561,N_14683,N_14292);
nand U15562 (N_15562,N_14942,N_14873);
nand U15563 (N_15563,N_13834,N_13854);
and U15564 (N_15564,N_14752,N_14496);
xor U15565 (N_15565,N_14662,N_13882);
nand U15566 (N_15566,N_14830,N_13773);
or U15567 (N_15567,N_13943,N_14458);
and U15568 (N_15568,N_14205,N_13829);
nor U15569 (N_15569,N_14824,N_14947);
or U15570 (N_15570,N_14403,N_13883);
and U15571 (N_15571,N_14587,N_14075);
and U15572 (N_15572,N_14229,N_13920);
or U15573 (N_15573,N_14226,N_13896);
or U15574 (N_15574,N_14032,N_14553);
xor U15575 (N_15575,N_14899,N_14639);
nand U15576 (N_15576,N_13927,N_14140);
and U15577 (N_15577,N_14767,N_14396);
xor U15578 (N_15578,N_13987,N_14196);
and U15579 (N_15579,N_14857,N_14650);
and U15580 (N_15580,N_14632,N_14725);
nand U15581 (N_15581,N_14357,N_14474);
or U15582 (N_15582,N_14307,N_14319);
and U15583 (N_15583,N_14442,N_13955);
xnor U15584 (N_15584,N_13785,N_14490);
xor U15585 (N_15585,N_13820,N_14372);
and U15586 (N_15586,N_14604,N_14907);
or U15587 (N_15587,N_13828,N_14613);
nor U15588 (N_15588,N_14797,N_14642);
or U15589 (N_15589,N_14321,N_14792);
nor U15590 (N_15590,N_14676,N_13786);
nor U15591 (N_15591,N_14839,N_14039);
nor U15592 (N_15592,N_14042,N_14518);
or U15593 (N_15593,N_14959,N_14082);
xor U15594 (N_15594,N_14052,N_14338);
nor U15595 (N_15595,N_14688,N_14800);
and U15596 (N_15596,N_14044,N_14626);
and U15597 (N_15597,N_14913,N_14500);
and U15598 (N_15598,N_14228,N_13856);
or U15599 (N_15599,N_14954,N_14979);
and U15600 (N_15600,N_14326,N_14168);
or U15601 (N_15601,N_13901,N_14628);
and U15602 (N_15602,N_14999,N_14706);
nor U15603 (N_15603,N_14278,N_14466);
xor U15604 (N_15604,N_14368,N_14004);
and U15605 (N_15605,N_13826,N_14190);
nor U15606 (N_15606,N_14894,N_14255);
and U15607 (N_15607,N_14811,N_14366);
nand U15608 (N_15608,N_14175,N_14275);
and U15609 (N_15609,N_14027,N_14392);
or U15610 (N_15610,N_14340,N_14143);
xor U15611 (N_15611,N_14768,N_13823);
nand U15612 (N_15612,N_14348,N_14978);
xnor U15613 (N_15613,N_14745,N_14629);
nor U15614 (N_15614,N_13767,N_14610);
xor U15615 (N_15615,N_13832,N_13966);
xor U15616 (N_15616,N_14801,N_13864);
nand U15617 (N_15617,N_14930,N_13894);
and U15618 (N_15618,N_14169,N_14106);
or U15619 (N_15619,N_13752,N_13903);
nor U15620 (N_15620,N_14498,N_14180);
or U15621 (N_15621,N_14809,N_14865);
and U15622 (N_15622,N_14805,N_14341);
nand U15623 (N_15623,N_14698,N_14686);
nand U15624 (N_15624,N_14739,N_13782);
xor U15625 (N_15625,N_13858,N_14325);
or U15626 (N_15626,N_13901,N_13767);
nand U15627 (N_15627,N_14721,N_13883);
nor U15628 (N_15628,N_14644,N_14189);
and U15629 (N_15629,N_14743,N_14798);
xor U15630 (N_15630,N_13794,N_14462);
xnor U15631 (N_15631,N_14477,N_13981);
nor U15632 (N_15632,N_14356,N_13793);
xor U15633 (N_15633,N_14401,N_13857);
nor U15634 (N_15634,N_14747,N_13832);
nor U15635 (N_15635,N_14734,N_13780);
xor U15636 (N_15636,N_13889,N_14275);
and U15637 (N_15637,N_13793,N_14307);
xnor U15638 (N_15638,N_14354,N_14356);
nand U15639 (N_15639,N_14345,N_13919);
and U15640 (N_15640,N_14698,N_13872);
or U15641 (N_15641,N_14930,N_14422);
xnor U15642 (N_15642,N_14731,N_14533);
nor U15643 (N_15643,N_14417,N_14889);
or U15644 (N_15644,N_14159,N_14097);
nor U15645 (N_15645,N_14857,N_14688);
xor U15646 (N_15646,N_14843,N_14014);
nor U15647 (N_15647,N_14968,N_13885);
and U15648 (N_15648,N_14918,N_13825);
or U15649 (N_15649,N_14657,N_14058);
xor U15650 (N_15650,N_14231,N_13984);
xor U15651 (N_15651,N_14768,N_13775);
and U15652 (N_15652,N_13892,N_14873);
nand U15653 (N_15653,N_14220,N_14598);
and U15654 (N_15654,N_14039,N_14504);
nand U15655 (N_15655,N_14129,N_13761);
and U15656 (N_15656,N_14286,N_13830);
nand U15657 (N_15657,N_14332,N_14312);
nor U15658 (N_15658,N_14232,N_14315);
nor U15659 (N_15659,N_14625,N_14243);
nor U15660 (N_15660,N_14048,N_14676);
nand U15661 (N_15661,N_14484,N_14984);
nor U15662 (N_15662,N_13832,N_14084);
and U15663 (N_15663,N_13752,N_14542);
or U15664 (N_15664,N_13924,N_14454);
or U15665 (N_15665,N_14548,N_14660);
nand U15666 (N_15666,N_14080,N_14175);
nor U15667 (N_15667,N_14251,N_14446);
nand U15668 (N_15668,N_13819,N_14360);
or U15669 (N_15669,N_14439,N_13936);
and U15670 (N_15670,N_14602,N_14457);
and U15671 (N_15671,N_13969,N_13919);
nand U15672 (N_15672,N_14867,N_14170);
xnor U15673 (N_15673,N_14938,N_14018);
xnor U15674 (N_15674,N_14427,N_14429);
and U15675 (N_15675,N_13960,N_14178);
xnor U15676 (N_15676,N_14313,N_14469);
or U15677 (N_15677,N_14704,N_13791);
or U15678 (N_15678,N_14279,N_14063);
or U15679 (N_15679,N_14026,N_14294);
nor U15680 (N_15680,N_13961,N_14800);
or U15681 (N_15681,N_13924,N_14891);
xor U15682 (N_15682,N_14471,N_14123);
nand U15683 (N_15683,N_14508,N_13998);
nand U15684 (N_15684,N_14864,N_14592);
and U15685 (N_15685,N_14297,N_13882);
nand U15686 (N_15686,N_14229,N_14001);
or U15687 (N_15687,N_13890,N_14311);
xnor U15688 (N_15688,N_14031,N_14199);
nor U15689 (N_15689,N_14347,N_13890);
or U15690 (N_15690,N_14193,N_13998);
xor U15691 (N_15691,N_13969,N_13865);
and U15692 (N_15692,N_14230,N_14795);
or U15693 (N_15693,N_14418,N_14992);
and U15694 (N_15694,N_14703,N_14232);
or U15695 (N_15695,N_14003,N_14801);
or U15696 (N_15696,N_14287,N_13929);
nand U15697 (N_15697,N_14089,N_14593);
nor U15698 (N_15698,N_13833,N_13866);
or U15699 (N_15699,N_14266,N_13911);
and U15700 (N_15700,N_13976,N_14430);
nor U15701 (N_15701,N_14861,N_13994);
xor U15702 (N_15702,N_14470,N_14363);
xnor U15703 (N_15703,N_14914,N_14968);
nand U15704 (N_15704,N_14629,N_13799);
or U15705 (N_15705,N_14239,N_13908);
nand U15706 (N_15706,N_14167,N_13896);
xor U15707 (N_15707,N_13781,N_14857);
and U15708 (N_15708,N_14320,N_13828);
xnor U15709 (N_15709,N_14475,N_14926);
and U15710 (N_15710,N_14739,N_14736);
or U15711 (N_15711,N_14271,N_14641);
and U15712 (N_15712,N_14966,N_14293);
nand U15713 (N_15713,N_14816,N_14396);
or U15714 (N_15714,N_14671,N_14622);
xnor U15715 (N_15715,N_13868,N_14760);
and U15716 (N_15716,N_14431,N_14986);
xor U15717 (N_15717,N_14203,N_13970);
nand U15718 (N_15718,N_14562,N_13999);
and U15719 (N_15719,N_14502,N_14210);
or U15720 (N_15720,N_13993,N_13750);
or U15721 (N_15721,N_14024,N_14759);
and U15722 (N_15722,N_14878,N_14951);
xnor U15723 (N_15723,N_13765,N_14617);
and U15724 (N_15724,N_13905,N_14291);
nor U15725 (N_15725,N_14556,N_14063);
or U15726 (N_15726,N_14589,N_14578);
nor U15727 (N_15727,N_14134,N_14245);
nor U15728 (N_15728,N_13992,N_14399);
or U15729 (N_15729,N_14812,N_14685);
nor U15730 (N_15730,N_14411,N_14091);
and U15731 (N_15731,N_14990,N_14049);
xnor U15732 (N_15732,N_13826,N_14614);
nand U15733 (N_15733,N_13975,N_14753);
xor U15734 (N_15734,N_14762,N_14749);
nor U15735 (N_15735,N_14175,N_14319);
nand U15736 (N_15736,N_14297,N_13804);
nand U15737 (N_15737,N_14424,N_14620);
nand U15738 (N_15738,N_14730,N_14255);
or U15739 (N_15739,N_14444,N_13887);
nand U15740 (N_15740,N_14441,N_14337);
nor U15741 (N_15741,N_14270,N_14121);
xor U15742 (N_15742,N_14299,N_14487);
and U15743 (N_15743,N_13897,N_13767);
and U15744 (N_15744,N_14430,N_14327);
nor U15745 (N_15745,N_14987,N_14656);
and U15746 (N_15746,N_14862,N_14587);
and U15747 (N_15747,N_14374,N_14381);
nand U15748 (N_15748,N_14267,N_13981);
xor U15749 (N_15749,N_13766,N_14033);
or U15750 (N_15750,N_14945,N_14329);
nor U15751 (N_15751,N_14834,N_14140);
or U15752 (N_15752,N_14183,N_13953);
xor U15753 (N_15753,N_14039,N_14674);
nand U15754 (N_15754,N_14277,N_13851);
and U15755 (N_15755,N_14123,N_14158);
or U15756 (N_15756,N_14260,N_14070);
xor U15757 (N_15757,N_14327,N_14539);
or U15758 (N_15758,N_14931,N_14145);
nand U15759 (N_15759,N_14858,N_14505);
nor U15760 (N_15760,N_14615,N_14549);
nor U15761 (N_15761,N_14832,N_14057);
or U15762 (N_15762,N_14032,N_14506);
and U15763 (N_15763,N_14444,N_14382);
and U15764 (N_15764,N_14489,N_13800);
nor U15765 (N_15765,N_14629,N_14815);
and U15766 (N_15766,N_14411,N_14151);
nand U15767 (N_15767,N_14768,N_14444);
xnor U15768 (N_15768,N_13893,N_14390);
nand U15769 (N_15769,N_13894,N_14971);
or U15770 (N_15770,N_14673,N_14257);
nor U15771 (N_15771,N_14682,N_14236);
and U15772 (N_15772,N_14693,N_14949);
nand U15773 (N_15773,N_13861,N_13846);
nand U15774 (N_15774,N_14804,N_14696);
nor U15775 (N_15775,N_14485,N_14765);
xnor U15776 (N_15776,N_13944,N_14311);
and U15777 (N_15777,N_14869,N_14510);
and U15778 (N_15778,N_14742,N_14021);
nand U15779 (N_15779,N_13843,N_14839);
and U15780 (N_15780,N_14327,N_13762);
nand U15781 (N_15781,N_14814,N_13790);
xnor U15782 (N_15782,N_14328,N_14253);
nand U15783 (N_15783,N_14808,N_14796);
nor U15784 (N_15784,N_13991,N_13778);
xor U15785 (N_15785,N_14118,N_14138);
or U15786 (N_15786,N_14525,N_14632);
and U15787 (N_15787,N_13996,N_14349);
or U15788 (N_15788,N_14533,N_14827);
and U15789 (N_15789,N_13839,N_14971);
nor U15790 (N_15790,N_14868,N_14599);
nand U15791 (N_15791,N_14985,N_14687);
or U15792 (N_15792,N_14828,N_14124);
nor U15793 (N_15793,N_14366,N_14317);
xor U15794 (N_15794,N_13966,N_14124);
nand U15795 (N_15795,N_14548,N_14610);
nand U15796 (N_15796,N_14941,N_13842);
nor U15797 (N_15797,N_14597,N_14546);
and U15798 (N_15798,N_14706,N_13863);
or U15799 (N_15799,N_14095,N_14803);
xor U15800 (N_15800,N_14854,N_14545);
xor U15801 (N_15801,N_13760,N_14439);
or U15802 (N_15802,N_14893,N_14488);
xnor U15803 (N_15803,N_14160,N_13761);
nor U15804 (N_15804,N_14291,N_13753);
and U15805 (N_15805,N_14297,N_14042);
and U15806 (N_15806,N_14886,N_14882);
nor U15807 (N_15807,N_13857,N_13953);
nand U15808 (N_15808,N_14531,N_13762);
and U15809 (N_15809,N_14567,N_13926);
nand U15810 (N_15810,N_14950,N_14369);
and U15811 (N_15811,N_14732,N_14366);
and U15812 (N_15812,N_14931,N_14354);
nor U15813 (N_15813,N_13894,N_14504);
nand U15814 (N_15814,N_13914,N_13912);
nand U15815 (N_15815,N_14476,N_13840);
nand U15816 (N_15816,N_14461,N_14802);
nor U15817 (N_15817,N_14739,N_14807);
and U15818 (N_15818,N_14788,N_14545);
nand U15819 (N_15819,N_14557,N_14067);
nor U15820 (N_15820,N_14504,N_14771);
nor U15821 (N_15821,N_13801,N_14863);
nand U15822 (N_15822,N_14097,N_13754);
nor U15823 (N_15823,N_14037,N_14616);
xnor U15824 (N_15824,N_14330,N_14654);
xnor U15825 (N_15825,N_14555,N_13943);
and U15826 (N_15826,N_14402,N_14515);
xor U15827 (N_15827,N_14294,N_14141);
and U15828 (N_15828,N_14122,N_13775);
and U15829 (N_15829,N_14973,N_14810);
nor U15830 (N_15830,N_14791,N_14770);
and U15831 (N_15831,N_14150,N_14125);
nor U15832 (N_15832,N_13996,N_14447);
xor U15833 (N_15833,N_13949,N_14109);
or U15834 (N_15834,N_14185,N_14838);
xnor U15835 (N_15835,N_14657,N_14113);
and U15836 (N_15836,N_14890,N_14853);
nand U15837 (N_15837,N_13859,N_13799);
nand U15838 (N_15838,N_14602,N_13881);
nor U15839 (N_15839,N_14106,N_14347);
or U15840 (N_15840,N_14518,N_14069);
xor U15841 (N_15841,N_14617,N_14116);
nor U15842 (N_15842,N_13923,N_14756);
nand U15843 (N_15843,N_14667,N_14761);
and U15844 (N_15844,N_14892,N_14213);
and U15845 (N_15845,N_14622,N_14045);
or U15846 (N_15846,N_13789,N_14955);
and U15847 (N_15847,N_14880,N_13981);
nand U15848 (N_15848,N_14122,N_13764);
nand U15849 (N_15849,N_14699,N_14073);
nor U15850 (N_15850,N_14971,N_13999);
nand U15851 (N_15851,N_14533,N_14086);
xor U15852 (N_15852,N_14996,N_14407);
and U15853 (N_15853,N_13753,N_14986);
or U15854 (N_15854,N_14432,N_14272);
nor U15855 (N_15855,N_14066,N_13893);
xnor U15856 (N_15856,N_14242,N_14260);
or U15857 (N_15857,N_14583,N_14780);
nand U15858 (N_15858,N_14131,N_14032);
nand U15859 (N_15859,N_14321,N_14521);
or U15860 (N_15860,N_13990,N_14990);
xnor U15861 (N_15861,N_14805,N_13946);
nand U15862 (N_15862,N_14352,N_14757);
xnor U15863 (N_15863,N_13819,N_14271);
xor U15864 (N_15864,N_14988,N_14658);
xnor U15865 (N_15865,N_14856,N_14074);
or U15866 (N_15866,N_14000,N_14102);
nor U15867 (N_15867,N_14892,N_14762);
or U15868 (N_15868,N_13752,N_14673);
nand U15869 (N_15869,N_14586,N_14411);
xor U15870 (N_15870,N_14874,N_13795);
nand U15871 (N_15871,N_14647,N_14589);
nor U15872 (N_15872,N_13871,N_14501);
or U15873 (N_15873,N_13897,N_13756);
nand U15874 (N_15874,N_14608,N_14094);
nor U15875 (N_15875,N_13840,N_13926);
nor U15876 (N_15876,N_14467,N_14443);
nand U15877 (N_15877,N_14561,N_14072);
xor U15878 (N_15878,N_13919,N_14175);
and U15879 (N_15879,N_14536,N_13783);
nand U15880 (N_15880,N_14597,N_14652);
xnor U15881 (N_15881,N_13936,N_13966);
nand U15882 (N_15882,N_14616,N_14170);
nor U15883 (N_15883,N_14033,N_14655);
nor U15884 (N_15884,N_14626,N_14661);
and U15885 (N_15885,N_13852,N_13776);
xnor U15886 (N_15886,N_13783,N_14863);
xnor U15887 (N_15887,N_14829,N_14920);
nand U15888 (N_15888,N_14500,N_14056);
nand U15889 (N_15889,N_13816,N_13822);
and U15890 (N_15890,N_13860,N_13965);
nor U15891 (N_15891,N_14619,N_14898);
nand U15892 (N_15892,N_14007,N_14545);
nor U15893 (N_15893,N_14406,N_14231);
xnor U15894 (N_15894,N_14435,N_14523);
nor U15895 (N_15895,N_14071,N_14327);
or U15896 (N_15896,N_14565,N_14391);
or U15897 (N_15897,N_14736,N_13858);
or U15898 (N_15898,N_14753,N_13928);
or U15899 (N_15899,N_13776,N_14033);
or U15900 (N_15900,N_14322,N_14146);
nor U15901 (N_15901,N_13886,N_13952);
xor U15902 (N_15902,N_14256,N_14482);
and U15903 (N_15903,N_14334,N_14907);
and U15904 (N_15904,N_14418,N_13953);
nor U15905 (N_15905,N_14435,N_14045);
and U15906 (N_15906,N_14453,N_14065);
xnor U15907 (N_15907,N_14323,N_14637);
xnor U15908 (N_15908,N_14162,N_14564);
or U15909 (N_15909,N_14419,N_14662);
xnor U15910 (N_15910,N_14716,N_14195);
or U15911 (N_15911,N_14657,N_13832);
nand U15912 (N_15912,N_13785,N_14988);
nand U15913 (N_15913,N_14691,N_13835);
xor U15914 (N_15914,N_14113,N_14122);
nand U15915 (N_15915,N_14796,N_13800);
nand U15916 (N_15916,N_14099,N_14076);
xnor U15917 (N_15917,N_14562,N_14893);
xor U15918 (N_15918,N_14708,N_14027);
nor U15919 (N_15919,N_14652,N_14266);
or U15920 (N_15920,N_13930,N_14212);
or U15921 (N_15921,N_14972,N_14169);
xnor U15922 (N_15922,N_13982,N_14040);
and U15923 (N_15923,N_13773,N_14530);
nand U15924 (N_15924,N_14496,N_13958);
and U15925 (N_15925,N_14799,N_14765);
xnor U15926 (N_15926,N_14460,N_14620);
nand U15927 (N_15927,N_14304,N_14561);
or U15928 (N_15928,N_13927,N_14851);
and U15929 (N_15929,N_14015,N_14461);
or U15930 (N_15930,N_13972,N_14859);
xnor U15931 (N_15931,N_13925,N_14967);
xor U15932 (N_15932,N_14674,N_14725);
nand U15933 (N_15933,N_14563,N_14808);
nand U15934 (N_15934,N_14906,N_14937);
nor U15935 (N_15935,N_14048,N_14592);
nand U15936 (N_15936,N_14989,N_14534);
nand U15937 (N_15937,N_14144,N_14056);
nor U15938 (N_15938,N_14887,N_13768);
nor U15939 (N_15939,N_14807,N_14865);
nand U15940 (N_15940,N_14410,N_14530);
nand U15941 (N_15941,N_14849,N_14915);
xnor U15942 (N_15942,N_14072,N_13776);
and U15943 (N_15943,N_13885,N_14479);
and U15944 (N_15944,N_14345,N_14952);
nand U15945 (N_15945,N_14907,N_14351);
nand U15946 (N_15946,N_13892,N_14039);
xnor U15947 (N_15947,N_14620,N_14018);
or U15948 (N_15948,N_14852,N_14821);
nand U15949 (N_15949,N_13984,N_14282);
or U15950 (N_15950,N_14070,N_13937);
or U15951 (N_15951,N_14075,N_13854);
xnor U15952 (N_15952,N_14213,N_14212);
and U15953 (N_15953,N_14764,N_14700);
and U15954 (N_15954,N_14628,N_14399);
xor U15955 (N_15955,N_14436,N_14547);
nand U15956 (N_15956,N_14548,N_14606);
nand U15957 (N_15957,N_14491,N_14720);
nor U15958 (N_15958,N_13798,N_14793);
nor U15959 (N_15959,N_14821,N_14655);
nor U15960 (N_15960,N_14440,N_14839);
nand U15961 (N_15961,N_14053,N_14356);
or U15962 (N_15962,N_14499,N_14097);
nand U15963 (N_15963,N_14576,N_14331);
nor U15964 (N_15964,N_14998,N_14838);
nor U15965 (N_15965,N_13867,N_14128);
and U15966 (N_15966,N_14426,N_14107);
and U15967 (N_15967,N_14973,N_14994);
nor U15968 (N_15968,N_14571,N_14188);
and U15969 (N_15969,N_14325,N_14906);
xnor U15970 (N_15970,N_13900,N_14908);
nand U15971 (N_15971,N_14847,N_14472);
nand U15972 (N_15972,N_13979,N_14270);
nand U15973 (N_15973,N_13795,N_13938);
xnor U15974 (N_15974,N_14199,N_14906);
nand U15975 (N_15975,N_14950,N_14777);
and U15976 (N_15976,N_14861,N_14250);
nor U15977 (N_15977,N_14201,N_14891);
nand U15978 (N_15978,N_14906,N_14708);
xnor U15979 (N_15979,N_13786,N_13891);
and U15980 (N_15980,N_14720,N_14389);
nor U15981 (N_15981,N_14277,N_14540);
xnor U15982 (N_15982,N_14253,N_14778);
xor U15983 (N_15983,N_14461,N_14299);
and U15984 (N_15984,N_14225,N_14175);
nand U15985 (N_15985,N_14792,N_13783);
nor U15986 (N_15986,N_14617,N_14262);
xor U15987 (N_15987,N_14709,N_13857);
or U15988 (N_15988,N_13948,N_14658);
nand U15989 (N_15989,N_14882,N_14892);
nor U15990 (N_15990,N_14168,N_14446);
and U15991 (N_15991,N_13792,N_14638);
nor U15992 (N_15992,N_14714,N_13968);
xor U15993 (N_15993,N_14277,N_14080);
and U15994 (N_15994,N_14133,N_14878);
and U15995 (N_15995,N_14380,N_13965);
or U15996 (N_15996,N_14210,N_14670);
or U15997 (N_15997,N_14317,N_14292);
and U15998 (N_15998,N_14747,N_14423);
or U15999 (N_15999,N_14370,N_13801);
and U16000 (N_16000,N_14558,N_14018);
or U16001 (N_16001,N_14690,N_14027);
xnor U16002 (N_16002,N_13845,N_13761);
nor U16003 (N_16003,N_13823,N_13810);
nand U16004 (N_16004,N_14855,N_13760);
nand U16005 (N_16005,N_13924,N_14088);
xnor U16006 (N_16006,N_14645,N_14795);
nand U16007 (N_16007,N_14688,N_14856);
and U16008 (N_16008,N_14584,N_14667);
nor U16009 (N_16009,N_14025,N_14235);
xnor U16010 (N_16010,N_13893,N_14927);
nor U16011 (N_16011,N_14619,N_14464);
xnor U16012 (N_16012,N_14442,N_14004);
or U16013 (N_16013,N_13889,N_14587);
nor U16014 (N_16014,N_14433,N_13984);
nor U16015 (N_16015,N_14840,N_13957);
and U16016 (N_16016,N_14739,N_14932);
and U16017 (N_16017,N_14862,N_14383);
nand U16018 (N_16018,N_14150,N_14596);
nor U16019 (N_16019,N_13814,N_14690);
nor U16020 (N_16020,N_14199,N_14996);
or U16021 (N_16021,N_14357,N_14453);
or U16022 (N_16022,N_14527,N_14089);
and U16023 (N_16023,N_14655,N_13771);
and U16024 (N_16024,N_13819,N_14433);
xnor U16025 (N_16025,N_14701,N_14903);
nand U16026 (N_16026,N_14509,N_14714);
xor U16027 (N_16027,N_14181,N_14115);
and U16028 (N_16028,N_14909,N_14600);
and U16029 (N_16029,N_14024,N_14916);
and U16030 (N_16030,N_14900,N_13809);
and U16031 (N_16031,N_14190,N_14144);
nand U16032 (N_16032,N_14234,N_14758);
nand U16033 (N_16033,N_14251,N_14019);
or U16034 (N_16034,N_13944,N_14509);
xor U16035 (N_16035,N_13822,N_14421);
nand U16036 (N_16036,N_14979,N_14625);
xnor U16037 (N_16037,N_14026,N_13916);
and U16038 (N_16038,N_14647,N_13913);
xor U16039 (N_16039,N_14672,N_14542);
nand U16040 (N_16040,N_14573,N_14411);
and U16041 (N_16041,N_14958,N_14708);
xnor U16042 (N_16042,N_14311,N_13876);
nor U16043 (N_16043,N_14407,N_14104);
and U16044 (N_16044,N_14765,N_13998);
xnor U16045 (N_16045,N_14056,N_13910);
xor U16046 (N_16046,N_14884,N_14782);
and U16047 (N_16047,N_14740,N_14812);
xnor U16048 (N_16048,N_13809,N_14494);
nor U16049 (N_16049,N_14424,N_14863);
nand U16050 (N_16050,N_14262,N_14134);
nand U16051 (N_16051,N_14597,N_14857);
and U16052 (N_16052,N_14170,N_14998);
nand U16053 (N_16053,N_14764,N_14644);
xnor U16054 (N_16054,N_14498,N_14323);
nor U16055 (N_16055,N_14967,N_13820);
nand U16056 (N_16056,N_14214,N_14185);
xnor U16057 (N_16057,N_14497,N_13852);
nor U16058 (N_16058,N_13800,N_14650);
or U16059 (N_16059,N_14244,N_14206);
or U16060 (N_16060,N_13993,N_13909);
xnor U16061 (N_16061,N_14826,N_14681);
nor U16062 (N_16062,N_14892,N_14653);
nand U16063 (N_16063,N_13907,N_14838);
nor U16064 (N_16064,N_13976,N_14249);
or U16065 (N_16065,N_14901,N_14643);
or U16066 (N_16066,N_14512,N_14438);
or U16067 (N_16067,N_13850,N_13766);
or U16068 (N_16068,N_13929,N_14987);
and U16069 (N_16069,N_14360,N_14409);
xor U16070 (N_16070,N_13866,N_14846);
and U16071 (N_16071,N_14558,N_14584);
nand U16072 (N_16072,N_13837,N_14214);
nand U16073 (N_16073,N_13862,N_14593);
or U16074 (N_16074,N_14995,N_14913);
and U16075 (N_16075,N_14947,N_14287);
and U16076 (N_16076,N_14781,N_14895);
and U16077 (N_16077,N_14287,N_13998);
nand U16078 (N_16078,N_14831,N_14173);
nor U16079 (N_16079,N_14587,N_14299);
nand U16080 (N_16080,N_14399,N_14177);
and U16081 (N_16081,N_14693,N_14452);
nand U16082 (N_16082,N_14718,N_14423);
nor U16083 (N_16083,N_14615,N_13942);
and U16084 (N_16084,N_14387,N_14406);
and U16085 (N_16085,N_14658,N_14432);
nand U16086 (N_16086,N_14975,N_14570);
xor U16087 (N_16087,N_14593,N_14862);
xor U16088 (N_16088,N_14635,N_13759);
and U16089 (N_16089,N_14583,N_14578);
xor U16090 (N_16090,N_13842,N_14851);
and U16091 (N_16091,N_14744,N_14968);
nor U16092 (N_16092,N_13759,N_14122);
nor U16093 (N_16093,N_13837,N_14887);
xnor U16094 (N_16094,N_14703,N_13798);
or U16095 (N_16095,N_14822,N_14261);
xor U16096 (N_16096,N_13851,N_14294);
and U16097 (N_16097,N_14641,N_14143);
and U16098 (N_16098,N_14739,N_14568);
and U16099 (N_16099,N_14923,N_14906);
or U16100 (N_16100,N_14239,N_14390);
xnor U16101 (N_16101,N_14968,N_14729);
nor U16102 (N_16102,N_14352,N_14656);
nor U16103 (N_16103,N_14775,N_14416);
and U16104 (N_16104,N_14803,N_14084);
nor U16105 (N_16105,N_14041,N_14152);
and U16106 (N_16106,N_14407,N_14398);
nand U16107 (N_16107,N_14230,N_14481);
xnor U16108 (N_16108,N_13760,N_13827);
nor U16109 (N_16109,N_14286,N_14877);
xor U16110 (N_16110,N_14844,N_14027);
xnor U16111 (N_16111,N_14138,N_14361);
and U16112 (N_16112,N_14020,N_14225);
xor U16113 (N_16113,N_14918,N_14956);
nand U16114 (N_16114,N_14303,N_14616);
nor U16115 (N_16115,N_14569,N_14735);
xnor U16116 (N_16116,N_14608,N_13866);
xor U16117 (N_16117,N_14765,N_14187);
or U16118 (N_16118,N_13957,N_14182);
and U16119 (N_16119,N_14383,N_14189);
nor U16120 (N_16120,N_14278,N_14807);
nand U16121 (N_16121,N_14857,N_14356);
and U16122 (N_16122,N_14255,N_13849);
xnor U16123 (N_16123,N_13910,N_14997);
nor U16124 (N_16124,N_14579,N_13963);
nand U16125 (N_16125,N_14527,N_14641);
or U16126 (N_16126,N_14471,N_13792);
xor U16127 (N_16127,N_13904,N_14954);
nand U16128 (N_16128,N_14212,N_13854);
xor U16129 (N_16129,N_13979,N_14521);
and U16130 (N_16130,N_14787,N_14868);
nand U16131 (N_16131,N_14069,N_14655);
nand U16132 (N_16132,N_14043,N_14042);
xor U16133 (N_16133,N_14398,N_14432);
nor U16134 (N_16134,N_13899,N_13859);
xor U16135 (N_16135,N_14314,N_14357);
xnor U16136 (N_16136,N_14835,N_14777);
nor U16137 (N_16137,N_13797,N_14662);
xnor U16138 (N_16138,N_14024,N_14540);
xnor U16139 (N_16139,N_14037,N_14051);
xnor U16140 (N_16140,N_14038,N_14265);
or U16141 (N_16141,N_14561,N_13967);
or U16142 (N_16142,N_14589,N_14021);
or U16143 (N_16143,N_14112,N_14351);
and U16144 (N_16144,N_14277,N_14874);
and U16145 (N_16145,N_14859,N_14257);
xor U16146 (N_16146,N_14193,N_14477);
nand U16147 (N_16147,N_14587,N_13916);
or U16148 (N_16148,N_14981,N_14692);
nand U16149 (N_16149,N_14814,N_14244);
and U16150 (N_16150,N_14281,N_14576);
nand U16151 (N_16151,N_14784,N_14872);
xnor U16152 (N_16152,N_13810,N_14555);
and U16153 (N_16153,N_14967,N_14529);
nand U16154 (N_16154,N_14474,N_14504);
nand U16155 (N_16155,N_13904,N_14795);
nand U16156 (N_16156,N_14126,N_14811);
or U16157 (N_16157,N_14455,N_14623);
nor U16158 (N_16158,N_14274,N_14115);
or U16159 (N_16159,N_14058,N_14734);
nor U16160 (N_16160,N_14835,N_14560);
nand U16161 (N_16161,N_14274,N_14398);
or U16162 (N_16162,N_13845,N_14520);
nor U16163 (N_16163,N_13808,N_14613);
xnor U16164 (N_16164,N_13965,N_13925);
nand U16165 (N_16165,N_13964,N_14450);
xnor U16166 (N_16166,N_14646,N_14986);
nor U16167 (N_16167,N_14816,N_14254);
nor U16168 (N_16168,N_14243,N_14186);
nor U16169 (N_16169,N_14915,N_14064);
nor U16170 (N_16170,N_14610,N_13820);
xor U16171 (N_16171,N_14488,N_14100);
xor U16172 (N_16172,N_14326,N_14591);
nor U16173 (N_16173,N_13974,N_14032);
or U16174 (N_16174,N_14535,N_13966);
nor U16175 (N_16175,N_14067,N_14140);
xnor U16176 (N_16176,N_14756,N_14759);
or U16177 (N_16177,N_13933,N_14974);
nor U16178 (N_16178,N_14733,N_14074);
nor U16179 (N_16179,N_14749,N_14322);
xnor U16180 (N_16180,N_14593,N_14547);
or U16181 (N_16181,N_14628,N_14671);
nor U16182 (N_16182,N_14514,N_14466);
and U16183 (N_16183,N_14162,N_13893);
nor U16184 (N_16184,N_14222,N_14022);
nand U16185 (N_16185,N_14390,N_14817);
or U16186 (N_16186,N_14926,N_14911);
nor U16187 (N_16187,N_13963,N_14809);
nor U16188 (N_16188,N_14743,N_14267);
nand U16189 (N_16189,N_14267,N_13781);
nor U16190 (N_16190,N_14901,N_14117);
or U16191 (N_16191,N_13946,N_14331);
xnor U16192 (N_16192,N_14204,N_13832);
and U16193 (N_16193,N_14328,N_14320);
nor U16194 (N_16194,N_14703,N_14353);
nand U16195 (N_16195,N_14729,N_14289);
xor U16196 (N_16196,N_14473,N_14371);
xnor U16197 (N_16197,N_14339,N_14170);
nor U16198 (N_16198,N_13948,N_14288);
nand U16199 (N_16199,N_14037,N_13893);
or U16200 (N_16200,N_14149,N_14529);
or U16201 (N_16201,N_14494,N_13873);
and U16202 (N_16202,N_14547,N_14971);
nor U16203 (N_16203,N_14483,N_14109);
nor U16204 (N_16204,N_14667,N_14266);
and U16205 (N_16205,N_14153,N_13974);
xor U16206 (N_16206,N_14221,N_14475);
nand U16207 (N_16207,N_13941,N_13961);
or U16208 (N_16208,N_14242,N_13770);
xnor U16209 (N_16209,N_14251,N_14653);
nand U16210 (N_16210,N_14249,N_13804);
xor U16211 (N_16211,N_14591,N_14093);
nand U16212 (N_16212,N_14874,N_14878);
and U16213 (N_16213,N_14294,N_14054);
nor U16214 (N_16214,N_13883,N_14715);
nor U16215 (N_16215,N_14784,N_14375);
or U16216 (N_16216,N_14606,N_14751);
and U16217 (N_16217,N_14745,N_14972);
or U16218 (N_16218,N_14708,N_14523);
nand U16219 (N_16219,N_14306,N_14956);
and U16220 (N_16220,N_13869,N_14757);
nor U16221 (N_16221,N_13899,N_14656);
nand U16222 (N_16222,N_14982,N_14064);
or U16223 (N_16223,N_14057,N_14134);
nor U16224 (N_16224,N_14219,N_14072);
or U16225 (N_16225,N_14057,N_14355);
or U16226 (N_16226,N_14855,N_14774);
xor U16227 (N_16227,N_13934,N_14271);
xnor U16228 (N_16228,N_14665,N_14282);
nor U16229 (N_16229,N_14918,N_13939);
nor U16230 (N_16230,N_14495,N_14786);
nor U16231 (N_16231,N_14597,N_14812);
xnor U16232 (N_16232,N_14108,N_14008);
nor U16233 (N_16233,N_14248,N_13828);
nand U16234 (N_16234,N_14340,N_14091);
and U16235 (N_16235,N_13908,N_14728);
nor U16236 (N_16236,N_14238,N_14015);
nand U16237 (N_16237,N_13796,N_14449);
xor U16238 (N_16238,N_13850,N_14071);
or U16239 (N_16239,N_14264,N_14874);
nor U16240 (N_16240,N_14483,N_14208);
or U16241 (N_16241,N_14756,N_14144);
nor U16242 (N_16242,N_14644,N_14122);
xor U16243 (N_16243,N_14708,N_14184);
nand U16244 (N_16244,N_14427,N_14436);
xor U16245 (N_16245,N_13942,N_14606);
or U16246 (N_16246,N_14973,N_14168);
and U16247 (N_16247,N_14052,N_14499);
nand U16248 (N_16248,N_13978,N_14573);
and U16249 (N_16249,N_13779,N_14866);
nor U16250 (N_16250,N_15236,N_15902);
nand U16251 (N_16251,N_16241,N_15838);
or U16252 (N_16252,N_15230,N_16134);
nor U16253 (N_16253,N_15713,N_16091);
and U16254 (N_16254,N_15849,N_15256);
xor U16255 (N_16255,N_15963,N_15916);
and U16256 (N_16256,N_16023,N_15299);
or U16257 (N_16257,N_15453,N_15495);
nor U16258 (N_16258,N_16239,N_15504);
xor U16259 (N_16259,N_15582,N_15008);
nand U16260 (N_16260,N_15531,N_15327);
and U16261 (N_16261,N_16149,N_15288);
nor U16262 (N_16262,N_15900,N_15124);
nor U16263 (N_16263,N_15325,N_15659);
or U16264 (N_16264,N_15723,N_15592);
xor U16265 (N_16265,N_15978,N_15593);
nand U16266 (N_16266,N_15852,N_15743);
and U16267 (N_16267,N_15228,N_15154);
xnor U16268 (N_16268,N_15729,N_15215);
nand U16269 (N_16269,N_15316,N_15808);
nand U16270 (N_16270,N_15158,N_15542);
or U16271 (N_16271,N_15745,N_16081);
nor U16272 (N_16272,N_15436,N_15605);
nand U16273 (N_16273,N_15002,N_15380);
nor U16274 (N_16274,N_15939,N_16128);
and U16275 (N_16275,N_15837,N_15586);
nand U16276 (N_16276,N_15570,N_15575);
nand U16277 (N_16277,N_15132,N_15526);
nor U16278 (N_16278,N_16164,N_16066);
nor U16279 (N_16279,N_15600,N_15049);
nand U16280 (N_16280,N_16244,N_15110);
xor U16281 (N_16281,N_15704,N_15927);
and U16282 (N_16282,N_16133,N_16040);
or U16283 (N_16283,N_15411,N_15553);
xor U16284 (N_16284,N_15076,N_16130);
and U16285 (N_16285,N_15482,N_16015);
and U16286 (N_16286,N_15468,N_15823);
nor U16287 (N_16287,N_16142,N_16162);
nand U16288 (N_16288,N_16000,N_15198);
or U16289 (N_16289,N_16160,N_16191);
nor U16290 (N_16290,N_15375,N_15845);
nor U16291 (N_16291,N_16017,N_15555);
xor U16292 (N_16292,N_15620,N_15752);
or U16293 (N_16293,N_15131,N_16152);
nand U16294 (N_16294,N_15298,N_16069);
or U16295 (N_16295,N_15185,N_15194);
nand U16296 (N_16296,N_15192,N_15233);
xor U16297 (N_16297,N_15767,N_15707);
or U16298 (N_16298,N_15874,N_15948);
or U16299 (N_16299,N_15412,N_15933);
or U16300 (N_16300,N_15832,N_15165);
nand U16301 (N_16301,N_15969,N_15274);
xor U16302 (N_16302,N_15027,N_16112);
nor U16303 (N_16303,N_15547,N_15287);
xor U16304 (N_16304,N_15277,N_15981);
or U16305 (N_16305,N_15078,N_15416);
or U16306 (N_16306,N_16094,N_15003);
xor U16307 (N_16307,N_15691,N_15182);
xnor U16308 (N_16308,N_15720,N_16020);
nor U16309 (N_16309,N_15738,N_15793);
or U16310 (N_16310,N_15394,N_15730);
nor U16311 (N_16311,N_15063,N_16217);
nand U16312 (N_16312,N_15992,N_15237);
or U16313 (N_16313,N_16246,N_15397);
or U16314 (N_16314,N_15535,N_15769);
and U16315 (N_16315,N_16001,N_15544);
xor U16316 (N_16316,N_15284,N_15410);
nor U16317 (N_16317,N_15034,N_16031);
and U16318 (N_16318,N_15486,N_15273);
xor U16319 (N_16319,N_15694,N_16054);
nand U16320 (N_16320,N_15561,N_15322);
nor U16321 (N_16321,N_16087,N_16170);
xor U16322 (N_16322,N_15150,N_15117);
nand U16323 (N_16323,N_15096,N_16126);
nor U16324 (N_16324,N_16182,N_16041);
nand U16325 (N_16325,N_15636,N_15760);
and U16326 (N_16326,N_15655,N_16093);
xnor U16327 (N_16327,N_16095,N_15431);
nand U16328 (N_16328,N_15229,N_16119);
xnor U16329 (N_16329,N_16228,N_15688);
nor U16330 (N_16330,N_15021,N_16127);
xnor U16331 (N_16331,N_15490,N_16120);
nor U16332 (N_16332,N_16079,N_15731);
nor U16333 (N_16333,N_16238,N_15275);
and U16334 (N_16334,N_15855,N_15227);
nand U16335 (N_16335,N_16064,N_15827);
or U16336 (N_16336,N_15303,N_16099);
and U16337 (N_16337,N_15762,N_15664);
or U16338 (N_16338,N_15595,N_16083);
or U16339 (N_16339,N_15304,N_15011);
nand U16340 (N_16340,N_15755,N_15498);
nand U16341 (N_16341,N_15653,N_15448);
nor U16342 (N_16342,N_16161,N_15678);
and U16343 (N_16343,N_15450,N_16145);
and U16344 (N_16344,N_16086,N_16240);
xor U16345 (N_16345,N_16200,N_15365);
and U16346 (N_16346,N_15732,N_16005);
or U16347 (N_16347,N_15953,N_15496);
and U16348 (N_16348,N_15965,N_15754);
nand U16349 (N_16349,N_15220,N_15751);
nor U16350 (N_16350,N_15590,N_15577);
xor U16351 (N_16351,N_15534,N_16062);
xnor U16352 (N_16352,N_15884,N_15536);
or U16353 (N_16353,N_15623,N_15982);
xor U16354 (N_16354,N_15455,N_15168);
and U16355 (N_16355,N_15301,N_15446);
nor U16356 (N_16356,N_15515,N_15193);
nand U16357 (N_16357,N_15361,N_15028);
xnor U16358 (N_16358,N_15666,N_16051);
xnor U16359 (N_16359,N_15148,N_16059);
and U16360 (N_16360,N_15947,N_16058);
xor U16361 (N_16361,N_15356,N_15216);
xnor U16362 (N_16362,N_15033,N_16024);
nor U16363 (N_16363,N_16010,N_16021);
and U16364 (N_16364,N_15006,N_15626);
nand U16365 (N_16365,N_15911,N_16146);
and U16366 (N_16366,N_15803,N_15784);
and U16367 (N_16367,N_15173,N_15646);
and U16368 (N_16368,N_15153,N_15259);
or U16369 (N_16369,N_15378,N_15061);
or U16370 (N_16370,N_15675,N_15300);
xor U16371 (N_16371,N_15766,N_15867);
nor U16372 (N_16372,N_15342,N_15866);
nor U16373 (N_16373,N_15499,N_15449);
or U16374 (N_16374,N_15782,N_15833);
or U16375 (N_16375,N_15726,N_15239);
or U16376 (N_16376,N_15095,N_15106);
nand U16377 (N_16377,N_15128,N_15210);
or U16378 (N_16378,N_15476,N_16063);
or U16379 (N_16379,N_15311,N_15541);
or U16380 (N_16380,N_15562,N_15140);
and U16381 (N_16381,N_16018,N_15090);
xor U16382 (N_16382,N_16205,N_15462);
and U16383 (N_16383,N_16019,N_16122);
nand U16384 (N_16384,N_15587,N_15251);
nor U16385 (N_16385,N_15960,N_15657);
or U16386 (N_16386,N_15088,N_15171);
xnor U16387 (N_16387,N_15614,N_15891);
and U16388 (N_16388,N_15355,N_15286);
nor U16389 (N_16389,N_15031,N_15332);
xnor U16390 (N_16390,N_15360,N_15494);
nand U16391 (N_16391,N_15492,N_15077);
xnor U16392 (N_16392,N_15177,N_15628);
nand U16393 (N_16393,N_15873,N_15371);
nand U16394 (N_16394,N_16074,N_15668);
or U16395 (N_16395,N_15379,N_15799);
or U16396 (N_16396,N_15501,N_15157);
and U16397 (N_16397,N_15041,N_15898);
and U16398 (N_16398,N_15139,N_15324);
nand U16399 (N_16399,N_15750,N_16103);
or U16400 (N_16400,N_15059,N_15554);
or U16401 (N_16401,N_16147,N_15924);
or U16402 (N_16402,N_15260,N_15125);
nand U16403 (N_16403,N_15114,N_16107);
or U16404 (N_16404,N_15334,N_15761);
nand U16405 (N_16405,N_15596,N_15432);
nor U16406 (N_16406,N_15143,N_15529);
or U16407 (N_16407,N_15406,N_15697);
nor U16408 (N_16408,N_15434,N_15004);
nand U16409 (N_16409,N_15999,N_15903);
nor U16410 (N_16410,N_15962,N_16016);
nor U16411 (N_16411,N_15607,N_15368);
nor U16412 (N_16412,N_15568,N_15170);
and U16413 (N_16413,N_15703,N_15997);
and U16414 (N_16414,N_15543,N_16221);
and U16415 (N_16415,N_15976,N_15692);
xnor U16416 (N_16416,N_15441,N_15885);
or U16417 (N_16417,N_15975,N_15527);
nor U16418 (N_16418,N_15429,N_15047);
nor U16419 (N_16419,N_16124,N_15439);
nor U16420 (N_16420,N_15112,N_15700);
nand U16421 (N_16421,N_16176,N_15961);
nand U16422 (N_16422,N_15471,N_15734);
or U16423 (N_16423,N_16140,N_15879);
or U16424 (N_16424,N_15856,N_15159);
and U16425 (N_16425,N_16012,N_15169);
xor U16426 (N_16426,N_15581,N_15461);
nor U16427 (N_16427,N_15661,N_15973);
xor U16428 (N_16428,N_16111,N_15865);
or U16429 (N_16429,N_15705,N_15557);
xnor U16430 (N_16430,N_15493,N_15142);
or U16431 (N_16431,N_15801,N_15224);
and U16432 (N_16432,N_16190,N_15306);
nand U16433 (N_16433,N_15000,N_15912);
and U16434 (N_16434,N_15042,N_16209);
nand U16435 (N_16435,N_15127,N_15934);
or U16436 (N_16436,N_15672,N_15176);
and U16437 (N_16437,N_15525,N_15359);
or U16438 (N_16438,N_15860,N_15815);
or U16439 (N_16439,N_15156,N_16245);
and U16440 (N_16440,N_16136,N_15331);
xor U16441 (N_16441,N_15319,N_15155);
nor U16442 (N_16442,N_15389,N_15980);
and U16443 (N_16443,N_15094,N_15473);
nand U16444 (N_16444,N_16036,N_16150);
nand U16445 (N_16445,N_15971,N_15853);
xnor U16446 (N_16446,N_15777,N_15813);
xor U16447 (N_16447,N_15100,N_15072);
xor U16448 (N_16448,N_15348,N_15179);
or U16449 (N_16449,N_15715,N_16044);
xor U16450 (N_16450,N_16218,N_15460);
nand U16451 (N_16451,N_15388,N_15787);
and U16452 (N_16452,N_15591,N_15321);
nand U16453 (N_16453,N_15172,N_16236);
nor U16454 (N_16454,N_15249,N_16177);
or U16455 (N_16455,N_15017,N_16039);
nand U16456 (N_16456,N_15282,N_15790);
xor U16457 (N_16457,N_15305,N_15187);
or U16458 (N_16458,N_15479,N_15617);
and U16459 (N_16459,N_15346,N_15573);
and U16460 (N_16460,N_15403,N_15611);
nor U16461 (N_16461,N_15421,N_15597);
nor U16462 (N_16462,N_15888,N_16233);
and U16463 (N_16463,N_15794,N_16193);
or U16464 (N_16464,N_16199,N_15753);
nor U16465 (N_16465,N_15503,N_15015);
nand U16466 (N_16466,N_15645,N_15010);
nand U16467 (N_16467,N_15444,N_15551);
or U16468 (N_16468,N_15629,N_15818);
nor U16469 (N_16469,N_16060,N_15550);
nand U16470 (N_16470,N_15013,N_16214);
nand U16471 (N_16471,N_15181,N_15069);
xnor U16472 (N_16472,N_15682,N_15056);
nand U16473 (N_16473,N_15101,N_15291);
and U16474 (N_16474,N_16050,N_15484);
nand U16475 (N_16475,N_15510,N_15763);
or U16476 (N_16476,N_16156,N_15895);
nand U16477 (N_16477,N_15477,N_15684);
nand U16478 (N_16478,N_16135,N_15062);
and U16479 (N_16479,N_15968,N_15716);
or U16480 (N_16480,N_15549,N_15950);
xnor U16481 (N_16481,N_15598,N_16154);
nor U16482 (N_16482,N_15910,N_15285);
nor U16483 (N_16483,N_16030,N_15202);
or U16484 (N_16484,N_15307,N_16148);
nand U16485 (N_16485,N_15647,N_15018);
and U16486 (N_16486,N_15424,N_15580);
nand U16487 (N_16487,N_15086,N_15023);
and U16488 (N_16488,N_15612,N_15201);
nor U16489 (N_16489,N_15774,N_15907);
nor U16490 (N_16490,N_15454,N_16027);
nor U16491 (N_16491,N_15826,N_15556);
and U16492 (N_16492,N_15560,N_15464);
or U16493 (N_16493,N_15292,N_15383);
xor U16494 (N_16494,N_16139,N_15757);
xnor U16495 (N_16495,N_15613,N_16115);
and U16496 (N_16496,N_15835,N_15868);
nand U16497 (N_16497,N_16098,N_15650);
xor U16498 (N_16498,N_15245,N_15806);
xor U16499 (N_16499,N_15875,N_15632);
and U16500 (N_16500,N_16029,N_15886);
xor U16501 (N_16501,N_15708,N_15058);
or U16502 (N_16502,N_15399,N_15578);
or U16503 (N_16503,N_15807,N_15830);
xnor U16504 (N_16504,N_15308,N_15872);
nand U16505 (N_16505,N_16195,N_15392);
and U16506 (N_16506,N_15213,N_15052);
and U16507 (N_16507,N_15706,N_15522);
xnor U16508 (N_16508,N_15564,N_15931);
xor U16509 (N_16509,N_15641,N_16125);
xnor U16510 (N_16510,N_15518,N_15656);
nand U16511 (N_16511,N_16025,N_15152);
nand U16512 (N_16512,N_16121,N_15337);
nor U16513 (N_16513,N_15548,N_15180);
and U16514 (N_16514,N_15068,N_15539);
xnor U16515 (N_16515,N_15054,N_16151);
xor U16516 (N_16516,N_16057,N_15797);
xor U16517 (N_16517,N_15111,N_15070);
and U16518 (N_16518,N_15205,N_16065);
xnor U16519 (N_16519,N_15988,N_15333);
nor U16520 (N_16520,N_15218,N_15524);
or U16521 (N_16521,N_15407,N_16208);
nor U16522 (N_16522,N_15133,N_16243);
nor U16523 (N_16523,N_15167,N_15391);
or U16524 (N_16524,N_15297,N_15440);
or U16525 (N_16525,N_15087,N_15798);
and U16526 (N_16526,N_16206,N_15478);
nor U16527 (N_16527,N_15913,N_15974);
nand U16528 (N_16528,N_15084,N_15926);
xor U16529 (N_16529,N_15350,N_15858);
and U16530 (N_16530,N_15340,N_15906);
nand U16531 (N_16531,N_16110,N_16034);
and U16532 (N_16532,N_15147,N_15433);
nand U16533 (N_16533,N_15733,N_15505);
nand U16534 (N_16534,N_15384,N_15386);
nor U16535 (N_16535,N_15579,N_15212);
or U16536 (N_16536,N_15022,N_15057);
xnor U16537 (N_16537,N_15458,N_15426);
xor U16538 (N_16538,N_16224,N_16222);
xnor U16539 (N_16539,N_15417,N_15373);
xor U16540 (N_16540,N_15475,N_15343);
and U16541 (N_16541,N_15309,N_15690);
xnor U16542 (N_16542,N_15622,N_15569);
or U16543 (N_16543,N_16068,N_15243);
nor U16544 (N_16544,N_15938,N_15451);
or U16545 (N_16545,N_16075,N_16032);
xor U16546 (N_16546,N_16009,N_15442);
nor U16547 (N_16547,N_15747,N_15588);
nand U16548 (N_16548,N_16226,N_15558);
nand U16549 (N_16549,N_15235,N_15639);
nor U16550 (N_16550,N_15401,N_15074);
xor U16551 (N_16551,N_15918,N_15480);
or U16552 (N_16552,N_15120,N_15402);
nand U16553 (N_16553,N_15899,N_15877);
or U16554 (N_16554,N_15178,N_15130);
xor U16555 (N_16555,N_15257,N_15897);
nor U16556 (N_16556,N_15651,N_15776);
nand U16557 (N_16557,N_15942,N_16229);
nor U16558 (N_16558,N_16207,N_16102);
and U16559 (N_16559,N_15116,N_15466);
nand U16560 (N_16560,N_15315,N_15634);
or U16561 (N_16561,N_16104,N_16237);
and U16562 (N_16562,N_16197,N_15294);
or U16563 (N_16563,N_15633,N_15817);
or U16564 (N_16564,N_16159,N_15265);
nand U16565 (N_16565,N_15370,N_15618);
xnor U16566 (N_16566,N_16178,N_15785);
nor U16567 (N_16567,N_15323,N_15644);
or U16568 (N_16568,N_16223,N_16037);
or U16569 (N_16569,N_15876,N_15437);
and U16570 (N_16570,N_15687,N_15184);
nand U16571 (N_16571,N_16076,N_15909);
xor U16572 (N_16572,N_16056,N_15452);
nor U16573 (N_16573,N_15080,N_15354);
and U16574 (N_16574,N_15940,N_16163);
nor U16575 (N_16575,N_15583,N_15843);
nand U16576 (N_16576,N_15396,N_15242);
xor U16577 (N_16577,N_15630,N_15850);
nor U16578 (N_16578,N_15363,N_16166);
or U16579 (N_16579,N_15024,N_15834);
xor U16580 (N_16580,N_16234,N_16210);
xnor U16581 (N_16581,N_15338,N_15721);
and U16582 (N_16582,N_15864,N_16042);
xnor U16583 (N_16583,N_15983,N_15418);
or U16584 (N_16584,N_16138,N_16108);
xnor U16585 (N_16585,N_15930,N_16035);
nor U16586 (N_16586,N_16049,N_15532);
nand U16587 (N_16587,N_15722,N_15296);
nor U16588 (N_16588,N_15162,N_15400);
xor U16589 (N_16589,N_15984,N_15221);
nor U16590 (N_16590,N_15563,N_15079);
xor U16591 (N_16591,N_15064,N_16132);
nor U16592 (N_16592,N_15161,N_16196);
or U16593 (N_16593,N_15105,N_15811);
nor U16594 (N_16594,N_15805,N_15883);
xor U16595 (N_16595,N_15280,N_15067);
nor U16596 (N_16596,N_15122,N_15698);
nand U16597 (N_16597,N_15851,N_15398);
nand U16598 (N_16598,N_15163,N_15796);
or U16599 (N_16599,N_15538,N_15483);
nor U16600 (N_16600,N_15472,N_15053);
or U16601 (N_16601,N_15863,N_15414);
xnor U16602 (N_16602,N_15904,N_15673);
or U16603 (N_16603,N_15804,N_15572);
and U16604 (N_16604,N_15206,N_15344);
and U16605 (N_16605,N_15737,N_15358);
nand U16606 (N_16606,N_15367,N_15075);
or U16607 (N_16607,N_15748,N_15624);
nor U16608 (N_16608,N_15328,N_15736);
xnor U16609 (N_16609,N_15727,N_15270);
and U16610 (N_16610,N_15941,N_15928);
nor U16611 (N_16611,N_15685,N_16113);
or U16612 (N_16612,N_16022,N_15840);
nor U16613 (N_16613,N_16184,N_15993);
xnor U16614 (N_16614,N_16203,N_15151);
nor U16615 (N_16615,N_15290,N_15862);
nand U16616 (N_16616,N_15841,N_15276);
and U16617 (N_16617,N_15469,N_16003);
nand U16618 (N_16618,N_15648,N_15638);
or U16619 (N_16619,N_16109,N_15995);
and U16620 (N_16620,N_15998,N_15640);
xnor U16621 (N_16621,N_15741,N_15728);
nand U16622 (N_16622,N_15362,N_16072);
and U16623 (N_16623,N_15289,N_15520);
nor U16624 (N_16624,N_15642,N_15264);
and U16625 (N_16625,N_15196,N_15966);
nor U16626 (N_16626,N_15822,N_15295);
and U16627 (N_16627,N_15739,N_16077);
or U16628 (N_16628,N_15791,N_16189);
and U16629 (N_16629,N_15020,N_15474);
nor U16630 (N_16630,N_16230,N_15467);
nand U16631 (N_16631,N_15514,N_15093);
nand U16632 (N_16632,N_15889,N_16084);
nor U16633 (N_16633,N_15714,N_15374);
or U16634 (N_16634,N_15652,N_15339);
nand U16635 (N_16635,N_16198,N_15552);
nand U16636 (N_16636,N_16061,N_15559);
nand U16637 (N_16637,N_16201,N_16212);
or U16638 (N_16638,N_15517,N_16179);
nand U16639 (N_16639,N_15395,N_15263);
xor U16640 (N_16640,N_15134,N_16007);
or U16641 (N_16641,N_15066,N_15244);
and U16642 (N_16642,N_16047,N_15985);
nor U16643 (N_16643,N_16100,N_16004);
nor U16644 (N_16644,N_16137,N_15415);
xnor U16645 (N_16645,N_15326,N_15943);
nor U16646 (N_16646,N_15330,N_15589);
nand U16647 (N_16647,N_16174,N_15857);
nor U16648 (N_16648,N_15922,N_15413);
xnor U16649 (N_16649,N_15487,N_15035);
nor U16650 (N_16650,N_16080,N_15232);
xor U16651 (N_16651,N_16073,N_15954);
or U16652 (N_16652,N_15248,N_16192);
or U16653 (N_16653,N_15677,N_15566);
or U16654 (N_16654,N_16131,N_15001);
and U16655 (N_16655,N_15238,N_15341);
nor U16656 (N_16656,N_15681,N_15625);
or U16657 (N_16657,N_16101,N_15491);
nand U16658 (N_16658,N_15621,N_15204);
nor U16659 (N_16659,N_15765,N_15457);
nor U16660 (N_16660,N_15771,N_15081);
xnor U16661 (N_16661,N_16204,N_15660);
and U16662 (N_16662,N_15183,N_15091);
nor U16663 (N_16663,N_15585,N_16185);
and U16664 (N_16664,N_15252,N_15914);
and U16665 (N_16665,N_15082,N_15576);
nand U16666 (N_16666,N_15956,N_15919);
nand U16667 (N_16667,N_15099,N_15654);
xnor U16668 (N_16668,N_15209,N_15702);
and U16669 (N_16669,N_15829,N_15369);
or U16670 (N_16670,N_15423,N_16143);
and U16671 (N_16671,N_15606,N_15207);
nor U16672 (N_16672,N_15281,N_15701);
xor U16673 (N_16673,N_15250,N_15045);
nand U16674 (N_16674,N_15693,N_15387);
or U16675 (N_16675,N_15537,N_15390);
nor U16676 (N_16676,N_15565,N_15459);
nor U16677 (N_16677,N_15773,N_16046);
or U16678 (N_16678,N_15637,N_15443);
or U16679 (N_16679,N_15724,N_15896);
nand U16680 (N_16680,N_15108,N_15967);
nor U16681 (N_16681,N_15508,N_15445);
or U16682 (N_16682,N_15226,N_15456);
xor U16683 (N_16683,N_15347,N_15335);
and U16684 (N_16684,N_15219,N_15255);
and U16685 (N_16685,N_15481,N_16096);
xnor U16686 (N_16686,N_15955,N_15658);
nor U16687 (N_16687,N_15073,N_16171);
nor U16688 (N_16688,N_15842,N_16242);
and U16689 (N_16689,N_16067,N_16188);
nand U16690 (N_16690,N_16053,N_15037);
nor U16691 (N_16691,N_15601,N_15254);
xnor U16692 (N_16692,N_15783,N_15279);
nor U16693 (N_16693,N_15145,N_15113);
xor U16694 (N_16694,N_16011,N_15144);
xor U16695 (N_16695,N_15816,N_15521);
nor U16696 (N_16696,N_16078,N_15861);
nand U16697 (N_16697,N_15602,N_16129);
xor U16698 (N_16698,N_15293,N_15759);
or U16699 (N_16699,N_16173,N_15241);
or U16700 (N_16700,N_15749,N_16168);
nor U16701 (N_16701,N_15772,N_15908);
or U16702 (N_16702,N_15507,N_15329);
and U16703 (N_16703,N_15836,N_15894);
and U16704 (N_16704,N_15141,N_15744);
xor U16705 (N_16705,N_15302,N_15717);
xor U16706 (N_16706,N_16092,N_15372);
xnor U16707 (N_16707,N_16155,N_15946);
nand U16708 (N_16708,N_15085,N_15200);
nand U16709 (N_16709,N_16167,N_15905);
and U16710 (N_16710,N_15065,N_15349);
or U16711 (N_16711,N_15878,N_15419);
nor U16712 (N_16712,N_15103,N_15115);
or U16713 (N_16713,N_15994,N_15137);
nor U16714 (N_16714,N_15121,N_15318);
nand U16715 (N_16715,N_16219,N_15032);
or U16716 (N_16716,N_15214,N_16117);
and U16717 (N_16717,N_15599,N_15970);
or U16718 (N_16718,N_16248,N_15846);
nor U16719 (N_16719,N_15788,N_15936);
or U16720 (N_16720,N_15014,N_15663);
and U16721 (N_16721,N_16158,N_16123);
xnor U16722 (N_16722,N_15509,N_15317);
nor U16723 (N_16723,N_15262,N_15314);
nor U16724 (N_16724,N_15977,N_16028);
xor U16725 (N_16725,N_15050,N_15921);
and U16726 (N_16726,N_16070,N_16114);
or U16727 (N_16727,N_15854,N_15408);
or U16728 (N_16728,N_15048,N_15915);
and U16729 (N_16729,N_16225,N_16105);
nor U16730 (N_16730,N_15175,N_16175);
nor U16731 (N_16731,N_15533,N_15880);
xnor U16732 (N_16732,N_16085,N_16216);
nor U16733 (N_16733,N_15005,N_16183);
nand U16734 (N_16734,N_15951,N_15792);
or U16735 (N_16735,N_16220,N_15670);
and U16736 (N_16736,N_15166,N_15820);
and U16737 (N_16737,N_15019,N_15420);
or U16738 (N_16738,N_15695,N_15012);
nand U16739 (N_16739,N_15381,N_15944);
or U16740 (N_16740,N_15699,N_15545);
xnor U16741 (N_16741,N_15800,N_15310);
nand U16742 (N_16742,N_15118,N_15674);
nor U16743 (N_16743,N_15887,N_15038);
and U16744 (N_16744,N_15186,N_15513);
or U16745 (N_16745,N_15470,N_15871);
or U16746 (N_16746,N_15528,N_15136);
or U16747 (N_16747,N_15126,N_15267);
or U16748 (N_16748,N_15044,N_15683);
xor U16749 (N_16749,N_16181,N_16211);
xor U16750 (N_16750,N_15199,N_15071);
and U16751 (N_16751,N_15631,N_15404);
and U16752 (N_16752,N_15571,N_15710);
xor U16753 (N_16753,N_15635,N_15725);
nor U16754 (N_16754,N_15506,N_15385);
and U16755 (N_16755,N_15990,N_15923);
and U16756 (N_16756,N_15979,N_16215);
and U16757 (N_16757,N_15352,N_15901);
nor U16758 (N_16758,N_16141,N_15203);
nand U16759 (N_16759,N_16213,N_16165);
xnor U16760 (N_16760,N_15283,N_15812);
xnor U16761 (N_16761,N_15123,N_15786);
nor U16762 (N_16762,N_15246,N_15223);
and U16763 (N_16763,N_16045,N_15511);
nand U16764 (N_16764,N_15320,N_15669);
nor U16765 (N_16765,N_16097,N_15119);
or U16766 (N_16766,N_15364,N_16227);
and U16767 (N_16767,N_15366,N_16082);
or U16768 (N_16768,N_15208,N_15351);
xnor U16769 (N_16769,N_15831,N_15463);
and U16770 (N_16770,N_15135,N_16247);
or U16771 (N_16771,N_15949,N_15425);
xor U16772 (N_16772,N_15098,N_15430);
or U16773 (N_16773,N_15809,N_15146);
and U16774 (N_16774,N_15217,N_15719);
nor U16775 (N_16775,N_15574,N_15882);
or U16776 (N_16776,N_15848,N_16180);
and U16777 (N_16777,N_16144,N_15272);
or U16778 (N_16778,N_15996,N_16071);
nor U16779 (N_16779,N_16008,N_15546);
and U16780 (N_16780,N_15735,N_15195);
or U16781 (N_16781,N_15060,N_15540);
nand U16782 (N_16782,N_15485,N_15775);
nor U16783 (N_16783,N_15662,N_15844);
nand U16784 (N_16784,N_15802,N_15502);
xor U16785 (N_16785,N_15746,N_16090);
and U16786 (N_16786,N_15129,N_16038);
nand U16787 (N_16787,N_15989,N_15040);
and U16788 (N_16788,N_15488,N_15190);
nand U16789 (N_16789,N_15007,N_15438);
xor U16790 (N_16790,N_15952,N_15089);
or U16791 (N_16791,N_15376,N_16187);
nand U16792 (N_16792,N_16118,N_15959);
or U16793 (N_16793,N_15758,N_15377);
nor U16794 (N_16794,N_16231,N_15211);
and U16795 (N_16795,N_15353,N_15711);
nand U16796 (N_16796,N_15819,N_15269);
and U16797 (N_16797,N_15188,N_15109);
xnor U16798 (N_16798,N_15197,N_15957);
nor U16799 (N_16799,N_15357,N_15519);
nand U16800 (N_16800,N_15869,N_15742);
and U16801 (N_16801,N_15920,N_15925);
and U16802 (N_16802,N_15770,N_16006);
nor U16803 (N_16803,N_15051,N_15881);
or U16804 (N_16804,N_15604,N_15810);
nand U16805 (N_16805,N_15917,N_15972);
or U16806 (N_16806,N_15680,N_15405);
xnor U16807 (N_16807,N_15261,N_16157);
nand U16808 (N_16808,N_15258,N_15029);
and U16809 (N_16809,N_15097,N_15313);
and U16810 (N_16810,N_15253,N_15083);
and U16811 (N_16811,N_16026,N_16089);
and U16812 (N_16812,N_15649,N_15046);
xor U16813 (N_16813,N_16169,N_16153);
and U16814 (N_16814,N_16232,N_16055);
or U16815 (N_16815,N_15500,N_16014);
nor U16816 (N_16816,N_15039,N_15932);
nand U16817 (N_16817,N_15712,N_15986);
and U16818 (N_16818,N_15686,N_15189);
or U16819 (N_16819,N_16116,N_15643);
or U16820 (N_16820,N_15234,N_15676);
and U16821 (N_16821,N_15336,N_15225);
or U16822 (N_16822,N_15756,N_15779);
nand U16823 (N_16823,N_15497,N_15382);
xnor U16824 (N_16824,N_16013,N_15240);
and U16825 (N_16825,N_15107,N_15102);
and U16826 (N_16826,N_15615,N_15679);
nor U16827 (N_16827,N_15393,N_15278);
xnor U16828 (N_16828,N_15104,N_15271);
or U16829 (N_16829,N_15824,N_15043);
nor U16830 (N_16830,N_16033,N_15821);
nand U16831 (N_16831,N_15016,N_15780);
or U16832 (N_16832,N_15627,N_16186);
and U16833 (N_16833,N_15764,N_15523);
xnor U16834 (N_16834,N_15958,N_15665);
nor U16835 (N_16835,N_15345,N_15191);
xnor U16836 (N_16836,N_15567,N_15929);
and U16837 (N_16837,N_15594,N_15026);
and U16838 (N_16838,N_16235,N_15828);
or U16839 (N_16839,N_15991,N_15839);
or U16840 (N_16840,N_15164,N_15937);
and U16841 (N_16841,N_15781,N_15709);
and U16842 (N_16842,N_15036,N_15778);
xor U16843 (N_16843,N_15671,N_15610);
or U16844 (N_16844,N_15247,N_15892);
or U16845 (N_16845,N_15435,N_15667);
or U16846 (N_16846,N_15222,N_15814);
xor U16847 (N_16847,N_15055,N_15847);
nor U16848 (N_16848,N_15266,N_15689);
or U16849 (N_16849,N_15530,N_16043);
nor U16850 (N_16850,N_15768,N_15945);
nor U16851 (N_16851,N_15025,N_16172);
nor U16852 (N_16852,N_16194,N_16202);
nand U16853 (N_16853,N_15789,N_15512);
nand U16854 (N_16854,N_15312,N_15935);
nand U16855 (N_16855,N_15696,N_15149);
nor U16856 (N_16856,N_16088,N_15030);
nand U16857 (N_16857,N_15870,N_15859);
and U16858 (N_16858,N_15174,N_15465);
and U16859 (N_16859,N_15516,N_16106);
nand U16860 (N_16860,N_15795,N_16002);
and U16861 (N_16861,N_15489,N_15160);
or U16862 (N_16862,N_15609,N_15893);
nand U16863 (N_16863,N_15422,N_15616);
or U16864 (N_16864,N_15009,N_15138);
nor U16865 (N_16865,N_15584,N_15603);
or U16866 (N_16866,N_15427,N_16052);
or U16867 (N_16867,N_15825,N_15409);
and U16868 (N_16868,N_15987,N_15608);
xor U16869 (N_16869,N_15428,N_15718);
nor U16870 (N_16870,N_15092,N_15619);
xor U16871 (N_16871,N_15740,N_15268);
and U16872 (N_16872,N_15447,N_15231);
xnor U16873 (N_16873,N_16048,N_15890);
and U16874 (N_16874,N_16249,N_15964);
and U16875 (N_16875,N_15359,N_15252);
or U16876 (N_16876,N_15440,N_16042);
or U16877 (N_16877,N_16066,N_16105);
xor U16878 (N_16878,N_15099,N_15538);
and U16879 (N_16879,N_15393,N_15591);
nand U16880 (N_16880,N_15592,N_15330);
nor U16881 (N_16881,N_15760,N_16019);
nor U16882 (N_16882,N_15878,N_16138);
nor U16883 (N_16883,N_16197,N_16154);
and U16884 (N_16884,N_15420,N_15401);
nand U16885 (N_16885,N_15228,N_15203);
nand U16886 (N_16886,N_15176,N_15252);
nor U16887 (N_16887,N_15138,N_16040);
and U16888 (N_16888,N_16032,N_15147);
xor U16889 (N_16889,N_15230,N_16156);
and U16890 (N_16890,N_15303,N_15123);
xnor U16891 (N_16891,N_15720,N_15015);
and U16892 (N_16892,N_15135,N_15401);
nor U16893 (N_16893,N_15345,N_15538);
xnor U16894 (N_16894,N_15436,N_15991);
xor U16895 (N_16895,N_15083,N_15017);
or U16896 (N_16896,N_15042,N_15907);
nor U16897 (N_16897,N_15978,N_15187);
or U16898 (N_16898,N_16228,N_15906);
xnor U16899 (N_16899,N_15630,N_16027);
nand U16900 (N_16900,N_16136,N_15833);
or U16901 (N_16901,N_15670,N_15497);
and U16902 (N_16902,N_15090,N_16114);
or U16903 (N_16903,N_15181,N_15095);
nor U16904 (N_16904,N_15302,N_15981);
nor U16905 (N_16905,N_16168,N_15612);
nand U16906 (N_16906,N_15415,N_16085);
and U16907 (N_16907,N_15955,N_15729);
or U16908 (N_16908,N_15287,N_15352);
or U16909 (N_16909,N_15519,N_16022);
nor U16910 (N_16910,N_16199,N_15579);
or U16911 (N_16911,N_15931,N_15683);
xor U16912 (N_16912,N_15923,N_16114);
and U16913 (N_16913,N_15684,N_15180);
nand U16914 (N_16914,N_15367,N_15445);
xor U16915 (N_16915,N_16077,N_15828);
nand U16916 (N_16916,N_16007,N_15380);
and U16917 (N_16917,N_15014,N_16086);
and U16918 (N_16918,N_15078,N_16025);
xor U16919 (N_16919,N_16197,N_15648);
or U16920 (N_16920,N_15174,N_15991);
nor U16921 (N_16921,N_15062,N_15625);
nor U16922 (N_16922,N_15934,N_16040);
nand U16923 (N_16923,N_15763,N_15917);
or U16924 (N_16924,N_16192,N_15829);
or U16925 (N_16925,N_15097,N_15471);
or U16926 (N_16926,N_15804,N_16112);
xor U16927 (N_16927,N_15785,N_15666);
and U16928 (N_16928,N_16127,N_15813);
or U16929 (N_16929,N_15546,N_15825);
nand U16930 (N_16930,N_15301,N_16195);
or U16931 (N_16931,N_16242,N_16004);
and U16932 (N_16932,N_15056,N_16220);
xor U16933 (N_16933,N_15765,N_16119);
xor U16934 (N_16934,N_15992,N_15436);
nand U16935 (N_16935,N_15941,N_15521);
and U16936 (N_16936,N_16060,N_15876);
nand U16937 (N_16937,N_15760,N_15620);
nor U16938 (N_16938,N_15337,N_16070);
xnor U16939 (N_16939,N_15618,N_15960);
nand U16940 (N_16940,N_15402,N_15622);
and U16941 (N_16941,N_15483,N_16232);
and U16942 (N_16942,N_15548,N_15257);
or U16943 (N_16943,N_15283,N_15469);
and U16944 (N_16944,N_15951,N_15973);
and U16945 (N_16945,N_15255,N_15888);
or U16946 (N_16946,N_16042,N_15730);
xor U16947 (N_16947,N_15903,N_15248);
nor U16948 (N_16948,N_15708,N_15889);
nand U16949 (N_16949,N_15498,N_16222);
or U16950 (N_16950,N_15265,N_15922);
nor U16951 (N_16951,N_15865,N_15278);
nor U16952 (N_16952,N_16079,N_16147);
or U16953 (N_16953,N_16152,N_15282);
nor U16954 (N_16954,N_15762,N_15257);
xnor U16955 (N_16955,N_15651,N_15214);
and U16956 (N_16956,N_15067,N_15852);
nor U16957 (N_16957,N_16102,N_15438);
xor U16958 (N_16958,N_15776,N_16194);
xor U16959 (N_16959,N_15868,N_15852);
or U16960 (N_16960,N_15870,N_15516);
and U16961 (N_16961,N_15867,N_16145);
or U16962 (N_16962,N_15440,N_15656);
nor U16963 (N_16963,N_15554,N_15547);
and U16964 (N_16964,N_15472,N_15753);
nor U16965 (N_16965,N_16196,N_15000);
or U16966 (N_16966,N_16036,N_15360);
nand U16967 (N_16967,N_15991,N_15498);
or U16968 (N_16968,N_15449,N_15382);
nand U16969 (N_16969,N_16117,N_15712);
xor U16970 (N_16970,N_15098,N_15359);
or U16971 (N_16971,N_16044,N_15465);
nand U16972 (N_16972,N_15454,N_15601);
and U16973 (N_16973,N_15480,N_15976);
xnor U16974 (N_16974,N_16110,N_15862);
xnor U16975 (N_16975,N_15730,N_15528);
and U16976 (N_16976,N_15154,N_15477);
or U16977 (N_16977,N_16178,N_15526);
and U16978 (N_16978,N_16018,N_15086);
xor U16979 (N_16979,N_16015,N_15214);
nand U16980 (N_16980,N_15952,N_15062);
xnor U16981 (N_16981,N_16045,N_16040);
nand U16982 (N_16982,N_15482,N_15997);
xor U16983 (N_16983,N_15124,N_15938);
nand U16984 (N_16984,N_16088,N_15731);
and U16985 (N_16985,N_15332,N_15539);
xor U16986 (N_16986,N_15069,N_16067);
xor U16987 (N_16987,N_15105,N_15795);
nor U16988 (N_16988,N_16116,N_16105);
xor U16989 (N_16989,N_15783,N_15701);
nor U16990 (N_16990,N_15803,N_15429);
nand U16991 (N_16991,N_15344,N_16119);
or U16992 (N_16992,N_15016,N_16166);
nor U16993 (N_16993,N_16152,N_15821);
nor U16994 (N_16994,N_15969,N_15720);
nand U16995 (N_16995,N_15641,N_15870);
nor U16996 (N_16996,N_15563,N_15223);
nor U16997 (N_16997,N_16036,N_15753);
and U16998 (N_16998,N_16011,N_15054);
nand U16999 (N_16999,N_15215,N_15444);
xor U17000 (N_17000,N_15582,N_15740);
xor U17001 (N_17001,N_15440,N_15356);
nor U17002 (N_17002,N_16121,N_16230);
nand U17003 (N_17003,N_15470,N_15045);
nand U17004 (N_17004,N_16094,N_15672);
xor U17005 (N_17005,N_16077,N_15348);
or U17006 (N_17006,N_15288,N_15379);
and U17007 (N_17007,N_15887,N_15128);
or U17008 (N_17008,N_16229,N_15753);
nand U17009 (N_17009,N_15547,N_15637);
and U17010 (N_17010,N_16235,N_15359);
or U17011 (N_17011,N_16227,N_15068);
and U17012 (N_17012,N_15931,N_15979);
nand U17013 (N_17013,N_15388,N_15663);
nand U17014 (N_17014,N_15884,N_15679);
and U17015 (N_17015,N_15385,N_15374);
xor U17016 (N_17016,N_16245,N_15117);
xor U17017 (N_17017,N_15454,N_15173);
nor U17018 (N_17018,N_15354,N_15667);
xnor U17019 (N_17019,N_15056,N_15723);
and U17020 (N_17020,N_15578,N_15176);
nor U17021 (N_17021,N_16137,N_15484);
or U17022 (N_17022,N_16234,N_15202);
xor U17023 (N_17023,N_15074,N_15292);
or U17024 (N_17024,N_15386,N_16058);
nand U17025 (N_17025,N_15842,N_16181);
nor U17026 (N_17026,N_15434,N_15614);
or U17027 (N_17027,N_15767,N_15899);
xor U17028 (N_17028,N_15169,N_15705);
and U17029 (N_17029,N_15013,N_15017);
nand U17030 (N_17030,N_16198,N_15334);
nand U17031 (N_17031,N_15878,N_15870);
xor U17032 (N_17032,N_16136,N_15809);
and U17033 (N_17033,N_15079,N_16188);
nor U17034 (N_17034,N_15533,N_15840);
nor U17035 (N_17035,N_15437,N_15173);
nand U17036 (N_17036,N_16156,N_15152);
or U17037 (N_17037,N_15743,N_15440);
nor U17038 (N_17038,N_15978,N_15185);
nor U17039 (N_17039,N_15938,N_15183);
xor U17040 (N_17040,N_15659,N_15645);
nand U17041 (N_17041,N_15552,N_16165);
nand U17042 (N_17042,N_16233,N_15950);
or U17043 (N_17043,N_15347,N_16185);
xor U17044 (N_17044,N_15548,N_15250);
nor U17045 (N_17045,N_15235,N_15102);
and U17046 (N_17046,N_15995,N_15794);
and U17047 (N_17047,N_15696,N_16029);
nand U17048 (N_17048,N_15946,N_15934);
nor U17049 (N_17049,N_15490,N_15055);
nand U17050 (N_17050,N_15194,N_15976);
nand U17051 (N_17051,N_15980,N_15705);
or U17052 (N_17052,N_15324,N_15551);
nand U17053 (N_17053,N_15074,N_15461);
or U17054 (N_17054,N_15067,N_16007);
nand U17055 (N_17055,N_15042,N_15961);
or U17056 (N_17056,N_15317,N_15364);
or U17057 (N_17057,N_15417,N_15565);
xnor U17058 (N_17058,N_15829,N_15259);
nand U17059 (N_17059,N_15235,N_15763);
nand U17060 (N_17060,N_15329,N_15472);
xnor U17061 (N_17061,N_15617,N_15940);
xnor U17062 (N_17062,N_16035,N_15000);
or U17063 (N_17063,N_15316,N_15337);
xor U17064 (N_17064,N_15007,N_16175);
xnor U17065 (N_17065,N_15279,N_15301);
nand U17066 (N_17066,N_15886,N_16212);
or U17067 (N_17067,N_15410,N_15755);
and U17068 (N_17068,N_15320,N_15929);
nand U17069 (N_17069,N_15997,N_15161);
nor U17070 (N_17070,N_15434,N_15540);
or U17071 (N_17071,N_15925,N_16177);
xnor U17072 (N_17072,N_15936,N_15287);
xor U17073 (N_17073,N_16211,N_15522);
or U17074 (N_17074,N_16157,N_16082);
and U17075 (N_17075,N_15426,N_15632);
or U17076 (N_17076,N_16024,N_15411);
and U17077 (N_17077,N_16196,N_16142);
nand U17078 (N_17078,N_15038,N_15740);
nand U17079 (N_17079,N_15103,N_15987);
or U17080 (N_17080,N_15802,N_15493);
and U17081 (N_17081,N_15193,N_15350);
and U17082 (N_17082,N_15715,N_15085);
xor U17083 (N_17083,N_16073,N_15421);
nand U17084 (N_17084,N_15408,N_16031);
xor U17085 (N_17085,N_15681,N_15317);
nor U17086 (N_17086,N_15927,N_15953);
nand U17087 (N_17087,N_15911,N_15019);
nor U17088 (N_17088,N_15098,N_15495);
nand U17089 (N_17089,N_15659,N_15825);
and U17090 (N_17090,N_15572,N_15289);
nand U17091 (N_17091,N_15922,N_16121);
or U17092 (N_17092,N_15470,N_16139);
nand U17093 (N_17093,N_15263,N_15239);
or U17094 (N_17094,N_16076,N_15179);
and U17095 (N_17095,N_15457,N_15741);
xor U17096 (N_17096,N_16056,N_15195);
xnor U17097 (N_17097,N_15069,N_16238);
nor U17098 (N_17098,N_15796,N_15607);
nand U17099 (N_17099,N_15627,N_15941);
or U17100 (N_17100,N_15368,N_15552);
nor U17101 (N_17101,N_16039,N_15235);
nor U17102 (N_17102,N_16219,N_15483);
nand U17103 (N_17103,N_15897,N_15838);
nor U17104 (N_17104,N_15826,N_15924);
or U17105 (N_17105,N_15896,N_15334);
nand U17106 (N_17106,N_15970,N_15674);
nand U17107 (N_17107,N_16058,N_16045);
nand U17108 (N_17108,N_15284,N_15156);
xor U17109 (N_17109,N_15147,N_15580);
or U17110 (N_17110,N_16041,N_15024);
xnor U17111 (N_17111,N_15953,N_15000);
nor U17112 (N_17112,N_15406,N_15209);
nand U17113 (N_17113,N_15758,N_15983);
xor U17114 (N_17114,N_15327,N_16237);
or U17115 (N_17115,N_15508,N_15696);
xor U17116 (N_17116,N_15335,N_16157);
xor U17117 (N_17117,N_15736,N_15446);
nor U17118 (N_17118,N_15583,N_15364);
nor U17119 (N_17119,N_16226,N_16054);
and U17120 (N_17120,N_15908,N_15495);
nor U17121 (N_17121,N_15661,N_15723);
xor U17122 (N_17122,N_15768,N_15170);
nand U17123 (N_17123,N_16122,N_15388);
or U17124 (N_17124,N_15649,N_16128);
nor U17125 (N_17125,N_15910,N_15413);
nand U17126 (N_17126,N_15846,N_16129);
or U17127 (N_17127,N_15929,N_15002);
nor U17128 (N_17128,N_15062,N_15420);
or U17129 (N_17129,N_16233,N_15552);
xor U17130 (N_17130,N_16075,N_15709);
and U17131 (N_17131,N_15923,N_15396);
nor U17132 (N_17132,N_16063,N_15147);
xnor U17133 (N_17133,N_16163,N_15035);
and U17134 (N_17134,N_15873,N_15878);
xnor U17135 (N_17135,N_15437,N_15194);
and U17136 (N_17136,N_15725,N_15578);
and U17137 (N_17137,N_15226,N_15532);
nand U17138 (N_17138,N_16008,N_15076);
or U17139 (N_17139,N_15322,N_15829);
and U17140 (N_17140,N_15866,N_15464);
or U17141 (N_17141,N_15955,N_15744);
and U17142 (N_17142,N_15160,N_15636);
nor U17143 (N_17143,N_16205,N_16004);
xnor U17144 (N_17144,N_15206,N_16236);
nand U17145 (N_17145,N_15644,N_15276);
nand U17146 (N_17146,N_15846,N_15000);
nand U17147 (N_17147,N_15373,N_15854);
xor U17148 (N_17148,N_15016,N_16097);
nand U17149 (N_17149,N_15750,N_15418);
xor U17150 (N_17150,N_15553,N_15982);
and U17151 (N_17151,N_15420,N_15637);
nor U17152 (N_17152,N_15939,N_16067);
xor U17153 (N_17153,N_15708,N_15658);
or U17154 (N_17154,N_16058,N_15536);
nand U17155 (N_17155,N_15990,N_16173);
and U17156 (N_17156,N_16086,N_15857);
nand U17157 (N_17157,N_15415,N_15497);
nand U17158 (N_17158,N_15032,N_15794);
or U17159 (N_17159,N_15164,N_15838);
xor U17160 (N_17160,N_15685,N_15528);
and U17161 (N_17161,N_15061,N_15539);
and U17162 (N_17162,N_15341,N_15572);
or U17163 (N_17163,N_15982,N_15791);
nor U17164 (N_17164,N_15420,N_15572);
nand U17165 (N_17165,N_15529,N_15621);
nand U17166 (N_17166,N_15789,N_15094);
xor U17167 (N_17167,N_15991,N_15221);
xor U17168 (N_17168,N_15135,N_16241);
nor U17169 (N_17169,N_15846,N_15699);
nor U17170 (N_17170,N_15434,N_15243);
xor U17171 (N_17171,N_15136,N_15984);
or U17172 (N_17172,N_15012,N_16062);
and U17173 (N_17173,N_15362,N_15699);
nand U17174 (N_17174,N_15494,N_15306);
xnor U17175 (N_17175,N_15822,N_15714);
nor U17176 (N_17176,N_15072,N_15146);
xor U17177 (N_17177,N_15912,N_16113);
nor U17178 (N_17178,N_15072,N_15604);
nand U17179 (N_17179,N_15958,N_16003);
or U17180 (N_17180,N_16238,N_15405);
nor U17181 (N_17181,N_15362,N_15914);
or U17182 (N_17182,N_15159,N_16221);
nor U17183 (N_17183,N_15016,N_15447);
xor U17184 (N_17184,N_15658,N_16194);
and U17185 (N_17185,N_15514,N_15377);
or U17186 (N_17186,N_15983,N_15384);
nor U17187 (N_17187,N_16111,N_16205);
or U17188 (N_17188,N_15216,N_15869);
nand U17189 (N_17189,N_15807,N_16076);
and U17190 (N_17190,N_15286,N_15922);
nor U17191 (N_17191,N_15363,N_15327);
xnor U17192 (N_17192,N_15446,N_15122);
nor U17193 (N_17193,N_16198,N_15557);
nand U17194 (N_17194,N_15480,N_15938);
nand U17195 (N_17195,N_15213,N_15764);
nand U17196 (N_17196,N_15140,N_15536);
and U17197 (N_17197,N_15173,N_15881);
nand U17198 (N_17198,N_15323,N_15452);
nand U17199 (N_17199,N_15043,N_15929);
xor U17200 (N_17200,N_15123,N_16086);
or U17201 (N_17201,N_15015,N_15700);
xnor U17202 (N_17202,N_15686,N_15288);
xnor U17203 (N_17203,N_15340,N_16116);
nand U17204 (N_17204,N_16005,N_15317);
xor U17205 (N_17205,N_16181,N_15136);
xnor U17206 (N_17206,N_15839,N_15675);
or U17207 (N_17207,N_15056,N_16071);
and U17208 (N_17208,N_15808,N_15172);
or U17209 (N_17209,N_15563,N_16091);
xor U17210 (N_17210,N_15995,N_15325);
nand U17211 (N_17211,N_15638,N_15788);
or U17212 (N_17212,N_16209,N_15333);
xor U17213 (N_17213,N_15026,N_15988);
xor U17214 (N_17214,N_15373,N_15153);
nand U17215 (N_17215,N_15352,N_15063);
nand U17216 (N_17216,N_15612,N_15039);
or U17217 (N_17217,N_15635,N_15625);
xor U17218 (N_17218,N_15832,N_15517);
nor U17219 (N_17219,N_16068,N_15580);
or U17220 (N_17220,N_15382,N_15833);
nor U17221 (N_17221,N_15646,N_16021);
xnor U17222 (N_17222,N_15838,N_15865);
xnor U17223 (N_17223,N_15028,N_15521);
and U17224 (N_17224,N_16241,N_15223);
and U17225 (N_17225,N_15094,N_16130);
xnor U17226 (N_17226,N_16241,N_15225);
xor U17227 (N_17227,N_16168,N_15738);
and U17228 (N_17228,N_15748,N_15709);
or U17229 (N_17229,N_15169,N_15596);
and U17230 (N_17230,N_16132,N_16244);
xor U17231 (N_17231,N_15551,N_15615);
nor U17232 (N_17232,N_15123,N_15738);
nand U17233 (N_17233,N_15801,N_16058);
and U17234 (N_17234,N_15008,N_16171);
nand U17235 (N_17235,N_15901,N_16140);
nor U17236 (N_17236,N_15197,N_16135);
nor U17237 (N_17237,N_15835,N_15062);
xnor U17238 (N_17238,N_15099,N_15097);
or U17239 (N_17239,N_16148,N_15785);
or U17240 (N_17240,N_15136,N_16052);
nand U17241 (N_17241,N_15437,N_16020);
nand U17242 (N_17242,N_15237,N_16049);
or U17243 (N_17243,N_15278,N_15324);
nand U17244 (N_17244,N_15762,N_16093);
nand U17245 (N_17245,N_15166,N_15388);
or U17246 (N_17246,N_15952,N_16212);
nand U17247 (N_17247,N_15424,N_15055);
xor U17248 (N_17248,N_15117,N_16061);
nand U17249 (N_17249,N_16004,N_15892);
xor U17250 (N_17250,N_15703,N_15435);
or U17251 (N_17251,N_15586,N_15997);
nor U17252 (N_17252,N_15648,N_15726);
xnor U17253 (N_17253,N_15533,N_15160);
or U17254 (N_17254,N_15664,N_15842);
or U17255 (N_17255,N_16085,N_15806);
and U17256 (N_17256,N_15345,N_15034);
nor U17257 (N_17257,N_15112,N_15561);
nor U17258 (N_17258,N_16032,N_15171);
and U17259 (N_17259,N_16238,N_15188);
nand U17260 (N_17260,N_16226,N_15636);
nand U17261 (N_17261,N_16156,N_16119);
or U17262 (N_17262,N_16202,N_15903);
xor U17263 (N_17263,N_15183,N_15471);
nor U17264 (N_17264,N_15772,N_15341);
and U17265 (N_17265,N_15542,N_15422);
and U17266 (N_17266,N_15910,N_15012);
xnor U17267 (N_17267,N_15080,N_15542);
and U17268 (N_17268,N_15270,N_15792);
xor U17269 (N_17269,N_16013,N_16034);
xor U17270 (N_17270,N_15412,N_15913);
or U17271 (N_17271,N_15030,N_15157);
nand U17272 (N_17272,N_16155,N_15304);
and U17273 (N_17273,N_16048,N_15953);
and U17274 (N_17274,N_15096,N_15418);
xnor U17275 (N_17275,N_15358,N_15775);
xnor U17276 (N_17276,N_15595,N_15761);
nand U17277 (N_17277,N_15527,N_15659);
nor U17278 (N_17278,N_15619,N_15580);
nor U17279 (N_17279,N_15072,N_15833);
or U17280 (N_17280,N_15527,N_15403);
nor U17281 (N_17281,N_15455,N_16202);
or U17282 (N_17282,N_15045,N_15594);
or U17283 (N_17283,N_15696,N_15210);
nor U17284 (N_17284,N_15628,N_15780);
xor U17285 (N_17285,N_16142,N_15773);
or U17286 (N_17286,N_15723,N_15847);
nor U17287 (N_17287,N_16011,N_15815);
nand U17288 (N_17288,N_15508,N_16026);
or U17289 (N_17289,N_15168,N_15197);
nand U17290 (N_17290,N_16147,N_15016);
or U17291 (N_17291,N_15828,N_15994);
xor U17292 (N_17292,N_15359,N_15883);
and U17293 (N_17293,N_15131,N_16067);
and U17294 (N_17294,N_16114,N_15021);
nand U17295 (N_17295,N_15225,N_15001);
nand U17296 (N_17296,N_16172,N_16242);
and U17297 (N_17297,N_15611,N_15602);
xor U17298 (N_17298,N_15282,N_15177);
nand U17299 (N_17299,N_15743,N_15040);
nor U17300 (N_17300,N_15278,N_16237);
xnor U17301 (N_17301,N_15043,N_15499);
nand U17302 (N_17302,N_15406,N_15486);
nor U17303 (N_17303,N_15493,N_15843);
xnor U17304 (N_17304,N_15092,N_15941);
or U17305 (N_17305,N_16128,N_16059);
and U17306 (N_17306,N_15401,N_15791);
xnor U17307 (N_17307,N_16148,N_15264);
xnor U17308 (N_17308,N_15217,N_15343);
or U17309 (N_17309,N_15813,N_16056);
nor U17310 (N_17310,N_15525,N_15339);
xnor U17311 (N_17311,N_15523,N_15846);
nand U17312 (N_17312,N_15489,N_15052);
and U17313 (N_17313,N_15311,N_16076);
or U17314 (N_17314,N_16105,N_15161);
nand U17315 (N_17315,N_16186,N_16057);
xnor U17316 (N_17316,N_15645,N_15817);
nor U17317 (N_17317,N_15225,N_15050);
nand U17318 (N_17318,N_15886,N_15405);
or U17319 (N_17319,N_15786,N_15049);
nor U17320 (N_17320,N_15138,N_15146);
and U17321 (N_17321,N_15289,N_15508);
nor U17322 (N_17322,N_15506,N_15916);
nor U17323 (N_17323,N_15059,N_15956);
or U17324 (N_17324,N_16025,N_16050);
xor U17325 (N_17325,N_15527,N_15512);
nor U17326 (N_17326,N_15597,N_15836);
or U17327 (N_17327,N_15576,N_15352);
or U17328 (N_17328,N_15683,N_15330);
or U17329 (N_17329,N_16060,N_15930);
or U17330 (N_17330,N_15413,N_15373);
nor U17331 (N_17331,N_15463,N_16165);
nand U17332 (N_17332,N_15986,N_15446);
and U17333 (N_17333,N_15324,N_15177);
nor U17334 (N_17334,N_15308,N_16017);
xnor U17335 (N_17335,N_15213,N_15892);
xor U17336 (N_17336,N_15371,N_16127);
nor U17337 (N_17337,N_15035,N_15210);
xnor U17338 (N_17338,N_15712,N_15380);
nand U17339 (N_17339,N_15515,N_15899);
xor U17340 (N_17340,N_15788,N_15429);
nor U17341 (N_17341,N_15067,N_15172);
or U17342 (N_17342,N_15814,N_15429);
xor U17343 (N_17343,N_15268,N_15307);
and U17344 (N_17344,N_15589,N_15187);
and U17345 (N_17345,N_16114,N_15028);
and U17346 (N_17346,N_15495,N_15822);
nor U17347 (N_17347,N_15869,N_15667);
nor U17348 (N_17348,N_15288,N_15048);
nor U17349 (N_17349,N_15012,N_15519);
xnor U17350 (N_17350,N_15549,N_15225);
xor U17351 (N_17351,N_15093,N_15665);
xnor U17352 (N_17352,N_16022,N_15799);
and U17353 (N_17353,N_15002,N_15257);
and U17354 (N_17354,N_15692,N_15575);
and U17355 (N_17355,N_15589,N_15643);
xor U17356 (N_17356,N_15342,N_15466);
nor U17357 (N_17357,N_15008,N_15891);
and U17358 (N_17358,N_15179,N_15993);
nor U17359 (N_17359,N_15461,N_15142);
nand U17360 (N_17360,N_15283,N_16230);
or U17361 (N_17361,N_15306,N_15907);
or U17362 (N_17362,N_15172,N_15001);
and U17363 (N_17363,N_16006,N_15797);
or U17364 (N_17364,N_16157,N_15849);
xnor U17365 (N_17365,N_15006,N_16239);
nor U17366 (N_17366,N_16193,N_16133);
nor U17367 (N_17367,N_15524,N_15758);
nor U17368 (N_17368,N_15200,N_15802);
or U17369 (N_17369,N_15851,N_15751);
nand U17370 (N_17370,N_15747,N_15964);
nor U17371 (N_17371,N_15967,N_15259);
or U17372 (N_17372,N_16187,N_15520);
nand U17373 (N_17373,N_16215,N_15736);
nor U17374 (N_17374,N_16045,N_15930);
or U17375 (N_17375,N_15706,N_15815);
xnor U17376 (N_17376,N_15509,N_15979);
nand U17377 (N_17377,N_16201,N_16037);
nor U17378 (N_17378,N_15602,N_16016);
or U17379 (N_17379,N_15839,N_16021);
xor U17380 (N_17380,N_15647,N_15383);
nor U17381 (N_17381,N_15039,N_15295);
xor U17382 (N_17382,N_15628,N_15975);
or U17383 (N_17383,N_15490,N_15567);
or U17384 (N_17384,N_15618,N_16099);
or U17385 (N_17385,N_16242,N_15195);
xnor U17386 (N_17386,N_16147,N_15552);
and U17387 (N_17387,N_15232,N_16231);
or U17388 (N_17388,N_15396,N_16024);
or U17389 (N_17389,N_15136,N_15032);
and U17390 (N_17390,N_15958,N_15037);
or U17391 (N_17391,N_15958,N_15095);
nand U17392 (N_17392,N_15920,N_15372);
or U17393 (N_17393,N_15665,N_16046);
nand U17394 (N_17394,N_15366,N_15671);
nand U17395 (N_17395,N_15578,N_15150);
nor U17396 (N_17396,N_15775,N_15494);
or U17397 (N_17397,N_16117,N_15590);
nand U17398 (N_17398,N_15314,N_16247);
xor U17399 (N_17399,N_15491,N_15036);
nor U17400 (N_17400,N_15563,N_16041);
nand U17401 (N_17401,N_15797,N_16200);
nor U17402 (N_17402,N_16019,N_15035);
nand U17403 (N_17403,N_16181,N_15014);
and U17404 (N_17404,N_15036,N_15511);
or U17405 (N_17405,N_15659,N_15397);
and U17406 (N_17406,N_15868,N_15075);
xnor U17407 (N_17407,N_15694,N_15312);
nor U17408 (N_17408,N_15745,N_16070);
nor U17409 (N_17409,N_15615,N_15844);
and U17410 (N_17410,N_15200,N_15845);
nand U17411 (N_17411,N_16044,N_15521);
and U17412 (N_17412,N_15598,N_15558);
or U17413 (N_17413,N_15139,N_15235);
or U17414 (N_17414,N_15307,N_16050);
nand U17415 (N_17415,N_15569,N_15013);
and U17416 (N_17416,N_16168,N_15957);
nor U17417 (N_17417,N_15157,N_15060);
xor U17418 (N_17418,N_15689,N_15277);
and U17419 (N_17419,N_15964,N_15333);
or U17420 (N_17420,N_15436,N_15674);
nor U17421 (N_17421,N_15080,N_16092);
nand U17422 (N_17422,N_16148,N_16061);
or U17423 (N_17423,N_16112,N_15086);
and U17424 (N_17424,N_15132,N_15710);
nor U17425 (N_17425,N_15574,N_15932);
xnor U17426 (N_17426,N_16161,N_15517);
nand U17427 (N_17427,N_15307,N_15767);
nand U17428 (N_17428,N_15314,N_15640);
and U17429 (N_17429,N_15406,N_16194);
and U17430 (N_17430,N_16033,N_16083);
and U17431 (N_17431,N_15723,N_15805);
nor U17432 (N_17432,N_15039,N_15117);
nor U17433 (N_17433,N_15522,N_16209);
or U17434 (N_17434,N_16244,N_15809);
nand U17435 (N_17435,N_15012,N_16140);
nor U17436 (N_17436,N_15091,N_15092);
and U17437 (N_17437,N_15735,N_16040);
nor U17438 (N_17438,N_15533,N_15348);
nand U17439 (N_17439,N_16098,N_15653);
nand U17440 (N_17440,N_15934,N_15047);
or U17441 (N_17441,N_16188,N_15761);
and U17442 (N_17442,N_15964,N_16200);
or U17443 (N_17443,N_15006,N_15745);
or U17444 (N_17444,N_15930,N_15030);
nand U17445 (N_17445,N_16171,N_16021);
xnor U17446 (N_17446,N_15514,N_15848);
nand U17447 (N_17447,N_16159,N_16113);
or U17448 (N_17448,N_15962,N_15600);
nor U17449 (N_17449,N_15713,N_15575);
and U17450 (N_17450,N_15935,N_15287);
xnor U17451 (N_17451,N_15981,N_15950);
nor U17452 (N_17452,N_15581,N_15482);
or U17453 (N_17453,N_16220,N_15891);
xnor U17454 (N_17454,N_16067,N_15166);
or U17455 (N_17455,N_15112,N_15416);
nor U17456 (N_17456,N_15468,N_15819);
or U17457 (N_17457,N_15168,N_15037);
nand U17458 (N_17458,N_16142,N_16191);
nand U17459 (N_17459,N_15404,N_15572);
and U17460 (N_17460,N_15846,N_15298);
nand U17461 (N_17461,N_16118,N_15439);
and U17462 (N_17462,N_15165,N_15769);
nor U17463 (N_17463,N_15846,N_15038);
nand U17464 (N_17464,N_15811,N_15790);
xnor U17465 (N_17465,N_15245,N_15799);
nand U17466 (N_17466,N_15295,N_15443);
nor U17467 (N_17467,N_15171,N_16201);
nand U17468 (N_17468,N_15201,N_15542);
xor U17469 (N_17469,N_16035,N_15145);
nor U17470 (N_17470,N_15166,N_15863);
nor U17471 (N_17471,N_15640,N_16117);
and U17472 (N_17472,N_15341,N_15618);
nand U17473 (N_17473,N_15958,N_15345);
nor U17474 (N_17474,N_16155,N_15114);
nand U17475 (N_17475,N_15866,N_16010);
or U17476 (N_17476,N_15768,N_15974);
nor U17477 (N_17477,N_15865,N_16135);
nand U17478 (N_17478,N_15934,N_15595);
nand U17479 (N_17479,N_15374,N_15909);
or U17480 (N_17480,N_15441,N_16226);
or U17481 (N_17481,N_15437,N_15462);
and U17482 (N_17482,N_15732,N_15425);
xor U17483 (N_17483,N_15681,N_15123);
nand U17484 (N_17484,N_15060,N_15154);
or U17485 (N_17485,N_16199,N_15809);
or U17486 (N_17486,N_15504,N_16153);
nor U17487 (N_17487,N_15555,N_15534);
or U17488 (N_17488,N_16012,N_15504);
or U17489 (N_17489,N_15309,N_15459);
and U17490 (N_17490,N_15407,N_15692);
nor U17491 (N_17491,N_15896,N_15542);
nor U17492 (N_17492,N_16185,N_15655);
nor U17493 (N_17493,N_15986,N_15359);
or U17494 (N_17494,N_15663,N_15018);
xnor U17495 (N_17495,N_15873,N_16147);
nor U17496 (N_17496,N_15330,N_15072);
nand U17497 (N_17497,N_15490,N_15421);
nor U17498 (N_17498,N_15398,N_15304);
and U17499 (N_17499,N_15683,N_15302);
and U17500 (N_17500,N_17479,N_16473);
nand U17501 (N_17501,N_17312,N_17043);
nand U17502 (N_17502,N_17143,N_17217);
nor U17503 (N_17503,N_17122,N_17068);
nor U17504 (N_17504,N_16831,N_17450);
and U17505 (N_17505,N_17069,N_16954);
xnor U17506 (N_17506,N_16577,N_17200);
nor U17507 (N_17507,N_17047,N_17014);
nand U17508 (N_17508,N_16888,N_17152);
nor U17509 (N_17509,N_17289,N_17250);
and U17510 (N_17510,N_17121,N_16523);
or U17511 (N_17511,N_16754,N_17347);
nand U17512 (N_17512,N_17215,N_17193);
and U17513 (N_17513,N_16460,N_16886);
nor U17514 (N_17514,N_16753,N_16876);
and U17515 (N_17515,N_17209,N_16775);
and U17516 (N_17516,N_16379,N_17073);
nand U17517 (N_17517,N_17429,N_16450);
and U17518 (N_17518,N_16591,N_16275);
nor U17519 (N_17519,N_17054,N_16397);
or U17520 (N_17520,N_17346,N_16571);
nor U17521 (N_17521,N_17452,N_17461);
nor U17522 (N_17522,N_16688,N_16630);
xor U17523 (N_17523,N_16493,N_16663);
and U17524 (N_17524,N_17168,N_16426);
nor U17525 (N_17525,N_16913,N_17368);
or U17526 (N_17526,N_16525,N_16385);
and U17527 (N_17527,N_17344,N_16787);
nand U17528 (N_17528,N_16905,N_16367);
and U17529 (N_17529,N_17225,N_16323);
nor U17530 (N_17530,N_16497,N_16603);
or U17531 (N_17531,N_16281,N_16760);
xnor U17532 (N_17532,N_17363,N_16793);
or U17533 (N_17533,N_17166,N_17196);
nor U17534 (N_17534,N_16767,N_16916);
or U17535 (N_17535,N_16956,N_17300);
xor U17536 (N_17536,N_16866,N_17383);
nor U17537 (N_17537,N_16666,N_16797);
nand U17538 (N_17538,N_16352,N_17324);
xnor U17539 (N_17539,N_16692,N_17431);
and U17540 (N_17540,N_17293,N_16257);
or U17541 (N_17541,N_17449,N_16803);
nand U17542 (N_17542,N_16883,N_16477);
nor U17543 (N_17543,N_16683,N_16621);
or U17544 (N_17544,N_17058,N_16359);
or U17545 (N_17545,N_17208,N_17007);
nor U17546 (N_17546,N_17235,N_16463);
and U17547 (N_17547,N_16798,N_17485);
and U17548 (N_17548,N_17448,N_17171);
xor U17549 (N_17549,N_17309,N_16826);
and U17550 (N_17550,N_16972,N_16776);
xnor U17551 (N_17551,N_16759,N_17318);
and U17552 (N_17552,N_17146,N_17160);
nand U17553 (N_17553,N_17304,N_17343);
nor U17554 (N_17554,N_16755,N_16900);
and U17555 (N_17555,N_16847,N_16893);
nand U17556 (N_17556,N_17302,N_17101);
xnor U17557 (N_17557,N_17236,N_16739);
and U17558 (N_17558,N_17157,N_16836);
nand U17559 (N_17559,N_17028,N_16895);
xnor U17560 (N_17560,N_16504,N_17335);
or U17561 (N_17561,N_16652,N_16838);
or U17562 (N_17562,N_16469,N_17412);
nand U17563 (N_17563,N_16973,N_16277);
and U17564 (N_17564,N_16537,N_16413);
xnor U17565 (N_17565,N_17390,N_16583);
xnor U17566 (N_17566,N_16660,N_16909);
xor U17567 (N_17567,N_17469,N_16619);
xor U17568 (N_17568,N_17388,N_17084);
or U17569 (N_17569,N_17252,N_16821);
nand U17570 (N_17570,N_16865,N_16773);
nor U17571 (N_17571,N_16606,N_16509);
or U17572 (N_17572,N_17366,N_17264);
nor U17573 (N_17573,N_16453,N_16500);
nand U17574 (N_17574,N_16890,N_17443);
and U17575 (N_17575,N_17331,N_17391);
or U17576 (N_17576,N_17371,N_16542);
nor U17577 (N_17577,N_17267,N_16372);
or U17578 (N_17578,N_16270,N_16943);
and U17579 (N_17579,N_16696,N_16851);
and U17580 (N_17580,N_17222,N_16837);
nand U17581 (N_17581,N_16333,N_16917);
or U17582 (N_17582,N_16875,N_16348);
nand U17583 (N_17583,N_17440,N_17389);
xor U17584 (N_17584,N_16977,N_17078);
and U17585 (N_17585,N_17308,N_17317);
and U17586 (N_17586,N_17032,N_16748);
and U17587 (N_17587,N_17133,N_16626);
xnor U17588 (N_17588,N_17057,N_16908);
xor U17589 (N_17589,N_16302,N_16639);
and U17590 (N_17590,N_17367,N_17397);
or U17591 (N_17591,N_16991,N_16314);
xor U17592 (N_17592,N_16356,N_16564);
nor U17593 (N_17593,N_16827,N_17056);
or U17594 (N_17594,N_16967,N_16587);
or U17595 (N_17595,N_16350,N_16378);
xor U17596 (N_17596,N_17240,N_17123);
and U17597 (N_17597,N_16613,N_17188);
xnor U17598 (N_17598,N_16769,N_16915);
and U17599 (N_17599,N_16365,N_17021);
and U17600 (N_17600,N_16389,N_16854);
nor U17601 (N_17601,N_16297,N_16830);
and U17602 (N_17602,N_16300,N_16870);
xor U17603 (N_17603,N_16633,N_16774);
xnor U17604 (N_17604,N_16730,N_17134);
and U17605 (N_17605,N_17035,N_17045);
nor U17606 (N_17606,N_16404,N_16716);
nor U17607 (N_17607,N_16501,N_17059);
nor U17608 (N_17608,N_17190,N_16993);
nor U17609 (N_17609,N_16401,N_16510);
or U17610 (N_17610,N_17067,N_16641);
xnor U17611 (N_17611,N_16702,N_16261);
nand U17612 (N_17612,N_16332,N_17170);
xnor U17613 (N_17613,N_17065,N_17341);
and U17614 (N_17614,N_16573,N_16354);
and U17615 (N_17615,N_16648,N_17204);
and U17616 (N_17616,N_16659,N_16313);
nand U17617 (N_17617,N_17219,N_16394);
nor U17618 (N_17618,N_16963,N_16996);
xnor U17619 (N_17619,N_16853,N_17287);
nand U17620 (N_17620,N_16757,N_17182);
nor U17621 (N_17621,N_17083,N_17022);
and U17622 (N_17622,N_17336,N_17223);
or U17623 (N_17623,N_17462,N_17072);
nor U17624 (N_17624,N_16299,N_16346);
or U17625 (N_17625,N_16285,N_17475);
and U17626 (N_17626,N_16945,N_17255);
xnor U17627 (N_17627,N_16693,N_16914);
or U17628 (N_17628,N_16391,N_17256);
or U17629 (N_17629,N_16687,N_17292);
and U17630 (N_17630,N_16650,N_17418);
nor U17631 (N_17631,N_16799,N_17307);
nor U17632 (N_17632,N_16265,N_16263);
or U17633 (N_17633,N_17420,N_16843);
and U17634 (N_17634,N_17147,N_16358);
nor U17635 (N_17635,N_16530,N_16428);
nor U17636 (N_17636,N_17115,N_16985);
and U17637 (N_17637,N_16361,N_16982);
nor U17638 (N_17638,N_16825,N_16946);
nor U17639 (N_17639,N_16386,N_16872);
nand U17640 (N_17640,N_16927,N_16910);
nand U17641 (N_17641,N_17135,N_16321);
nand U17642 (N_17642,N_17494,N_16536);
nor U17643 (N_17643,N_16325,N_17338);
or U17644 (N_17644,N_17424,N_17203);
xnor U17645 (N_17645,N_16283,N_17254);
or U17646 (N_17646,N_16515,N_16535);
nand U17647 (N_17647,N_16834,N_17176);
and U17648 (N_17648,N_16654,N_16483);
xnor U17649 (N_17649,N_16809,N_16360);
xnor U17650 (N_17650,N_16820,N_16408);
nor U17651 (N_17651,N_17109,N_16789);
nand U17652 (N_17652,N_16912,N_16565);
nor U17653 (N_17653,N_16474,N_16745);
and U17654 (N_17654,N_17098,N_17396);
nor U17655 (N_17655,N_16522,N_16835);
nand U17656 (N_17656,N_17298,N_16676);
nand U17657 (N_17657,N_16715,N_17149);
xor U17658 (N_17658,N_16637,N_17474);
nand U17659 (N_17659,N_16980,N_16792);
or U17660 (N_17660,N_16618,N_17359);
or U17661 (N_17661,N_16863,N_16423);
xor U17662 (N_17662,N_17386,N_16287);
or U17663 (N_17663,N_16289,N_17230);
xor U17664 (N_17664,N_16976,N_16988);
xnor U17665 (N_17665,N_16488,N_17159);
xor U17666 (N_17666,N_17144,N_16387);
xnor U17667 (N_17667,N_17198,N_17185);
and U17668 (N_17668,N_17046,N_17408);
xnor U17669 (N_17669,N_17114,N_16364);
xor U17670 (N_17670,N_17333,N_16327);
and U17671 (N_17671,N_16725,N_16464);
nand U17672 (N_17672,N_17273,N_16765);
or U17673 (N_17673,N_16925,N_16931);
nor U17674 (N_17674,N_16407,N_16955);
nand U17675 (N_17675,N_17457,N_16860);
or U17676 (N_17676,N_16766,N_16528);
nand U17677 (N_17677,N_16881,N_16567);
and U17678 (N_17678,N_16429,N_17214);
or U17679 (N_17679,N_16832,N_16778);
nand U17680 (N_17680,N_16944,N_16761);
or U17681 (N_17681,N_17179,N_16329);
nand U17682 (N_17682,N_16402,N_17361);
and U17683 (N_17683,N_17053,N_16324);
or U17684 (N_17684,N_17194,N_17498);
nand U17685 (N_17685,N_17232,N_17097);
nor U17686 (N_17686,N_16458,N_17374);
nand U17687 (N_17687,N_17082,N_16627);
nand U17688 (N_17688,N_16740,N_17216);
and U17689 (N_17689,N_16952,N_17493);
nor U17690 (N_17690,N_16703,N_16783);
nand U17691 (N_17691,N_16309,N_16634);
nand U17692 (N_17692,N_17484,N_16884);
nand U17693 (N_17693,N_17294,N_16852);
nor U17694 (N_17694,N_16625,N_17093);
and U17695 (N_17695,N_16801,N_16431);
and U17696 (N_17696,N_16635,N_16343);
and U17697 (N_17697,N_16370,N_16505);
xor U17698 (N_17698,N_16710,N_17476);
or U17699 (N_17699,N_16345,N_16588);
or U17700 (N_17700,N_17370,N_16709);
or U17701 (N_17701,N_17112,N_16294);
nor U17702 (N_17702,N_16719,N_16507);
nand U17703 (N_17703,N_16494,N_16472);
or U17704 (N_17704,N_17221,N_16484);
or U17705 (N_17705,N_17076,N_17410);
nor U17706 (N_17706,N_16341,N_17094);
nand U17707 (N_17707,N_16903,N_16490);
or U17708 (N_17708,N_16369,N_16572);
or U17709 (N_17709,N_16264,N_16858);
nor U17710 (N_17710,N_16975,N_16540);
and U17711 (N_17711,N_16434,N_16651);
and U17712 (N_17712,N_16878,N_16492);
nand U17713 (N_17713,N_16962,N_16561);
or U17714 (N_17714,N_17062,N_17434);
nand U17715 (N_17715,N_16935,N_16259);
xnor U17716 (N_17716,N_16254,N_17055);
and U17717 (N_17717,N_17274,N_17316);
and U17718 (N_17718,N_17070,N_16796);
xor U17719 (N_17719,N_16738,N_16506);
xor U17720 (N_17720,N_16411,N_16271);
xnor U17721 (N_17721,N_17445,N_16595);
xnor U17722 (N_17722,N_16258,N_16547);
xnor U17723 (N_17723,N_17174,N_16871);
nand U17724 (N_17724,N_16318,N_17422);
and U17725 (N_17725,N_17402,N_17348);
nand U17726 (N_17726,N_16701,N_17413);
or U17727 (N_17727,N_16602,N_17224);
or U17728 (N_17728,N_16685,N_17245);
nand U17729 (N_17729,N_16758,N_17407);
xor U17730 (N_17730,N_16462,N_16657);
or U17731 (N_17731,N_16815,N_16763);
nor U17732 (N_17732,N_16310,N_16780);
and U17733 (N_17733,N_17088,N_17118);
and U17734 (N_17734,N_17387,N_16449);
and U17735 (N_17735,N_17433,N_16427);
or U17736 (N_17736,N_17125,N_16785);
nand U17737 (N_17737,N_16622,N_16467);
nand U17738 (N_17738,N_16942,N_16316);
xor U17739 (N_17739,N_16276,N_17460);
and U17740 (N_17740,N_16723,N_16608);
nand U17741 (N_17741,N_16384,N_17148);
xor U17742 (N_17742,N_16339,N_16959);
nor U17743 (N_17743,N_16303,N_17169);
xor U17744 (N_17744,N_16999,N_16322);
nor U17745 (N_17745,N_16713,N_17063);
xor U17746 (N_17746,N_17323,N_16274);
and U17747 (N_17747,N_17427,N_16861);
and U17748 (N_17748,N_16779,N_17036);
xnor U17749 (N_17749,N_17016,N_16312);
nand U17750 (N_17750,N_17442,N_16777);
nand U17751 (N_17751,N_16711,N_17353);
and U17752 (N_17752,N_16425,N_16894);
or U17753 (N_17753,N_17282,N_16272);
nand U17754 (N_17754,N_16373,N_16306);
or U17755 (N_17755,N_16400,N_17326);
xnor U17756 (N_17756,N_16447,N_17131);
nand U17757 (N_17757,N_16947,N_16308);
xnor U17758 (N_17758,N_16794,N_16415);
xor U17759 (N_17759,N_16278,N_17002);
and U17760 (N_17760,N_16568,N_16670);
xnor U17761 (N_17761,N_17241,N_16465);
and U17762 (N_17762,N_17436,N_16502);
or U17763 (N_17763,N_17465,N_17154);
xnor U17764 (N_17764,N_16867,N_17111);
nor U17765 (N_17765,N_17438,N_17291);
nand U17766 (N_17766,N_16614,N_16690);
and U17767 (N_17767,N_17401,N_16563);
xor U17768 (N_17768,N_17364,N_17334);
or U17769 (N_17769,N_16526,N_16399);
nand U17770 (N_17770,N_17044,N_17048);
xor U17771 (N_17771,N_17419,N_16416);
nor U17772 (N_17772,N_16933,N_16366);
nor U17773 (N_17773,N_16390,N_17080);
nor U17774 (N_17774,N_16279,N_17471);
or U17775 (N_17775,N_17261,N_17126);
or U17776 (N_17776,N_16601,N_16856);
and U17777 (N_17777,N_16700,N_16335);
xnor U17778 (N_17778,N_16623,N_17060);
nand U17779 (N_17779,N_16694,N_17150);
and U17780 (N_17780,N_17011,N_16266);
nor U17781 (N_17781,N_16684,N_17173);
nand U17782 (N_17782,N_17310,N_16554);
nor U17783 (N_17783,N_16818,N_17000);
nand U17784 (N_17784,N_16849,N_17253);
nand U17785 (N_17785,N_17033,N_16334);
and U17786 (N_17786,N_17066,N_16291);
nor U17787 (N_17787,N_17142,N_17330);
nand U17788 (N_17788,N_16786,N_16788);
or U17789 (N_17789,N_16671,N_16732);
nor U17790 (N_17790,N_17180,N_17006);
nand U17791 (N_17791,N_16337,N_16848);
xnor U17792 (N_17792,N_16901,N_17362);
xor U17793 (N_17793,N_17453,N_16610);
and U17794 (N_17794,N_17244,N_17089);
nor U17795 (N_17795,N_16560,N_17064);
and U17796 (N_17796,N_17491,N_17435);
and U17797 (N_17797,N_16969,N_16879);
xnor U17798 (N_17798,N_16841,N_17195);
nand U17799 (N_17799,N_16586,N_17394);
nand U17800 (N_17800,N_16989,N_17092);
nor U17801 (N_17801,N_16664,N_17430);
nor U17802 (N_17802,N_16482,N_17266);
nand U17803 (N_17803,N_16669,N_16422);
nand U17804 (N_17804,N_17151,N_16363);
nor U17805 (N_17805,N_17480,N_16470);
or U17806 (N_17806,N_16548,N_17399);
nand U17807 (N_17807,N_17263,N_16344);
and U17808 (N_17808,N_17315,N_16673);
xnor U17809 (N_17809,N_16771,N_17466);
nand U17810 (N_17810,N_17459,N_17275);
nand U17811 (N_17811,N_17458,N_16762);
nor U17812 (N_17812,N_16668,N_16691);
and U17813 (N_17813,N_17379,N_17329);
nor U17814 (N_17814,N_16770,N_16403);
and U17815 (N_17815,N_16288,N_16877);
or U17816 (N_17816,N_17237,N_17246);
xnor U17817 (N_17817,N_16612,N_16398);
nor U17818 (N_17818,N_16442,N_17400);
xor U17819 (N_17819,N_17117,N_17417);
xnor U17820 (N_17820,N_16708,N_17226);
or U17821 (N_17821,N_17110,N_16750);
nor U17822 (N_17822,N_16672,N_16508);
nor U17823 (N_17823,N_17153,N_16459);
or U17824 (N_17824,N_16937,N_17488);
xnor U17825 (N_17825,N_17155,N_17280);
nor U17826 (N_17826,N_17482,N_17281);
nand U17827 (N_17827,N_16987,N_16896);
or U17828 (N_17828,N_17050,N_16282);
nor U17829 (N_17829,N_17013,N_17186);
nand U17830 (N_17830,N_17325,N_17385);
nand U17831 (N_17831,N_17103,N_17259);
or U17832 (N_17832,N_16751,N_17052);
nand U17833 (N_17833,N_16496,N_16349);
or U17834 (N_17834,N_17249,N_16475);
xor U17835 (N_17835,N_17130,N_16628);
xor U17836 (N_17836,N_16643,N_17439);
xnor U17837 (N_17837,N_16468,N_16791);
xor U17838 (N_17838,N_17243,N_17376);
xor U17839 (N_17839,N_16889,N_16768);
nor U17840 (N_17840,N_16461,N_17090);
or U17841 (N_17841,N_16374,N_16533);
xnor U17842 (N_17842,N_16534,N_16524);
nor U17843 (N_17843,N_16706,N_17455);
xnor U17844 (N_17844,N_16380,N_16499);
and U17845 (N_17845,N_17020,N_16966);
nand U17846 (N_17846,N_16772,N_16727);
and U17847 (N_17847,N_17004,N_16897);
xor U17848 (N_17848,N_17119,N_16882);
nand U17849 (N_17849,N_16305,N_17276);
nand U17850 (N_17850,N_17290,N_16436);
nor U17851 (N_17851,N_16457,N_17034);
and U17852 (N_17852,N_16992,N_16412);
xor U17853 (N_17853,N_17463,N_16326);
and U17854 (N_17854,N_17297,N_16418);
nor U17855 (N_17855,N_16932,N_17113);
xor U17856 (N_17856,N_17349,N_16414);
or U17857 (N_17857,N_16581,N_17178);
or U17858 (N_17858,N_17495,N_17358);
or U17859 (N_17859,N_16292,N_17165);
and U17860 (N_17860,N_17128,N_16377);
and U17861 (N_17861,N_17025,N_16924);
nand U17862 (N_17862,N_17392,N_16580);
nor U17863 (N_17863,N_16336,N_17105);
and U17864 (N_17864,N_17061,N_17345);
or U17865 (N_17865,N_16647,N_16911);
xor U17866 (N_17866,N_16998,N_17187);
nor U17867 (N_17867,N_16576,N_16950);
or U17868 (N_17868,N_16790,N_16728);
nand U17869 (N_17869,N_16656,N_16569);
and U17870 (N_17870,N_16938,N_16615);
xor U17871 (N_17871,N_17156,N_16986);
nand U17872 (N_17872,N_16317,N_17369);
nor U17873 (N_17873,N_16655,N_17238);
nor U17874 (N_17874,N_16511,N_16828);
xor U17875 (N_17875,N_17029,N_17191);
or U17876 (N_17876,N_16984,N_16632);
nand U17877 (N_17877,N_16640,N_17247);
nand U17878 (N_17878,N_17478,N_17406);
or U17879 (N_17879,N_16466,N_16448);
nand U17880 (N_17880,N_17177,N_17271);
nand U17881 (N_17881,N_16964,N_16440);
xnor U17882 (N_17882,N_16679,N_17099);
xnor U17883 (N_17883,N_16644,N_17183);
nand U17884 (N_17884,N_17486,N_16810);
xor U17885 (N_17885,N_16438,N_16579);
or U17886 (N_17886,N_17031,N_16819);
xnor U17887 (N_17887,N_16782,N_17205);
xnor U17888 (N_17888,N_16295,N_17199);
xor U17889 (N_17889,N_16990,N_16296);
nand U17890 (N_17890,N_16347,N_17295);
and U17891 (N_17891,N_17081,N_17432);
nand U17892 (N_17892,N_16868,N_16487);
or U17893 (N_17893,N_16405,N_16743);
and U17894 (N_17894,N_17023,N_16362);
nor U17895 (N_17895,N_16741,N_17306);
xor U17896 (N_17896,N_17161,N_17421);
or U17897 (N_17897,N_17039,N_17041);
or U17898 (N_17898,N_17409,N_17124);
or U17899 (N_17899,N_16607,N_17415);
or U17900 (N_17900,N_17030,N_16965);
or U17901 (N_17901,N_17136,N_17079);
xor U17902 (N_17902,N_17251,N_16646);
xnor U17903 (N_17903,N_16697,N_16752);
xnor U17904 (N_17904,N_16551,N_16922);
xnor U17905 (N_17905,N_17220,N_16546);
nor U17906 (N_17906,N_16558,N_16262);
and U17907 (N_17907,N_16566,N_16611);
nor U17908 (N_17908,N_16939,N_16355);
and U17909 (N_17909,N_17210,N_16631);
or U17910 (N_17910,N_16539,N_16953);
nor U17911 (N_17911,N_16517,N_16814);
nor U17912 (N_17912,N_17116,N_17139);
xor U17913 (N_17913,N_16455,N_17437);
or U17914 (N_17914,N_16845,N_16550);
nand U17915 (N_17915,N_16452,N_17423);
or U17916 (N_17916,N_17071,N_17145);
and U17917 (N_17917,N_17140,N_16503);
xnor U17918 (N_17918,N_17218,N_16340);
nand U17919 (N_17919,N_16891,N_16971);
and U17920 (N_17920,N_17472,N_16273);
and U17921 (N_17921,N_17311,N_16744);
or U17922 (N_17922,N_16395,N_16960);
nor U17923 (N_17923,N_16353,N_16961);
nor U17924 (N_17924,N_17017,N_17380);
nor U17925 (N_17925,N_16873,N_17189);
nand U17926 (N_17926,N_16444,N_16616);
nand U17927 (N_17927,N_17248,N_16978);
nand U17928 (N_17928,N_16562,N_16594);
xnor U17929 (N_17929,N_16979,N_16410);
or U17930 (N_17930,N_16553,N_16734);
nor U17931 (N_17931,N_16513,N_16747);
xnor U17932 (N_17932,N_17085,N_17239);
nor U17933 (N_17933,N_16735,N_16880);
nand U17934 (N_17934,N_17229,N_16286);
xnor U17935 (N_17935,N_16393,N_16549);
nor U17936 (N_17936,N_16806,N_17301);
nor U17937 (N_17937,N_17272,N_17354);
xnor U17938 (N_17938,N_16629,N_16948);
xnor U17939 (N_17939,N_16280,N_17051);
xnor U17940 (N_17940,N_16293,N_16529);
or U17941 (N_17941,N_16409,N_16476);
nand U17942 (N_17942,N_16839,N_16342);
and U17943 (N_17943,N_16957,N_16311);
xnor U17944 (N_17944,N_16816,N_16538);
nor U17945 (N_17945,N_17327,N_16645);
nor U17946 (N_17946,N_17319,N_16638);
nand U17947 (N_17947,N_16307,N_16904);
xor U17948 (N_17948,N_16592,N_16590);
or U17949 (N_17949,N_16717,N_17242);
xor U17950 (N_17950,N_17257,N_16514);
nor U17951 (N_17951,N_16812,N_16328);
nand U17952 (N_17952,N_16584,N_17285);
or U17953 (N_17953,N_17227,N_17024);
and U17954 (N_17954,N_16857,N_17350);
nand U17955 (N_17955,N_16736,N_16519);
xnor U17956 (N_17956,N_16267,N_16330);
nor U17957 (N_17957,N_16489,N_16813);
nand U17958 (N_17958,N_17477,N_17278);
or U17959 (N_17959,N_17001,N_17497);
nand U17960 (N_17960,N_16667,N_16923);
nor U17961 (N_17961,N_16874,N_16480);
nor U17962 (N_17962,N_16892,N_17077);
or U17963 (N_17963,N_17372,N_17003);
nor U17964 (N_17964,N_16545,N_16445);
nor U17965 (N_17965,N_16609,N_17087);
and U17966 (N_17966,N_17164,N_17481);
xor U17967 (N_17967,N_17100,N_16485);
nor U17968 (N_17968,N_17162,N_17132);
nor U17969 (N_17969,N_17137,N_17403);
xor U17970 (N_17970,N_17342,N_17382);
or U17971 (N_17971,N_16437,N_17129);
or U17972 (N_17972,N_16605,N_16593);
nand U17973 (N_17973,N_17228,N_17231);
or U17974 (N_17974,N_17393,N_17284);
or U17975 (N_17975,N_16833,N_16695);
xor U17976 (N_17976,N_16720,N_16800);
and U17977 (N_17977,N_17197,N_17473);
nand U17978 (N_17978,N_17405,N_17213);
xnor U17979 (N_17979,N_16681,N_16850);
nand U17980 (N_17980,N_17499,N_17012);
xnor U17981 (N_17981,N_17120,N_17258);
xnor U17982 (N_17982,N_16304,N_17106);
xor U17983 (N_17983,N_17095,N_17005);
and U17984 (N_17984,N_16855,N_16516);
nand U17985 (N_17985,N_17026,N_17260);
nand U17986 (N_17986,N_17288,N_16811);
or U17987 (N_17987,N_16682,N_16698);
nand U17988 (N_17988,N_17352,N_16704);
xnor U17989 (N_17989,N_16406,N_16570);
nor U17990 (N_17990,N_16443,N_16958);
nor U17991 (N_17991,N_17234,N_16712);
or U17992 (N_17992,N_16658,N_16435);
nand U17993 (N_17993,N_16357,N_16381);
and U17994 (N_17994,N_16662,N_16557);
nand U17995 (N_17995,N_17038,N_16869);
nor U17996 (N_17996,N_17384,N_16887);
nor U17997 (N_17997,N_17019,N_16899);
xnor U17998 (N_17998,N_16906,N_17163);
nand U17999 (N_17999,N_16624,N_17127);
nor U18000 (N_18000,N_16726,N_16729);
nor U18001 (N_18001,N_16995,N_16559);
and U18002 (N_18002,N_17269,N_16941);
and U18003 (N_18003,N_16926,N_16319);
nor U18004 (N_18004,N_16430,N_16665);
nand U18005 (N_18005,N_16268,N_17464);
xnor U18006 (N_18006,N_17305,N_16844);
and U18007 (N_18007,N_16250,N_16951);
nand U18008 (N_18008,N_16521,N_16898);
or U18009 (N_18009,N_17015,N_16320);
nor U18010 (N_18010,N_16351,N_16375);
and U18011 (N_18011,N_17355,N_16589);
xnor U18012 (N_18012,N_16582,N_16388);
xnor U18013 (N_18013,N_16968,N_17428);
and U18014 (N_18014,N_16620,N_17441);
xnor U18015 (N_18015,N_17373,N_16543);
or U18016 (N_18016,N_16859,N_16252);
and U18017 (N_18017,N_17212,N_16420);
xnor U18018 (N_18018,N_16678,N_16556);
nor U18019 (N_18019,N_16807,N_17086);
and U18020 (N_18020,N_16575,N_17299);
xor U18021 (N_18021,N_16290,N_17262);
or U18022 (N_18022,N_16804,N_17270);
and U18023 (N_18023,N_16677,N_16531);
nand U18024 (N_18024,N_16456,N_16921);
and U18025 (N_18025,N_16371,N_16376);
nand U18026 (N_18026,N_16929,N_17425);
xnor U18027 (N_18027,N_16756,N_16907);
nand U18028 (N_18028,N_17268,N_17365);
nand U18029 (N_18029,N_17108,N_17340);
or U18030 (N_18030,N_17496,N_17451);
or U18031 (N_18031,N_16368,N_16338);
nand U18032 (N_18032,N_16846,N_16298);
or U18033 (N_18033,N_16823,N_16260);
and U18034 (N_18034,N_17265,N_17360);
or U18035 (N_18035,N_17049,N_16392);
xnor U18036 (N_18036,N_16518,N_16721);
and U18037 (N_18037,N_17192,N_17158);
and U18038 (N_18038,N_16974,N_16382);
nand U18039 (N_18039,N_17201,N_16498);
or U18040 (N_18040,N_16599,N_17375);
or U18041 (N_18041,N_17211,N_16454);
and U18042 (N_18042,N_16862,N_16424);
and U18043 (N_18043,N_16936,N_17283);
and U18044 (N_18044,N_17104,N_16731);
xnor U18045 (N_18045,N_16596,N_17328);
nor U18046 (N_18046,N_16802,N_16808);
or U18047 (N_18047,N_17175,N_17018);
and U18048 (N_18048,N_17206,N_16781);
nor U18049 (N_18049,N_16902,N_16661);
and U18050 (N_18050,N_16544,N_16733);
or U18051 (N_18051,N_16940,N_17138);
xor U18052 (N_18052,N_17172,N_17042);
nor U18053 (N_18053,N_16805,N_16396);
nor U18054 (N_18054,N_16724,N_17414);
or U18055 (N_18055,N_17411,N_16994);
nor U18056 (N_18056,N_17446,N_16585);
nand U18057 (N_18057,N_16479,N_16930);
nand U18058 (N_18058,N_17404,N_17426);
xnor U18059 (N_18059,N_16829,N_17320);
nor U18060 (N_18060,N_17381,N_17356);
or U18061 (N_18061,N_17470,N_17107);
nand U18062 (N_18062,N_16742,N_16486);
nor U18063 (N_18063,N_16284,N_16680);
and U18064 (N_18064,N_16689,N_16532);
xor U18065 (N_18065,N_16949,N_16714);
nor U18066 (N_18066,N_17444,N_16842);
nor U18067 (N_18067,N_16441,N_16981);
nand U18068 (N_18068,N_16600,N_16578);
nor U18069 (N_18069,N_16269,N_17207);
and U18070 (N_18070,N_16520,N_17233);
nor U18071 (N_18071,N_17337,N_16495);
nand U18072 (N_18072,N_16527,N_16315);
nand U18073 (N_18073,N_16636,N_16417);
nand U18074 (N_18074,N_17314,N_16255);
and U18075 (N_18075,N_16481,N_17447);
nor U18076 (N_18076,N_17489,N_16446);
and U18077 (N_18077,N_16552,N_16433);
xnor U18078 (N_18078,N_16598,N_16478);
xor U18079 (N_18079,N_17416,N_16997);
nand U18080 (N_18080,N_16983,N_16642);
and U18081 (N_18081,N_16604,N_17492);
and U18082 (N_18082,N_16597,N_17483);
xnor U18083 (N_18083,N_17102,N_16432);
xnor U18084 (N_18084,N_16541,N_16256);
xor U18085 (N_18085,N_17321,N_17277);
or U18086 (N_18086,N_17167,N_16885);
nand U18087 (N_18087,N_17141,N_16512);
or U18088 (N_18088,N_17279,N_17037);
nand U18089 (N_18089,N_16722,N_17010);
or U18090 (N_18090,N_16746,N_17357);
nand U18091 (N_18091,N_16920,N_17181);
and U18092 (N_18092,N_16419,N_16686);
and U18093 (N_18093,N_17467,N_17351);
or U18094 (N_18094,N_16928,N_17322);
nand U18095 (N_18095,N_17009,N_16674);
nand U18096 (N_18096,N_17074,N_16649);
nor U18097 (N_18097,N_16675,N_17339);
nand U18098 (N_18098,N_17027,N_16301);
and U18099 (N_18099,N_16331,N_16784);
nand U18100 (N_18100,N_17202,N_16737);
nand U18101 (N_18101,N_17303,N_16383);
xor U18102 (N_18102,N_16471,N_16705);
nand U18103 (N_18103,N_17096,N_16764);
and U18104 (N_18104,N_16918,N_17468);
nor U18105 (N_18105,N_16795,N_17091);
nand U18106 (N_18106,N_16718,N_16251);
xnor U18107 (N_18107,N_16749,N_16491);
nor U18108 (N_18108,N_16555,N_17332);
and U18109 (N_18109,N_16934,N_16864);
xor U18110 (N_18110,N_16653,N_17454);
nand U18111 (N_18111,N_17313,N_16253);
or U18112 (N_18112,N_16970,N_17286);
xor U18113 (N_18113,N_16421,N_16439);
or U18114 (N_18114,N_16451,N_17398);
or U18115 (N_18115,N_17377,N_17008);
xor U18116 (N_18116,N_17490,N_17487);
or U18117 (N_18117,N_16824,N_17456);
nor U18118 (N_18118,N_16699,N_16574);
nor U18119 (N_18119,N_16919,N_17075);
nand U18120 (N_18120,N_17184,N_17040);
and U18121 (N_18121,N_17378,N_16822);
nor U18122 (N_18122,N_17395,N_17296);
or U18123 (N_18123,N_16617,N_16707);
or U18124 (N_18124,N_16817,N_16840);
nor U18125 (N_18125,N_16327,N_17106);
nand U18126 (N_18126,N_17145,N_16558);
or U18127 (N_18127,N_16981,N_17347);
nand U18128 (N_18128,N_17362,N_16787);
or U18129 (N_18129,N_17342,N_16438);
nor U18130 (N_18130,N_16674,N_17265);
xnor U18131 (N_18131,N_17233,N_16898);
nand U18132 (N_18132,N_17006,N_16707);
or U18133 (N_18133,N_16381,N_16500);
nor U18134 (N_18134,N_16481,N_17341);
nand U18135 (N_18135,N_16287,N_16686);
or U18136 (N_18136,N_16352,N_16620);
xor U18137 (N_18137,N_16730,N_16654);
nand U18138 (N_18138,N_16765,N_16602);
xor U18139 (N_18139,N_16680,N_17412);
and U18140 (N_18140,N_16676,N_17437);
or U18141 (N_18141,N_17185,N_16796);
and U18142 (N_18142,N_16685,N_17195);
xnor U18143 (N_18143,N_16984,N_17065);
and U18144 (N_18144,N_16359,N_17120);
or U18145 (N_18145,N_17400,N_16551);
xnor U18146 (N_18146,N_16790,N_17127);
nand U18147 (N_18147,N_16815,N_16705);
and U18148 (N_18148,N_16971,N_17005);
and U18149 (N_18149,N_17100,N_17380);
nor U18150 (N_18150,N_17366,N_16301);
xor U18151 (N_18151,N_17431,N_16532);
and U18152 (N_18152,N_16800,N_17381);
nand U18153 (N_18153,N_16500,N_16593);
or U18154 (N_18154,N_16813,N_17429);
xor U18155 (N_18155,N_17111,N_16491);
nor U18156 (N_18156,N_16701,N_16750);
nand U18157 (N_18157,N_16346,N_17296);
and U18158 (N_18158,N_17354,N_17313);
nand U18159 (N_18159,N_17090,N_17445);
xnor U18160 (N_18160,N_17400,N_17149);
and U18161 (N_18161,N_17433,N_16314);
xor U18162 (N_18162,N_17304,N_16822);
nor U18163 (N_18163,N_16766,N_17001);
xor U18164 (N_18164,N_16755,N_16341);
or U18165 (N_18165,N_17175,N_16359);
nor U18166 (N_18166,N_16903,N_17051);
nor U18167 (N_18167,N_16267,N_17267);
or U18168 (N_18168,N_16448,N_16339);
or U18169 (N_18169,N_17316,N_17444);
nand U18170 (N_18170,N_17440,N_17012);
xor U18171 (N_18171,N_17318,N_16864);
xor U18172 (N_18172,N_16708,N_16646);
and U18173 (N_18173,N_17454,N_16253);
and U18174 (N_18174,N_16515,N_17032);
nand U18175 (N_18175,N_17208,N_17089);
nand U18176 (N_18176,N_16953,N_17479);
or U18177 (N_18177,N_16733,N_16798);
or U18178 (N_18178,N_16318,N_16754);
nand U18179 (N_18179,N_17367,N_16892);
nand U18180 (N_18180,N_17405,N_16627);
nor U18181 (N_18181,N_16624,N_16379);
nor U18182 (N_18182,N_17130,N_17296);
nor U18183 (N_18183,N_17264,N_16322);
xor U18184 (N_18184,N_17222,N_16589);
and U18185 (N_18185,N_16353,N_17335);
xnor U18186 (N_18186,N_17088,N_16357);
and U18187 (N_18187,N_17274,N_17028);
nand U18188 (N_18188,N_17334,N_16943);
nor U18189 (N_18189,N_16784,N_16574);
xor U18190 (N_18190,N_16560,N_16626);
nand U18191 (N_18191,N_17397,N_16723);
and U18192 (N_18192,N_16775,N_16930);
and U18193 (N_18193,N_17196,N_16354);
nand U18194 (N_18194,N_16975,N_16892);
and U18195 (N_18195,N_17169,N_16762);
or U18196 (N_18196,N_17111,N_17329);
nor U18197 (N_18197,N_16538,N_16443);
or U18198 (N_18198,N_17160,N_17326);
xnor U18199 (N_18199,N_16375,N_17197);
or U18200 (N_18200,N_17125,N_16912);
nor U18201 (N_18201,N_16483,N_17020);
xor U18202 (N_18202,N_17196,N_16349);
and U18203 (N_18203,N_16797,N_17106);
xnor U18204 (N_18204,N_17414,N_16723);
nand U18205 (N_18205,N_17418,N_16828);
nor U18206 (N_18206,N_17354,N_16481);
xnor U18207 (N_18207,N_16572,N_16383);
and U18208 (N_18208,N_17326,N_16485);
or U18209 (N_18209,N_17261,N_16818);
nor U18210 (N_18210,N_16391,N_16707);
or U18211 (N_18211,N_16730,N_16438);
nand U18212 (N_18212,N_16297,N_17496);
nor U18213 (N_18213,N_17281,N_16601);
xor U18214 (N_18214,N_17044,N_16489);
nand U18215 (N_18215,N_17418,N_16357);
xnor U18216 (N_18216,N_17371,N_17006);
nor U18217 (N_18217,N_17153,N_17254);
nor U18218 (N_18218,N_17111,N_16981);
or U18219 (N_18219,N_17466,N_16674);
nand U18220 (N_18220,N_16376,N_16777);
nor U18221 (N_18221,N_16873,N_16407);
nor U18222 (N_18222,N_16266,N_17306);
and U18223 (N_18223,N_16523,N_17029);
nand U18224 (N_18224,N_16918,N_16706);
or U18225 (N_18225,N_16327,N_16719);
xnor U18226 (N_18226,N_17371,N_17308);
nand U18227 (N_18227,N_17105,N_16318);
xnor U18228 (N_18228,N_16670,N_16818);
nand U18229 (N_18229,N_16337,N_16787);
nor U18230 (N_18230,N_17086,N_16638);
nand U18231 (N_18231,N_17371,N_16298);
nand U18232 (N_18232,N_16819,N_17063);
or U18233 (N_18233,N_17266,N_16604);
xor U18234 (N_18234,N_16368,N_16726);
nor U18235 (N_18235,N_17435,N_16805);
and U18236 (N_18236,N_16681,N_16466);
or U18237 (N_18237,N_16415,N_16948);
nand U18238 (N_18238,N_16748,N_17374);
nor U18239 (N_18239,N_16266,N_16864);
xor U18240 (N_18240,N_16534,N_17431);
nor U18241 (N_18241,N_16701,N_16575);
nor U18242 (N_18242,N_16469,N_16506);
nor U18243 (N_18243,N_16310,N_17433);
nor U18244 (N_18244,N_16286,N_16913);
and U18245 (N_18245,N_16563,N_16456);
nand U18246 (N_18246,N_17246,N_16326);
or U18247 (N_18247,N_17437,N_17355);
nor U18248 (N_18248,N_16668,N_17380);
xnor U18249 (N_18249,N_16276,N_16537);
or U18250 (N_18250,N_16748,N_17137);
nand U18251 (N_18251,N_16839,N_17281);
and U18252 (N_18252,N_17106,N_16425);
nor U18253 (N_18253,N_16887,N_17170);
and U18254 (N_18254,N_16940,N_17131);
or U18255 (N_18255,N_17076,N_16960);
xor U18256 (N_18256,N_16421,N_16967);
nand U18257 (N_18257,N_17209,N_17212);
and U18258 (N_18258,N_16928,N_16268);
and U18259 (N_18259,N_16343,N_17316);
xor U18260 (N_18260,N_16439,N_17441);
or U18261 (N_18261,N_16303,N_16988);
nor U18262 (N_18262,N_16526,N_16815);
xor U18263 (N_18263,N_16309,N_16708);
and U18264 (N_18264,N_16801,N_16298);
xor U18265 (N_18265,N_17210,N_17365);
xor U18266 (N_18266,N_17050,N_16550);
and U18267 (N_18267,N_16667,N_16991);
nand U18268 (N_18268,N_17058,N_16520);
xor U18269 (N_18269,N_17114,N_17428);
nand U18270 (N_18270,N_17254,N_16547);
xnor U18271 (N_18271,N_16725,N_16724);
xnor U18272 (N_18272,N_16763,N_17405);
xor U18273 (N_18273,N_17241,N_16741);
nor U18274 (N_18274,N_16745,N_17367);
nand U18275 (N_18275,N_17471,N_16261);
and U18276 (N_18276,N_16812,N_16708);
nand U18277 (N_18277,N_16814,N_17364);
nand U18278 (N_18278,N_17012,N_16723);
and U18279 (N_18279,N_17248,N_17204);
xnor U18280 (N_18280,N_17105,N_16709);
xnor U18281 (N_18281,N_16676,N_16987);
nor U18282 (N_18282,N_16432,N_17439);
and U18283 (N_18283,N_16322,N_16843);
nor U18284 (N_18284,N_16384,N_17257);
or U18285 (N_18285,N_16950,N_17354);
or U18286 (N_18286,N_16922,N_17381);
xor U18287 (N_18287,N_17397,N_16713);
xor U18288 (N_18288,N_16960,N_16604);
nand U18289 (N_18289,N_16438,N_16903);
or U18290 (N_18290,N_16955,N_16920);
xnor U18291 (N_18291,N_17152,N_17190);
or U18292 (N_18292,N_17091,N_16262);
xnor U18293 (N_18293,N_16529,N_16857);
nand U18294 (N_18294,N_16295,N_16282);
nand U18295 (N_18295,N_16491,N_17401);
and U18296 (N_18296,N_16274,N_17027);
nand U18297 (N_18297,N_16269,N_16302);
nor U18298 (N_18298,N_17399,N_16393);
or U18299 (N_18299,N_16810,N_16589);
or U18300 (N_18300,N_17259,N_16798);
or U18301 (N_18301,N_17239,N_16294);
or U18302 (N_18302,N_16843,N_16439);
or U18303 (N_18303,N_17040,N_17272);
or U18304 (N_18304,N_17396,N_16919);
and U18305 (N_18305,N_16599,N_17040);
or U18306 (N_18306,N_16587,N_16811);
nand U18307 (N_18307,N_16607,N_16735);
xor U18308 (N_18308,N_16960,N_17381);
or U18309 (N_18309,N_17195,N_16720);
or U18310 (N_18310,N_17203,N_17109);
xor U18311 (N_18311,N_16571,N_16959);
nor U18312 (N_18312,N_16291,N_17090);
or U18313 (N_18313,N_17331,N_17461);
xnor U18314 (N_18314,N_16874,N_16674);
nand U18315 (N_18315,N_16386,N_16289);
or U18316 (N_18316,N_16831,N_16567);
nand U18317 (N_18317,N_17218,N_16571);
xor U18318 (N_18318,N_17310,N_17322);
xor U18319 (N_18319,N_17488,N_16349);
xor U18320 (N_18320,N_16712,N_17477);
and U18321 (N_18321,N_16909,N_16504);
nor U18322 (N_18322,N_17261,N_16665);
nor U18323 (N_18323,N_17081,N_16458);
xor U18324 (N_18324,N_17453,N_17038);
or U18325 (N_18325,N_17064,N_16927);
nor U18326 (N_18326,N_17376,N_17391);
and U18327 (N_18327,N_17302,N_17128);
and U18328 (N_18328,N_17405,N_17134);
or U18329 (N_18329,N_17161,N_16763);
and U18330 (N_18330,N_16759,N_17403);
nor U18331 (N_18331,N_16510,N_17364);
or U18332 (N_18332,N_16820,N_17175);
nor U18333 (N_18333,N_16549,N_16724);
and U18334 (N_18334,N_17082,N_16287);
xnor U18335 (N_18335,N_16927,N_16640);
nor U18336 (N_18336,N_16558,N_17074);
xnor U18337 (N_18337,N_16306,N_17301);
nand U18338 (N_18338,N_17427,N_16520);
xnor U18339 (N_18339,N_16517,N_16699);
and U18340 (N_18340,N_16334,N_16840);
nor U18341 (N_18341,N_17428,N_17090);
xnor U18342 (N_18342,N_17255,N_16499);
or U18343 (N_18343,N_16600,N_17298);
and U18344 (N_18344,N_17403,N_17462);
and U18345 (N_18345,N_16409,N_16952);
nor U18346 (N_18346,N_16948,N_17283);
and U18347 (N_18347,N_17136,N_16670);
or U18348 (N_18348,N_16851,N_16771);
xor U18349 (N_18349,N_17421,N_16439);
nand U18350 (N_18350,N_16408,N_17147);
xnor U18351 (N_18351,N_16364,N_17099);
nand U18352 (N_18352,N_17493,N_16414);
and U18353 (N_18353,N_16482,N_17362);
nor U18354 (N_18354,N_17124,N_16644);
nand U18355 (N_18355,N_17375,N_16633);
nor U18356 (N_18356,N_16512,N_17451);
and U18357 (N_18357,N_16781,N_16883);
nand U18358 (N_18358,N_17251,N_16377);
and U18359 (N_18359,N_17141,N_17002);
nor U18360 (N_18360,N_16472,N_17470);
xor U18361 (N_18361,N_17486,N_16534);
or U18362 (N_18362,N_16253,N_17180);
and U18363 (N_18363,N_17345,N_17125);
and U18364 (N_18364,N_16826,N_17347);
and U18365 (N_18365,N_16944,N_16397);
xnor U18366 (N_18366,N_17423,N_17264);
or U18367 (N_18367,N_16490,N_17452);
nor U18368 (N_18368,N_16967,N_16560);
xnor U18369 (N_18369,N_16541,N_16388);
xor U18370 (N_18370,N_16418,N_17038);
or U18371 (N_18371,N_16327,N_16767);
and U18372 (N_18372,N_17274,N_16742);
nor U18373 (N_18373,N_16362,N_16405);
xor U18374 (N_18374,N_16348,N_16485);
nor U18375 (N_18375,N_16692,N_16995);
nand U18376 (N_18376,N_16312,N_16273);
or U18377 (N_18377,N_16861,N_16969);
nor U18378 (N_18378,N_16640,N_17223);
or U18379 (N_18379,N_16799,N_17476);
nand U18380 (N_18380,N_17334,N_16599);
and U18381 (N_18381,N_17381,N_17075);
nand U18382 (N_18382,N_16907,N_17274);
nor U18383 (N_18383,N_17296,N_16553);
xor U18384 (N_18384,N_16647,N_17347);
nand U18385 (N_18385,N_17106,N_17224);
or U18386 (N_18386,N_16766,N_16443);
xor U18387 (N_18387,N_16348,N_16351);
nand U18388 (N_18388,N_16330,N_17108);
xor U18389 (N_18389,N_17430,N_17145);
xor U18390 (N_18390,N_16412,N_16705);
or U18391 (N_18391,N_17057,N_16599);
or U18392 (N_18392,N_17059,N_16911);
and U18393 (N_18393,N_17209,N_17411);
nor U18394 (N_18394,N_17441,N_17056);
nor U18395 (N_18395,N_16692,N_16893);
xnor U18396 (N_18396,N_17161,N_17046);
xor U18397 (N_18397,N_16397,N_16615);
nor U18398 (N_18398,N_16710,N_17426);
or U18399 (N_18399,N_17353,N_17419);
xor U18400 (N_18400,N_17338,N_16308);
and U18401 (N_18401,N_16978,N_17283);
or U18402 (N_18402,N_17160,N_16490);
or U18403 (N_18403,N_17392,N_17102);
xnor U18404 (N_18404,N_17260,N_17313);
xnor U18405 (N_18405,N_16949,N_16703);
nand U18406 (N_18406,N_17367,N_17023);
nand U18407 (N_18407,N_16712,N_16601);
xnor U18408 (N_18408,N_16867,N_16647);
nor U18409 (N_18409,N_16343,N_16652);
nand U18410 (N_18410,N_16337,N_16807);
nor U18411 (N_18411,N_17103,N_16727);
nand U18412 (N_18412,N_16585,N_16916);
and U18413 (N_18413,N_16486,N_17365);
nand U18414 (N_18414,N_17205,N_17058);
nor U18415 (N_18415,N_16618,N_17070);
and U18416 (N_18416,N_16510,N_16298);
and U18417 (N_18417,N_16355,N_16365);
xnor U18418 (N_18418,N_16893,N_16310);
nand U18419 (N_18419,N_17042,N_17226);
or U18420 (N_18420,N_16547,N_16516);
and U18421 (N_18421,N_17142,N_17034);
or U18422 (N_18422,N_17137,N_16989);
or U18423 (N_18423,N_17495,N_16992);
and U18424 (N_18424,N_16396,N_17119);
nand U18425 (N_18425,N_17457,N_16535);
and U18426 (N_18426,N_17446,N_17172);
xor U18427 (N_18427,N_17302,N_16983);
xnor U18428 (N_18428,N_17254,N_17148);
nand U18429 (N_18429,N_16645,N_17034);
or U18430 (N_18430,N_17045,N_16764);
xor U18431 (N_18431,N_16965,N_17201);
nor U18432 (N_18432,N_17413,N_17084);
or U18433 (N_18433,N_16638,N_16331);
xnor U18434 (N_18434,N_16958,N_17474);
nor U18435 (N_18435,N_16752,N_16755);
nand U18436 (N_18436,N_16569,N_17335);
or U18437 (N_18437,N_17206,N_16267);
xor U18438 (N_18438,N_17112,N_16613);
nand U18439 (N_18439,N_16611,N_16436);
nand U18440 (N_18440,N_16552,N_16891);
or U18441 (N_18441,N_16947,N_16757);
nand U18442 (N_18442,N_17115,N_16907);
and U18443 (N_18443,N_17285,N_16263);
nor U18444 (N_18444,N_16699,N_16391);
and U18445 (N_18445,N_16790,N_17072);
and U18446 (N_18446,N_16601,N_16390);
nor U18447 (N_18447,N_16460,N_17090);
nand U18448 (N_18448,N_17302,N_17122);
or U18449 (N_18449,N_16321,N_16336);
nand U18450 (N_18450,N_17493,N_17477);
and U18451 (N_18451,N_16856,N_17151);
xnor U18452 (N_18452,N_16642,N_17302);
nor U18453 (N_18453,N_17006,N_16831);
nand U18454 (N_18454,N_16485,N_17019);
nand U18455 (N_18455,N_16769,N_17018);
xor U18456 (N_18456,N_16263,N_16418);
and U18457 (N_18457,N_16508,N_16648);
xor U18458 (N_18458,N_17411,N_16258);
nor U18459 (N_18459,N_17106,N_17044);
nand U18460 (N_18460,N_17078,N_17277);
nor U18461 (N_18461,N_17360,N_16546);
or U18462 (N_18462,N_17196,N_16934);
nor U18463 (N_18463,N_16453,N_16640);
xor U18464 (N_18464,N_17128,N_17371);
and U18465 (N_18465,N_16590,N_16259);
nand U18466 (N_18466,N_16613,N_17045);
or U18467 (N_18467,N_16420,N_17356);
xnor U18468 (N_18468,N_16975,N_16971);
nand U18469 (N_18469,N_16934,N_16781);
nand U18470 (N_18470,N_16750,N_16608);
or U18471 (N_18471,N_17360,N_17132);
and U18472 (N_18472,N_16690,N_17069);
and U18473 (N_18473,N_16729,N_16945);
xnor U18474 (N_18474,N_16547,N_17438);
xor U18475 (N_18475,N_16830,N_17479);
and U18476 (N_18476,N_16629,N_16536);
xnor U18477 (N_18477,N_17075,N_16626);
nor U18478 (N_18478,N_17426,N_17083);
nand U18479 (N_18479,N_16888,N_17388);
and U18480 (N_18480,N_16822,N_17490);
nor U18481 (N_18481,N_17266,N_17376);
nor U18482 (N_18482,N_16998,N_16984);
or U18483 (N_18483,N_16672,N_16911);
or U18484 (N_18484,N_17359,N_16846);
nand U18485 (N_18485,N_16662,N_16709);
xor U18486 (N_18486,N_17441,N_16391);
xor U18487 (N_18487,N_16680,N_16407);
nor U18488 (N_18488,N_16960,N_16404);
nand U18489 (N_18489,N_16770,N_16916);
xor U18490 (N_18490,N_17302,N_17307);
nor U18491 (N_18491,N_17191,N_16480);
nor U18492 (N_18492,N_17120,N_16406);
and U18493 (N_18493,N_17141,N_16603);
nor U18494 (N_18494,N_16563,N_17060);
or U18495 (N_18495,N_17365,N_16427);
xor U18496 (N_18496,N_16753,N_17340);
xnor U18497 (N_18497,N_17467,N_16813);
and U18498 (N_18498,N_16908,N_17336);
nand U18499 (N_18499,N_17360,N_16843);
xnor U18500 (N_18500,N_16975,N_16554);
and U18501 (N_18501,N_17086,N_16318);
and U18502 (N_18502,N_16802,N_16832);
or U18503 (N_18503,N_16414,N_17069);
nand U18504 (N_18504,N_17484,N_16925);
or U18505 (N_18505,N_16778,N_16908);
or U18506 (N_18506,N_16416,N_16470);
nor U18507 (N_18507,N_16761,N_17475);
nand U18508 (N_18508,N_16488,N_16882);
xnor U18509 (N_18509,N_16628,N_16354);
and U18510 (N_18510,N_17031,N_16444);
xor U18511 (N_18511,N_16856,N_16540);
nand U18512 (N_18512,N_16635,N_16960);
and U18513 (N_18513,N_16386,N_16667);
xor U18514 (N_18514,N_16764,N_16894);
nor U18515 (N_18515,N_17213,N_17475);
nor U18516 (N_18516,N_17107,N_17099);
and U18517 (N_18517,N_16796,N_16323);
nor U18518 (N_18518,N_16492,N_16266);
nand U18519 (N_18519,N_16795,N_16454);
and U18520 (N_18520,N_16937,N_17179);
nor U18521 (N_18521,N_17466,N_16624);
nand U18522 (N_18522,N_16939,N_16445);
nor U18523 (N_18523,N_17300,N_17067);
or U18524 (N_18524,N_17239,N_17207);
and U18525 (N_18525,N_16889,N_16950);
nor U18526 (N_18526,N_16448,N_16436);
nand U18527 (N_18527,N_17305,N_17441);
or U18528 (N_18528,N_16949,N_17159);
nand U18529 (N_18529,N_16878,N_17288);
nor U18530 (N_18530,N_16861,N_17191);
or U18531 (N_18531,N_16687,N_17226);
or U18532 (N_18532,N_17280,N_17456);
nor U18533 (N_18533,N_16297,N_17452);
nand U18534 (N_18534,N_16661,N_16913);
and U18535 (N_18535,N_17002,N_16380);
xor U18536 (N_18536,N_17044,N_17043);
nor U18537 (N_18537,N_16251,N_16254);
nor U18538 (N_18538,N_17265,N_17221);
nand U18539 (N_18539,N_16788,N_17188);
nor U18540 (N_18540,N_16722,N_17416);
xor U18541 (N_18541,N_16643,N_16740);
nand U18542 (N_18542,N_17209,N_17254);
and U18543 (N_18543,N_16586,N_16317);
nand U18544 (N_18544,N_16482,N_16826);
nor U18545 (N_18545,N_17323,N_16660);
and U18546 (N_18546,N_17051,N_16379);
nor U18547 (N_18547,N_17370,N_16759);
and U18548 (N_18548,N_16687,N_16790);
nand U18549 (N_18549,N_16337,N_16881);
xor U18550 (N_18550,N_16467,N_17382);
xor U18551 (N_18551,N_16937,N_16450);
xnor U18552 (N_18552,N_17001,N_16742);
xnor U18553 (N_18553,N_17263,N_16811);
nand U18554 (N_18554,N_16462,N_16273);
or U18555 (N_18555,N_16996,N_16890);
nor U18556 (N_18556,N_17124,N_16380);
nand U18557 (N_18557,N_16910,N_17448);
or U18558 (N_18558,N_17337,N_16651);
or U18559 (N_18559,N_16338,N_16790);
xor U18560 (N_18560,N_16674,N_17116);
or U18561 (N_18561,N_16735,N_17007);
nor U18562 (N_18562,N_16334,N_16701);
nor U18563 (N_18563,N_17103,N_16470);
or U18564 (N_18564,N_16299,N_16520);
nand U18565 (N_18565,N_17044,N_16513);
nor U18566 (N_18566,N_17081,N_17074);
xor U18567 (N_18567,N_17454,N_16430);
nor U18568 (N_18568,N_16937,N_17093);
xor U18569 (N_18569,N_17194,N_17346);
and U18570 (N_18570,N_16759,N_16722);
nor U18571 (N_18571,N_16890,N_16572);
nand U18572 (N_18572,N_16843,N_16735);
and U18573 (N_18573,N_16705,N_17175);
and U18574 (N_18574,N_17253,N_16450);
nand U18575 (N_18575,N_16855,N_16761);
and U18576 (N_18576,N_16323,N_16908);
nor U18577 (N_18577,N_16514,N_17147);
or U18578 (N_18578,N_16612,N_16591);
and U18579 (N_18579,N_16456,N_17436);
xor U18580 (N_18580,N_16862,N_16568);
and U18581 (N_18581,N_17413,N_16494);
and U18582 (N_18582,N_17440,N_17161);
or U18583 (N_18583,N_17051,N_16985);
and U18584 (N_18584,N_16505,N_16304);
nor U18585 (N_18585,N_16258,N_17399);
nor U18586 (N_18586,N_16403,N_17419);
nor U18587 (N_18587,N_16404,N_16746);
and U18588 (N_18588,N_16850,N_17207);
nand U18589 (N_18589,N_16515,N_16451);
xor U18590 (N_18590,N_17320,N_17128);
nand U18591 (N_18591,N_16716,N_16929);
nand U18592 (N_18592,N_17279,N_16346);
nor U18593 (N_18593,N_17448,N_16766);
nand U18594 (N_18594,N_16338,N_16729);
or U18595 (N_18595,N_16513,N_17060);
nor U18596 (N_18596,N_16322,N_16520);
nor U18597 (N_18597,N_16544,N_16663);
nand U18598 (N_18598,N_17429,N_17396);
and U18599 (N_18599,N_16674,N_17289);
nand U18600 (N_18600,N_17139,N_17287);
nor U18601 (N_18601,N_16467,N_16440);
nand U18602 (N_18602,N_16959,N_17354);
xnor U18603 (N_18603,N_16664,N_16558);
xnor U18604 (N_18604,N_16992,N_16572);
nand U18605 (N_18605,N_17104,N_16258);
xnor U18606 (N_18606,N_17442,N_16277);
xnor U18607 (N_18607,N_16274,N_16865);
xnor U18608 (N_18608,N_16980,N_17053);
nor U18609 (N_18609,N_16329,N_16749);
nor U18610 (N_18610,N_17406,N_16300);
or U18611 (N_18611,N_17134,N_16813);
xnor U18612 (N_18612,N_17305,N_17358);
xnor U18613 (N_18613,N_17387,N_16744);
or U18614 (N_18614,N_17053,N_17062);
xor U18615 (N_18615,N_17033,N_16434);
nand U18616 (N_18616,N_17425,N_16796);
nand U18617 (N_18617,N_17058,N_16350);
and U18618 (N_18618,N_16828,N_16267);
nand U18619 (N_18619,N_16484,N_16545);
xnor U18620 (N_18620,N_16745,N_16592);
xor U18621 (N_18621,N_16462,N_16560);
and U18622 (N_18622,N_16919,N_17186);
or U18623 (N_18623,N_16420,N_16336);
nand U18624 (N_18624,N_17430,N_17380);
nand U18625 (N_18625,N_17379,N_16558);
nor U18626 (N_18626,N_16641,N_16705);
nor U18627 (N_18627,N_16337,N_16948);
and U18628 (N_18628,N_16900,N_16419);
or U18629 (N_18629,N_17178,N_16726);
xor U18630 (N_18630,N_17094,N_17099);
nor U18631 (N_18631,N_17059,N_16313);
and U18632 (N_18632,N_16316,N_16829);
xnor U18633 (N_18633,N_16585,N_16484);
nor U18634 (N_18634,N_17265,N_16882);
or U18635 (N_18635,N_16962,N_16687);
nor U18636 (N_18636,N_17289,N_16270);
nand U18637 (N_18637,N_16880,N_17316);
and U18638 (N_18638,N_16946,N_16350);
nor U18639 (N_18639,N_16555,N_16576);
or U18640 (N_18640,N_16463,N_16497);
and U18641 (N_18641,N_17134,N_16837);
nand U18642 (N_18642,N_16622,N_16623);
or U18643 (N_18643,N_16977,N_16845);
xnor U18644 (N_18644,N_16947,N_16421);
or U18645 (N_18645,N_16385,N_16257);
xor U18646 (N_18646,N_17483,N_16394);
or U18647 (N_18647,N_16590,N_17320);
xor U18648 (N_18648,N_17239,N_16661);
and U18649 (N_18649,N_17353,N_17374);
nand U18650 (N_18650,N_17183,N_17156);
nor U18651 (N_18651,N_16708,N_16905);
xor U18652 (N_18652,N_16350,N_16766);
nor U18653 (N_18653,N_16733,N_16370);
nand U18654 (N_18654,N_16747,N_17480);
nand U18655 (N_18655,N_17459,N_17072);
and U18656 (N_18656,N_16628,N_17056);
nor U18657 (N_18657,N_16386,N_16854);
nor U18658 (N_18658,N_17348,N_16518);
nor U18659 (N_18659,N_16913,N_16700);
xor U18660 (N_18660,N_17030,N_17456);
nor U18661 (N_18661,N_16955,N_16622);
and U18662 (N_18662,N_17363,N_16740);
and U18663 (N_18663,N_17357,N_17396);
or U18664 (N_18664,N_16529,N_17391);
nand U18665 (N_18665,N_16626,N_17286);
nand U18666 (N_18666,N_16312,N_16332);
and U18667 (N_18667,N_16977,N_17462);
nor U18668 (N_18668,N_16833,N_16787);
nor U18669 (N_18669,N_16380,N_16931);
and U18670 (N_18670,N_17141,N_16852);
and U18671 (N_18671,N_16473,N_17332);
nor U18672 (N_18672,N_16939,N_17068);
or U18673 (N_18673,N_16435,N_16973);
nor U18674 (N_18674,N_16678,N_16411);
xor U18675 (N_18675,N_17161,N_16977);
and U18676 (N_18676,N_16453,N_17279);
nand U18677 (N_18677,N_17000,N_17394);
nand U18678 (N_18678,N_17010,N_16570);
or U18679 (N_18679,N_16623,N_16510);
and U18680 (N_18680,N_16402,N_16588);
xor U18681 (N_18681,N_17006,N_17218);
xnor U18682 (N_18682,N_17145,N_16704);
or U18683 (N_18683,N_16934,N_16914);
xor U18684 (N_18684,N_16857,N_17210);
or U18685 (N_18685,N_16251,N_16388);
xor U18686 (N_18686,N_17352,N_16974);
xnor U18687 (N_18687,N_17235,N_16326);
xnor U18688 (N_18688,N_16566,N_17461);
xor U18689 (N_18689,N_17481,N_16621);
or U18690 (N_18690,N_17069,N_16911);
or U18691 (N_18691,N_16618,N_16372);
nor U18692 (N_18692,N_17175,N_16281);
nor U18693 (N_18693,N_17390,N_17225);
nand U18694 (N_18694,N_17199,N_17409);
or U18695 (N_18695,N_16663,N_16913);
or U18696 (N_18696,N_17026,N_17484);
nand U18697 (N_18697,N_17049,N_16255);
or U18698 (N_18698,N_16260,N_17265);
nand U18699 (N_18699,N_17457,N_16701);
or U18700 (N_18700,N_17034,N_17013);
nand U18701 (N_18701,N_17117,N_17449);
and U18702 (N_18702,N_16459,N_16743);
nand U18703 (N_18703,N_17219,N_17353);
and U18704 (N_18704,N_17093,N_17279);
xor U18705 (N_18705,N_16898,N_16766);
nor U18706 (N_18706,N_16729,N_16649);
xor U18707 (N_18707,N_17235,N_16896);
and U18708 (N_18708,N_16388,N_17188);
or U18709 (N_18709,N_16593,N_17099);
nor U18710 (N_18710,N_16929,N_17494);
and U18711 (N_18711,N_17147,N_17326);
nand U18712 (N_18712,N_17437,N_16634);
or U18713 (N_18713,N_16834,N_16395);
and U18714 (N_18714,N_16531,N_16635);
xor U18715 (N_18715,N_16784,N_17496);
nor U18716 (N_18716,N_16690,N_16372);
nand U18717 (N_18717,N_17499,N_17233);
and U18718 (N_18718,N_17277,N_16623);
nand U18719 (N_18719,N_17319,N_17051);
and U18720 (N_18720,N_16611,N_16876);
or U18721 (N_18721,N_17162,N_16713);
and U18722 (N_18722,N_16440,N_16989);
nand U18723 (N_18723,N_17455,N_17421);
nand U18724 (N_18724,N_17383,N_16886);
or U18725 (N_18725,N_16855,N_16682);
xnor U18726 (N_18726,N_17140,N_17166);
or U18727 (N_18727,N_16550,N_17106);
nor U18728 (N_18728,N_16641,N_16567);
nor U18729 (N_18729,N_16466,N_16514);
xnor U18730 (N_18730,N_17105,N_17310);
nor U18731 (N_18731,N_17350,N_17132);
nand U18732 (N_18732,N_17469,N_16744);
and U18733 (N_18733,N_17457,N_16988);
nand U18734 (N_18734,N_16668,N_16394);
and U18735 (N_18735,N_16994,N_17285);
xnor U18736 (N_18736,N_16899,N_16722);
nand U18737 (N_18737,N_16343,N_17348);
and U18738 (N_18738,N_16752,N_17099);
xor U18739 (N_18739,N_17118,N_17062);
nor U18740 (N_18740,N_16755,N_17117);
nor U18741 (N_18741,N_16751,N_16652);
nor U18742 (N_18742,N_17029,N_17410);
and U18743 (N_18743,N_16657,N_17304);
xnor U18744 (N_18744,N_16895,N_17431);
nor U18745 (N_18745,N_17304,N_16353);
xnor U18746 (N_18746,N_17236,N_16530);
xnor U18747 (N_18747,N_16470,N_16512);
nor U18748 (N_18748,N_16521,N_16817);
nand U18749 (N_18749,N_16689,N_16253);
nor U18750 (N_18750,N_18464,N_18007);
or U18751 (N_18751,N_18140,N_18501);
or U18752 (N_18752,N_17635,N_18317);
and U18753 (N_18753,N_18193,N_18234);
or U18754 (N_18754,N_18264,N_17680);
and U18755 (N_18755,N_18242,N_17810);
nor U18756 (N_18756,N_17505,N_18456);
and U18757 (N_18757,N_18228,N_17684);
and U18758 (N_18758,N_17817,N_17881);
xnor U18759 (N_18759,N_18164,N_18408);
xnor U18760 (N_18760,N_18575,N_18612);
and U18761 (N_18761,N_17794,N_17627);
or U18762 (N_18762,N_18025,N_17690);
or U18763 (N_18763,N_18513,N_17622);
and U18764 (N_18764,N_18411,N_18555);
and U18765 (N_18765,N_18515,N_18433);
nor U18766 (N_18766,N_18064,N_18202);
nor U18767 (N_18767,N_17616,N_17509);
or U18768 (N_18768,N_18271,N_17702);
or U18769 (N_18769,N_17954,N_18578);
nor U18770 (N_18770,N_17758,N_18167);
and U18771 (N_18771,N_18090,N_18546);
nand U18772 (N_18772,N_17695,N_17527);
nand U18773 (N_18773,N_17503,N_17745);
or U18774 (N_18774,N_17528,N_18061);
and U18775 (N_18775,N_17538,N_18142);
nand U18776 (N_18776,N_18582,N_18051);
nor U18777 (N_18777,N_17923,N_17928);
nor U18778 (N_18778,N_18650,N_18223);
or U18779 (N_18779,N_17589,N_17671);
or U18780 (N_18780,N_17991,N_17831);
xor U18781 (N_18781,N_18625,N_17956);
nor U18782 (N_18782,N_17526,N_18360);
or U18783 (N_18783,N_18545,N_18727);
xnor U18784 (N_18784,N_17813,N_18648);
nand U18785 (N_18785,N_17851,N_17681);
nor U18786 (N_18786,N_17919,N_18010);
and U18787 (N_18787,N_17763,N_17764);
nand U18788 (N_18788,N_17677,N_18425);
nor U18789 (N_18789,N_17696,N_17988);
and U18790 (N_18790,N_18141,N_18044);
or U18791 (N_18791,N_18337,N_18079);
xnor U18792 (N_18792,N_18574,N_18748);
or U18793 (N_18793,N_18628,N_17512);
and U18794 (N_18794,N_17762,N_18112);
nor U18795 (N_18795,N_17872,N_18399);
nor U18796 (N_18796,N_18221,N_18267);
nand U18797 (N_18797,N_17520,N_18571);
or U18798 (N_18798,N_18063,N_18346);
nand U18799 (N_18799,N_18700,N_18060);
or U18800 (N_18800,N_17768,N_18354);
nand U18801 (N_18801,N_18481,N_18101);
nor U18802 (N_18802,N_18418,N_17893);
xor U18803 (N_18803,N_18486,N_17782);
or U18804 (N_18804,N_18633,N_17734);
nor U18805 (N_18805,N_18181,N_18632);
xnor U18806 (N_18806,N_17746,N_18531);
xor U18807 (N_18807,N_18056,N_17701);
xor U18808 (N_18808,N_18716,N_18472);
xor U18809 (N_18809,N_18547,N_17897);
nor U18810 (N_18810,N_18459,N_18284);
xor U18811 (N_18811,N_17668,N_18527);
or U18812 (N_18812,N_18341,N_18324);
and U18813 (N_18813,N_17900,N_18718);
nor U18814 (N_18814,N_18173,N_17926);
or U18815 (N_18815,N_18130,N_18244);
nand U18816 (N_18816,N_18589,N_18435);
nand U18817 (N_18817,N_17652,N_18713);
nand U18818 (N_18818,N_17916,N_17580);
nor U18819 (N_18819,N_17973,N_18232);
xor U18820 (N_18820,N_17947,N_18094);
nor U18821 (N_18821,N_18370,N_17638);
or U18822 (N_18822,N_18380,N_17769);
or U18823 (N_18823,N_18092,N_17549);
xor U18824 (N_18824,N_17508,N_17921);
xor U18825 (N_18825,N_18504,N_17590);
xor U18826 (N_18826,N_18676,N_18148);
or U18827 (N_18827,N_18630,N_18562);
nor U18828 (N_18828,N_18375,N_17883);
nor U18829 (N_18829,N_18514,N_18033);
or U18830 (N_18830,N_17952,N_17812);
nor U18831 (N_18831,N_18484,N_18200);
xor U18832 (N_18832,N_18474,N_18576);
or U18833 (N_18833,N_17726,N_18157);
or U18834 (N_18834,N_17833,N_17826);
and U18835 (N_18835,N_18078,N_18693);
xor U18836 (N_18836,N_17890,N_18155);
xor U18837 (N_18837,N_17927,N_17785);
xor U18838 (N_18838,N_17767,N_17755);
xnor U18839 (N_18839,N_17687,N_18478);
xor U18840 (N_18840,N_18607,N_18672);
nand U18841 (N_18841,N_18196,N_18381);
nand U18842 (N_18842,N_17725,N_17649);
nor U18843 (N_18843,N_17686,N_17678);
or U18844 (N_18844,N_17800,N_18490);
nand U18845 (N_18845,N_18583,N_17710);
nor U18846 (N_18846,N_18454,N_18421);
nand U18847 (N_18847,N_17732,N_17797);
and U18848 (N_18848,N_17539,N_17636);
nand U18849 (N_18849,N_18150,N_18175);
and U18850 (N_18850,N_18037,N_18054);
nor U18851 (N_18851,N_18369,N_18241);
and U18852 (N_18852,N_17946,N_18134);
nor U18853 (N_18853,N_18506,N_18445);
or U18854 (N_18854,N_18736,N_18059);
nand U18855 (N_18855,N_18641,N_18251);
or U18856 (N_18856,N_18351,N_18505);
or U18857 (N_18857,N_17516,N_18172);
nor U18858 (N_18858,N_17752,N_18032);
and U18859 (N_18859,N_18365,N_18143);
or U18860 (N_18860,N_18388,N_18372);
nor U18861 (N_18861,N_18055,N_17601);
and U18862 (N_18862,N_17811,N_18534);
xnor U18863 (N_18863,N_18208,N_17859);
and U18864 (N_18864,N_18177,N_18584);
and U18865 (N_18865,N_17847,N_18746);
or U18866 (N_18866,N_17896,N_17941);
nand U18867 (N_18867,N_18133,N_18410);
nor U18868 (N_18868,N_18678,N_18338);
xor U18869 (N_18869,N_18734,N_18020);
nor U18870 (N_18870,N_17662,N_17554);
and U18871 (N_18871,N_18116,N_18248);
xnor U18872 (N_18872,N_18414,N_18384);
nor U18873 (N_18873,N_17550,N_17808);
and U18874 (N_18874,N_18247,N_18170);
or U18875 (N_18875,N_17888,N_17541);
or U18876 (N_18876,N_18668,N_17802);
or U18877 (N_18877,N_18488,N_18580);
or U18878 (N_18878,N_17587,N_18136);
nor U18879 (N_18879,N_18691,N_17880);
xor U18880 (N_18880,N_17663,N_17978);
and U18881 (N_18881,N_18739,N_18126);
or U18882 (N_18882,N_18715,N_18413);
or U18883 (N_18883,N_17836,N_18619);
and U18884 (N_18884,N_17868,N_18110);
and U18885 (N_18885,N_17532,N_18500);
nand U18886 (N_18886,N_18249,N_18246);
and U18887 (N_18887,N_17674,N_17524);
xnor U18888 (N_18888,N_18238,N_17693);
nand U18889 (N_18889,N_18460,N_18696);
and U18890 (N_18890,N_18254,N_18266);
xor U18891 (N_18891,N_18226,N_18186);
nor U18892 (N_18892,N_18396,N_18053);
nand U18893 (N_18893,N_18269,N_17694);
nor U18894 (N_18894,N_17892,N_17595);
nand U18895 (N_18895,N_18307,N_18541);
xnor U18896 (N_18896,N_18189,N_18685);
xnor U18897 (N_18897,N_18635,N_18458);
xnor U18898 (N_18898,N_17980,N_17940);
xnor U18899 (N_18899,N_17992,N_17700);
nand U18900 (N_18900,N_17856,N_18400);
nand U18901 (N_18901,N_18732,N_17865);
xor U18902 (N_18902,N_18294,N_18694);
nor U18903 (N_18903,N_18675,N_17560);
nor U18904 (N_18904,N_17559,N_18482);
xnor U18905 (N_18905,N_18533,N_17898);
nand U18906 (N_18906,N_18398,N_17912);
and U18907 (N_18907,N_18364,N_18469);
nand U18908 (N_18908,N_17637,N_17722);
or U18909 (N_18909,N_18543,N_17536);
xor U18910 (N_18910,N_17564,N_18397);
nand U18911 (N_18911,N_18253,N_18636);
nor U18912 (N_18912,N_18525,N_17670);
xor U18913 (N_18913,N_18551,N_18376);
and U18914 (N_18914,N_18345,N_18273);
nand U18915 (N_18915,N_17879,N_17739);
xor U18916 (N_18916,N_18479,N_17593);
xor U18917 (N_18917,N_18024,N_18227);
nand U18918 (N_18918,N_18156,N_17712);
and U18919 (N_18919,N_18282,N_17709);
and U18920 (N_18920,N_18076,N_18520);
nand U18921 (N_18921,N_17567,N_18434);
xnor U18922 (N_18922,N_17777,N_18074);
nor U18923 (N_18923,N_18035,N_18538);
and U18924 (N_18924,N_18080,N_18424);
xnor U18925 (N_18925,N_17644,N_18412);
nand U18926 (N_18926,N_18461,N_18688);
or U18927 (N_18927,N_17704,N_18496);
nor U18928 (N_18928,N_18611,N_18508);
nand U18929 (N_18929,N_17801,N_18334);
nand U18930 (N_18930,N_17982,N_17976);
xnor U18931 (N_18931,N_18431,N_17962);
nor U18932 (N_18932,N_18489,N_17787);
nor U18933 (N_18933,N_18509,N_17965);
or U18934 (N_18934,N_18644,N_18728);
nor U18935 (N_18935,N_17798,N_18415);
nand U18936 (N_18936,N_18596,N_17786);
xor U18937 (N_18937,N_18296,N_17740);
and U18938 (N_18938,N_17791,N_18093);
nand U18939 (N_18939,N_18406,N_18297);
nor U18940 (N_18940,N_18326,N_18483);
or U18941 (N_18941,N_17773,N_18503);
nand U18942 (N_18942,N_18724,N_18211);
nand U18943 (N_18943,N_18229,N_18096);
or U18944 (N_18944,N_17805,N_18194);
nor U18945 (N_18945,N_17850,N_17818);
nor U18946 (N_18946,N_17544,N_18091);
nor U18947 (N_18947,N_18213,N_17876);
and U18948 (N_18948,N_18595,N_18058);
nand U18949 (N_18949,N_17972,N_17819);
xnor U18950 (N_18950,N_18599,N_18615);
or U18951 (N_18951,N_18068,N_18717);
nor U18952 (N_18952,N_17789,N_17737);
nor U18953 (N_18953,N_17967,N_18304);
xor U18954 (N_18954,N_18220,N_18327);
nand U18955 (N_18955,N_18627,N_17578);
nand U18956 (N_18956,N_18480,N_17906);
and U18957 (N_18957,N_17860,N_18475);
nor U18958 (N_18958,N_18066,N_17943);
and U18959 (N_18959,N_18419,N_17568);
and U18960 (N_18960,N_17611,N_17625);
nor U18961 (N_18961,N_17873,N_17821);
or U18962 (N_18962,N_17552,N_17957);
nor U18963 (N_18963,N_18390,N_18147);
nand U18964 (N_18964,N_18437,N_18686);
nor U18965 (N_18965,N_17910,N_18394);
nand U18966 (N_18966,N_18322,N_17672);
nor U18967 (N_18967,N_18030,N_18250);
and U18968 (N_18968,N_18203,N_17588);
or U18969 (N_18969,N_18107,N_18653);
xnor U18970 (N_18970,N_18318,N_17891);
nand U18971 (N_18971,N_18477,N_17698);
xor U18972 (N_18972,N_17929,N_18152);
nand U18973 (N_18973,N_18707,N_17842);
and U18974 (N_18974,N_18522,N_17853);
nand U18975 (N_18975,N_17983,N_17718);
nor U18976 (N_18976,N_18233,N_18314);
xor U18977 (N_18977,N_17529,N_17780);
nand U18978 (N_18978,N_18385,N_17996);
and U18979 (N_18979,N_18467,N_17753);
nand U18980 (N_18980,N_18403,N_17632);
xor U18981 (N_18981,N_17735,N_18013);
nor U18982 (N_18982,N_18492,N_18018);
xor U18983 (N_18983,N_17615,N_18183);
nor U18984 (N_18984,N_18048,N_17731);
xnor U18985 (N_18985,N_18111,N_17829);
nand U18986 (N_18986,N_17760,N_18295);
and U18987 (N_18987,N_17609,N_18682);
and U18988 (N_18988,N_18377,N_18119);
and U18989 (N_18989,N_17660,N_17922);
nor U18990 (N_18990,N_18401,N_18290);
or U18991 (N_18991,N_18146,N_18023);
and U18992 (N_18992,N_18714,N_18237);
nand U18993 (N_18993,N_17815,N_18311);
and U18994 (N_18994,N_18039,N_17665);
or U18995 (N_18995,N_18163,N_18298);
xor U18996 (N_18996,N_17573,N_18335);
or U18997 (N_18997,N_18100,N_17598);
and U18998 (N_18998,N_18620,N_18182);
nor U18999 (N_18999,N_18590,N_18587);
nor U19000 (N_19000,N_17515,N_17523);
nor U19001 (N_19001,N_17707,N_17729);
and U19002 (N_19002,N_18586,N_18701);
or U19003 (N_19003,N_18663,N_18206);
and U19004 (N_19004,N_17548,N_18639);
or U19005 (N_19005,N_17986,N_18276);
and U19006 (N_19006,N_18499,N_18255);
xor U19007 (N_19007,N_17518,N_17669);
nor U19008 (N_19008,N_18214,N_18428);
nor U19009 (N_19009,N_17793,N_17570);
or U19010 (N_19010,N_18529,N_18559);
nand U19011 (N_19011,N_17933,N_18521);
xor U19012 (N_19012,N_17691,N_18745);
nand U19013 (N_19013,N_18512,N_18149);
xor U19014 (N_19014,N_17531,N_17506);
nor U19015 (N_19015,N_17581,N_17779);
and U19016 (N_19016,N_18315,N_18216);
xor U19017 (N_19017,N_18448,N_18174);
nor U19018 (N_19018,N_18613,N_18444);
or U19019 (N_19019,N_17820,N_17855);
xor U19020 (N_19020,N_18260,N_17866);
nor U19021 (N_19021,N_18165,N_18601);
nand U19022 (N_19022,N_18017,N_17594);
nand U19023 (N_19023,N_17838,N_17903);
nor U19024 (N_19024,N_18108,N_18540);
nand U19025 (N_19025,N_18617,N_18550);
and U19026 (N_19026,N_18683,N_18669);
or U19027 (N_19027,N_18702,N_18359);
xnor U19028 (N_19028,N_17641,N_18288);
nor U19029 (N_19029,N_18537,N_17736);
or U19030 (N_19030,N_18446,N_18191);
nor U19031 (N_19031,N_18022,N_17931);
or U19032 (N_19032,N_17809,N_17602);
or U19033 (N_19033,N_18123,N_17562);
nor U19034 (N_19034,N_18319,N_17938);
and U19035 (N_19035,N_17653,N_17708);
nor U19036 (N_19036,N_17751,N_18239);
nor U19037 (N_19037,N_17924,N_18643);
nor U19038 (N_19038,N_18045,N_17711);
or U19039 (N_19039,N_17543,N_17667);
nor U19040 (N_19040,N_18677,N_18352);
and U19041 (N_19041,N_18106,N_18602);
nand U19042 (N_19042,N_18452,N_18333);
nand U19043 (N_19043,N_17985,N_18634);
nor U19044 (N_19044,N_18081,N_18692);
and U19045 (N_19045,N_18006,N_17519);
nor U19046 (N_19046,N_17871,N_18673);
nor U19047 (N_19047,N_17864,N_17781);
or U19048 (N_19048,N_17617,N_18357);
nor U19049 (N_19049,N_18160,N_17828);
and U19050 (N_19050,N_18552,N_18569);
xnor U19051 (N_19051,N_17547,N_18187);
xor U19052 (N_19052,N_18706,N_18511);
and U19053 (N_19053,N_17688,N_17950);
nor U19054 (N_19054,N_17959,N_17534);
xor U19055 (N_19055,N_17948,N_18002);
nor U19056 (N_19056,N_17981,N_17844);
nor U19057 (N_19057,N_18358,N_18363);
nor U19058 (N_19058,N_18217,N_17823);
or U19059 (N_19059,N_17766,N_18417);
or U19060 (N_19060,N_17877,N_17997);
and U19061 (N_19061,N_18657,N_17626);
xnor U19062 (N_19062,N_18117,N_18272);
or U19063 (N_19063,N_18651,N_18470);
or U19064 (N_19064,N_17803,N_18642);
nand U19065 (N_19065,N_18145,N_18622);
nand U19066 (N_19066,N_17806,N_18258);
and U19067 (N_19067,N_18563,N_18197);
xnor U19068 (N_19068,N_18243,N_17630);
nor U19069 (N_19069,N_17754,N_17841);
and U19070 (N_19070,N_18299,N_18095);
or U19071 (N_19071,N_18593,N_18703);
nor U19072 (N_19072,N_17995,N_17999);
or U19073 (N_19073,N_17676,N_18084);
nor U19074 (N_19074,N_18218,N_18313);
or U19075 (N_19075,N_17655,N_18199);
and U19076 (N_19076,N_18270,N_18518);
nand U19077 (N_19077,N_18286,N_17790);
nor U19078 (N_19078,N_17723,N_18626);
nor U19079 (N_19079,N_17683,N_18158);
xor U19080 (N_19080,N_18339,N_17792);
and U19081 (N_19081,N_18553,N_17631);
xnor U19082 (N_19082,N_18179,N_18350);
or U19083 (N_19083,N_18067,N_18618);
nor U19084 (N_19084,N_17827,N_17643);
xnor U19085 (N_19085,N_18349,N_18741);
nand U19086 (N_19086,N_17507,N_18287);
or U19087 (N_19087,N_17908,N_17591);
nand U19088 (N_19088,N_17642,N_18664);
or U19089 (N_19089,N_17650,N_18436);
and U19090 (N_19090,N_17994,N_17807);
or U19091 (N_19091,N_18698,N_17942);
and U19092 (N_19092,N_18524,N_17500);
xnor U19093 (N_19093,N_17744,N_18494);
or U19094 (N_19094,N_18723,N_17998);
xor U19095 (N_19095,N_17861,N_18325);
nand U19096 (N_19096,N_17867,N_17743);
and U19097 (N_19097,N_17504,N_18449);
nor U19098 (N_19098,N_18029,N_18050);
nor U19099 (N_19099,N_18422,N_18329);
nand U19100 (N_19100,N_18560,N_18679);
xnor U19101 (N_19101,N_18747,N_17553);
or U19102 (N_19102,N_18262,N_18684);
xnor U19103 (N_19103,N_18062,N_18120);
nor U19104 (N_19104,N_17721,N_18231);
xor U19105 (N_19105,N_17837,N_18426);
xor U19106 (N_19106,N_17621,N_18631);
or U19107 (N_19107,N_18565,N_18485);
or U19108 (N_19108,N_18104,N_17961);
nor U19109 (N_19109,N_18001,N_17964);
nand U19110 (N_19110,N_18274,N_18608);
or U19111 (N_19111,N_17756,N_17825);
nor U19112 (N_19112,N_18451,N_18252);
or U19113 (N_19113,N_17612,N_17832);
nand U19114 (N_19114,N_17555,N_18275);
and U19115 (N_19115,N_18131,N_18647);
nor U19116 (N_19116,N_17822,N_18749);
and U19117 (N_19117,N_18070,N_18402);
or U19118 (N_19118,N_18212,N_17592);
nor U19119 (N_19119,N_18528,N_18502);
xnor U19120 (N_19120,N_17585,N_18222);
nand U19121 (N_19121,N_18305,N_18000);
or U19122 (N_19122,N_18331,N_17535);
nand U19123 (N_19123,N_18621,N_17738);
xnor U19124 (N_19124,N_18564,N_17648);
xnor U19125 (N_19125,N_18124,N_17989);
or U19126 (N_19126,N_17920,N_17606);
nand U19127 (N_19127,N_18666,N_18277);
and U19128 (N_19128,N_18105,N_17596);
nor U19129 (N_19129,N_18405,N_17511);
nor U19130 (N_19130,N_18725,N_17584);
nor U19131 (N_19131,N_17974,N_17514);
nor U19132 (N_19132,N_17963,N_18256);
xnor U19133 (N_19133,N_18498,N_18443);
xor U19134 (N_19134,N_18236,N_17848);
xor U19135 (N_19135,N_18473,N_18086);
xnor U19136 (N_19136,N_18077,N_18597);
xor U19137 (N_19137,N_18278,N_18071);
xnor U19138 (N_19138,N_18153,N_17843);
xor U19139 (N_19139,N_17870,N_18088);
nor U19140 (N_19140,N_18115,N_17608);
nor U19141 (N_19141,N_17628,N_18052);
or U19142 (N_19142,N_17716,N_18516);
nand U19143 (N_19143,N_18047,N_17761);
xor U19144 (N_19144,N_18671,N_18371);
xor U19145 (N_19145,N_17706,N_17955);
nor U19146 (N_19146,N_17915,N_18738);
or U19147 (N_19147,N_18014,N_17566);
and U19148 (N_19148,N_18566,N_18209);
xor U19149 (N_19149,N_17658,N_18535);
xor U19150 (N_19150,N_18204,N_17741);
nor U19151 (N_19151,N_18378,N_18159);
or U19152 (N_19152,N_17692,N_18487);
and U19153 (N_19153,N_17968,N_18423);
nor U19154 (N_19154,N_17750,N_18442);
xnor U19155 (N_19155,N_17936,N_17576);
nand U19156 (N_19156,N_18122,N_18429);
or U19157 (N_19157,N_18015,N_18409);
and U19158 (N_19158,N_18468,N_17623);
or U19159 (N_19159,N_18103,N_17525);
or U19160 (N_19160,N_17977,N_18661);
and U19161 (N_19161,N_17887,N_18720);
xor U19162 (N_19162,N_17607,N_18034);
or U19163 (N_19163,N_18289,N_17937);
xor U19164 (N_19164,N_17501,N_17858);
xnor U19165 (N_19165,N_17730,N_18348);
or U19166 (N_19166,N_18730,N_18558);
nor U19167 (N_19167,N_17824,N_17558);
xnor U19168 (N_19168,N_18530,N_17697);
nand U19169 (N_19169,N_17640,N_17816);
or U19170 (N_19170,N_18336,N_17774);
nand U19171 (N_19171,N_17522,N_18235);
nor U19172 (N_19172,N_17857,N_17902);
nand U19173 (N_19173,N_18735,N_18466);
or U19174 (N_19174,N_18450,N_18215);
nand U19175 (N_19175,N_18114,N_18623);
xnor U19176 (N_19176,N_18667,N_17788);
or U19177 (N_19177,N_18285,N_18729);
or U19178 (N_19178,N_18554,N_17517);
xor U19179 (N_19179,N_18603,N_18162);
and U19180 (N_19180,N_18393,N_17878);
nor U19181 (N_19181,N_18347,N_18151);
and U19182 (N_19182,N_17899,N_18323);
nor U19183 (N_19183,N_18659,N_17682);
or U19184 (N_19184,N_18009,N_17571);
nand U19185 (N_19185,N_18328,N_17835);
nand U19186 (N_19186,N_17904,N_18645);
xor U19187 (N_19187,N_17664,N_18026);
or U19188 (N_19188,N_17699,N_17685);
xor U19189 (N_19189,N_18008,N_18665);
nor U19190 (N_19190,N_18557,N_18711);
nand U19191 (N_19191,N_17759,N_17561);
nor U19192 (N_19192,N_17513,N_17645);
or U19193 (N_19193,N_18302,N_18646);
nor U19194 (N_19194,N_17778,N_18447);
xnor U19195 (N_19195,N_17849,N_18395);
nand U19196 (N_19196,N_18709,N_18561);
or U19197 (N_19197,N_18031,N_18169);
and U19198 (N_19198,N_18240,N_17799);
or U19199 (N_19199,N_18308,N_18268);
xor U19200 (N_19200,N_18737,N_17909);
xnor U19201 (N_19201,N_18649,N_18176);
xnor U19202 (N_19202,N_17770,N_18043);
nor U19203 (N_19203,N_18330,N_18344);
or U19204 (N_19204,N_18462,N_17533);
or U19205 (N_19205,N_17804,N_17604);
nand U19206 (N_19206,N_18144,N_18379);
nor U19207 (N_19207,N_18089,N_18689);
nor U19208 (N_19208,N_18366,N_18733);
xnor U19209 (N_19209,N_18510,N_18740);
nand U19210 (N_19210,N_17783,N_17618);
xnor U19211 (N_19211,N_18279,N_18263);
nand U19212 (N_19212,N_18310,N_18392);
nand U19213 (N_19213,N_18532,N_18629);
xor U19214 (N_19214,N_17563,N_17993);
nor U19215 (N_19215,N_18057,N_18332);
nor U19216 (N_19216,N_18710,N_17510);
nand U19217 (N_19217,N_18343,N_18073);
nand U19218 (N_19218,N_17796,N_18493);
nor U19219 (N_19219,N_18201,N_18656);
xor U19220 (N_19220,N_18726,N_17582);
or U19221 (N_19221,N_18517,N_17945);
nor U19222 (N_19222,N_18687,N_18742);
and U19223 (N_19223,N_18606,N_17586);
nor U19224 (N_19224,N_17556,N_18291);
nand U19225 (N_19225,N_17661,N_17689);
and U19226 (N_19226,N_18438,N_17624);
xnor U19227 (N_19227,N_18577,N_18072);
nor U19228 (N_19228,N_18362,N_18662);
xor U19229 (N_19229,N_17875,N_17530);
nand U19230 (N_19230,N_17545,N_18526);
nor U19231 (N_19231,N_18265,N_17884);
nand U19232 (N_19232,N_18019,N_17679);
or U19233 (N_19233,N_17666,N_18190);
xnor U19234 (N_19234,N_17895,N_18476);
nor U19235 (N_19235,N_17905,N_17979);
nand U19236 (N_19236,N_17600,N_17747);
or U19237 (N_19237,N_17749,N_18135);
nor U19238 (N_19238,N_17565,N_17720);
and U19239 (N_19239,N_17715,N_17619);
xor U19240 (N_19240,N_17834,N_17830);
xnor U19241 (N_19241,N_17932,N_17886);
nor U19242 (N_19242,N_17869,N_18041);
nand U19243 (N_19243,N_18281,N_17572);
or U19244 (N_19244,N_17633,N_18604);
nor U19245 (N_19245,N_18556,N_18610);
nand U19246 (N_19246,N_17882,N_17975);
xor U19247 (N_19247,N_18098,N_18430);
nor U19248 (N_19248,N_18549,N_18519);
xnor U19249 (N_19249,N_18722,N_18420);
or U19250 (N_19250,N_18439,N_18128);
or U19251 (N_19251,N_18320,N_17724);
or U19252 (N_19252,N_17634,N_17949);
or U19253 (N_19253,N_18383,N_18523);
xnor U19254 (N_19254,N_18257,N_17757);
or U19255 (N_19255,N_17597,N_17918);
and U19256 (N_19256,N_18065,N_17639);
nor U19257 (N_19257,N_18581,N_18161);
and U19258 (N_19258,N_18674,N_18658);
and U19259 (N_19259,N_18138,N_17537);
xnor U19260 (N_19260,N_18404,N_18592);
or U19261 (N_19261,N_18536,N_18374);
and U19262 (N_19262,N_18624,N_18049);
or U19263 (N_19263,N_18188,N_18300);
nor U19264 (N_19264,N_18591,N_18708);
nor U19265 (N_19265,N_18261,N_17614);
and U19266 (N_19266,N_17894,N_17657);
nand U19267 (N_19267,N_17577,N_18230);
nor U19268 (N_19268,N_18036,N_17874);
and U19269 (N_19269,N_17728,N_17795);
xor U19270 (N_19270,N_17654,N_18386);
or U19271 (N_19271,N_17733,N_18573);
or U19272 (N_19272,N_17647,N_18637);
and U19273 (N_19273,N_17599,N_18712);
nand U19274 (N_19274,N_17971,N_18605);
and U19275 (N_19275,N_18699,N_18028);
nand U19276 (N_19276,N_17613,N_18594);
and U19277 (N_19277,N_17840,N_18453);
and U19278 (N_19278,N_18180,N_17620);
nand U19279 (N_19279,N_18491,N_18207);
nand U19280 (N_19280,N_17656,N_17925);
and U19281 (N_19281,N_17727,N_18042);
or U19282 (N_19282,N_17574,N_18353);
xnor U19283 (N_19283,N_17960,N_17970);
xor U19284 (N_19284,N_17605,N_17542);
and U19285 (N_19285,N_17901,N_18416);
and U19286 (N_19286,N_18640,N_18245);
xor U19287 (N_19287,N_18570,N_18121);
nand U19288 (N_19288,N_18132,N_18012);
or U19289 (N_19289,N_17673,N_18638);
nand U19290 (N_19290,N_17583,N_18118);
xnor U19291 (N_19291,N_18660,N_18139);
xor U19292 (N_19292,N_17839,N_18011);
or U19293 (N_19293,N_18040,N_18109);
nand U19294 (N_19294,N_18497,N_17889);
nand U19295 (N_19295,N_18016,N_18312);
and U19296 (N_19296,N_17575,N_17814);
and U19297 (N_19297,N_18355,N_17784);
xor U19298 (N_19298,N_18495,N_17719);
nor U19299 (N_19299,N_18387,N_18027);
xnor U19300 (N_19300,N_18280,N_17765);
xor U19301 (N_19301,N_18192,N_18038);
nand U19302 (N_19302,N_18306,N_18259);
nand U19303 (N_19303,N_17502,N_18609);
nor U19304 (N_19304,N_18588,N_17603);
xor U19305 (N_19305,N_18382,N_18507);
or U19306 (N_19306,N_18654,N_18705);
xnor U19307 (N_19307,N_18719,N_18389);
and U19308 (N_19308,N_18166,N_18083);
xnor U19309 (N_19309,N_18198,N_17772);
nand U19310 (N_19310,N_18368,N_18342);
nor U19311 (N_19311,N_18224,N_17569);
or U19312 (N_19312,N_18168,N_18455);
xnor U19313 (N_19313,N_17930,N_17629);
xnor U19314 (N_19314,N_18113,N_17540);
and U19315 (N_19315,N_17987,N_18046);
and U19316 (N_19316,N_18695,N_17659);
xor U19317 (N_19317,N_18171,N_18004);
and U19318 (N_19318,N_17546,N_18655);
nand U19319 (N_19319,N_17863,N_17944);
and U19320 (N_19320,N_18069,N_17984);
or U19321 (N_19321,N_17911,N_18731);
nor U19322 (N_19322,N_18129,N_18614);
and U19323 (N_19323,N_18219,N_17966);
nor U19324 (N_19324,N_18744,N_17776);
or U19325 (N_19325,N_18021,N_18210);
or U19326 (N_19326,N_18178,N_17703);
or U19327 (N_19327,N_17969,N_17557);
or U19328 (N_19328,N_17846,N_18572);
xnor U19329 (N_19329,N_18427,N_18184);
and U19330 (N_19330,N_17748,N_17714);
or U19331 (N_19331,N_18361,N_18082);
nor U19332 (N_19332,N_18283,N_18185);
or U19333 (N_19333,N_18087,N_18097);
nor U19334 (N_19334,N_17913,N_17958);
xnor U19335 (N_19335,N_18441,N_17885);
nand U19336 (N_19336,N_18407,N_18137);
xnor U19337 (N_19337,N_18585,N_18356);
and U19338 (N_19338,N_17951,N_18471);
nor U19339 (N_19339,N_17845,N_17939);
and U19340 (N_19340,N_18303,N_18743);
nor U19341 (N_19341,N_18154,N_17742);
and U19342 (N_19342,N_17579,N_17907);
nand U19343 (N_19343,N_18690,N_17717);
and U19344 (N_19344,N_18579,N_18391);
nand U19345 (N_19345,N_18681,N_18099);
or U19346 (N_19346,N_18367,N_18373);
nor U19347 (N_19347,N_17914,N_18127);
or U19348 (N_19348,N_17775,N_17771);
nand U19349 (N_19349,N_18463,N_18457);
nand U19350 (N_19350,N_18440,N_17917);
nor U19351 (N_19351,N_18003,N_18225);
nand U19352 (N_19352,N_17713,N_18721);
or U19353 (N_19353,N_18321,N_18567);
or U19354 (N_19354,N_17953,N_18316);
nor U19355 (N_19355,N_18616,N_18340);
nor U19356 (N_19356,N_17705,N_18598);
xor U19357 (N_19357,N_18697,N_17854);
and U19358 (N_19358,N_18309,N_17551);
or U19359 (N_19359,N_18005,N_17646);
nor U19360 (N_19360,N_18075,N_17521);
xnor U19361 (N_19361,N_18542,N_17675);
nand U19362 (N_19362,N_18301,N_18680);
xor U19363 (N_19363,N_18195,N_18102);
or U19364 (N_19364,N_18293,N_17935);
nor U19365 (N_19365,N_17862,N_18600);
and U19366 (N_19366,N_18432,N_17852);
xnor U19367 (N_19367,N_17990,N_18292);
xor U19368 (N_19368,N_17651,N_18568);
nor U19369 (N_19369,N_17934,N_18544);
and U19370 (N_19370,N_18205,N_18085);
nand U19371 (N_19371,N_18125,N_18539);
nor U19372 (N_19372,N_18465,N_18704);
nor U19373 (N_19373,N_17610,N_18670);
nand U19374 (N_19374,N_18548,N_18652);
nor U19375 (N_19375,N_18352,N_17701);
nand U19376 (N_19376,N_18000,N_18633);
xnor U19377 (N_19377,N_18594,N_18601);
nor U19378 (N_19378,N_18388,N_17949);
nand U19379 (N_19379,N_18555,N_18354);
and U19380 (N_19380,N_17780,N_17579);
nor U19381 (N_19381,N_17639,N_17846);
and U19382 (N_19382,N_18382,N_18194);
nor U19383 (N_19383,N_17719,N_17622);
xnor U19384 (N_19384,N_18097,N_18391);
nand U19385 (N_19385,N_18248,N_18098);
xnor U19386 (N_19386,N_18124,N_18640);
xor U19387 (N_19387,N_18590,N_17922);
nand U19388 (N_19388,N_18652,N_17807);
nor U19389 (N_19389,N_18068,N_17888);
or U19390 (N_19390,N_17673,N_18063);
nor U19391 (N_19391,N_18039,N_17904);
xor U19392 (N_19392,N_17919,N_18734);
and U19393 (N_19393,N_18745,N_18137);
or U19394 (N_19394,N_17579,N_18441);
nand U19395 (N_19395,N_18391,N_18517);
nand U19396 (N_19396,N_18665,N_18074);
or U19397 (N_19397,N_17988,N_18000);
xnor U19398 (N_19398,N_17847,N_17822);
nor U19399 (N_19399,N_17617,N_18696);
xor U19400 (N_19400,N_18535,N_18254);
nor U19401 (N_19401,N_18050,N_18742);
nor U19402 (N_19402,N_18491,N_18026);
or U19403 (N_19403,N_18409,N_18063);
or U19404 (N_19404,N_18338,N_17697);
and U19405 (N_19405,N_18564,N_18167);
nor U19406 (N_19406,N_18388,N_18086);
nor U19407 (N_19407,N_17831,N_18698);
xor U19408 (N_19408,N_17677,N_18383);
or U19409 (N_19409,N_18257,N_18569);
nand U19410 (N_19410,N_18369,N_17595);
or U19411 (N_19411,N_18459,N_18056);
and U19412 (N_19412,N_17904,N_18481);
xor U19413 (N_19413,N_17705,N_18111);
nor U19414 (N_19414,N_17789,N_18063);
xnor U19415 (N_19415,N_17851,N_18065);
and U19416 (N_19416,N_18322,N_17805);
nor U19417 (N_19417,N_17882,N_18286);
xor U19418 (N_19418,N_18486,N_18515);
or U19419 (N_19419,N_17710,N_17846);
or U19420 (N_19420,N_18718,N_17658);
and U19421 (N_19421,N_18722,N_17961);
xnor U19422 (N_19422,N_18571,N_18068);
nor U19423 (N_19423,N_18507,N_18019);
nor U19424 (N_19424,N_18154,N_18526);
xnor U19425 (N_19425,N_18421,N_18553);
nor U19426 (N_19426,N_17811,N_17787);
nand U19427 (N_19427,N_18746,N_17665);
or U19428 (N_19428,N_18374,N_17892);
nand U19429 (N_19429,N_17992,N_17907);
xnor U19430 (N_19430,N_17759,N_18345);
xnor U19431 (N_19431,N_17637,N_18477);
and U19432 (N_19432,N_18391,N_17983);
and U19433 (N_19433,N_17965,N_18388);
xnor U19434 (N_19434,N_17779,N_18224);
or U19435 (N_19435,N_18216,N_18558);
xor U19436 (N_19436,N_18464,N_18186);
and U19437 (N_19437,N_17780,N_18139);
nand U19438 (N_19438,N_17874,N_18233);
nor U19439 (N_19439,N_18101,N_18515);
nor U19440 (N_19440,N_18469,N_18136);
and U19441 (N_19441,N_18206,N_18420);
or U19442 (N_19442,N_18316,N_18258);
xnor U19443 (N_19443,N_17519,N_17633);
and U19444 (N_19444,N_18283,N_18092);
xnor U19445 (N_19445,N_17530,N_18573);
nor U19446 (N_19446,N_18275,N_18078);
xor U19447 (N_19447,N_18370,N_17903);
and U19448 (N_19448,N_18659,N_18714);
nand U19449 (N_19449,N_18177,N_17508);
and U19450 (N_19450,N_18732,N_17674);
xnor U19451 (N_19451,N_18197,N_17905);
or U19452 (N_19452,N_18531,N_18626);
and U19453 (N_19453,N_17846,N_17766);
nor U19454 (N_19454,N_17560,N_18364);
nor U19455 (N_19455,N_17521,N_18070);
nand U19456 (N_19456,N_18746,N_17629);
xnor U19457 (N_19457,N_18628,N_18507);
nand U19458 (N_19458,N_18485,N_17869);
and U19459 (N_19459,N_17543,N_17690);
and U19460 (N_19460,N_17744,N_18663);
or U19461 (N_19461,N_17626,N_18284);
and U19462 (N_19462,N_18325,N_17806);
xor U19463 (N_19463,N_18017,N_17697);
or U19464 (N_19464,N_18213,N_18458);
nand U19465 (N_19465,N_18489,N_17588);
xnor U19466 (N_19466,N_18741,N_17918);
nand U19467 (N_19467,N_18505,N_17993);
and U19468 (N_19468,N_18611,N_17821);
or U19469 (N_19469,N_17577,N_17545);
nand U19470 (N_19470,N_18250,N_17814);
nand U19471 (N_19471,N_18392,N_18571);
or U19472 (N_19472,N_17988,N_18299);
nor U19473 (N_19473,N_18244,N_18006);
nand U19474 (N_19474,N_18569,N_18094);
nor U19475 (N_19475,N_18389,N_18180);
xor U19476 (N_19476,N_17613,N_17719);
xnor U19477 (N_19477,N_18429,N_18330);
xor U19478 (N_19478,N_17872,N_17530);
nand U19479 (N_19479,N_17873,N_17810);
and U19480 (N_19480,N_18343,N_17763);
and U19481 (N_19481,N_18405,N_18656);
nor U19482 (N_19482,N_17914,N_17743);
nor U19483 (N_19483,N_17976,N_18542);
or U19484 (N_19484,N_17761,N_18273);
nor U19485 (N_19485,N_17916,N_17765);
and U19486 (N_19486,N_17851,N_18426);
or U19487 (N_19487,N_18432,N_17926);
and U19488 (N_19488,N_17756,N_17873);
or U19489 (N_19489,N_18064,N_18700);
and U19490 (N_19490,N_17556,N_18708);
nand U19491 (N_19491,N_18368,N_18268);
xnor U19492 (N_19492,N_17980,N_18511);
nand U19493 (N_19493,N_17519,N_17813);
nor U19494 (N_19494,N_18597,N_17726);
and U19495 (N_19495,N_17675,N_18052);
nand U19496 (N_19496,N_17612,N_18564);
nand U19497 (N_19497,N_18266,N_17924);
nand U19498 (N_19498,N_17575,N_18270);
nor U19499 (N_19499,N_17912,N_18249);
xnor U19500 (N_19500,N_17964,N_17984);
and U19501 (N_19501,N_18377,N_17751);
xnor U19502 (N_19502,N_18300,N_18293);
nor U19503 (N_19503,N_17964,N_17735);
or U19504 (N_19504,N_18286,N_18717);
nor U19505 (N_19505,N_17612,N_18243);
or U19506 (N_19506,N_18105,N_17733);
xor U19507 (N_19507,N_18247,N_17819);
xnor U19508 (N_19508,N_17705,N_18715);
nor U19509 (N_19509,N_17883,N_17817);
and U19510 (N_19510,N_18333,N_18704);
xnor U19511 (N_19511,N_17624,N_18546);
nand U19512 (N_19512,N_17968,N_17572);
and U19513 (N_19513,N_18442,N_18734);
and U19514 (N_19514,N_18258,N_17714);
nand U19515 (N_19515,N_17728,N_17504);
and U19516 (N_19516,N_18405,N_17535);
and U19517 (N_19517,N_17776,N_18717);
nand U19518 (N_19518,N_18158,N_18172);
or U19519 (N_19519,N_18732,N_18379);
and U19520 (N_19520,N_17790,N_18405);
xor U19521 (N_19521,N_18298,N_18322);
nor U19522 (N_19522,N_18685,N_17564);
and U19523 (N_19523,N_18294,N_17505);
xnor U19524 (N_19524,N_18501,N_18345);
or U19525 (N_19525,N_17787,N_17899);
nand U19526 (N_19526,N_17841,N_17525);
or U19527 (N_19527,N_18470,N_18490);
or U19528 (N_19528,N_18198,N_17514);
xor U19529 (N_19529,N_17924,N_18334);
or U19530 (N_19530,N_18078,N_17522);
and U19531 (N_19531,N_18695,N_18481);
nand U19532 (N_19532,N_18650,N_17810);
nand U19533 (N_19533,N_18035,N_18421);
xor U19534 (N_19534,N_17795,N_18061);
nor U19535 (N_19535,N_18684,N_17926);
or U19536 (N_19536,N_17748,N_18556);
xnor U19537 (N_19537,N_18090,N_17619);
nor U19538 (N_19538,N_18702,N_18497);
or U19539 (N_19539,N_18542,N_17910);
and U19540 (N_19540,N_17917,N_18141);
and U19541 (N_19541,N_17939,N_18259);
or U19542 (N_19542,N_18449,N_18024);
nand U19543 (N_19543,N_18275,N_17524);
nor U19544 (N_19544,N_18126,N_17569);
xor U19545 (N_19545,N_18143,N_18220);
nand U19546 (N_19546,N_18748,N_18362);
nand U19547 (N_19547,N_18166,N_17717);
xor U19548 (N_19548,N_17954,N_17609);
xnor U19549 (N_19549,N_18546,N_18541);
xnor U19550 (N_19550,N_18256,N_18425);
xnor U19551 (N_19551,N_18288,N_18670);
nor U19552 (N_19552,N_18508,N_18123);
nor U19553 (N_19553,N_18105,N_18531);
and U19554 (N_19554,N_17604,N_17718);
and U19555 (N_19555,N_18082,N_18290);
nor U19556 (N_19556,N_17667,N_18115);
or U19557 (N_19557,N_17811,N_18574);
or U19558 (N_19558,N_17997,N_18202);
or U19559 (N_19559,N_18102,N_18706);
or U19560 (N_19560,N_18371,N_18465);
xnor U19561 (N_19561,N_18568,N_17913);
nand U19562 (N_19562,N_18245,N_17956);
or U19563 (N_19563,N_18165,N_18583);
nor U19564 (N_19564,N_18309,N_18522);
xnor U19565 (N_19565,N_18175,N_17760);
nor U19566 (N_19566,N_18571,N_18297);
nor U19567 (N_19567,N_17682,N_17547);
and U19568 (N_19568,N_18157,N_18526);
nor U19569 (N_19569,N_18461,N_18178);
or U19570 (N_19570,N_17586,N_17925);
nand U19571 (N_19571,N_18547,N_17851);
and U19572 (N_19572,N_18221,N_17531);
nand U19573 (N_19573,N_18363,N_17839);
xor U19574 (N_19574,N_17561,N_17581);
or U19575 (N_19575,N_18388,N_18146);
nor U19576 (N_19576,N_18650,N_18319);
and U19577 (N_19577,N_18519,N_18368);
nand U19578 (N_19578,N_17917,N_18724);
xor U19579 (N_19579,N_17556,N_18530);
xor U19580 (N_19580,N_17647,N_17818);
nor U19581 (N_19581,N_18020,N_18345);
or U19582 (N_19582,N_18039,N_18201);
and U19583 (N_19583,N_17700,N_18094);
nor U19584 (N_19584,N_18528,N_18123);
xor U19585 (N_19585,N_18643,N_17585);
nor U19586 (N_19586,N_18019,N_18364);
or U19587 (N_19587,N_18360,N_18074);
and U19588 (N_19588,N_17927,N_18445);
and U19589 (N_19589,N_17610,N_18171);
xor U19590 (N_19590,N_18451,N_17819);
nor U19591 (N_19591,N_17919,N_17629);
xnor U19592 (N_19592,N_17990,N_17997);
nand U19593 (N_19593,N_17629,N_18128);
nor U19594 (N_19594,N_18683,N_17573);
xor U19595 (N_19595,N_18083,N_18316);
xnor U19596 (N_19596,N_17688,N_18105);
nand U19597 (N_19597,N_17507,N_18564);
nand U19598 (N_19598,N_17572,N_18085);
and U19599 (N_19599,N_17887,N_18509);
nor U19600 (N_19600,N_17543,N_17692);
xnor U19601 (N_19601,N_17544,N_18725);
nor U19602 (N_19602,N_17573,N_18067);
xor U19603 (N_19603,N_18155,N_18137);
or U19604 (N_19604,N_18080,N_17762);
or U19605 (N_19605,N_18016,N_18371);
nor U19606 (N_19606,N_17529,N_18200);
nor U19607 (N_19607,N_17930,N_18318);
xnor U19608 (N_19608,N_18199,N_17787);
nand U19609 (N_19609,N_18436,N_18669);
nand U19610 (N_19610,N_17865,N_18707);
nor U19611 (N_19611,N_18741,N_18604);
or U19612 (N_19612,N_18256,N_17997);
nand U19613 (N_19613,N_17634,N_18383);
xnor U19614 (N_19614,N_18483,N_18258);
and U19615 (N_19615,N_18611,N_18663);
xor U19616 (N_19616,N_17680,N_17802);
nand U19617 (N_19617,N_18257,N_17639);
xnor U19618 (N_19618,N_18262,N_17500);
nor U19619 (N_19619,N_18713,N_18124);
nand U19620 (N_19620,N_18571,N_17652);
xnor U19621 (N_19621,N_18322,N_17956);
nor U19622 (N_19622,N_18705,N_18748);
xor U19623 (N_19623,N_17900,N_18295);
and U19624 (N_19624,N_17710,N_18144);
xor U19625 (N_19625,N_17526,N_17842);
or U19626 (N_19626,N_18566,N_18642);
xor U19627 (N_19627,N_18385,N_18570);
and U19628 (N_19628,N_18479,N_18445);
nor U19629 (N_19629,N_17834,N_18577);
or U19630 (N_19630,N_17798,N_18373);
nor U19631 (N_19631,N_18010,N_18607);
or U19632 (N_19632,N_17804,N_18400);
or U19633 (N_19633,N_18686,N_17531);
xor U19634 (N_19634,N_18303,N_18413);
and U19635 (N_19635,N_17550,N_18425);
and U19636 (N_19636,N_18315,N_17862);
nand U19637 (N_19637,N_18603,N_18468);
and U19638 (N_19638,N_17612,N_17953);
or U19639 (N_19639,N_17694,N_18674);
nand U19640 (N_19640,N_17665,N_18406);
xor U19641 (N_19641,N_18583,N_17877);
or U19642 (N_19642,N_17794,N_18154);
nand U19643 (N_19643,N_17768,N_17809);
nand U19644 (N_19644,N_17765,N_18268);
or U19645 (N_19645,N_18486,N_17671);
and U19646 (N_19646,N_18038,N_17794);
and U19647 (N_19647,N_17888,N_18130);
and U19648 (N_19648,N_18207,N_17576);
xor U19649 (N_19649,N_18469,N_18715);
and U19650 (N_19650,N_18559,N_18114);
and U19651 (N_19651,N_18532,N_18699);
nor U19652 (N_19652,N_17655,N_18107);
or U19653 (N_19653,N_17938,N_18531);
and U19654 (N_19654,N_18517,N_18192);
nand U19655 (N_19655,N_18102,N_18521);
and U19656 (N_19656,N_17814,N_17996);
xnor U19657 (N_19657,N_18609,N_18344);
nand U19658 (N_19658,N_18152,N_18469);
nand U19659 (N_19659,N_17624,N_17574);
and U19660 (N_19660,N_18448,N_18111);
and U19661 (N_19661,N_17503,N_18540);
xor U19662 (N_19662,N_18115,N_17998);
xor U19663 (N_19663,N_17764,N_18314);
and U19664 (N_19664,N_18147,N_18249);
and U19665 (N_19665,N_18266,N_18361);
or U19666 (N_19666,N_17773,N_18401);
nand U19667 (N_19667,N_18639,N_17988);
and U19668 (N_19668,N_18334,N_17879);
nor U19669 (N_19669,N_18272,N_17903);
nand U19670 (N_19670,N_17983,N_18389);
and U19671 (N_19671,N_17531,N_18454);
nand U19672 (N_19672,N_18707,N_18386);
and U19673 (N_19673,N_18312,N_17763);
xor U19674 (N_19674,N_18117,N_17704);
nor U19675 (N_19675,N_18178,N_17734);
nor U19676 (N_19676,N_17839,N_18740);
xor U19677 (N_19677,N_18315,N_18518);
nand U19678 (N_19678,N_18242,N_18596);
and U19679 (N_19679,N_17912,N_18303);
and U19680 (N_19680,N_18650,N_17868);
nor U19681 (N_19681,N_17965,N_18079);
and U19682 (N_19682,N_17843,N_18694);
nor U19683 (N_19683,N_18056,N_17675);
nor U19684 (N_19684,N_18713,N_18042);
and U19685 (N_19685,N_18102,N_18393);
xor U19686 (N_19686,N_18474,N_18575);
nor U19687 (N_19687,N_18665,N_18392);
nor U19688 (N_19688,N_17632,N_18084);
nand U19689 (N_19689,N_17511,N_18299);
xor U19690 (N_19690,N_18730,N_18290);
or U19691 (N_19691,N_18423,N_18393);
xor U19692 (N_19692,N_17624,N_18441);
or U19693 (N_19693,N_18337,N_18606);
nor U19694 (N_19694,N_17540,N_17868);
nor U19695 (N_19695,N_18372,N_18267);
and U19696 (N_19696,N_17871,N_18072);
and U19697 (N_19697,N_17735,N_18090);
and U19698 (N_19698,N_18548,N_17986);
xor U19699 (N_19699,N_17848,N_18649);
or U19700 (N_19700,N_18302,N_18583);
xor U19701 (N_19701,N_17972,N_18654);
nand U19702 (N_19702,N_17721,N_18600);
and U19703 (N_19703,N_18132,N_18734);
nand U19704 (N_19704,N_18074,N_17597);
or U19705 (N_19705,N_18450,N_18594);
nand U19706 (N_19706,N_18082,N_18135);
nand U19707 (N_19707,N_18019,N_18223);
nor U19708 (N_19708,N_18522,N_18555);
xnor U19709 (N_19709,N_17683,N_17824);
nor U19710 (N_19710,N_18658,N_17718);
and U19711 (N_19711,N_18174,N_17704);
and U19712 (N_19712,N_18647,N_17739);
or U19713 (N_19713,N_18591,N_18235);
or U19714 (N_19714,N_18417,N_18497);
nand U19715 (N_19715,N_17922,N_18271);
nor U19716 (N_19716,N_18693,N_18545);
nand U19717 (N_19717,N_17540,N_17543);
xnor U19718 (N_19718,N_18071,N_17648);
and U19719 (N_19719,N_17649,N_18648);
nand U19720 (N_19720,N_17694,N_18622);
nand U19721 (N_19721,N_18652,N_17602);
xor U19722 (N_19722,N_18222,N_18248);
xor U19723 (N_19723,N_18059,N_17708);
and U19724 (N_19724,N_17526,N_18271);
xnor U19725 (N_19725,N_18722,N_18314);
and U19726 (N_19726,N_18021,N_18638);
nand U19727 (N_19727,N_18429,N_17701);
and U19728 (N_19728,N_17743,N_18363);
xnor U19729 (N_19729,N_17887,N_18675);
xnor U19730 (N_19730,N_18388,N_18258);
xor U19731 (N_19731,N_18550,N_18440);
and U19732 (N_19732,N_18727,N_17592);
xor U19733 (N_19733,N_17610,N_18471);
and U19734 (N_19734,N_18285,N_18152);
nor U19735 (N_19735,N_18747,N_17694);
nor U19736 (N_19736,N_17904,N_18042);
and U19737 (N_19737,N_17728,N_17917);
nor U19738 (N_19738,N_18181,N_17696);
xnor U19739 (N_19739,N_18657,N_18342);
nor U19740 (N_19740,N_17500,N_18446);
or U19741 (N_19741,N_18387,N_18202);
nand U19742 (N_19742,N_18710,N_17618);
nand U19743 (N_19743,N_18260,N_18334);
and U19744 (N_19744,N_18190,N_18427);
xor U19745 (N_19745,N_17974,N_18496);
nor U19746 (N_19746,N_17735,N_17909);
or U19747 (N_19747,N_17944,N_18229);
and U19748 (N_19748,N_17578,N_18661);
and U19749 (N_19749,N_17535,N_17978);
nor U19750 (N_19750,N_18635,N_18375);
nand U19751 (N_19751,N_17999,N_17557);
nand U19752 (N_19752,N_18636,N_18368);
xor U19753 (N_19753,N_17965,N_18685);
xnor U19754 (N_19754,N_17762,N_18318);
nand U19755 (N_19755,N_17530,N_17662);
nand U19756 (N_19756,N_17690,N_17620);
and U19757 (N_19757,N_18569,N_17940);
or U19758 (N_19758,N_18305,N_18415);
or U19759 (N_19759,N_17537,N_18303);
and U19760 (N_19760,N_18743,N_18308);
nand U19761 (N_19761,N_18584,N_18611);
nand U19762 (N_19762,N_17507,N_18137);
or U19763 (N_19763,N_17544,N_18397);
or U19764 (N_19764,N_17668,N_17538);
nand U19765 (N_19765,N_18031,N_18112);
xor U19766 (N_19766,N_17588,N_18526);
nor U19767 (N_19767,N_18121,N_18344);
or U19768 (N_19768,N_17524,N_18676);
and U19769 (N_19769,N_18346,N_18121);
or U19770 (N_19770,N_18028,N_17970);
and U19771 (N_19771,N_18088,N_18485);
or U19772 (N_19772,N_18635,N_18522);
nor U19773 (N_19773,N_17697,N_17992);
nand U19774 (N_19774,N_18390,N_17822);
or U19775 (N_19775,N_18062,N_17642);
nor U19776 (N_19776,N_18744,N_17995);
nand U19777 (N_19777,N_17869,N_17774);
or U19778 (N_19778,N_17606,N_18239);
or U19779 (N_19779,N_17630,N_18609);
or U19780 (N_19780,N_17830,N_17645);
nor U19781 (N_19781,N_17957,N_18029);
nor U19782 (N_19782,N_17868,N_17808);
and U19783 (N_19783,N_17509,N_18736);
nand U19784 (N_19784,N_17540,N_18737);
and U19785 (N_19785,N_17998,N_18259);
nor U19786 (N_19786,N_18248,N_18555);
and U19787 (N_19787,N_17748,N_17596);
or U19788 (N_19788,N_18332,N_18036);
nor U19789 (N_19789,N_18033,N_18162);
nand U19790 (N_19790,N_17937,N_18258);
and U19791 (N_19791,N_17535,N_18259);
nand U19792 (N_19792,N_18116,N_17527);
and U19793 (N_19793,N_18313,N_17961);
or U19794 (N_19794,N_18679,N_17654);
nand U19795 (N_19795,N_18059,N_18333);
or U19796 (N_19796,N_18736,N_18452);
or U19797 (N_19797,N_18421,N_18237);
nor U19798 (N_19798,N_17949,N_18339);
or U19799 (N_19799,N_17729,N_18027);
or U19800 (N_19800,N_18116,N_18065);
xor U19801 (N_19801,N_17558,N_18255);
and U19802 (N_19802,N_18334,N_18667);
or U19803 (N_19803,N_18217,N_18322);
or U19804 (N_19804,N_17800,N_18675);
and U19805 (N_19805,N_17921,N_18082);
xor U19806 (N_19806,N_18162,N_18034);
nor U19807 (N_19807,N_17506,N_17638);
nand U19808 (N_19808,N_18312,N_18035);
or U19809 (N_19809,N_17853,N_18501);
or U19810 (N_19810,N_17839,N_17922);
or U19811 (N_19811,N_18004,N_17521);
nand U19812 (N_19812,N_17726,N_18176);
or U19813 (N_19813,N_18230,N_17795);
or U19814 (N_19814,N_17903,N_17928);
xnor U19815 (N_19815,N_17717,N_18259);
xor U19816 (N_19816,N_17832,N_18058);
nand U19817 (N_19817,N_18033,N_18570);
nor U19818 (N_19818,N_18397,N_17537);
and U19819 (N_19819,N_17891,N_18592);
xor U19820 (N_19820,N_18637,N_17580);
or U19821 (N_19821,N_18075,N_17738);
nor U19822 (N_19822,N_17554,N_17647);
xnor U19823 (N_19823,N_18331,N_17836);
nor U19824 (N_19824,N_18272,N_17909);
nor U19825 (N_19825,N_18472,N_18687);
and U19826 (N_19826,N_17746,N_18198);
and U19827 (N_19827,N_18224,N_17938);
nand U19828 (N_19828,N_17634,N_18014);
nor U19829 (N_19829,N_18004,N_18680);
or U19830 (N_19830,N_17574,N_18440);
and U19831 (N_19831,N_18661,N_18454);
nor U19832 (N_19832,N_18180,N_18308);
and U19833 (N_19833,N_18262,N_17799);
and U19834 (N_19834,N_18524,N_18066);
nand U19835 (N_19835,N_18054,N_18465);
or U19836 (N_19836,N_18507,N_18556);
nand U19837 (N_19837,N_17535,N_18710);
xnor U19838 (N_19838,N_17822,N_17919);
nor U19839 (N_19839,N_17528,N_18151);
nand U19840 (N_19840,N_17702,N_18473);
nand U19841 (N_19841,N_17517,N_18377);
nor U19842 (N_19842,N_17935,N_17939);
or U19843 (N_19843,N_17614,N_18590);
nor U19844 (N_19844,N_18649,N_17803);
nor U19845 (N_19845,N_18033,N_18465);
xor U19846 (N_19846,N_17936,N_17825);
nand U19847 (N_19847,N_17801,N_18043);
or U19848 (N_19848,N_18166,N_18051);
and U19849 (N_19849,N_18168,N_18393);
nor U19850 (N_19850,N_18344,N_17791);
nand U19851 (N_19851,N_18510,N_18143);
nor U19852 (N_19852,N_17615,N_18419);
nand U19853 (N_19853,N_18030,N_18378);
nor U19854 (N_19854,N_17851,N_17609);
nand U19855 (N_19855,N_17550,N_17927);
xnor U19856 (N_19856,N_18607,N_18353);
or U19857 (N_19857,N_18392,N_18166);
or U19858 (N_19858,N_18478,N_17860);
nor U19859 (N_19859,N_17828,N_17801);
and U19860 (N_19860,N_18395,N_17756);
xor U19861 (N_19861,N_18004,N_17861);
nor U19862 (N_19862,N_18607,N_18680);
xnor U19863 (N_19863,N_17665,N_17583);
or U19864 (N_19864,N_18006,N_17694);
nor U19865 (N_19865,N_18024,N_18278);
or U19866 (N_19866,N_18035,N_18179);
nand U19867 (N_19867,N_18610,N_17636);
and U19868 (N_19868,N_18747,N_17528);
xnor U19869 (N_19869,N_18644,N_17836);
or U19870 (N_19870,N_17802,N_18132);
or U19871 (N_19871,N_18590,N_18410);
or U19872 (N_19872,N_17645,N_17632);
and U19873 (N_19873,N_17842,N_18222);
and U19874 (N_19874,N_17640,N_18556);
and U19875 (N_19875,N_17720,N_18093);
nand U19876 (N_19876,N_17984,N_18127);
xnor U19877 (N_19877,N_18196,N_17709);
and U19878 (N_19878,N_17554,N_17790);
and U19879 (N_19879,N_18459,N_17926);
and U19880 (N_19880,N_18029,N_17620);
xor U19881 (N_19881,N_17543,N_18670);
xor U19882 (N_19882,N_18568,N_17690);
nor U19883 (N_19883,N_17568,N_18013);
xnor U19884 (N_19884,N_18447,N_18670);
and U19885 (N_19885,N_17880,N_18081);
xnor U19886 (N_19886,N_17925,N_18604);
and U19887 (N_19887,N_17996,N_18728);
and U19888 (N_19888,N_17856,N_18300);
nor U19889 (N_19889,N_17927,N_18686);
nand U19890 (N_19890,N_17968,N_18665);
nor U19891 (N_19891,N_17728,N_17534);
nand U19892 (N_19892,N_18071,N_18398);
nor U19893 (N_19893,N_18566,N_18620);
and U19894 (N_19894,N_18531,N_18202);
nand U19895 (N_19895,N_18186,N_18328);
xnor U19896 (N_19896,N_18007,N_18584);
nor U19897 (N_19897,N_17779,N_18188);
xnor U19898 (N_19898,N_17508,N_17960);
xor U19899 (N_19899,N_18031,N_18680);
xnor U19900 (N_19900,N_18544,N_17628);
xor U19901 (N_19901,N_17558,N_17662);
or U19902 (N_19902,N_18057,N_17587);
nor U19903 (N_19903,N_17937,N_17800);
nor U19904 (N_19904,N_17689,N_18267);
nor U19905 (N_19905,N_18420,N_18236);
xor U19906 (N_19906,N_17626,N_18072);
xor U19907 (N_19907,N_17559,N_18093);
nand U19908 (N_19908,N_18343,N_17664);
nor U19909 (N_19909,N_18590,N_17895);
nand U19910 (N_19910,N_18473,N_17870);
and U19911 (N_19911,N_18119,N_17906);
or U19912 (N_19912,N_18215,N_18099);
nor U19913 (N_19913,N_18675,N_18056);
and U19914 (N_19914,N_18234,N_17914);
or U19915 (N_19915,N_17823,N_17908);
nand U19916 (N_19916,N_18157,N_18201);
and U19917 (N_19917,N_17698,N_18394);
xor U19918 (N_19918,N_18115,N_18546);
and U19919 (N_19919,N_17590,N_17625);
nor U19920 (N_19920,N_17603,N_18443);
nor U19921 (N_19921,N_18095,N_17846);
or U19922 (N_19922,N_18512,N_18444);
xor U19923 (N_19923,N_18509,N_17954);
or U19924 (N_19924,N_17600,N_18135);
nand U19925 (N_19925,N_18330,N_17848);
or U19926 (N_19926,N_18192,N_17878);
and U19927 (N_19927,N_17852,N_17814);
xor U19928 (N_19928,N_18297,N_18304);
xnor U19929 (N_19929,N_18381,N_17778);
nand U19930 (N_19930,N_18714,N_18567);
or U19931 (N_19931,N_17917,N_17707);
and U19932 (N_19932,N_17670,N_17820);
and U19933 (N_19933,N_17705,N_18135);
nor U19934 (N_19934,N_18361,N_18066);
nand U19935 (N_19935,N_17780,N_18546);
or U19936 (N_19936,N_18233,N_18687);
or U19937 (N_19937,N_18389,N_18233);
nor U19938 (N_19938,N_17747,N_18124);
xnor U19939 (N_19939,N_18730,N_18647);
xnor U19940 (N_19940,N_18611,N_17996);
nand U19941 (N_19941,N_17745,N_17779);
nor U19942 (N_19942,N_17529,N_18261);
or U19943 (N_19943,N_18284,N_18044);
nor U19944 (N_19944,N_18198,N_18451);
nand U19945 (N_19945,N_18396,N_17945);
nand U19946 (N_19946,N_18724,N_17827);
nand U19947 (N_19947,N_18622,N_17988);
and U19948 (N_19948,N_18709,N_18223);
nor U19949 (N_19949,N_17535,N_18212);
and U19950 (N_19950,N_18204,N_18169);
or U19951 (N_19951,N_17749,N_17950);
and U19952 (N_19952,N_17968,N_18016);
xnor U19953 (N_19953,N_18682,N_18442);
or U19954 (N_19954,N_18351,N_18210);
nand U19955 (N_19955,N_17885,N_18630);
nor U19956 (N_19956,N_18527,N_18331);
or U19957 (N_19957,N_18314,N_18038);
nand U19958 (N_19958,N_18566,N_18407);
nand U19959 (N_19959,N_18619,N_17587);
nand U19960 (N_19960,N_17850,N_17523);
xnor U19961 (N_19961,N_18696,N_17685);
xnor U19962 (N_19962,N_18319,N_18652);
xnor U19963 (N_19963,N_17768,N_17765);
nand U19964 (N_19964,N_17989,N_18150);
xor U19965 (N_19965,N_17536,N_18202);
or U19966 (N_19966,N_17640,N_17963);
or U19967 (N_19967,N_17789,N_18168);
or U19968 (N_19968,N_18171,N_17786);
nand U19969 (N_19969,N_18673,N_17688);
nand U19970 (N_19970,N_18350,N_18371);
and U19971 (N_19971,N_18348,N_18059);
and U19972 (N_19972,N_18067,N_18196);
and U19973 (N_19973,N_17885,N_18204);
nor U19974 (N_19974,N_18432,N_17557);
and U19975 (N_19975,N_18019,N_17878);
nor U19976 (N_19976,N_18666,N_18003);
nand U19977 (N_19977,N_17893,N_18157);
and U19978 (N_19978,N_18214,N_18692);
and U19979 (N_19979,N_17941,N_18207);
nor U19980 (N_19980,N_18480,N_18412);
xor U19981 (N_19981,N_18306,N_18434);
or U19982 (N_19982,N_17996,N_17605);
nand U19983 (N_19983,N_17929,N_17741);
nor U19984 (N_19984,N_18728,N_18317);
nor U19985 (N_19985,N_18119,N_18473);
xor U19986 (N_19986,N_17865,N_18191);
nand U19987 (N_19987,N_18644,N_17922);
or U19988 (N_19988,N_18382,N_18197);
xor U19989 (N_19989,N_18358,N_18357);
xor U19990 (N_19990,N_18039,N_18415);
or U19991 (N_19991,N_18696,N_18633);
nand U19992 (N_19992,N_17715,N_17702);
or U19993 (N_19993,N_17610,N_18704);
xnor U19994 (N_19994,N_17946,N_17666);
or U19995 (N_19995,N_17503,N_18305);
nand U19996 (N_19996,N_17838,N_18307);
or U19997 (N_19997,N_18175,N_18540);
nand U19998 (N_19998,N_18696,N_17822);
or U19999 (N_19999,N_17543,N_18730);
or U20000 (N_20000,N_19666,N_19959);
or U20001 (N_20001,N_19095,N_19688);
and U20002 (N_20002,N_19555,N_19043);
nand U20003 (N_20003,N_18824,N_19971);
nor U20004 (N_20004,N_19753,N_19827);
nand U20005 (N_20005,N_18788,N_19149);
nor U20006 (N_20006,N_19842,N_19854);
nand U20007 (N_20007,N_18910,N_19157);
nand U20008 (N_20008,N_19447,N_18841);
and U20009 (N_20009,N_19075,N_19328);
and U20010 (N_20010,N_19796,N_19798);
or U20011 (N_20011,N_19805,N_19445);
xnor U20012 (N_20012,N_18805,N_19623);
and U20013 (N_20013,N_19893,N_18772);
xnor U20014 (N_20014,N_19776,N_19803);
nand U20015 (N_20015,N_19984,N_19215);
xnor U20016 (N_20016,N_19271,N_19812);
and U20017 (N_20017,N_19383,N_19404);
xnor U20018 (N_20018,N_19579,N_19491);
nor U20019 (N_20019,N_18804,N_19477);
and U20020 (N_20020,N_19542,N_19539);
or U20021 (N_20021,N_19218,N_19444);
nor U20022 (N_20022,N_19018,N_19860);
nand U20023 (N_20023,N_19127,N_19394);
and U20024 (N_20024,N_19606,N_19918);
or U20025 (N_20025,N_19686,N_19137);
or U20026 (N_20026,N_19675,N_19158);
and U20027 (N_20027,N_19638,N_19933);
or U20028 (N_20028,N_19395,N_18792);
nand U20029 (N_20029,N_19020,N_19295);
xnor U20030 (N_20030,N_19829,N_19197);
xor U20031 (N_20031,N_19389,N_19219);
and U20032 (N_20032,N_19924,N_19031);
and U20033 (N_20033,N_18818,N_18832);
xor U20034 (N_20034,N_19713,N_19000);
and U20035 (N_20035,N_19265,N_18908);
and U20036 (N_20036,N_19093,N_19490);
and U20037 (N_20037,N_19493,N_19278);
nor U20038 (N_20038,N_19844,N_19837);
nand U20039 (N_20039,N_18996,N_19501);
xnor U20040 (N_20040,N_19706,N_19629);
nor U20041 (N_20041,N_19177,N_19474);
nor U20042 (N_20042,N_19921,N_19572);
or U20043 (N_20043,N_18813,N_19712);
or U20044 (N_20044,N_19139,N_19225);
nand U20045 (N_20045,N_18885,N_19014);
nand U20046 (N_20046,N_18790,N_19125);
nand U20047 (N_20047,N_18958,N_19897);
and U20048 (N_20048,N_19355,N_19274);
nor U20049 (N_20049,N_19323,N_19154);
nor U20050 (N_20050,N_19305,N_19524);
nor U20051 (N_20051,N_18897,N_19540);
xnor U20052 (N_20052,N_19636,N_19815);
nand U20053 (N_20053,N_18859,N_19683);
nor U20054 (N_20054,N_19207,N_19496);
or U20055 (N_20055,N_19202,N_19301);
xnor U20056 (N_20056,N_19546,N_19859);
nor U20057 (N_20057,N_19864,N_19588);
and U20058 (N_20058,N_19571,N_18932);
and U20059 (N_20059,N_19168,N_19567);
nor U20060 (N_20060,N_19169,N_19433);
xnor U20061 (N_20061,N_19724,N_19267);
and U20062 (N_20062,N_19610,N_19104);
or U20063 (N_20063,N_19242,N_18839);
or U20064 (N_20064,N_19845,N_19819);
xnor U20065 (N_20065,N_19049,N_18759);
nand U20066 (N_20066,N_19699,N_19937);
nor U20067 (N_20067,N_18942,N_19377);
nand U20068 (N_20068,N_19966,N_19160);
nor U20069 (N_20069,N_19528,N_19547);
and U20070 (N_20070,N_19254,N_19703);
or U20071 (N_20071,N_18887,N_18921);
or U20072 (N_20072,N_18969,N_19998);
xor U20073 (N_20073,N_19601,N_19633);
or U20074 (N_20074,N_19064,N_19578);
or U20075 (N_20075,N_18871,N_19269);
nand U20076 (N_20076,N_19044,N_19804);
xor U20077 (N_20077,N_19670,N_19485);
nor U20078 (N_20078,N_18778,N_19058);
or U20079 (N_20079,N_19416,N_19928);
nor U20080 (N_20080,N_19917,N_19153);
nand U20081 (N_20081,N_19620,N_19194);
and U20082 (N_20082,N_19236,N_19308);
nand U20083 (N_20083,N_19521,N_19660);
or U20084 (N_20084,N_19087,N_19599);
or U20085 (N_20085,N_19658,N_19942);
and U20086 (N_20086,N_19584,N_18856);
nand U20087 (N_20087,N_19604,N_19347);
or U20088 (N_20088,N_18828,N_18931);
nor U20089 (N_20089,N_19861,N_18909);
xnor U20090 (N_20090,N_19936,N_18926);
nand U20091 (N_20091,N_19988,N_19097);
nand U20092 (N_20092,N_19920,N_18893);
xnor U20093 (N_20093,N_19339,N_19500);
nand U20094 (N_20094,N_19820,N_18928);
or U20095 (N_20095,N_18999,N_19028);
nand U20096 (N_20096,N_18806,N_19226);
nand U20097 (N_20097,N_18915,N_19009);
xnor U20098 (N_20098,N_19774,N_19392);
nand U20099 (N_20099,N_18853,N_18929);
nor U20100 (N_20100,N_19746,N_19237);
nand U20101 (N_20101,N_19553,N_18793);
nor U20102 (N_20102,N_18950,N_19007);
nand U20103 (N_20103,N_19905,N_18782);
nor U20104 (N_20104,N_19580,N_19507);
nor U20105 (N_20105,N_18940,N_19786);
nand U20106 (N_20106,N_19078,N_19875);
or U20107 (N_20107,N_19250,N_19630);
nor U20108 (N_20108,N_19109,N_19212);
nand U20109 (N_20109,N_18982,N_19282);
or U20110 (N_20110,N_18970,N_19489);
xor U20111 (N_20111,N_19256,N_19784);
nand U20112 (N_20112,N_19129,N_19431);
or U20113 (N_20113,N_18924,N_19393);
and U20114 (N_20114,N_19639,N_19053);
nand U20115 (N_20115,N_19478,N_18811);
and U20116 (N_20116,N_19895,N_18923);
or U20117 (N_20117,N_19674,N_19464);
and U20118 (N_20118,N_18937,N_19326);
nor U20119 (N_20119,N_19742,N_19340);
xnor U20120 (N_20120,N_19557,N_18842);
and U20121 (N_20121,N_19698,N_18765);
nor U20122 (N_20122,N_19626,N_19329);
and U20123 (N_20123,N_19082,N_19611);
nand U20124 (N_20124,N_19946,N_19901);
nand U20125 (N_20125,N_19608,N_18836);
nor U20126 (N_20126,N_19065,N_19973);
nor U20127 (N_20127,N_18868,N_18873);
or U20128 (N_20128,N_19963,N_19899);
or U20129 (N_20129,N_19067,N_19843);
xnor U20130 (N_20130,N_19915,N_18878);
and U20131 (N_20131,N_19165,N_19307);
and U20132 (N_20132,N_19051,N_19298);
xnor U20133 (N_20133,N_19642,N_19126);
xor U20134 (N_20134,N_19766,N_19440);
or U20135 (N_20135,N_19970,N_19257);
or U20136 (N_20136,N_19791,N_19617);
and U20137 (N_20137,N_19881,N_19775);
nor U20138 (N_20138,N_19759,N_19175);
or U20139 (N_20139,N_19529,N_19909);
nand U20140 (N_20140,N_19371,N_19330);
xnor U20141 (N_20141,N_19927,N_19132);
nor U20142 (N_20142,N_19466,N_18852);
xnor U20143 (N_20143,N_19799,N_18976);
nand U20144 (N_20144,N_19955,N_19726);
or U20145 (N_20145,N_18857,N_19982);
or U20146 (N_20146,N_19613,N_19284);
nand U20147 (N_20147,N_19084,N_19332);
and U20148 (N_20148,N_19600,N_19564);
or U20149 (N_20149,N_18860,N_19554);
nor U20150 (N_20150,N_19708,N_18957);
nand U20151 (N_20151,N_19645,N_19164);
or U20152 (N_20152,N_19400,N_19846);
xnor U20153 (N_20153,N_19516,N_19076);
and U20154 (N_20154,N_19107,N_19460);
or U20155 (N_20155,N_19072,N_19193);
nor U20156 (N_20156,N_19628,N_19956);
nand U20157 (N_20157,N_19800,N_19593);
nor U20158 (N_20158,N_19213,N_19810);
or U20159 (N_20159,N_19720,N_18762);
nand U20160 (N_20160,N_19890,N_19405);
or U20161 (N_20161,N_19381,N_19052);
xor U20162 (N_20162,N_19693,N_19309);
and U20163 (N_20163,N_19446,N_19756);
and U20164 (N_20164,N_19740,N_19372);
and U20165 (N_20165,N_19866,N_19480);
nand U20166 (N_20166,N_18858,N_18954);
nand U20167 (N_20167,N_19867,N_18851);
nor U20168 (N_20168,N_19731,N_19486);
or U20169 (N_20169,N_19525,N_19981);
nor U20170 (N_20170,N_18930,N_19352);
xnor U20171 (N_20171,N_19575,N_19430);
and U20172 (N_20172,N_19426,N_19935);
xor U20173 (N_20173,N_18833,N_19681);
xor U20174 (N_20174,N_19908,N_19987);
nor U20175 (N_20175,N_18819,N_19417);
and U20176 (N_20176,N_19481,N_18879);
xnor U20177 (N_20177,N_19900,N_18994);
or U20178 (N_20178,N_19318,N_18768);
xor U20179 (N_20179,N_19163,N_19989);
and U20180 (N_20180,N_18964,N_18935);
xnor U20181 (N_20181,N_18927,N_18773);
nand U20182 (N_20182,N_19378,N_19025);
or U20183 (N_20183,N_19437,N_19889);
or U20184 (N_20184,N_19527,N_18870);
or U20185 (N_20185,N_18945,N_18801);
nor U20186 (N_20186,N_19349,N_19513);
xnor U20187 (N_20187,N_18803,N_19824);
and U20188 (N_20188,N_18980,N_19131);
nor U20189 (N_20189,N_19559,N_19316);
and U20190 (N_20190,N_19427,N_19865);
and U20191 (N_20191,N_18786,N_19324);
and U20192 (N_20192,N_19607,N_19229);
xor U20193 (N_20193,N_19035,N_19596);
nor U20194 (N_20194,N_18830,N_19764);
or U20195 (N_20195,N_19632,N_19692);
nand U20196 (N_20196,N_19855,N_19128);
nand U20197 (N_20197,N_19336,N_19133);
nand U20198 (N_20198,N_19587,N_19190);
nor U20199 (N_20199,N_18750,N_19813);
nand U20200 (N_20200,N_18906,N_19839);
and U20201 (N_20201,N_19090,N_19765);
or U20202 (N_20202,N_19678,N_19958);
or U20203 (N_20203,N_19353,N_19522);
nand U20204 (N_20204,N_19105,N_19436);
and U20205 (N_20205,N_19398,N_19047);
nor U20206 (N_20206,N_18877,N_19577);
or U20207 (N_20207,N_19360,N_18884);
nand U20208 (N_20208,N_19003,N_19231);
or U20209 (N_20209,N_18767,N_18962);
nor U20210 (N_20210,N_19022,N_19291);
xor U20211 (N_20211,N_19173,N_19140);
nand U20212 (N_20212,N_19983,N_18952);
and U20213 (N_20213,N_18894,N_19010);
or U20214 (N_20214,N_19245,N_19871);
nand U20215 (N_20215,N_19004,N_18829);
xnor U20216 (N_20216,N_18876,N_19055);
xnor U20217 (N_20217,N_18796,N_19406);
nor U20218 (N_20218,N_18881,N_19467);
xor U20219 (N_20219,N_19710,N_19755);
or U20220 (N_20220,N_19648,N_19171);
nand U20221 (N_20221,N_19502,N_19411);
or U20222 (N_20222,N_19979,N_19618);
or U20223 (N_20223,N_18903,N_19880);
nor U20224 (N_20224,N_19985,N_19877);
and U20225 (N_20225,N_19365,N_19359);
and U20226 (N_20226,N_19387,N_19224);
nor U20227 (N_20227,N_18874,N_18752);
nand U20228 (N_20228,N_19705,N_19672);
xnor U20229 (N_20229,N_18972,N_19509);
nor U20230 (N_20230,N_18902,N_19566);
nand U20231 (N_20231,N_19120,N_19299);
or U20232 (N_20232,N_19386,N_19719);
nor U20233 (N_20233,N_19422,N_19376);
nand U20234 (N_20234,N_19576,N_19621);
nand U20235 (N_20235,N_19399,N_19801);
or U20236 (N_20236,N_19814,N_19530);
or U20237 (N_20237,N_19325,N_19272);
nor U20238 (N_20238,N_19320,N_19993);
or U20239 (N_20239,N_19156,N_18785);
xor U20240 (N_20240,N_19737,N_19066);
xnor U20241 (N_20241,N_19828,N_18948);
nand U20242 (N_20242,N_19694,N_19531);
nor U20243 (N_20243,N_19655,N_19954);
nor U20244 (N_20244,N_18986,N_19721);
nand U20245 (N_20245,N_19362,N_19734);
nor U20246 (N_20246,N_19421,N_19255);
xor U20247 (N_20247,N_19735,N_19147);
and U20248 (N_20248,N_18889,N_19709);
nor U20249 (N_20249,N_19560,N_19410);
and U20250 (N_20250,N_19117,N_18774);
xnor U20251 (N_20251,N_18783,N_19728);
nand U20252 (N_20252,N_19045,N_19586);
nor U20253 (N_20253,N_19170,N_19281);
nor U20254 (N_20254,N_18934,N_19488);
or U20255 (N_20255,N_19263,N_19034);
xnor U20256 (N_20256,N_18872,N_19906);
nor U20257 (N_20257,N_19960,N_18900);
nor U20258 (N_20258,N_19641,N_19346);
xor U20259 (N_20259,N_19515,N_19184);
or U20260 (N_20260,N_19779,N_18760);
and U20261 (N_20261,N_19382,N_19280);
nor U20262 (N_20262,N_19196,N_19852);
nor U20263 (N_20263,N_18892,N_19614);
or U20264 (N_20264,N_19057,N_19634);
nor U20265 (N_20265,N_19858,N_19585);
xor U20266 (N_20266,N_18985,N_19419);
and U20267 (N_20267,N_18754,N_18867);
nand U20268 (N_20268,N_18770,N_19101);
and U20269 (N_20269,N_18941,N_19150);
nor U20270 (N_20270,N_19717,N_19294);
or U20271 (N_20271,N_19304,N_19931);
or U20272 (N_20272,N_18756,N_19873);
and U20273 (N_20273,N_19220,N_18864);
nor U20274 (N_20274,N_19646,N_19403);
and U20275 (N_20275,N_19733,N_18763);
xor U20276 (N_20276,N_19947,N_19391);
xor U20277 (N_20277,N_19050,N_19448);
nand U20278 (N_20278,N_19006,N_19402);
xnor U20279 (N_20279,N_19762,N_19874);
nor U20280 (N_20280,N_19232,N_19943);
xor U20281 (N_20281,N_19870,N_19950);
xnor U20282 (N_20282,N_19597,N_19505);
nor U20283 (N_20283,N_19697,N_19754);
nor U20284 (N_20284,N_19289,N_19741);
or U20285 (N_20285,N_19206,N_19130);
nor U20286 (N_20286,N_19806,N_19653);
nor U20287 (N_20287,N_19195,N_19744);
xnor U20288 (N_20288,N_19777,N_19696);
and U20289 (N_20289,N_19707,N_19986);
nor U20290 (N_20290,N_18998,N_19743);
and U20291 (N_20291,N_19227,N_19262);
or U20292 (N_20292,N_19470,N_19913);
nor U20293 (N_20293,N_19757,N_19968);
nand U20294 (N_20294,N_19663,N_19487);
and U20295 (N_20295,N_19100,N_18826);
xnor U20296 (N_20296,N_19583,N_18820);
nor U20297 (N_20297,N_19662,N_18850);
or U20298 (N_20298,N_19081,N_19676);
nor U20299 (N_20299,N_18775,N_19356);
xor U20300 (N_20300,N_19367,N_18978);
xnor U20301 (N_20301,N_18914,N_19518);
or U20302 (N_20302,N_18955,N_19079);
and U20303 (N_20303,N_19322,N_19119);
or U20304 (N_20304,N_18827,N_18837);
nor U20305 (N_20305,N_19581,N_19283);
xnor U20306 (N_20306,N_19181,N_19342);
xnor U20307 (N_20307,N_19241,N_19450);
nand U20308 (N_20308,N_19162,N_19461);
nand U20309 (N_20309,N_19499,N_19974);
xnor U20310 (N_20310,N_19664,N_19545);
and U20311 (N_20311,N_19351,N_19136);
or U20312 (N_20312,N_19673,N_19514);
nand U20313 (N_20313,N_18863,N_19166);
nor U20314 (N_20314,N_19285,N_19551);
nand U20315 (N_20315,N_19135,N_19923);
and U20316 (N_20316,N_19767,N_19046);
and U20317 (N_20317,N_18875,N_19401);
or U20318 (N_20318,N_19040,N_19538);
or U20319 (N_20319,N_18771,N_19727);
and U20320 (N_20320,N_19335,N_19121);
nor U20321 (N_20321,N_19293,N_19725);
nor U20322 (N_20322,N_19159,N_18797);
nand U20323 (N_20323,N_19483,N_19442);
xnor U20324 (N_20324,N_18789,N_19103);
nor U20325 (N_20325,N_18944,N_19465);
and U20326 (N_20326,N_19822,N_18947);
or U20327 (N_20327,N_19114,N_18855);
nand U20328 (N_20328,N_19428,N_19615);
and U20329 (N_20329,N_19244,N_18917);
nor U20330 (N_20330,N_19124,N_19823);
xor U20331 (N_20331,N_19234,N_19223);
nand U20332 (N_20332,N_19957,N_18794);
nand U20333 (N_20333,N_19235,N_19826);
nor U20334 (N_20334,N_18854,N_19691);
nor U20335 (N_20335,N_19134,N_18835);
or U20336 (N_20336,N_19209,N_19690);
nand U20337 (N_20337,N_19669,N_19677);
nand U20338 (N_20338,N_19520,N_19408);
nand U20339 (N_20339,N_19992,N_19476);
nand U20340 (N_20340,N_19198,N_19102);
xnor U20341 (N_20341,N_19793,N_19005);
and U20342 (N_20342,N_19438,N_19296);
or U20343 (N_20343,N_19687,N_19167);
and U20344 (N_20344,N_18951,N_18791);
or U20345 (N_20345,N_19763,N_19965);
nor U20346 (N_20346,N_19747,N_19680);
or U20347 (N_20347,N_18844,N_19337);
and U20348 (N_20348,N_19882,N_19794);
nor U20349 (N_20349,N_19062,N_19785);
nand U20350 (N_20350,N_19247,N_18777);
and U20351 (N_20351,N_19178,N_19449);
and U20352 (N_20352,N_18987,N_18869);
or U20353 (N_20353,N_19385,N_19598);
or U20354 (N_20354,N_19185,N_19856);
or U20355 (N_20355,N_19217,N_19379);
nor U20356 (N_20356,N_19848,N_19469);
and U20357 (N_20357,N_18846,N_19056);
and U20358 (N_20358,N_18808,N_19013);
nand U20359 (N_20359,N_19199,N_19647);
and U20360 (N_20360,N_18848,N_19967);
xnor U20361 (N_20361,N_18784,N_18988);
nand U20362 (N_20362,N_19661,N_19659);
or U20363 (N_20363,N_19711,N_19919);
or U20364 (N_20364,N_19644,N_19825);
and U20365 (N_20365,N_18925,N_18973);
nand U20366 (N_20366,N_19484,N_19434);
nand U20367 (N_20367,N_18781,N_19701);
nand U20368 (N_20368,N_19457,N_19111);
and U20369 (N_20369,N_19768,N_19369);
nand U20370 (N_20370,N_19543,N_19907);
xor U20371 (N_20371,N_19068,N_19432);
xnor U20372 (N_20372,N_19652,N_19952);
nand U20373 (N_20373,N_19504,N_19695);
nand U20374 (N_20374,N_19038,N_19573);
nor U20375 (N_20375,N_19073,N_19321);
or U20376 (N_20376,N_18861,N_19962);
xor U20377 (N_20377,N_19344,N_19558);
xor U20378 (N_20378,N_19331,N_19668);
nand U20379 (N_20379,N_18912,N_19279);
nand U20380 (N_20380,N_18776,N_18907);
and U20381 (N_20381,N_19722,N_19074);
nor U20382 (N_20382,N_19667,N_19180);
xnor U20383 (N_20383,N_18769,N_19603);
nor U20384 (N_20384,N_19780,N_19561);
and U20385 (N_20385,N_19818,N_19210);
or U20386 (N_20386,N_19736,N_19704);
or U20387 (N_20387,N_19468,N_18966);
nor U20388 (N_20388,N_19758,N_19334);
or U20389 (N_20389,N_19083,N_19361);
nand U20390 (N_20390,N_19182,N_19495);
nand U20391 (N_20391,N_19769,N_19790);
nand U20392 (N_20392,N_19243,N_18898);
or U20393 (N_20393,N_18840,N_19650);
nor U20394 (N_20394,N_18822,N_19749);
nor U20395 (N_20395,N_18920,N_19789);
and U20396 (N_20396,N_19479,N_19788);
nor U20397 (N_20397,N_19418,N_18904);
nor U20398 (N_20398,N_19751,N_19266);
xnor U20399 (N_20399,N_19649,N_19685);
and U20400 (N_20400,N_18971,N_19904);
nor U20401 (N_20401,N_19302,N_19851);
or U20402 (N_20402,N_18938,N_18984);
nand U20403 (N_20403,N_19192,N_19876);
xor U20404 (N_20404,N_19635,N_18817);
and U20405 (N_20405,N_19951,N_19602);
xor U20406 (N_20406,N_19240,N_18891);
or U20407 (N_20407,N_19248,N_19214);
xnor U20408 (N_20408,N_19834,N_19333);
and U20409 (N_20409,N_18787,N_19016);
or U20410 (N_20410,N_19407,N_19783);
and U20411 (N_20411,N_19482,N_19995);
xor U20412 (N_20412,N_18816,N_19060);
nand U20413 (N_20413,N_19884,N_19930);
xnor U20414 (N_20414,N_19510,N_19397);
nand U20415 (N_20415,N_19143,N_19179);
nand U20416 (N_20416,N_19222,N_19589);
xnor U20417 (N_20417,N_19473,N_19249);
and U20418 (N_20418,N_19938,N_19413);
or U20419 (N_20419,N_19976,N_19868);
or U20420 (N_20420,N_19886,N_19463);
and U20421 (N_20421,N_18949,N_18758);
and U20422 (N_20422,N_19024,N_18896);
nor U20423 (N_20423,N_19141,N_19850);
and U20424 (N_20424,N_19435,N_19108);
nor U20425 (N_20425,N_19273,N_19089);
or U20426 (N_20426,N_19631,N_18974);
and U20427 (N_20427,N_18802,N_19570);
nor U20428 (N_20428,N_19781,N_19363);
or U20429 (N_20429,N_19714,N_19311);
and U20430 (N_20430,N_19679,N_19239);
nor U20431 (N_20431,N_19017,N_18753);
and U20432 (N_20432,N_19230,N_18899);
nor U20433 (N_20433,N_19991,N_19999);
or U20434 (N_20434,N_19021,N_19503);
xnor U20435 (N_20435,N_19903,N_18968);
or U20436 (N_20436,N_19452,N_19313);
nor U20437 (N_20437,N_19750,N_19552);
xor U20438 (N_20438,N_19816,N_19898);
nor U20439 (N_20439,N_19896,N_19723);
nor U20440 (N_20440,N_18809,N_19384);
and U20441 (N_20441,N_19287,N_19972);
xnor U20442 (N_20442,N_19412,N_19350);
nand U20443 (N_20443,N_19116,N_19071);
or U20444 (N_20444,N_19032,N_19787);
or U20445 (N_20445,N_19592,N_18866);
nand U20446 (N_20446,N_19745,N_19715);
or U20447 (N_20447,N_18779,N_18960);
and U20448 (N_20448,N_19145,N_19375);
or U20449 (N_20449,N_19259,N_19792);
nor U20450 (N_20450,N_19548,N_18849);
and U20451 (N_20451,N_19830,N_19425);
xnor U20452 (N_20452,N_18993,N_19811);
xor U20453 (N_20453,N_18933,N_19622);
nor U20454 (N_20454,N_19494,N_19569);
nor U20455 (N_20455,N_19926,N_19773);
nor U20456 (N_20456,N_19238,N_19625);
nand U20457 (N_20457,N_19080,N_19019);
or U20458 (N_20458,N_18800,N_18764);
or U20459 (N_20459,N_19315,N_19760);
xnor U20460 (N_20460,N_19700,N_19233);
and U20461 (N_20461,N_19290,N_19512);
and U20462 (N_20462,N_18901,N_19439);
or U20463 (N_20463,N_19535,N_19532);
or U20464 (N_20464,N_18834,N_19454);
or U20465 (N_20465,N_19471,N_18862);
nand U20466 (N_20466,N_19912,N_19037);
nand U20467 (N_20467,N_18943,N_19099);
nor U20468 (N_20468,N_18798,N_18843);
xor U20469 (N_20469,N_19497,N_18766);
and U20470 (N_20470,N_19069,N_19977);
nor U20471 (N_20471,N_19883,N_19261);
xor U20472 (N_20472,N_18936,N_18911);
xnor U20473 (N_20473,N_19029,N_19605);
or U20474 (N_20474,N_19894,N_19200);
and U20475 (N_20475,N_19782,N_19203);
and U20476 (N_20476,N_18888,N_19144);
or U20477 (N_20477,N_19831,N_19739);
nand U20478 (N_20478,N_18895,N_19821);
or U20479 (N_20479,N_19396,N_19187);
xor U20480 (N_20480,N_19092,N_19929);
and U20481 (N_20481,N_19511,N_18975);
or U20482 (N_20482,N_18815,N_19374);
nor U20483 (N_20483,N_19949,N_19373);
and U20484 (N_20484,N_19094,N_19012);
and U20485 (N_20485,N_19059,N_19590);
nor U20486 (N_20486,N_19770,N_19748);
nand U20487 (N_20487,N_19110,N_19802);
xnor U20488 (N_20488,N_19888,N_19969);
xnor U20489 (N_20489,N_19684,N_19506);
nor U20490 (N_20490,N_19183,N_19303);
or U20491 (N_20491,N_19341,N_19808);
xnor U20492 (N_20492,N_18946,N_18961);
xor U20493 (N_20493,N_19716,N_19940);
and U20494 (N_20494,N_19451,N_19997);
and U20495 (N_20495,N_19517,N_19380);
or U20496 (N_20496,N_19840,N_19390);
xnor U20497 (N_20497,N_19498,N_19934);
xor U20498 (N_20498,N_19002,N_19568);
nor U20499 (N_20499,N_19027,N_19310);
xnor U20500 (N_20500,N_19795,N_19978);
nor U20501 (N_20501,N_19063,N_19036);
nor U20502 (N_20502,N_19061,N_18865);
xnor U20503 (N_20503,N_18991,N_19809);
xnor U20504 (N_20504,N_19771,N_19549);
nor U20505 (N_20505,N_19211,N_19026);
nor U20506 (N_20506,N_19841,N_18807);
nor U20507 (N_20507,N_19252,N_18751);
nand U20508 (N_20508,N_19264,N_19508);
and U20509 (N_20509,N_19729,N_19188);
or U20510 (N_20510,N_19594,N_19718);
or U20511 (N_20511,N_18886,N_19008);
or U20512 (N_20512,N_19443,N_19533);
xor U20513 (N_20513,N_19441,N_19534);
or U20514 (N_20514,N_19916,N_19612);
or U20515 (N_20515,N_19327,N_19857);
nand U20516 (N_20516,N_19319,N_19702);
nor U20517 (N_20517,N_19085,N_19420);
xnor U20518 (N_20518,N_19033,N_19591);
nor U20519 (N_20519,N_19925,N_19541);
and U20520 (N_20520,N_19152,N_19536);
nor U20521 (N_20521,N_19996,N_19778);
or U20522 (N_20522,N_19562,N_19189);
or U20523 (N_20523,N_18812,N_19343);
nor U20524 (N_20524,N_18825,N_19878);
nand U20525 (N_20525,N_19519,N_19115);
xor U20526 (N_20526,N_19689,N_19458);
or U20527 (N_20527,N_19911,N_19297);
and U20528 (N_20528,N_18880,N_19654);
xnor U20529 (N_20529,N_19258,N_18965);
xnor U20530 (N_20530,N_19011,N_19205);
nand U20531 (N_20531,N_19932,N_18831);
nand U20532 (N_20532,N_19853,N_18977);
and U20533 (N_20533,N_19388,N_19348);
nor U20534 (N_20534,N_19994,N_19556);
and U20535 (N_20535,N_19086,N_18959);
and U20536 (N_20536,N_18956,N_19565);
or U20537 (N_20537,N_19944,N_19216);
xor U20538 (N_20538,N_19885,N_19582);
xnor U20539 (N_20539,N_19251,N_19651);
and U20540 (N_20540,N_19953,N_18823);
nand U20541 (N_20541,N_19948,N_19537);
or U20542 (N_20542,N_19041,N_19023);
nand U20543 (N_20543,N_18755,N_19106);
nand U20544 (N_20544,N_19368,N_19268);
xor U20545 (N_20545,N_18795,N_19836);
nand U20546 (N_20546,N_19155,N_19752);
or U20547 (N_20547,N_19914,N_18918);
xor U20548 (N_20548,N_19671,N_19077);
nand U20549 (N_20549,N_19366,N_18995);
and U20550 (N_20550,N_19370,N_18919);
nand U20551 (N_20551,N_19204,N_18916);
nand U20552 (N_20552,N_19286,N_18981);
and U20553 (N_20553,N_19682,N_19990);
nand U20554 (N_20554,N_19123,N_19472);
xor U20555 (N_20555,N_19253,N_19191);
nand U20556 (N_20556,N_18990,N_19098);
or U20557 (N_20557,N_19142,N_19260);
nor U20558 (N_20558,N_19964,N_19872);
nand U20559 (N_20559,N_19945,N_19902);
nand U20560 (N_20560,N_19277,N_19772);
nor U20561 (N_20561,N_19314,N_19312);
or U20562 (N_20562,N_19030,N_18939);
and U20563 (N_20563,N_19338,N_19208);
or U20564 (N_20564,N_18799,N_18821);
xnor U20565 (N_20565,N_18963,N_19665);
nand U20566 (N_20566,N_18992,N_19616);
nor U20567 (N_20567,N_19113,N_18979);
and U20568 (N_20568,N_18780,N_19414);
nor U20569 (N_20569,N_19892,N_19939);
nand U20570 (N_20570,N_18953,N_19492);
and U20571 (N_20571,N_19174,N_19345);
nor U20572 (N_20572,N_18989,N_19869);
and U20573 (N_20573,N_18997,N_19453);
nor U20574 (N_20574,N_19288,N_19563);
xor U20575 (N_20575,N_19980,N_19475);
xnor U20576 (N_20576,N_19276,N_19054);
nand U20577 (N_20577,N_18967,N_19148);
and U20578 (N_20578,N_18890,N_19112);
nand U20579 (N_20579,N_19039,N_19048);
nor U20580 (N_20580,N_19015,N_18883);
nor U20581 (N_20581,N_19817,N_19122);
or U20582 (N_20582,N_18847,N_19640);
and U20583 (N_20583,N_19270,N_19424);
nor U20584 (N_20584,N_19797,N_19643);
or U20585 (N_20585,N_18905,N_19730);
nor U20586 (N_20586,N_19462,N_19832);
nand U20587 (N_20587,N_19186,N_19001);
xor U20588 (N_20588,N_19357,N_19526);
xnor U20589 (N_20589,N_19091,N_19455);
and U20590 (N_20590,N_19172,N_19221);
and U20591 (N_20591,N_18814,N_19523);
nand U20592 (N_20592,N_19138,N_19409);
or U20593 (N_20593,N_19961,N_19429);
xnor U20594 (N_20594,N_19849,N_19292);
nor U20595 (N_20595,N_19246,N_19595);
nor U20596 (N_20596,N_18882,N_19910);
and U20597 (N_20597,N_19456,N_19364);
xnor U20598 (N_20598,N_18913,N_19151);
nor U20599 (N_20599,N_19941,N_19306);
xor U20600 (N_20600,N_19879,N_18810);
nor U20601 (N_20601,N_19738,N_18922);
nand U20602 (N_20602,N_18838,N_19887);
xnor U20603 (N_20603,N_19891,N_19096);
and U20604 (N_20604,N_19300,N_19146);
nor U20605 (N_20605,N_19835,N_18983);
or U20606 (N_20606,N_19459,N_19042);
nand U20607 (N_20607,N_19761,N_19609);
and U20608 (N_20608,N_19833,N_19228);
xor U20609 (N_20609,N_19201,N_19415);
or U20610 (N_20610,N_19838,N_18757);
nor U20611 (N_20611,N_19358,N_19574);
nand U20612 (N_20612,N_19275,N_19657);
nor U20613 (N_20613,N_18845,N_19423);
nor U20614 (N_20614,N_19922,N_19317);
xor U20615 (N_20615,N_19544,N_19624);
xnor U20616 (N_20616,N_19975,N_19070);
or U20617 (N_20617,N_19807,N_19863);
and U20618 (N_20618,N_19619,N_19354);
nand U20619 (N_20619,N_19627,N_19656);
xnor U20620 (N_20620,N_19118,N_19847);
nor U20621 (N_20621,N_19088,N_19161);
nor U20622 (N_20622,N_19862,N_19550);
and U20623 (N_20623,N_19637,N_19176);
nor U20624 (N_20624,N_18761,N_19732);
and U20625 (N_20625,N_19516,N_19866);
xnor U20626 (N_20626,N_19763,N_19238);
nand U20627 (N_20627,N_18973,N_18762);
nand U20628 (N_20628,N_19189,N_19220);
xor U20629 (N_20629,N_19931,N_19890);
xor U20630 (N_20630,N_19671,N_19905);
nor U20631 (N_20631,N_19613,N_19614);
and U20632 (N_20632,N_19803,N_19890);
or U20633 (N_20633,N_19113,N_19689);
nor U20634 (N_20634,N_19171,N_19803);
xor U20635 (N_20635,N_19037,N_19367);
or U20636 (N_20636,N_19498,N_19428);
or U20637 (N_20637,N_19640,N_19934);
nand U20638 (N_20638,N_19019,N_19820);
or U20639 (N_20639,N_19830,N_19625);
or U20640 (N_20640,N_19771,N_18842);
nor U20641 (N_20641,N_19019,N_19398);
or U20642 (N_20642,N_18993,N_19041);
nand U20643 (N_20643,N_19788,N_19596);
xnor U20644 (N_20644,N_18946,N_19149);
or U20645 (N_20645,N_19805,N_19421);
nor U20646 (N_20646,N_19453,N_19439);
and U20647 (N_20647,N_19545,N_19653);
or U20648 (N_20648,N_19304,N_19923);
or U20649 (N_20649,N_19073,N_19698);
and U20650 (N_20650,N_19995,N_19219);
or U20651 (N_20651,N_19315,N_19361);
or U20652 (N_20652,N_19704,N_18873);
xor U20653 (N_20653,N_19019,N_19758);
and U20654 (N_20654,N_19587,N_18767);
and U20655 (N_20655,N_19981,N_19222);
or U20656 (N_20656,N_19689,N_18793);
nor U20657 (N_20657,N_19404,N_18861);
xnor U20658 (N_20658,N_19136,N_19173);
nor U20659 (N_20659,N_18905,N_18969);
nand U20660 (N_20660,N_19475,N_19100);
nand U20661 (N_20661,N_19331,N_19906);
nor U20662 (N_20662,N_18803,N_18862);
xnor U20663 (N_20663,N_19207,N_19598);
xor U20664 (N_20664,N_19889,N_19859);
nand U20665 (N_20665,N_19430,N_19233);
or U20666 (N_20666,N_19800,N_19066);
or U20667 (N_20667,N_19640,N_18888);
nor U20668 (N_20668,N_19203,N_19126);
nand U20669 (N_20669,N_19292,N_19497);
and U20670 (N_20670,N_19017,N_19708);
or U20671 (N_20671,N_18804,N_19035);
nor U20672 (N_20672,N_19106,N_19630);
and U20673 (N_20673,N_19957,N_19883);
and U20674 (N_20674,N_18972,N_19295);
nor U20675 (N_20675,N_19466,N_19130);
and U20676 (N_20676,N_18940,N_19826);
nand U20677 (N_20677,N_19600,N_19926);
xnor U20678 (N_20678,N_19178,N_19296);
nand U20679 (N_20679,N_19908,N_19299);
xor U20680 (N_20680,N_19211,N_19390);
nand U20681 (N_20681,N_19867,N_19415);
nor U20682 (N_20682,N_19366,N_18763);
xor U20683 (N_20683,N_19204,N_19918);
xnor U20684 (N_20684,N_19155,N_19917);
xnor U20685 (N_20685,N_18941,N_18813);
or U20686 (N_20686,N_18831,N_18883);
and U20687 (N_20687,N_19477,N_19742);
or U20688 (N_20688,N_19084,N_18791);
xnor U20689 (N_20689,N_19921,N_19914);
nand U20690 (N_20690,N_19287,N_19970);
and U20691 (N_20691,N_19893,N_19589);
or U20692 (N_20692,N_19526,N_19397);
and U20693 (N_20693,N_19019,N_19621);
xor U20694 (N_20694,N_19872,N_19174);
nor U20695 (N_20695,N_19442,N_18788);
or U20696 (N_20696,N_19186,N_19465);
nor U20697 (N_20697,N_18938,N_18860);
or U20698 (N_20698,N_18994,N_19363);
xor U20699 (N_20699,N_19355,N_19996);
and U20700 (N_20700,N_19807,N_19221);
and U20701 (N_20701,N_19585,N_19487);
xnor U20702 (N_20702,N_18968,N_19559);
nor U20703 (N_20703,N_19330,N_19584);
nand U20704 (N_20704,N_19007,N_19398);
or U20705 (N_20705,N_18923,N_19295);
nor U20706 (N_20706,N_19889,N_19189);
nand U20707 (N_20707,N_19465,N_19540);
or U20708 (N_20708,N_19924,N_18837);
or U20709 (N_20709,N_19338,N_18968);
or U20710 (N_20710,N_19316,N_19889);
xor U20711 (N_20711,N_19949,N_19142);
or U20712 (N_20712,N_19029,N_19791);
nor U20713 (N_20713,N_19654,N_19410);
nand U20714 (N_20714,N_19405,N_18809);
nor U20715 (N_20715,N_19152,N_19793);
xor U20716 (N_20716,N_19548,N_18835);
nand U20717 (N_20717,N_19572,N_19562);
or U20718 (N_20718,N_19020,N_19419);
and U20719 (N_20719,N_19691,N_19715);
nor U20720 (N_20720,N_19668,N_19646);
xnor U20721 (N_20721,N_18886,N_19406);
or U20722 (N_20722,N_19094,N_19946);
xor U20723 (N_20723,N_19650,N_19713);
nand U20724 (N_20724,N_19311,N_19683);
or U20725 (N_20725,N_19191,N_19430);
and U20726 (N_20726,N_18928,N_19914);
nor U20727 (N_20727,N_18973,N_19565);
xor U20728 (N_20728,N_19078,N_19666);
xor U20729 (N_20729,N_19130,N_19910);
nand U20730 (N_20730,N_19306,N_19256);
nor U20731 (N_20731,N_19561,N_19497);
or U20732 (N_20732,N_19034,N_19873);
xnor U20733 (N_20733,N_19906,N_19437);
nor U20734 (N_20734,N_19236,N_19231);
nand U20735 (N_20735,N_18885,N_19728);
and U20736 (N_20736,N_19417,N_19815);
nor U20737 (N_20737,N_18904,N_19412);
and U20738 (N_20738,N_18992,N_19757);
nand U20739 (N_20739,N_18757,N_19687);
nor U20740 (N_20740,N_19468,N_19511);
nand U20741 (N_20741,N_19263,N_18853);
nand U20742 (N_20742,N_18794,N_18952);
or U20743 (N_20743,N_19942,N_19807);
xor U20744 (N_20744,N_19725,N_18995);
xnor U20745 (N_20745,N_19702,N_19447);
or U20746 (N_20746,N_19526,N_19243);
or U20747 (N_20747,N_18943,N_19841);
or U20748 (N_20748,N_19282,N_18818);
nor U20749 (N_20749,N_19849,N_19242);
nand U20750 (N_20750,N_19922,N_18999);
xnor U20751 (N_20751,N_19355,N_19163);
or U20752 (N_20752,N_19093,N_18753);
nor U20753 (N_20753,N_19912,N_18882);
nand U20754 (N_20754,N_18928,N_18759);
or U20755 (N_20755,N_19003,N_18881);
and U20756 (N_20756,N_18864,N_19966);
and U20757 (N_20757,N_19958,N_18850);
nand U20758 (N_20758,N_19700,N_19838);
nand U20759 (N_20759,N_18878,N_19793);
and U20760 (N_20760,N_19711,N_18819);
nor U20761 (N_20761,N_19662,N_19020);
nand U20762 (N_20762,N_19264,N_19646);
xor U20763 (N_20763,N_19433,N_19880);
xor U20764 (N_20764,N_19072,N_19731);
or U20765 (N_20765,N_19787,N_18800);
or U20766 (N_20766,N_18973,N_19838);
nand U20767 (N_20767,N_19752,N_19083);
nand U20768 (N_20768,N_19431,N_19347);
and U20769 (N_20769,N_19085,N_19861);
and U20770 (N_20770,N_19600,N_19585);
nand U20771 (N_20771,N_19289,N_18902);
or U20772 (N_20772,N_19602,N_19713);
nand U20773 (N_20773,N_19446,N_19204);
nor U20774 (N_20774,N_19166,N_19155);
or U20775 (N_20775,N_19462,N_19631);
xnor U20776 (N_20776,N_19289,N_19415);
nor U20777 (N_20777,N_18995,N_18770);
or U20778 (N_20778,N_19377,N_19250);
nand U20779 (N_20779,N_18827,N_19899);
or U20780 (N_20780,N_19700,N_19106);
nor U20781 (N_20781,N_19589,N_19687);
xnor U20782 (N_20782,N_19899,N_19522);
or U20783 (N_20783,N_19164,N_19423);
and U20784 (N_20784,N_18750,N_19600);
xnor U20785 (N_20785,N_19749,N_19969);
xnor U20786 (N_20786,N_19143,N_19405);
nand U20787 (N_20787,N_18951,N_19158);
and U20788 (N_20788,N_19466,N_19708);
and U20789 (N_20789,N_19246,N_19093);
xor U20790 (N_20790,N_19550,N_19688);
nand U20791 (N_20791,N_18874,N_19074);
xnor U20792 (N_20792,N_19211,N_19903);
nand U20793 (N_20793,N_19099,N_19345);
nor U20794 (N_20794,N_18883,N_19374);
nor U20795 (N_20795,N_19654,N_19972);
and U20796 (N_20796,N_19976,N_19008);
or U20797 (N_20797,N_19598,N_18893);
and U20798 (N_20798,N_19323,N_19860);
nor U20799 (N_20799,N_19933,N_19195);
nor U20800 (N_20800,N_19518,N_18829);
xor U20801 (N_20801,N_19188,N_19681);
nor U20802 (N_20802,N_19066,N_18993);
xnor U20803 (N_20803,N_19868,N_18878);
or U20804 (N_20804,N_19773,N_18960);
xor U20805 (N_20805,N_19468,N_19763);
or U20806 (N_20806,N_19917,N_19806);
nor U20807 (N_20807,N_19907,N_19565);
nor U20808 (N_20808,N_19533,N_19805);
xnor U20809 (N_20809,N_19768,N_19831);
and U20810 (N_20810,N_19892,N_19800);
or U20811 (N_20811,N_19027,N_19080);
xnor U20812 (N_20812,N_19671,N_19977);
or U20813 (N_20813,N_19039,N_19279);
xnor U20814 (N_20814,N_19438,N_18917);
nor U20815 (N_20815,N_18967,N_18916);
or U20816 (N_20816,N_19795,N_19008);
nor U20817 (N_20817,N_19709,N_19631);
nand U20818 (N_20818,N_19386,N_19541);
nor U20819 (N_20819,N_19811,N_18923);
nor U20820 (N_20820,N_19544,N_19573);
nor U20821 (N_20821,N_19521,N_19144);
nor U20822 (N_20822,N_19089,N_19766);
xnor U20823 (N_20823,N_18917,N_19074);
nand U20824 (N_20824,N_19927,N_19011);
xor U20825 (N_20825,N_19585,N_19074);
or U20826 (N_20826,N_19943,N_19250);
nand U20827 (N_20827,N_19207,N_19352);
xnor U20828 (N_20828,N_19786,N_19168);
nand U20829 (N_20829,N_19163,N_19636);
or U20830 (N_20830,N_19138,N_19573);
xnor U20831 (N_20831,N_19944,N_18994);
and U20832 (N_20832,N_18991,N_18982);
and U20833 (N_20833,N_19981,N_19124);
nor U20834 (N_20834,N_19560,N_19343);
nor U20835 (N_20835,N_19801,N_19785);
nand U20836 (N_20836,N_18987,N_19721);
nand U20837 (N_20837,N_18993,N_19825);
xor U20838 (N_20838,N_19572,N_19251);
and U20839 (N_20839,N_19093,N_19452);
and U20840 (N_20840,N_19262,N_18762);
nor U20841 (N_20841,N_19331,N_19445);
xor U20842 (N_20842,N_19292,N_19477);
xor U20843 (N_20843,N_18903,N_19538);
xnor U20844 (N_20844,N_19289,N_18757);
xnor U20845 (N_20845,N_19862,N_19428);
nor U20846 (N_20846,N_18874,N_19012);
nand U20847 (N_20847,N_18971,N_19308);
and U20848 (N_20848,N_19168,N_19303);
or U20849 (N_20849,N_18757,N_19137);
nand U20850 (N_20850,N_19726,N_19834);
nand U20851 (N_20851,N_19476,N_18837);
and U20852 (N_20852,N_18853,N_19558);
nand U20853 (N_20853,N_19545,N_19332);
nand U20854 (N_20854,N_19555,N_19723);
and U20855 (N_20855,N_19170,N_18914);
nor U20856 (N_20856,N_19352,N_19400);
nor U20857 (N_20857,N_18904,N_18878);
and U20858 (N_20858,N_19594,N_19066);
and U20859 (N_20859,N_19688,N_19666);
or U20860 (N_20860,N_19937,N_19465);
or U20861 (N_20861,N_19691,N_19811);
nand U20862 (N_20862,N_18979,N_18804);
nand U20863 (N_20863,N_19791,N_18974);
nand U20864 (N_20864,N_18861,N_19954);
xor U20865 (N_20865,N_19338,N_19921);
and U20866 (N_20866,N_19446,N_19906);
or U20867 (N_20867,N_18756,N_19689);
xor U20868 (N_20868,N_19097,N_19411);
and U20869 (N_20869,N_19427,N_19584);
nor U20870 (N_20870,N_19570,N_19397);
nor U20871 (N_20871,N_18874,N_19476);
and U20872 (N_20872,N_19412,N_19899);
nor U20873 (N_20873,N_19717,N_19403);
nand U20874 (N_20874,N_19793,N_18957);
nor U20875 (N_20875,N_19045,N_18843);
xor U20876 (N_20876,N_19534,N_19352);
nor U20877 (N_20877,N_18959,N_19649);
nor U20878 (N_20878,N_18941,N_19171);
or U20879 (N_20879,N_19740,N_19714);
nand U20880 (N_20880,N_19555,N_19768);
or U20881 (N_20881,N_19777,N_18962);
xnor U20882 (N_20882,N_19081,N_19415);
and U20883 (N_20883,N_18981,N_19182);
and U20884 (N_20884,N_18751,N_19600);
xor U20885 (N_20885,N_18875,N_19360);
nand U20886 (N_20886,N_19175,N_19945);
nand U20887 (N_20887,N_18949,N_19311);
nand U20888 (N_20888,N_19670,N_19498);
nand U20889 (N_20889,N_19995,N_19983);
xnor U20890 (N_20890,N_18793,N_19964);
or U20891 (N_20891,N_19862,N_19783);
xor U20892 (N_20892,N_18965,N_19617);
nand U20893 (N_20893,N_19773,N_19177);
nor U20894 (N_20894,N_19147,N_19871);
nor U20895 (N_20895,N_19814,N_19573);
nor U20896 (N_20896,N_18855,N_19367);
or U20897 (N_20897,N_18797,N_18858);
xnor U20898 (N_20898,N_19222,N_19218);
xnor U20899 (N_20899,N_19853,N_18870);
and U20900 (N_20900,N_19888,N_19802);
xor U20901 (N_20901,N_19756,N_19587);
nand U20902 (N_20902,N_19420,N_19287);
or U20903 (N_20903,N_19485,N_19954);
nor U20904 (N_20904,N_18961,N_19938);
nand U20905 (N_20905,N_18917,N_19550);
and U20906 (N_20906,N_19887,N_19709);
nand U20907 (N_20907,N_18811,N_19727);
xnor U20908 (N_20908,N_19008,N_19791);
and U20909 (N_20909,N_19231,N_18812);
and U20910 (N_20910,N_19356,N_19396);
and U20911 (N_20911,N_19179,N_18821);
and U20912 (N_20912,N_19502,N_18867);
xor U20913 (N_20913,N_18943,N_19748);
and U20914 (N_20914,N_19215,N_19057);
nand U20915 (N_20915,N_19964,N_19490);
xor U20916 (N_20916,N_18961,N_18952);
nor U20917 (N_20917,N_19256,N_19257);
or U20918 (N_20918,N_19911,N_19363);
or U20919 (N_20919,N_18952,N_19278);
or U20920 (N_20920,N_19998,N_19991);
xnor U20921 (N_20921,N_18817,N_19777);
xor U20922 (N_20922,N_19112,N_19313);
nand U20923 (N_20923,N_19333,N_19284);
or U20924 (N_20924,N_18869,N_19003);
nand U20925 (N_20925,N_19582,N_19595);
nand U20926 (N_20926,N_19464,N_19405);
xnor U20927 (N_20927,N_18971,N_18953);
xnor U20928 (N_20928,N_19631,N_19561);
nand U20929 (N_20929,N_19575,N_19898);
xor U20930 (N_20930,N_19200,N_19962);
xor U20931 (N_20931,N_19337,N_18935);
nor U20932 (N_20932,N_19987,N_18774);
or U20933 (N_20933,N_19951,N_19741);
or U20934 (N_20934,N_19599,N_19131);
nor U20935 (N_20935,N_19413,N_18894);
nand U20936 (N_20936,N_18978,N_19312);
nor U20937 (N_20937,N_19964,N_18923);
nand U20938 (N_20938,N_19455,N_19369);
or U20939 (N_20939,N_19972,N_18852);
xnor U20940 (N_20940,N_18940,N_19651);
nor U20941 (N_20941,N_19784,N_19428);
nand U20942 (N_20942,N_19187,N_19888);
or U20943 (N_20943,N_19962,N_19491);
or U20944 (N_20944,N_19962,N_19197);
and U20945 (N_20945,N_19252,N_19330);
nor U20946 (N_20946,N_19183,N_19710);
nand U20947 (N_20947,N_19757,N_18977);
xnor U20948 (N_20948,N_19921,N_19746);
nor U20949 (N_20949,N_19067,N_19224);
or U20950 (N_20950,N_18941,N_19674);
xnor U20951 (N_20951,N_19260,N_19099);
or U20952 (N_20952,N_19568,N_19402);
nor U20953 (N_20953,N_19906,N_19243);
xor U20954 (N_20954,N_19815,N_19613);
and U20955 (N_20955,N_19780,N_19642);
nand U20956 (N_20956,N_18832,N_19680);
and U20957 (N_20957,N_19230,N_19057);
nand U20958 (N_20958,N_19458,N_18950);
xor U20959 (N_20959,N_19799,N_19549);
and U20960 (N_20960,N_19195,N_19896);
and U20961 (N_20961,N_18858,N_19341);
or U20962 (N_20962,N_19752,N_19461);
nor U20963 (N_20963,N_19775,N_19560);
nor U20964 (N_20964,N_19781,N_19613);
and U20965 (N_20965,N_19056,N_18987);
and U20966 (N_20966,N_19774,N_18826);
xor U20967 (N_20967,N_18809,N_19674);
nor U20968 (N_20968,N_19637,N_19362);
or U20969 (N_20969,N_18790,N_19380);
or U20970 (N_20970,N_19591,N_19359);
and U20971 (N_20971,N_19377,N_19767);
or U20972 (N_20972,N_19062,N_19850);
nor U20973 (N_20973,N_18997,N_19738);
xnor U20974 (N_20974,N_19905,N_19482);
or U20975 (N_20975,N_19402,N_19508);
or U20976 (N_20976,N_19554,N_19383);
nor U20977 (N_20977,N_19585,N_19659);
nand U20978 (N_20978,N_19847,N_19294);
and U20979 (N_20979,N_19215,N_19807);
nor U20980 (N_20980,N_19639,N_19946);
or U20981 (N_20981,N_19352,N_18893);
xor U20982 (N_20982,N_19324,N_19082);
xor U20983 (N_20983,N_19445,N_19169);
and U20984 (N_20984,N_18879,N_19296);
and U20985 (N_20985,N_19696,N_19177);
nand U20986 (N_20986,N_18973,N_19583);
and U20987 (N_20987,N_19544,N_19476);
or U20988 (N_20988,N_19179,N_18801);
or U20989 (N_20989,N_19121,N_19384);
nand U20990 (N_20990,N_18862,N_19370);
and U20991 (N_20991,N_19952,N_18844);
and U20992 (N_20992,N_18865,N_18818);
or U20993 (N_20993,N_19530,N_19912);
or U20994 (N_20994,N_19894,N_19405);
nand U20995 (N_20995,N_19049,N_19925);
or U20996 (N_20996,N_19288,N_19459);
nand U20997 (N_20997,N_19257,N_19055);
nor U20998 (N_20998,N_18960,N_19003);
nor U20999 (N_20999,N_19535,N_19301);
nor U21000 (N_21000,N_18778,N_19739);
and U21001 (N_21001,N_19378,N_19004);
nand U21002 (N_21002,N_18827,N_18816);
nand U21003 (N_21003,N_19571,N_19250);
or U21004 (N_21004,N_19334,N_18770);
xnor U21005 (N_21005,N_19995,N_19351);
xnor U21006 (N_21006,N_19797,N_19546);
and U21007 (N_21007,N_19642,N_18945);
or U21008 (N_21008,N_18905,N_19709);
or U21009 (N_21009,N_18928,N_18816);
nor U21010 (N_21010,N_19000,N_18753);
nor U21011 (N_21011,N_19031,N_19462);
or U21012 (N_21012,N_19325,N_19529);
or U21013 (N_21013,N_19587,N_19391);
xor U21014 (N_21014,N_18756,N_19549);
xor U21015 (N_21015,N_19543,N_19400);
or U21016 (N_21016,N_19378,N_18928);
nand U21017 (N_21017,N_19318,N_18757);
and U21018 (N_21018,N_18793,N_19110);
nor U21019 (N_21019,N_18947,N_18925);
nor U21020 (N_21020,N_19792,N_19843);
nor U21021 (N_21021,N_19682,N_19750);
and U21022 (N_21022,N_18850,N_18811);
and U21023 (N_21023,N_18936,N_18861);
nand U21024 (N_21024,N_19394,N_18925);
xnor U21025 (N_21025,N_19327,N_19383);
nor U21026 (N_21026,N_19616,N_19479);
xor U21027 (N_21027,N_19222,N_18972);
xnor U21028 (N_21028,N_19923,N_19754);
xnor U21029 (N_21029,N_18830,N_19332);
nand U21030 (N_21030,N_19831,N_19648);
nand U21031 (N_21031,N_19841,N_19133);
xnor U21032 (N_21032,N_18950,N_19552);
nand U21033 (N_21033,N_19426,N_19384);
nor U21034 (N_21034,N_19547,N_19129);
and U21035 (N_21035,N_19220,N_18961);
or U21036 (N_21036,N_18822,N_19287);
nor U21037 (N_21037,N_19684,N_19144);
or U21038 (N_21038,N_19905,N_19199);
and U21039 (N_21039,N_18970,N_18798);
and U21040 (N_21040,N_19221,N_18766);
nand U21041 (N_21041,N_19817,N_19593);
nand U21042 (N_21042,N_19991,N_18980);
or U21043 (N_21043,N_19538,N_19074);
nand U21044 (N_21044,N_19045,N_19839);
nor U21045 (N_21045,N_19063,N_19745);
xnor U21046 (N_21046,N_19628,N_19324);
or U21047 (N_21047,N_19811,N_18762);
nand U21048 (N_21048,N_19231,N_19239);
nor U21049 (N_21049,N_18946,N_19742);
nand U21050 (N_21050,N_19339,N_19198);
or U21051 (N_21051,N_19521,N_19615);
and U21052 (N_21052,N_19438,N_18854);
or U21053 (N_21053,N_19255,N_19910);
xnor U21054 (N_21054,N_19249,N_19299);
and U21055 (N_21055,N_19142,N_19401);
and U21056 (N_21056,N_19386,N_18872);
nor U21057 (N_21057,N_19439,N_18962);
xor U21058 (N_21058,N_19423,N_19827);
nor U21059 (N_21059,N_19858,N_19097);
nor U21060 (N_21060,N_18959,N_19857);
or U21061 (N_21061,N_19782,N_19474);
xor U21062 (N_21062,N_19147,N_19336);
nand U21063 (N_21063,N_19302,N_19443);
nor U21064 (N_21064,N_19689,N_19006);
and U21065 (N_21065,N_19238,N_19747);
and U21066 (N_21066,N_18797,N_18854);
and U21067 (N_21067,N_19058,N_19332);
or U21068 (N_21068,N_18868,N_19123);
nand U21069 (N_21069,N_18761,N_18952);
nor U21070 (N_21070,N_19728,N_19099);
nand U21071 (N_21071,N_19843,N_19334);
xnor U21072 (N_21072,N_19625,N_19373);
nand U21073 (N_21073,N_19548,N_19497);
xor U21074 (N_21074,N_19360,N_18856);
xnor U21075 (N_21075,N_19726,N_19818);
nor U21076 (N_21076,N_19673,N_18884);
or U21077 (N_21077,N_19728,N_19742);
or U21078 (N_21078,N_19989,N_19147);
and U21079 (N_21079,N_19259,N_19684);
xnor U21080 (N_21080,N_19731,N_19041);
and U21081 (N_21081,N_18981,N_19453);
nor U21082 (N_21082,N_19296,N_19826);
and U21083 (N_21083,N_19728,N_19315);
nor U21084 (N_21084,N_19884,N_19799);
nand U21085 (N_21085,N_19636,N_19373);
xnor U21086 (N_21086,N_18998,N_19176);
or U21087 (N_21087,N_19654,N_19142);
nand U21088 (N_21088,N_18850,N_19779);
or U21089 (N_21089,N_19549,N_19864);
nand U21090 (N_21090,N_19143,N_19818);
nand U21091 (N_21091,N_19193,N_18762);
xnor U21092 (N_21092,N_19109,N_18996);
or U21093 (N_21093,N_19186,N_19148);
nor U21094 (N_21094,N_19912,N_19348);
nand U21095 (N_21095,N_19128,N_19485);
xor U21096 (N_21096,N_19312,N_19358);
and U21097 (N_21097,N_19922,N_18942);
nor U21098 (N_21098,N_19948,N_18857);
and U21099 (N_21099,N_18974,N_18792);
nand U21100 (N_21100,N_19985,N_19287);
nor U21101 (N_21101,N_18820,N_19493);
xor U21102 (N_21102,N_19501,N_18868);
or U21103 (N_21103,N_19135,N_19650);
or U21104 (N_21104,N_19718,N_19358);
nor U21105 (N_21105,N_19642,N_19395);
and U21106 (N_21106,N_19841,N_19750);
and U21107 (N_21107,N_19836,N_19841);
nand U21108 (N_21108,N_19182,N_19820);
nor U21109 (N_21109,N_19971,N_19134);
or U21110 (N_21110,N_19521,N_19229);
nand U21111 (N_21111,N_19297,N_19062);
or U21112 (N_21112,N_19411,N_19702);
and U21113 (N_21113,N_19386,N_19776);
xnor U21114 (N_21114,N_19923,N_19826);
nor U21115 (N_21115,N_18852,N_18993);
xnor U21116 (N_21116,N_18948,N_19175);
and U21117 (N_21117,N_19120,N_18847);
xor U21118 (N_21118,N_19320,N_18942);
xnor U21119 (N_21119,N_19408,N_19259);
and U21120 (N_21120,N_19587,N_19696);
or U21121 (N_21121,N_18954,N_19334);
nand U21122 (N_21122,N_18935,N_19757);
nand U21123 (N_21123,N_19991,N_19840);
xnor U21124 (N_21124,N_19258,N_19918);
and U21125 (N_21125,N_18751,N_19858);
and U21126 (N_21126,N_18902,N_19347);
xor U21127 (N_21127,N_19228,N_19129);
and U21128 (N_21128,N_19417,N_19356);
nand U21129 (N_21129,N_19872,N_19094);
or U21130 (N_21130,N_19309,N_19303);
xor U21131 (N_21131,N_19545,N_19303);
and U21132 (N_21132,N_18950,N_19100);
and U21133 (N_21133,N_19381,N_18874);
and U21134 (N_21134,N_19126,N_19544);
xor U21135 (N_21135,N_19513,N_19730);
and U21136 (N_21136,N_19598,N_19775);
nor U21137 (N_21137,N_19425,N_18946);
and U21138 (N_21138,N_18947,N_19599);
nand U21139 (N_21139,N_19054,N_19551);
nor U21140 (N_21140,N_19269,N_19560);
and U21141 (N_21141,N_19245,N_19677);
or U21142 (N_21142,N_19178,N_18944);
nor U21143 (N_21143,N_19209,N_19090);
nand U21144 (N_21144,N_19097,N_19840);
and U21145 (N_21145,N_19176,N_19872);
and U21146 (N_21146,N_18824,N_19561);
nor U21147 (N_21147,N_18976,N_19460);
or U21148 (N_21148,N_19003,N_19462);
nand U21149 (N_21149,N_19602,N_19224);
nor U21150 (N_21150,N_19581,N_19627);
nand U21151 (N_21151,N_19891,N_19933);
or U21152 (N_21152,N_19683,N_19261);
nor U21153 (N_21153,N_19962,N_18807);
xor U21154 (N_21154,N_19003,N_19075);
nor U21155 (N_21155,N_18842,N_19619);
nand U21156 (N_21156,N_19772,N_19846);
nor U21157 (N_21157,N_18852,N_19310);
and U21158 (N_21158,N_19759,N_19811);
xnor U21159 (N_21159,N_19579,N_19989);
and U21160 (N_21160,N_19834,N_19717);
and U21161 (N_21161,N_19572,N_19220);
nand U21162 (N_21162,N_19133,N_19132);
and U21163 (N_21163,N_19023,N_19063);
or U21164 (N_21164,N_19604,N_19772);
nor U21165 (N_21165,N_18889,N_18911);
nand U21166 (N_21166,N_18760,N_19583);
xor U21167 (N_21167,N_19595,N_18836);
or U21168 (N_21168,N_18938,N_19947);
and U21169 (N_21169,N_19057,N_19867);
xnor U21170 (N_21170,N_19523,N_19895);
and U21171 (N_21171,N_19545,N_18779);
nor U21172 (N_21172,N_19692,N_19866);
xor U21173 (N_21173,N_18852,N_19360);
or U21174 (N_21174,N_19212,N_19450);
nand U21175 (N_21175,N_19478,N_19953);
or U21176 (N_21176,N_19430,N_19170);
or U21177 (N_21177,N_19776,N_18929);
or U21178 (N_21178,N_19073,N_18998);
and U21179 (N_21179,N_19497,N_19204);
nand U21180 (N_21180,N_19710,N_19534);
and U21181 (N_21181,N_19474,N_19002);
nand U21182 (N_21182,N_19511,N_18906);
xnor U21183 (N_21183,N_19433,N_19787);
and U21184 (N_21184,N_19726,N_19792);
nor U21185 (N_21185,N_19843,N_19931);
and U21186 (N_21186,N_19924,N_19216);
and U21187 (N_21187,N_19687,N_19193);
xor U21188 (N_21188,N_19879,N_19173);
xor U21189 (N_21189,N_19039,N_19901);
nand U21190 (N_21190,N_19811,N_19426);
nor U21191 (N_21191,N_19408,N_19625);
or U21192 (N_21192,N_19288,N_18969);
and U21193 (N_21193,N_18927,N_19395);
or U21194 (N_21194,N_19371,N_19064);
and U21195 (N_21195,N_19651,N_19129);
nor U21196 (N_21196,N_19926,N_19886);
and U21197 (N_21197,N_19227,N_19698);
or U21198 (N_21198,N_19832,N_19809);
or U21199 (N_21199,N_19592,N_19640);
nand U21200 (N_21200,N_19588,N_19860);
or U21201 (N_21201,N_19060,N_19528);
xnor U21202 (N_21202,N_19765,N_19481);
nand U21203 (N_21203,N_18913,N_18940);
nor U21204 (N_21204,N_19028,N_19555);
or U21205 (N_21205,N_19471,N_18833);
and U21206 (N_21206,N_19066,N_19298);
nor U21207 (N_21207,N_19080,N_18784);
and U21208 (N_21208,N_19640,N_19702);
nor U21209 (N_21209,N_19181,N_19703);
xnor U21210 (N_21210,N_19618,N_19929);
nor U21211 (N_21211,N_19468,N_19479);
or U21212 (N_21212,N_19273,N_19030);
nor U21213 (N_21213,N_19786,N_19716);
and U21214 (N_21214,N_19679,N_18780);
or U21215 (N_21215,N_19346,N_19047);
xor U21216 (N_21216,N_19392,N_19189);
or U21217 (N_21217,N_19817,N_19941);
xor U21218 (N_21218,N_18760,N_19149);
xnor U21219 (N_21219,N_19403,N_19352);
or U21220 (N_21220,N_19270,N_19253);
and U21221 (N_21221,N_19481,N_19372);
or U21222 (N_21222,N_19406,N_19299);
nor U21223 (N_21223,N_19916,N_18813);
nor U21224 (N_21224,N_19114,N_18899);
nand U21225 (N_21225,N_19165,N_19603);
nand U21226 (N_21226,N_18908,N_18905);
nor U21227 (N_21227,N_19182,N_19050);
or U21228 (N_21228,N_19086,N_19444);
or U21229 (N_21229,N_19387,N_19475);
and U21230 (N_21230,N_19412,N_19189);
nand U21231 (N_21231,N_19312,N_19986);
nor U21232 (N_21232,N_18768,N_19642);
nand U21233 (N_21233,N_19103,N_19372);
or U21234 (N_21234,N_19834,N_19145);
xor U21235 (N_21235,N_18825,N_19815);
xnor U21236 (N_21236,N_19742,N_19795);
xor U21237 (N_21237,N_19650,N_19229);
or U21238 (N_21238,N_19043,N_19643);
and U21239 (N_21239,N_19579,N_19643);
or U21240 (N_21240,N_19484,N_19420);
and U21241 (N_21241,N_19712,N_19577);
nor U21242 (N_21242,N_19774,N_19898);
nand U21243 (N_21243,N_18920,N_19572);
xnor U21244 (N_21244,N_18943,N_18873);
and U21245 (N_21245,N_19802,N_19975);
nand U21246 (N_21246,N_18822,N_19217);
xor U21247 (N_21247,N_18944,N_19987);
nor U21248 (N_21248,N_19008,N_19029);
nand U21249 (N_21249,N_19690,N_19275);
nor U21250 (N_21250,N_20750,N_21096);
nor U21251 (N_21251,N_21120,N_20524);
or U21252 (N_21252,N_20166,N_21197);
nor U21253 (N_21253,N_20325,N_20417);
and U21254 (N_21254,N_21190,N_20774);
or U21255 (N_21255,N_20897,N_20021);
or U21256 (N_21256,N_20405,N_20557);
nand U21257 (N_21257,N_20331,N_20708);
and U21258 (N_21258,N_20099,N_20330);
nand U21259 (N_21259,N_20853,N_20544);
and U21260 (N_21260,N_21101,N_20333);
nand U21261 (N_21261,N_20630,N_20051);
nand U21262 (N_21262,N_20769,N_21174);
or U21263 (N_21263,N_20874,N_20757);
nor U21264 (N_21264,N_20679,N_20819);
and U21265 (N_21265,N_20680,N_20436);
nand U21266 (N_21266,N_20886,N_20985);
nand U21267 (N_21267,N_20908,N_20097);
nor U21268 (N_21268,N_20010,N_21032);
or U21269 (N_21269,N_20885,N_21110);
xor U21270 (N_21270,N_20268,N_20532);
or U21271 (N_21271,N_20872,N_20720);
and U21272 (N_21272,N_20512,N_20128);
nand U21273 (N_21273,N_20256,N_20996);
or U21274 (N_21274,N_20569,N_20786);
or U21275 (N_21275,N_20346,N_20339);
and U21276 (N_21276,N_20876,N_21220);
or U21277 (N_21277,N_21082,N_20471);
nor U21278 (N_21278,N_21076,N_20131);
nor U21279 (N_21279,N_20059,N_20558);
and U21280 (N_21280,N_20401,N_20929);
xor U21281 (N_21281,N_20984,N_20926);
or U21282 (N_21282,N_20954,N_20168);
xor U21283 (N_21283,N_21107,N_20006);
nand U21284 (N_21284,N_20434,N_20304);
xor U21285 (N_21285,N_20510,N_21182);
nor U21286 (N_21286,N_20081,N_20972);
nor U21287 (N_21287,N_20693,N_20347);
xor U21288 (N_21288,N_21170,N_20249);
nand U21289 (N_21289,N_20461,N_20554);
and U21290 (N_21290,N_20931,N_20751);
or U21291 (N_21291,N_20823,N_20525);
nor U21292 (N_21292,N_20445,N_21249);
or U21293 (N_21293,N_21022,N_20018);
or U21294 (N_21294,N_20592,N_20068);
and U21295 (N_21295,N_20211,N_20754);
nor U21296 (N_21296,N_21121,N_20190);
or U21297 (N_21297,N_20617,N_20384);
or U21298 (N_21298,N_21228,N_21067);
or U21299 (N_21299,N_21136,N_20807);
and U21300 (N_21300,N_20290,N_21088);
nand U21301 (N_21301,N_20517,N_20318);
nand U21302 (N_21302,N_20585,N_21070);
and U21303 (N_21303,N_21078,N_20838);
nor U21304 (N_21304,N_20988,N_20820);
nand U21305 (N_21305,N_20174,N_20079);
xor U21306 (N_21306,N_20618,N_20580);
and U21307 (N_21307,N_21181,N_20443);
nand U21308 (N_21308,N_20684,N_20343);
nand U21309 (N_21309,N_20121,N_21048);
nand U21310 (N_21310,N_21122,N_20199);
or U21311 (N_21311,N_20085,N_20639);
xor U21312 (N_21312,N_21105,N_20624);
xor U21313 (N_21313,N_20119,N_20701);
nand U21314 (N_21314,N_20578,N_20887);
xor U21315 (N_21315,N_21218,N_20016);
xnor U21316 (N_21316,N_20670,N_20899);
and U21317 (N_21317,N_20894,N_20740);
nand U21318 (N_21318,N_20251,N_20799);
and U21319 (N_21319,N_21116,N_20412);
and U21320 (N_21320,N_20400,N_20364);
nor U21321 (N_21321,N_20845,N_20194);
nor U21322 (N_21322,N_21104,N_20378);
nand U21323 (N_21323,N_21168,N_21213);
or U21324 (N_21324,N_20065,N_20977);
or U21325 (N_21325,N_20386,N_20044);
xnor U21326 (N_21326,N_21146,N_20735);
and U21327 (N_21327,N_20681,N_20348);
or U21328 (N_21328,N_20116,N_20429);
nand U21329 (N_21329,N_20257,N_20516);
or U21330 (N_21330,N_20748,N_20046);
or U21331 (N_21331,N_20489,N_21045);
nand U21332 (N_21332,N_20672,N_20396);
or U21333 (N_21333,N_20221,N_21207);
or U21334 (N_21334,N_20153,N_20547);
nand U21335 (N_21335,N_20289,N_20255);
xor U21336 (N_21336,N_20594,N_20125);
xor U21337 (N_21337,N_21030,N_20178);
nand U21338 (N_21338,N_20865,N_21231);
xnor U21339 (N_21339,N_20064,N_20635);
xnor U21340 (N_21340,N_20810,N_20784);
nand U21341 (N_21341,N_21149,N_20572);
nor U21342 (N_21342,N_20224,N_20969);
or U21343 (N_21343,N_20548,N_20531);
xnor U21344 (N_21344,N_20669,N_20599);
nand U21345 (N_21345,N_21156,N_20342);
or U21346 (N_21346,N_20056,N_20135);
xnor U21347 (N_21347,N_20582,N_20365);
or U21348 (N_21348,N_20832,N_20733);
and U21349 (N_21349,N_20377,N_20239);
or U21350 (N_21350,N_20738,N_21098);
nor U21351 (N_21351,N_21199,N_20511);
nor U21352 (N_21352,N_20614,N_20413);
nand U21353 (N_21353,N_21138,N_20546);
nand U21354 (N_21354,N_20833,N_20375);
nor U21355 (N_21355,N_21242,N_21196);
xor U21356 (N_21356,N_21083,N_20830);
nor U21357 (N_21357,N_20976,N_20514);
nand U21358 (N_21358,N_21113,N_20918);
and U21359 (N_21359,N_21123,N_20453);
and U21360 (N_21360,N_20593,N_21009);
or U21361 (N_21361,N_20382,N_20250);
and U21362 (N_21362,N_20392,N_20702);
and U21363 (N_21363,N_20629,N_20942);
or U21364 (N_21364,N_20816,N_20687);
nand U21365 (N_21365,N_21095,N_20328);
nor U21366 (N_21366,N_20998,N_20509);
and U21367 (N_21367,N_21198,N_20794);
and U21368 (N_21368,N_20004,N_20243);
nand U21369 (N_21369,N_21155,N_20835);
xnor U21370 (N_21370,N_20039,N_20898);
nand U21371 (N_21371,N_21239,N_20266);
and U21372 (N_21372,N_21084,N_21127);
or U21373 (N_21373,N_20092,N_20631);
and U21374 (N_21374,N_20465,N_20041);
and U21375 (N_21375,N_20123,N_20458);
and U21376 (N_21376,N_20207,N_20246);
or U21377 (N_21377,N_20462,N_20418);
or U21378 (N_21378,N_20965,N_20208);
and U21379 (N_21379,N_20351,N_20916);
or U21380 (N_21380,N_20966,N_20107);
or U21381 (N_21381,N_20612,N_20935);
and U21382 (N_21382,N_20692,N_20873);
and U21383 (N_21383,N_20235,N_20181);
nor U21384 (N_21384,N_21154,N_20924);
nor U21385 (N_21385,N_20999,N_20852);
and U21386 (N_21386,N_20504,N_20283);
nand U21387 (N_21387,N_20499,N_20619);
nand U21388 (N_21388,N_20219,N_20581);
nor U21389 (N_21389,N_20536,N_20076);
nor U21390 (N_21390,N_21038,N_20034);
xnor U21391 (N_21391,N_20451,N_20171);
nand U21392 (N_21392,N_20216,N_20476);
and U21393 (N_21393,N_21052,N_21069);
or U21394 (N_21394,N_20971,N_20848);
and U21395 (N_21395,N_20997,N_20490);
xor U21396 (N_21396,N_20668,N_21019);
or U21397 (N_21397,N_21180,N_20561);
nor U21398 (N_21398,N_20921,N_20053);
or U21399 (N_21399,N_20888,N_20473);
and U21400 (N_21400,N_20529,N_20310);
and U21401 (N_21401,N_20858,N_21039);
nand U21402 (N_21402,N_20498,N_20469);
xor U21403 (N_21403,N_20080,N_20608);
nand U21404 (N_21404,N_21109,N_20336);
nand U21405 (N_21405,N_20817,N_20744);
or U21406 (N_21406,N_20362,N_20430);
or U21407 (N_21407,N_20084,N_20045);
nand U21408 (N_21408,N_20588,N_20930);
xor U21409 (N_21409,N_21016,N_20063);
or U21410 (N_21410,N_20553,N_20800);
nand U21411 (N_21411,N_20066,N_20648);
or U21412 (N_21412,N_21074,N_20944);
and U21413 (N_21413,N_20882,N_20674);
nor U21414 (N_21414,N_20220,N_21046);
and U21415 (N_21415,N_21137,N_20460);
nand U21416 (N_21416,N_20366,N_20089);
and U21417 (N_21417,N_20940,N_20369);
nand U21418 (N_21418,N_21108,N_20513);
or U21419 (N_21419,N_21063,N_20978);
xnor U21420 (N_21420,N_20309,N_20111);
nand U21421 (N_21421,N_20160,N_20764);
xor U21422 (N_21422,N_21055,N_20454);
and U21423 (N_21423,N_21087,N_20301);
nor U21424 (N_21424,N_20154,N_20167);
or U21425 (N_21425,N_20227,N_20422);
nand U21426 (N_21426,N_20533,N_21172);
xor U21427 (N_21427,N_20566,N_20054);
and U21428 (N_21428,N_21077,N_21236);
nand U21429 (N_21429,N_20000,N_20613);
xnor U21430 (N_21430,N_20108,N_20156);
nand U21431 (N_21431,N_20537,N_20144);
or U21432 (N_21432,N_20716,N_20103);
xor U21433 (N_21433,N_20398,N_20974);
nand U21434 (N_21434,N_20542,N_20960);
xor U21435 (N_21435,N_20298,N_20270);
and U21436 (N_21436,N_20427,N_20201);
nand U21437 (N_21437,N_20431,N_20739);
or U21438 (N_21438,N_20410,N_21194);
nor U21439 (N_21439,N_20941,N_21235);
or U21440 (N_21440,N_21216,N_20657);
or U21441 (N_21441,N_20214,N_20688);
xor U21442 (N_21442,N_21102,N_21097);
nor U21443 (N_21443,N_20947,N_20003);
xor U21444 (N_21444,N_20552,N_21128);
and U21445 (N_21445,N_21100,N_21056);
or U21446 (N_21446,N_20851,N_20315);
nor U21447 (N_21447,N_20404,N_20633);
and U21448 (N_21448,N_20933,N_20082);
or U21449 (N_21449,N_21031,N_20397);
nor U21450 (N_21450,N_21191,N_20983);
nand U21451 (N_21451,N_20015,N_20903);
nor U21452 (N_21452,N_21215,N_20560);
nor U21453 (N_21453,N_20245,N_20914);
xor U21454 (N_21454,N_20615,N_21064);
nor U21455 (N_21455,N_20466,N_20905);
nor U21456 (N_21456,N_20213,N_21159);
or U21457 (N_21457,N_20381,N_20920);
nor U21458 (N_21458,N_20083,N_20264);
or U21459 (N_21459,N_20749,N_20008);
and U21460 (N_21460,N_20332,N_20137);
or U21461 (N_21461,N_20225,N_20959);
and U21462 (N_21462,N_20549,N_20487);
nand U21463 (N_21463,N_20936,N_20494);
xnor U21464 (N_21464,N_20587,N_20215);
or U21465 (N_21465,N_20822,N_20488);
nand U21466 (N_21466,N_20340,N_20326);
xor U21467 (N_21467,N_20598,N_20275);
nand U21468 (N_21468,N_20306,N_20191);
and U21469 (N_21469,N_20550,N_21153);
and U21470 (N_21470,N_20162,N_20062);
nor U21471 (N_21471,N_20906,N_20175);
xnor U21472 (N_21472,N_20987,N_20122);
xnor U21473 (N_21473,N_20372,N_21033);
xnor U21474 (N_21474,N_20379,N_20180);
nor U21475 (N_21475,N_20530,N_21021);
nand U21476 (N_21476,N_20651,N_20282);
xor U21477 (N_21477,N_21224,N_20100);
xor U21478 (N_21478,N_20927,N_20196);
or U21479 (N_21479,N_21246,N_20932);
xor U21480 (N_21480,N_20798,N_20258);
or U21481 (N_21481,N_20990,N_20409);
or U21482 (N_21482,N_20170,N_20995);
and U21483 (N_21483,N_20907,N_20895);
nor U21484 (N_21484,N_20611,N_20197);
xor U21485 (N_21485,N_20755,N_20269);
nand U21486 (N_21486,N_20742,N_20640);
nand U21487 (N_21487,N_20296,N_20142);
nand U21488 (N_21488,N_20857,N_21247);
nand U21489 (N_21489,N_20705,N_20272);
nand U21490 (N_21490,N_20446,N_20442);
and U21491 (N_21491,N_20109,N_20747);
nor U21492 (N_21492,N_20795,N_20535);
and U21493 (N_21493,N_20622,N_20112);
or U21494 (N_21494,N_20586,N_20715);
nand U21495 (N_21495,N_20893,N_20470);
nand U21496 (N_21496,N_20479,N_20871);
nand U21497 (N_21497,N_20049,N_20846);
and U21498 (N_21498,N_20945,N_20165);
nand U21499 (N_21499,N_20884,N_20609);
and U21500 (N_21500,N_21029,N_20038);
xor U21501 (N_21501,N_21002,N_20023);
nand U21502 (N_21502,N_20478,N_20299);
or U21503 (N_21503,N_20957,N_20424);
or U21504 (N_21504,N_20937,N_21189);
xnor U21505 (N_21505,N_20659,N_20238);
or U21506 (N_21506,N_21027,N_20236);
xor U21507 (N_21507,N_20013,N_20787);
and U21508 (N_21508,N_20939,N_20195);
xor U21509 (N_21509,N_20475,N_20145);
nor U21510 (N_21510,N_20603,N_20782);
nand U21511 (N_21511,N_20818,N_20877);
and U21512 (N_21512,N_20570,N_21144);
nand U21513 (N_21513,N_21011,N_21079);
nand U21514 (N_21514,N_20009,N_20237);
or U21515 (N_21515,N_20205,N_20295);
nor U21516 (N_21516,N_21050,N_20867);
nor U21517 (N_21517,N_20909,N_20344);
and U21518 (N_21518,N_20765,N_20277);
xnor U21519 (N_21519,N_20724,N_20105);
xor U21520 (N_21520,N_20928,N_20241);
xnor U21521 (N_21521,N_20649,N_20808);
nand U21522 (N_21522,N_20778,N_21192);
and U21523 (N_21523,N_20891,N_21240);
or U21524 (N_21524,N_20953,N_21068);
xnor U21525 (N_21525,N_20730,N_20130);
xor U21526 (N_21526,N_20441,N_20758);
nor U21527 (N_21527,N_20204,N_20706);
and U21528 (N_21528,N_20358,N_21061);
xnor U21529 (N_21529,N_20539,N_20452);
nor U21530 (N_21530,N_20970,N_20831);
and U21531 (N_21531,N_21162,N_20601);
nand U21532 (N_21532,N_21230,N_20883);
xnor U21533 (N_21533,N_20416,N_20047);
nand U21534 (N_21534,N_20228,N_21183);
and U21535 (N_21535,N_21217,N_20813);
nand U21536 (N_21536,N_20792,N_20634);
and U21537 (N_21537,N_20294,N_20809);
or U21538 (N_21538,N_20610,N_21177);
xnor U21539 (N_21539,N_20001,N_20012);
and U21540 (N_21540,N_20834,N_20002);
and U21541 (N_21541,N_20713,N_20158);
and U21542 (N_21542,N_20802,N_20164);
nor U21543 (N_21543,N_20568,N_20902);
xor U21544 (N_21544,N_20077,N_20373);
nand U21545 (N_21545,N_21072,N_21053);
nor U21546 (N_21546,N_21037,N_20091);
or U21547 (N_21547,N_20327,N_20133);
nand U21548 (N_21548,N_20623,N_20115);
nor U21549 (N_21549,N_20698,N_20380);
xor U21550 (N_21550,N_20663,N_21167);
nor U21551 (N_21551,N_20696,N_20638);
or U21552 (N_21552,N_20143,N_20850);
xor U21553 (N_21553,N_20480,N_21219);
xnor U21554 (N_21554,N_20334,N_20438);
and U21555 (N_21555,N_21018,N_20756);
nand U21556 (N_21556,N_20726,N_20420);
nand U21557 (N_21557,N_20789,N_21185);
or U21558 (N_21558,N_20485,N_20783);
and U21559 (N_21559,N_21111,N_20033);
nor U21560 (N_21560,N_21126,N_20704);
or U21561 (N_21561,N_20699,N_20811);
nand U21562 (N_21562,N_20341,N_21124);
and U21563 (N_21563,N_21035,N_21186);
nand U21564 (N_21564,N_20647,N_21203);
nor U21565 (N_21565,N_20360,N_20700);
nand U21566 (N_21566,N_20745,N_20703);
and U21567 (N_21567,N_20448,N_20654);
or U21568 (N_21568,N_20736,N_20423);
and U21569 (N_21569,N_20222,N_20632);
xor U21570 (N_21570,N_20048,N_20260);
or U21571 (N_21571,N_20956,N_20727);
nand U21572 (N_21572,N_20775,N_20415);
and U21573 (N_21573,N_20198,N_20564);
xnor U21574 (N_21574,N_20780,N_20685);
xnor U21575 (N_21575,N_20508,N_20114);
nor U21576 (N_21576,N_20913,N_20345);
xnor U21577 (N_21577,N_20989,N_20032);
xnor U21578 (N_21578,N_20433,N_20646);
or U21579 (N_21579,N_21041,N_20805);
and U21580 (N_21580,N_21161,N_20719);
xnor U21581 (N_21581,N_20875,N_20973);
nand U21582 (N_21582,N_20037,N_21178);
and U21583 (N_21583,N_21086,N_21143);
nand U21584 (N_21584,N_20312,N_20658);
nor U21585 (N_21585,N_20616,N_20506);
or U21586 (N_21586,N_20571,N_20011);
and U21587 (N_21587,N_20102,N_20551);
nor U21588 (N_21588,N_20991,N_21179);
xor U21589 (N_21589,N_20355,N_20484);
and U21590 (N_21590,N_20311,N_21085);
nand U21591 (N_21591,N_20094,N_20495);
xor U21592 (N_21592,N_21043,N_21129);
nor U21593 (N_21593,N_20661,N_20862);
nor U21594 (N_21594,N_20254,N_20291);
and U21595 (N_21595,N_20829,N_20286);
and U21596 (N_21596,N_21151,N_21007);
xnor U21597 (N_21597,N_21008,N_20760);
and U21598 (N_21598,N_20562,N_20050);
nand U21599 (N_21599,N_21040,N_20645);
nand U21600 (N_21600,N_20242,N_21119);
nand U21601 (N_21601,N_20767,N_20159);
and U21602 (N_21602,N_20743,N_20389);
nand U21603 (N_21603,N_21223,N_20234);
or U21604 (N_21604,N_20854,N_20644);
nand U21605 (N_21605,N_20722,N_20839);
nor U21606 (N_21606,N_20467,N_20093);
xor U21607 (N_21607,N_20172,N_20505);
and U21608 (N_21608,N_20652,N_20428);
or U21609 (N_21609,N_20151,N_21004);
xnor U21610 (N_21610,N_20126,N_20086);
nor U21611 (N_21611,N_20218,N_21062);
nor U21612 (N_21612,N_20797,N_20078);
or U21613 (N_21613,N_21047,N_21015);
or U21614 (N_21614,N_21209,N_20677);
nor U21615 (N_21615,N_20463,N_21243);
xnor U21616 (N_21616,N_20986,N_20481);
and U21617 (N_21617,N_20492,N_21075);
nor U21618 (N_21618,N_20911,N_20357);
or U21619 (N_21619,N_20161,N_20005);
or U21620 (N_21620,N_21001,N_20432);
and U21621 (N_21621,N_20855,N_20274);
nand U21622 (N_21622,N_20052,N_20859);
and U21623 (N_21623,N_20951,N_20889);
nand U21624 (N_21624,N_21103,N_20261);
nand U21625 (N_21625,N_21173,N_21065);
nand U21626 (N_21626,N_20024,N_20402);
or U21627 (N_21627,N_20671,N_21245);
xnor U21628 (N_21628,N_20025,N_20796);
or U21629 (N_21629,N_20752,N_20019);
and U21630 (N_21630,N_20098,N_20982);
and U21631 (N_21631,N_21057,N_20806);
nor U21632 (N_21632,N_21099,N_20714);
nor U21633 (N_21633,N_20140,N_20202);
nand U21634 (N_21634,N_20259,N_20522);
and U21635 (N_21635,N_21066,N_20335);
xnor U21636 (N_21636,N_20803,N_20324);
xnor U21637 (N_21637,N_20595,N_20781);
or U21638 (N_21638,N_20604,N_20528);
or U21639 (N_21639,N_21071,N_21013);
and U21640 (N_21640,N_20457,N_20840);
xnor U21641 (N_21641,N_20042,N_20814);
or U21642 (N_21642,N_20447,N_20545);
or U21643 (N_21643,N_20878,N_21034);
and U21644 (N_21644,N_20555,N_20248);
and U21645 (N_21645,N_21054,N_20147);
nor U21646 (N_21646,N_20421,N_20127);
nor U21647 (N_21647,N_20737,N_20709);
xor U21648 (N_21648,N_20496,N_20605);
nand U21649 (N_21649,N_20753,N_20027);
or U21650 (N_21650,N_20763,N_20253);
nor U21651 (N_21651,N_20187,N_20288);
xor U21652 (N_21652,N_20229,N_20950);
or U21653 (N_21653,N_20354,N_20917);
nand U21654 (N_21654,N_20507,N_21114);
or U21655 (N_21655,N_20919,N_20964);
or U21656 (N_21656,N_20790,N_20641);
nor U21657 (N_21657,N_20527,N_20625);
and U21658 (N_21658,N_21201,N_20673);
xnor U21659 (N_21659,N_20262,N_20643);
nand U21660 (N_21660,N_20329,N_20022);
or U21661 (N_21661,N_20090,N_20226);
xor U21662 (N_21662,N_20591,N_21000);
and U21663 (N_21663,N_21134,N_20028);
nand U21664 (N_21664,N_20824,N_21044);
xnor U21665 (N_21665,N_20665,N_20650);
nor U21666 (N_21666,N_20303,N_20826);
nand U21667 (N_21667,N_21005,N_20356);
nor U21668 (N_21668,N_20321,N_20203);
or U21669 (N_21669,N_20880,N_20148);
nand U21670 (N_21670,N_20801,N_20653);
nand U21671 (N_21671,N_20534,N_21152);
xnor U21672 (N_21672,N_20450,N_20169);
nor U21673 (N_21673,N_21006,N_21176);
nor U21674 (N_21674,N_20104,N_20192);
xnor U21675 (N_21675,N_20721,N_21028);
and U21676 (N_21676,N_20963,N_20391);
or U21677 (N_21677,N_20759,N_20771);
and U21678 (N_21678,N_20209,N_20276);
and U21679 (N_21679,N_21187,N_20761);
nor U21680 (N_21680,N_20182,N_20697);
nand U21681 (N_21681,N_21208,N_21145);
xnor U21682 (N_21682,N_20281,N_20020);
or U21683 (N_21683,N_20828,N_20732);
nor U21684 (N_21684,N_20029,N_21225);
and U21685 (N_21685,N_20955,N_20788);
and U21686 (N_21686,N_20136,N_20399);
nor U21687 (N_21687,N_20660,N_20762);
nor U21688 (N_21688,N_20584,N_20425);
and U21689 (N_21689,N_20305,N_20728);
xnor U21690 (N_21690,N_20731,N_20350);
or U21691 (N_21691,N_20746,N_20394);
nor U21692 (N_21692,N_20031,N_20293);
nand U21693 (N_21693,N_20177,N_20856);
xor U21694 (N_21694,N_20901,N_20439);
nor U21695 (N_21695,N_20992,N_20317);
or U21696 (N_21696,N_20777,N_20718);
xnor U21697 (N_21697,N_20287,N_20411);
xor U21698 (N_21698,N_20186,N_20695);
nand U21699 (N_21699,N_20879,N_20707);
or U21700 (N_21700,N_20860,N_20322);
and U21701 (N_21701,N_20390,N_21042);
or U21702 (N_21702,N_21092,N_20353);
xor U21703 (N_21703,N_20686,N_20847);
or U21704 (N_21704,N_20007,N_20184);
nand U21705 (N_21705,N_20993,N_21160);
nor U21706 (N_21706,N_20134,N_20271);
and U21707 (N_21707,N_20030,N_20656);
xor U21708 (N_21708,N_20923,N_20188);
nand U21709 (N_21709,N_20043,N_20503);
nand U21710 (N_21710,N_20675,N_20628);
nor U21711 (N_21711,N_20836,N_20337);
or U21712 (N_21712,N_20067,N_21195);
nor U21713 (N_21713,N_20866,N_20088);
xnor U21714 (N_21714,N_20231,N_21211);
nor U21715 (N_21715,N_21241,N_20385);
or U21716 (N_21716,N_20189,N_20414);
nor U21717 (N_21717,N_20278,N_21233);
or U21718 (N_21718,N_20662,N_20118);
or U21719 (N_21719,N_20300,N_20376);
nor U21720 (N_21720,N_20486,N_20626);
xor U21721 (N_21721,N_20212,N_20113);
or U21722 (N_21722,N_20904,N_21058);
and U21723 (N_21723,N_21147,N_20501);
nand U21724 (N_21724,N_20981,N_20596);
xor U21725 (N_21725,N_20812,N_20711);
or U21726 (N_21726,N_20636,N_20183);
nand U21727 (N_21727,N_20600,N_21133);
or U21728 (N_21728,N_20217,N_21073);
xnor U21729 (N_21729,N_21158,N_21229);
xnor U21730 (N_21730,N_20864,N_20233);
and U21731 (N_21731,N_20861,N_20338);
or U21732 (N_21732,N_21193,N_20383);
and U21733 (N_21733,N_20519,N_20141);
or U21734 (N_21734,N_20069,N_20682);
and U21735 (N_21735,N_20667,N_20607);
xnor U21736 (N_21736,N_20734,N_20120);
nand U21737 (N_21737,N_20961,N_20602);
nor U21738 (N_21738,N_20606,N_20779);
nor U21739 (N_21739,N_20565,N_20406);
or U21740 (N_21740,N_20247,N_20468);
or U21741 (N_21741,N_21106,N_20482);
and U21742 (N_21742,N_20210,N_20265);
xor U21743 (N_21743,N_20776,N_20284);
or U21744 (N_21744,N_20770,N_20437);
nand U21745 (N_21745,N_20320,N_20280);
or U21746 (N_21746,N_20459,N_21238);
xnor U21747 (N_21747,N_20152,N_20691);
nor U21748 (N_21748,N_20252,N_20408);
nor U21749 (N_21749,N_20323,N_20071);
nor U21750 (N_21750,N_21200,N_20407);
nor U21751 (N_21751,N_20302,N_20900);
nor U21752 (N_21752,N_20559,N_20308);
or U21753 (N_21753,N_20359,N_21169);
xor U21754 (N_21754,N_20576,N_20892);
nand U21755 (N_21755,N_21024,N_21222);
nand U21756 (N_21756,N_21164,N_20155);
nor U21757 (N_21757,N_20368,N_20967);
nor U21758 (N_21758,N_20979,N_20267);
xnor U21759 (N_21759,N_20642,N_21060);
xnor U21760 (N_21760,N_21141,N_20949);
nand U21761 (N_21761,N_20316,N_20477);
xnor U21762 (N_21762,N_20388,N_20741);
xor U21763 (N_21763,N_20627,N_20540);
or U21764 (N_21764,N_20768,N_20313);
xor U21765 (N_21765,N_20664,N_20793);
nor U21766 (N_21766,N_20193,N_20712);
nor U21767 (N_21767,N_20095,N_20725);
nand U21768 (N_21768,N_20870,N_20678);
xnor U21769 (N_21769,N_20837,N_20597);
and U21770 (N_21770,N_20073,N_21026);
and U21771 (N_21771,N_20403,N_20589);
nor U21772 (N_21772,N_20690,N_20502);
nand U21773 (N_21773,N_20230,N_20994);
nor U21774 (N_21774,N_21090,N_21184);
nor U21775 (N_21775,N_20943,N_20419);
xor U21776 (N_21776,N_21014,N_20474);
or U21777 (N_21777,N_20035,N_20117);
and U21778 (N_21778,N_20057,N_20101);
nor U21779 (N_21779,N_20521,N_21202);
or U21780 (N_21780,N_20124,N_20785);
xnor U21781 (N_21781,N_20567,N_20821);
nand U21782 (N_21782,N_20074,N_21248);
or U21783 (N_21783,N_20689,N_20868);
nand U21784 (N_21784,N_20577,N_20449);
nand U21785 (N_21785,N_20583,N_20526);
nor U21786 (N_21786,N_21115,N_21214);
xnor U21787 (N_21787,N_21142,N_20952);
nand U21788 (N_21788,N_21132,N_21125);
nand U21789 (N_21789,N_20058,N_20163);
and U21790 (N_21790,N_20263,N_21010);
and U21791 (N_21791,N_20842,N_21244);
and U21792 (N_21792,N_21051,N_20563);
or U21793 (N_21793,N_20223,N_20694);
xor U21794 (N_21794,N_20395,N_21117);
xor U21795 (N_21795,N_20292,N_20393);
nand U21796 (N_21796,N_20367,N_20149);
or U21797 (N_21797,N_21023,N_20520);
nand U21798 (N_21798,N_21012,N_20319);
xor U21799 (N_21799,N_20518,N_20244);
or U21800 (N_21800,N_20370,N_21080);
nand U21801 (N_21801,N_20841,N_21148);
and U21802 (N_21802,N_20500,N_20843);
and U21803 (N_21803,N_20717,N_20946);
xor U21804 (N_21804,N_20975,N_20579);
nor U21805 (N_21805,N_21175,N_21036);
xor U21806 (N_21806,N_20637,N_20014);
nor U21807 (N_21807,N_20556,N_20146);
or U21808 (N_21808,N_20980,N_20285);
xor U21809 (N_21809,N_20440,N_20472);
and U21810 (N_21810,N_20849,N_20574);
and U21811 (N_21811,N_20948,N_20361);
xor U21812 (N_21812,N_20444,N_20497);
or U21813 (N_21813,N_20110,N_21210);
or U21814 (N_21814,N_21140,N_20523);
nor U21815 (N_21815,N_20655,N_20922);
and U21816 (N_21816,N_21237,N_20017);
nand U21817 (N_21817,N_20232,N_21094);
or U21818 (N_21818,N_20139,N_21139);
nor U21819 (N_21819,N_20676,N_20129);
and U21820 (N_21820,N_20176,N_20157);
nor U21821 (N_21821,N_20869,N_21017);
nand U21822 (N_21822,N_20072,N_20374);
and U21823 (N_21823,N_20968,N_21232);
and U21824 (N_21824,N_20910,N_20387);
and U21825 (N_21825,N_20958,N_20363);
nand U21826 (N_21826,N_20683,N_21188);
or U21827 (N_21827,N_20962,N_21205);
nand U21828 (N_21828,N_21131,N_21093);
xnor U21829 (N_21829,N_20240,N_20132);
xor U21830 (N_21830,N_21118,N_21171);
nand U21831 (N_21831,N_20938,N_20825);
nand U21832 (N_21832,N_20150,N_20791);
and U21833 (N_21833,N_20349,N_21221);
or U21834 (N_21834,N_20456,N_20915);
nor U21835 (N_21835,N_20621,N_20055);
xnor U21836 (N_21836,N_20772,N_20620);
xor U21837 (N_21837,N_20106,N_21163);
or U21838 (N_21838,N_20096,N_20575);
or U21839 (N_21839,N_20307,N_21112);
xnor U21840 (N_21840,N_20491,N_21166);
nand U21841 (N_21841,N_20185,N_20075);
or U21842 (N_21842,N_21150,N_20666);
nor U21843 (N_21843,N_20061,N_20138);
nor U21844 (N_21844,N_20173,N_20352);
nand U21845 (N_21845,N_20279,N_20827);
nor U21846 (N_21846,N_20815,N_20297);
xnor U21847 (N_21847,N_21135,N_20590);
nand U21848 (N_21848,N_21091,N_20515);
nand U21849 (N_21849,N_20493,N_21003);
and U21850 (N_21850,N_20912,N_21130);
nor U21851 (N_21851,N_21089,N_21157);
xnor U21852 (N_21852,N_20483,N_20087);
nor U21853 (N_21853,N_20844,N_21212);
and U21854 (N_21854,N_21020,N_20543);
nor U21855 (N_21855,N_20179,N_21226);
xnor U21856 (N_21856,N_20729,N_21049);
xnor U21857 (N_21857,N_20314,N_20036);
xor U21858 (N_21858,N_20896,N_21204);
nand U21859 (N_21859,N_20273,N_20925);
nor U21860 (N_21860,N_21227,N_21025);
and U21861 (N_21861,N_20573,N_20206);
nand U21862 (N_21862,N_20890,N_20371);
nor U21863 (N_21863,N_20538,N_20200);
nand U21864 (N_21864,N_21234,N_20040);
and U21865 (N_21865,N_20766,N_21059);
nand U21866 (N_21866,N_21206,N_20710);
xor U21867 (N_21867,N_20426,N_20435);
and U21868 (N_21868,N_20723,N_20773);
nand U21869 (N_21869,N_20863,N_20060);
xor U21870 (N_21870,N_20026,N_20541);
and U21871 (N_21871,N_20455,N_21081);
xnor U21872 (N_21872,N_20804,N_20881);
nand U21873 (N_21873,N_20070,N_21165);
nand U21874 (N_21874,N_20934,N_20464);
nor U21875 (N_21875,N_20872,N_20771);
and U21876 (N_21876,N_20676,N_20543);
or U21877 (N_21877,N_20167,N_21127);
and U21878 (N_21878,N_20304,N_20773);
xnor U21879 (N_21879,N_20346,N_20084);
and U21880 (N_21880,N_20383,N_20242);
or U21881 (N_21881,N_20932,N_20347);
nor U21882 (N_21882,N_20648,N_20094);
or U21883 (N_21883,N_21060,N_20206);
nand U21884 (N_21884,N_20945,N_20376);
xor U21885 (N_21885,N_20359,N_20892);
or U21886 (N_21886,N_21171,N_20908);
nand U21887 (N_21887,N_21171,N_20030);
nand U21888 (N_21888,N_20574,N_20920);
or U21889 (N_21889,N_20712,N_20508);
or U21890 (N_21890,N_20928,N_20345);
and U21891 (N_21891,N_20323,N_20226);
nand U21892 (N_21892,N_21175,N_20032);
nor U21893 (N_21893,N_20884,N_20940);
nor U21894 (N_21894,N_20241,N_20276);
xor U21895 (N_21895,N_20765,N_20657);
xor U21896 (N_21896,N_20252,N_20881);
or U21897 (N_21897,N_20442,N_21130);
and U21898 (N_21898,N_20724,N_21081);
nor U21899 (N_21899,N_21200,N_20287);
nand U21900 (N_21900,N_20297,N_20762);
nand U21901 (N_21901,N_20972,N_21068);
xor U21902 (N_21902,N_20930,N_20774);
nand U21903 (N_21903,N_20741,N_20018);
nor U21904 (N_21904,N_21205,N_21202);
or U21905 (N_21905,N_20934,N_20663);
or U21906 (N_21906,N_20605,N_21105);
nor U21907 (N_21907,N_20604,N_21174);
and U21908 (N_21908,N_20345,N_20144);
nand U21909 (N_21909,N_20785,N_20879);
or U21910 (N_21910,N_20786,N_21167);
xnor U21911 (N_21911,N_20653,N_20094);
and U21912 (N_21912,N_20607,N_21103);
nand U21913 (N_21913,N_20946,N_20471);
or U21914 (N_21914,N_20956,N_20625);
nand U21915 (N_21915,N_20145,N_21092);
nor U21916 (N_21916,N_20785,N_20993);
and U21917 (N_21917,N_20656,N_20633);
or U21918 (N_21918,N_20726,N_20974);
or U21919 (N_21919,N_20324,N_20852);
xor U21920 (N_21920,N_20257,N_21080);
and U21921 (N_21921,N_20729,N_20382);
and U21922 (N_21922,N_20635,N_20678);
xnor U21923 (N_21923,N_21137,N_20584);
nor U21924 (N_21924,N_21013,N_20631);
nand U21925 (N_21925,N_20626,N_20927);
xor U21926 (N_21926,N_20558,N_20054);
nor U21927 (N_21927,N_21180,N_21109);
nand U21928 (N_21928,N_21093,N_20495);
nor U21929 (N_21929,N_20535,N_21063);
nor U21930 (N_21930,N_20951,N_20369);
or U21931 (N_21931,N_20852,N_20066);
or U21932 (N_21932,N_20352,N_20598);
nand U21933 (N_21933,N_21165,N_20848);
nand U21934 (N_21934,N_20948,N_20431);
nor U21935 (N_21935,N_20247,N_20764);
nand U21936 (N_21936,N_21186,N_21175);
and U21937 (N_21937,N_20518,N_20091);
and U21938 (N_21938,N_20716,N_20889);
nand U21939 (N_21939,N_20195,N_20359);
xor U21940 (N_21940,N_21135,N_20647);
and U21941 (N_21941,N_20986,N_20300);
xor U21942 (N_21942,N_20353,N_20203);
nand U21943 (N_21943,N_21054,N_20782);
and U21944 (N_21944,N_20589,N_21216);
nor U21945 (N_21945,N_20324,N_20624);
nand U21946 (N_21946,N_20384,N_21191);
xor U21947 (N_21947,N_20260,N_21244);
nand U21948 (N_21948,N_21021,N_20461);
xnor U21949 (N_21949,N_21023,N_20101);
xnor U21950 (N_21950,N_20793,N_20098);
or U21951 (N_21951,N_20201,N_20688);
xor U21952 (N_21952,N_21024,N_20329);
or U21953 (N_21953,N_20862,N_20520);
nor U21954 (N_21954,N_20070,N_20470);
or U21955 (N_21955,N_20523,N_21231);
and U21956 (N_21956,N_21063,N_21007);
nor U21957 (N_21957,N_21125,N_21205);
xnor U21958 (N_21958,N_20504,N_20090);
nand U21959 (N_21959,N_20175,N_20473);
nor U21960 (N_21960,N_21158,N_20510);
and U21961 (N_21961,N_20234,N_20224);
and U21962 (N_21962,N_20171,N_20772);
nand U21963 (N_21963,N_20168,N_20210);
nor U21964 (N_21964,N_20469,N_21086);
nand U21965 (N_21965,N_20207,N_20284);
nor U21966 (N_21966,N_20206,N_20273);
xor U21967 (N_21967,N_20027,N_20103);
nor U21968 (N_21968,N_20971,N_20797);
xnor U21969 (N_21969,N_21046,N_20275);
xnor U21970 (N_21970,N_21060,N_20139);
or U21971 (N_21971,N_21077,N_20230);
or U21972 (N_21972,N_21204,N_20157);
and U21973 (N_21973,N_20448,N_20291);
nand U21974 (N_21974,N_20864,N_20409);
nand U21975 (N_21975,N_20976,N_21146);
nand U21976 (N_21976,N_20125,N_20658);
and U21977 (N_21977,N_20765,N_20024);
and U21978 (N_21978,N_20272,N_20011);
xnor U21979 (N_21979,N_20134,N_21215);
nor U21980 (N_21980,N_20468,N_20802);
and U21981 (N_21981,N_20544,N_21194);
nor U21982 (N_21982,N_21105,N_20030);
xor U21983 (N_21983,N_21196,N_20439);
nor U21984 (N_21984,N_20922,N_20342);
or U21985 (N_21985,N_20568,N_21005);
nand U21986 (N_21986,N_20462,N_21075);
or U21987 (N_21987,N_20061,N_21238);
and U21988 (N_21988,N_20866,N_20376);
or U21989 (N_21989,N_20044,N_20875);
xor U21990 (N_21990,N_20080,N_20696);
and U21991 (N_21991,N_20668,N_20374);
or U21992 (N_21992,N_20662,N_20000);
xnor U21993 (N_21993,N_21202,N_20376);
xnor U21994 (N_21994,N_20433,N_21067);
xor U21995 (N_21995,N_20632,N_20503);
nand U21996 (N_21996,N_20166,N_20479);
nor U21997 (N_21997,N_20934,N_20773);
nor U21998 (N_21998,N_20615,N_20930);
nor U21999 (N_21999,N_20418,N_21109);
and U22000 (N_22000,N_20739,N_21075);
nand U22001 (N_22001,N_20117,N_21007);
and U22002 (N_22002,N_20991,N_21072);
nand U22003 (N_22003,N_20586,N_20702);
or U22004 (N_22004,N_20578,N_20057);
or U22005 (N_22005,N_20225,N_20684);
xor U22006 (N_22006,N_20417,N_20441);
or U22007 (N_22007,N_20801,N_20399);
and U22008 (N_22008,N_21131,N_21248);
nand U22009 (N_22009,N_20998,N_20445);
xnor U22010 (N_22010,N_20347,N_20999);
and U22011 (N_22011,N_20072,N_20985);
nor U22012 (N_22012,N_20269,N_21107);
and U22013 (N_22013,N_20717,N_21076);
and U22014 (N_22014,N_20676,N_20368);
xor U22015 (N_22015,N_20062,N_20786);
xor U22016 (N_22016,N_20986,N_20594);
or U22017 (N_22017,N_20669,N_20257);
and U22018 (N_22018,N_20931,N_20605);
nand U22019 (N_22019,N_20361,N_21244);
xor U22020 (N_22020,N_20091,N_20507);
nand U22021 (N_22021,N_21091,N_21067);
nand U22022 (N_22022,N_21075,N_20546);
nand U22023 (N_22023,N_20658,N_20331);
and U22024 (N_22024,N_20774,N_20474);
nor U22025 (N_22025,N_20904,N_20844);
xnor U22026 (N_22026,N_20419,N_20725);
xnor U22027 (N_22027,N_20450,N_20951);
or U22028 (N_22028,N_20490,N_20289);
or U22029 (N_22029,N_20975,N_20357);
nand U22030 (N_22030,N_20731,N_20710);
nor U22031 (N_22031,N_20646,N_20784);
xor U22032 (N_22032,N_20571,N_20199);
xor U22033 (N_22033,N_20339,N_20844);
xor U22034 (N_22034,N_21095,N_20448);
xor U22035 (N_22035,N_20141,N_20245);
xor U22036 (N_22036,N_20078,N_20147);
and U22037 (N_22037,N_20671,N_20563);
and U22038 (N_22038,N_21244,N_20957);
or U22039 (N_22039,N_20131,N_20763);
nor U22040 (N_22040,N_21238,N_21135);
nand U22041 (N_22041,N_20558,N_21078);
nand U22042 (N_22042,N_20700,N_21179);
xor U22043 (N_22043,N_21024,N_20277);
or U22044 (N_22044,N_20544,N_20690);
xor U22045 (N_22045,N_20550,N_20619);
nand U22046 (N_22046,N_20256,N_20501);
xor U22047 (N_22047,N_21050,N_20578);
or U22048 (N_22048,N_20044,N_20160);
nor U22049 (N_22049,N_20888,N_20982);
nor U22050 (N_22050,N_21219,N_20964);
or U22051 (N_22051,N_20864,N_20602);
nand U22052 (N_22052,N_20259,N_20066);
nand U22053 (N_22053,N_20284,N_20940);
nor U22054 (N_22054,N_20062,N_20183);
nor U22055 (N_22055,N_21230,N_20420);
nor U22056 (N_22056,N_20460,N_20363);
xnor U22057 (N_22057,N_21002,N_20626);
nand U22058 (N_22058,N_20714,N_21058);
and U22059 (N_22059,N_20754,N_20017);
nor U22060 (N_22060,N_21089,N_21133);
nor U22061 (N_22061,N_20539,N_20143);
or U22062 (N_22062,N_20564,N_21000);
or U22063 (N_22063,N_20384,N_20409);
and U22064 (N_22064,N_21177,N_20693);
xor U22065 (N_22065,N_20430,N_20082);
and U22066 (N_22066,N_20927,N_20816);
xnor U22067 (N_22067,N_20949,N_21084);
nor U22068 (N_22068,N_20189,N_20789);
xor U22069 (N_22069,N_20627,N_20285);
xnor U22070 (N_22070,N_20434,N_20566);
and U22071 (N_22071,N_21133,N_20471);
nor U22072 (N_22072,N_20859,N_20847);
or U22073 (N_22073,N_20277,N_21208);
nor U22074 (N_22074,N_20309,N_20582);
or U22075 (N_22075,N_20126,N_20985);
and U22076 (N_22076,N_20901,N_21091);
xnor U22077 (N_22077,N_20359,N_20822);
nand U22078 (N_22078,N_20438,N_20410);
nand U22079 (N_22079,N_20930,N_20660);
and U22080 (N_22080,N_20011,N_20994);
nor U22081 (N_22081,N_20222,N_21075);
and U22082 (N_22082,N_20803,N_20465);
nand U22083 (N_22083,N_20849,N_20679);
and U22084 (N_22084,N_20938,N_20530);
xnor U22085 (N_22085,N_20570,N_20807);
xnor U22086 (N_22086,N_20403,N_20415);
nand U22087 (N_22087,N_20650,N_20816);
and U22088 (N_22088,N_20869,N_20686);
nor U22089 (N_22089,N_21119,N_20602);
xor U22090 (N_22090,N_21004,N_20820);
or U22091 (N_22091,N_20298,N_20277);
xor U22092 (N_22092,N_20378,N_21070);
nor U22093 (N_22093,N_20747,N_21080);
or U22094 (N_22094,N_20317,N_20729);
and U22095 (N_22095,N_20481,N_21215);
xnor U22096 (N_22096,N_21058,N_21203);
xnor U22097 (N_22097,N_20996,N_20354);
xor U22098 (N_22098,N_20572,N_20331);
or U22099 (N_22099,N_21104,N_21199);
xor U22100 (N_22100,N_20998,N_21034);
nand U22101 (N_22101,N_20158,N_21126);
nor U22102 (N_22102,N_20815,N_21075);
and U22103 (N_22103,N_20698,N_20222);
and U22104 (N_22104,N_20265,N_20970);
nor U22105 (N_22105,N_20232,N_20638);
and U22106 (N_22106,N_20701,N_20185);
xor U22107 (N_22107,N_20281,N_20025);
nor U22108 (N_22108,N_20878,N_20695);
and U22109 (N_22109,N_20630,N_20133);
xnor U22110 (N_22110,N_20682,N_20984);
or U22111 (N_22111,N_21115,N_20810);
nand U22112 (N_22112,N_21032,N_21099);
nand U22113 (N_22113,N_20978,N_20613);
nand U22114 (N_22114,N_21124,N_20248);
and U22115 (N_22115,N_20926,N_20086);
nor U22116 (N_22116,N_20960,N_20403);
or U22117 (N_22117,N_20666,N_20070);
and U22118 (N_22118,N_21130,N_20301);
and U22119 (N_22119,N_20686,N_20137);
and U22120 (N_22120,N_20360,N_21007);
or U22121 (N_22121,N_20649,N_20348);
or U22122 (N_22122,N_20523,N_21175);
nor U22123 (N_22123,N_21021,N_21072);
and U22124 (N_22124,N_20623,N_20327);
or U22125 (N_22125,N_21103,N_21063);
xor U22126 (N_22126,N_21179,N_20836);
or U22127 (N_22127,N_20213,N_20512);
nor U22128 (N_22128,N_20175,N_21019);
xnor U22129 (N_22129,N_20529,N_20948);
nor U22130 (N_22130,N_20155,N_20329);
or U22131 (N_22131,N_20421,N_20779);
nor U22132 (N_22132,N_20432,N_21086);
nor U22133 (N_22133,N_20188,N_20184);
nand U22134 (N_22134,N_20741,N_20319);
xnor U22135 (N_22135,N_21052,N_20458);
nand U22136 (N_22136,N_21103,N_20092);
nand U22137 (N_22137,N_20221,N_20733);
nand U22138 (N_22138,N_20565,N_20026);
xnor U22139 (N_22139,N_20791,N_20525);
and U22140 (N_22140,N_20134,N_21061);
nand U22141 (N_22141,N_20958,N_20781);
or U22142 (N_22142,N_20535,N_20951);
nor U22143 (N_22143,N_20946,N_20307);
xnor U22144 (N_22144,N_20509,N_20233);
nand U22145 (N_22145,N_20782,N_20499);
and U22146 (N_22146,N_20575,N_21108);
and U22147 (N_22147,N_20146,N_20986);
xor U22148 (N_22148,N_20826,N_20512);
or U22149 (N_22149,N_20828,N_20065);
nand U22150 (N_22150,N_20254,N_20724);
nand U22151 (N_22151,N_20831,N_20019);
and U22152 (N_22152,N_21110,N_20916);
xnor U22153 (N_22153,N_21203,N_21121);
and U22154 (N_22154,N_21179,N_20051);
and U22155 (N_22155,N_21204,N_20805);
nand U22156 (N_22156,N_20510,N_20855);
or U22157 (N_22157,N_20753,N_20914);
nand U22158 (N_22158,N_20931,N_20626);
nor U22159 (N_22159,N_20309,N_20809);
nand U22160 (N_22160,N_20303,N_21060);
xnor U22161 (N_22161,N_21225,N_20277);
nand U22162 (N_22162,N_20533,N_20315);
nand U22163 (N_22163,N_20536,N_20059);
or U22164 (N_22164,N_21126,N_20210);
nand U22165 (N_22165,N_20688,N_21139);
xnor U22166 (N_22166,N_20987,N_20688);
xor U22167 (N_22167,N_20471,N_20985);
nand U22168 (N_22168,N_20854,N_20935);
and U22169 (N_22169,N_20695,N_20572);
nand U22170 (N_22170,N_20246,N_20620);
xnor U22171 (N_22171,N_20041,N_20535);
xor U22172 (N_22172,N_21195,N_20680);
xnor U22173 (N_22173,N_20461,N_21111);
and U22174 (N_22174,N_20584,N_20998);
nand U22175 (N_22175,N_20109,N_20203);
and U22176 (N_22176,N_20496,N_20220);
or U22177 (N_22177,N_20511,N_20334);
or U22178 (N_22178,N_21204,N_20048);
or U22179 (N_22179,N_20535,N_20182);
nor U22180 (N_22180,N_20978,N_20831);
xnor U22181 (N_22181,N_20671,N_20342);
or U22182 (N_22182,N_20303,N_20880);
or U22183 (N_22183,N_21086,N_20676);
and U22184 (N_22184,N_20339,N_20664);
nor U22185 (N_22185,N_20326,N_20724);
or U22186 (N_22186,N_20981,N_20911);
and U22187 (N_22187,N_20719,N_20372);
nand U22188 (N_22188,N_20637,N_20726);
nand U22189 (N_22189,N_20823,N_20162);
xnor U22190 (N_22190,N_20504,N_20007);
nand U22191 (N_22191,N_20684,N_20656);
nor U22192 (N_22192,N_20249,N_20883);
and U22193 (N_22193,N_20176,N_20935);
and U22194 (N_22194,N_20103,N_20373);
nor U22195 (N_22195,N_20951,N_21240);
and U22196 (N_22196,N_20140,N_20417);
or U22197 (N_22197,N_20712,N_20494);
xnor U22198 (N_22198,N_20371,N_20162);
and U22199 (N_22199,N_20916,N_20620);
or U22200 (N_22200,N_20753,N_20342);
xor U22201 (N_22201,N_20353,N_20908);
xor U22202 (N_22202,N_21023,N_20622);
xnor U22203 (N_22203,N_20415,N_20411);
or U22204 (N_22204,N_20968,N_20622);
and U22205 (N_22205,N_20244,N_20014);
nor U22206 (N_22206,N_20369,N_20751);
nor U22207 (N_22207,N_20361,N_20343);
or U22208 (N_22208,N_20239,N_20801);
nor U22209 (N_22209,N_21132,N_20153);
nand U22210 (N_22210,N_20150,N_20738);
nand U22211 (N_22211,N_20032,N_20542);
xor U22212 (N_22212,N_20401,N_20244);
nand U22213 (N_22213,N_20021,N_20628);
and U22214 (N_22214,N_20528,N_20072);
xnor U22215 (N_22215,N_20602,N_21009);
nor U22216 (N_22216,N_20676,N_20959);
nand U22217 (N_22217,N_20891,N_20666);
and U22218 (N_22218,N_20864,N_20321);
nand U22219 (N_22219,N_20073,N_20143);
xnor U22220 (N_22220,N_20631,N_20762);
or U22221 (N_22221,N_21001,N_20189);
and U22222 (N_22222,N_20881,N_20257);
nor U22223 (N_22223,N_20055,N_20648);
and U22224 (N_22224,N_20780,N_20261);
nand U22225 (N_22225,N_20483,N_21234);
xor U22226 (N_22226,N_20450,N_20255);
and U22227 (N_22227,N_20083,N_20781);
nor U22228 (N_22228,N_20781,N_21241);
xor U22229 (N_22229,N_20383,N_21048);
nor U22230 (N_22230,N_20415,N_20268);
nand U22231 (N_22231,N_20373,N_20145);
nor U22232 (N_22232,N_20866,N_20349);
nor U22233 (N_22233,N_20789,N_20539);
nor U22234 (N_22234,N_20620,N_20226);
or U22235 (N_22235,N_20963,N_20594);
nand U22236 (N_22236,N_20873,N_20563);
nand U22237 (N_22237,N_21049,N_20159);
or U22238 (N_22238,N_20283,N_20372);
xor U22239 (N_22239,N_20960,N_20897);
nand U22240 (N_22240,N_20306,N_21093);
nand U22241 (N_22241,N_21194,N_20431);
and U22242 (N_22242,N_20676,N_21109);
and U22243 (N_22243,N_20910,N_20224);
or U22244 (N_22244,N_20916,N_21201);
or U22245 (N_22245,N_20065,N_21070);
nand U22246 (N_22246,N_21058,N_20515);
xor U22247 (N_22247,N_20825,N_20470);
nand U22248 (N_22248,N_20788,N_20669);
and U22249 (N_22249,N_20469,N_20164);
xnor U22250 (N_22250,N_20168,N_20708);
or U22251 (N_22251,N_20069,N_21165);
or U22252 (N_22252,N_21037,N_21082);
xor U22253 (N_22253,N_20761,N_20576);
or U22254 (N_22254,N_21227,N_20359);
nand U22255 (N_22255,N_20696,N_20646);
nor U22256 (N_22256,N_20812,N_20084);
or U22257 (N_22257,N_21136,N_20232);
and U22258 (N_22258,N_20949,N_20574);
nand U22259 (N_22259,N_20333,N_20270);
or U22260 (N_22260,N_20347,N_20130);
or U22261 (N_22261,N_20578,N_20112);
and U22262 (N_22262,N_20690,N_20044);
or U22263 (N_22263,N_20357,N_20008);
xnor U22264 (N_22264,N_20802,N_20439);
or U22265 (N_22265,N_21086,N_20650);
xor U22266 (N_22266,N_20354,N_20680);
nor U22267 (N_22267,N_20025,N_20817);
nor U22268 (N_22268,N_21117,N_20054);
xnor U22269 (N_22269,N_20568,N_20727);
xnor U22270 (N_22270,N_20562,N_20012);
nor U22271 (N_22271,N_20973,N_20576);
nand U22272 (N_22272,N_20268,N_20033);
nor U22273 (N_22273,N_20233,N_20494);
nor U22274 (N_22274,N_20295,N_20116);
or U22275 (N_22275,N_21207,N_20676);
nand U22276 (N_22276,N_20043,N_20208);
nor U22277 (N_22277,N_20087,N_20783);
and U22278 (N_22278,N_20451,N_21109);
and U22279 (N_22279,N_20137,N_20864);
xnor U22280 (N_22280,N_20656,N_21218);
xor U22281 (N_22281,N_20603,N_20865);
xnor U22282 (N_22282,N_20442,N_20053);
and U22283 (N_22283,N_20809,N_20340);
nor U22284 (N_22284,N_20205,N_20253);
xnor U22285 (N_22285,N_21026,N_21193);
xnor U22286 (N_22286,N_21175,N_20173);
nand U22287 (N_22287,N_20644,N_20152);
nand U22288 (N_22288,N_20321,N_21061);
nor U22289 (N_22289,N_20366,N_21102);
or U22290 (N_22290,N_20359,N_20570);
and U22291 (N_22291,N_20034,N_20605);
nor U22292 (N_22292,N_20563,N_20978);
nor U22293 (N_22293,N_20801,N_20856);
and U22294 (N_22294,N_20368,N_20922);
or U22295 (N_22295,N_20605,N_20098);
xnor U22296 (N_22296,N_21026,N_20241);
nand U22297 (N_22297,N_20075,N_20428);
and U22298 (N_22298,N_21033,N_21175);
or U22299 (N_22299,N_20081,N_20284);
nor U22300 (N_22300,N_20642,N_20486);
xnor U22301 (N_22301,N_21248,N_20769);
and U22302 (N_22302,N_20227,N_20884);
and U22303 (N_22303,N_20510,N_20979);
or U22304 (N_22304,N_20437,N_20656);
and U22305 (N_22305,N_21227,N_21217);
nor U22306 (N_22306,N_20033,N_20951);
xnor U22307 (N_22307,N_20845,N_20373);
or U22308 (N_22308,N_20693,N_21206);
nor U22309 (N_22309,N_21132,N_20185);
nand U22310 (N_22310,N_20895,N_20276);
xor U22311 (N_22311,N_20309,N_21187);
nand U22312 (N_22312,N_21130,N_20399);
nor U22313 (N_22313,N_20397,N_20074);
nor U22314 (N_22314,N_20118,N_20420);
xor U22315 (N_22315,N_20010,N_20462);
and U22316 (N_22316,N_20562,N_20341);
nand U22317 (N_22317,N_20194,N_20569);
or U22318 (N_22318,N_21113,N_20642);
nand U22319 (N_22319,N_20874,N_20477);
and U22320 (N_22320,N_20254,N_20500);
nand U22321 (N_22321,N_21108,N_20156);
or U22322 (N_22322,N_20042,N_20121);
xnor U22323 (N_22323,N_21045,N_21061);
nand U22324 (N_22324,N_20886,N_20794);
nand U22325 (N_22325,N_20386,N_21086);
or U22326 (N_22326,N_21155,N_20076);
nand U22327 (N_22327,N_20573,N_20086);
nand U22328 (N_22328,N_21080,N_20363);
or U22329 (N_22329,N_21177,N_20371);
and U22330 (N_22330,N_21118,N_20801);
nor U22331 (N_22331,N_20384,N_20537);
nand U22332 (N_22332,N_20096,N_20197);
and U22333 (N_22333,N_20257,N_20838);
or U22334 (N_22334,N_21193,N_20121);
or U22335 (N_22335,N_20584,N_20662);
nand U22336 (N_22336,N_20555,N_20969);
nand U22337 (N_22337,N_20977,N_20724);
nand U22338 (N_22338,N_20916,N_20040);
xor U22339 (N_22339,N_20114,N_20116);
xnor U22340 (N_22340,N_20920,N_20536);
xnor U22341 (N_22341,N_20435,N_20508);
nor U22342 (N_22342,N_20834,N_20564);
xnor U22343 (N_22343,N_20919,N_20557);
and U22344 (N_22344,N_20165,N_20696);
or U22345 (N_22345,N_20685,N_21141);
nor U22346 (N_22346,N_21211,N_20887);
or U22347 (N_22347,N_20192,N_20423);
nor U22348 (N_22348,N_20462,N_20614);
nor U22349 (N_22349,N_20075,N_20514);
xor U22350 (N_22350,N_20650,N_20180);
nand U22351 (N_22351,N_20940,N_20791);
or U22352 (N_22352,N_20339,N_20967);
xnor U22353 (N_22353,N_21176,N_20892);
xnor U22354 (N_22354,N_20246,N_20762);
nand U22355 (N_22355,N_20846,N_20498);
and U22356 (N_22356,N_20555,N_20336);
nor U22357 (N_22357,N_20299,N_20928);
and U22358 (N_22358,N_21037,N_20679);
nand U22359 (N_22359,N_21121,N_20152);
nand U22360 (N_22360,N_21229,N_20471);
nor U22361 (N_22361,N_21120,N_20603);
nand U22362 (N_22362,N_20312,N_20317);
and U22363 (N_22363,N_20236,N_20812);
xor U22364 (N_22364,N_20721,N_20038);
nor U22365 (N_22365,N_20282,N_20315);
nor U22366 (N_22366,N_20331,N_20365);
xor U22367 (N_22367,N_21022,N_20689);
xnor U22368 (N_22368,N_20629,N_21116);
nor U22369 (N_22369,N_20039,N_20859);
or U22370 (N_22370,N_20076,N_20224);
or U22371 (N_22371,N_20791,N_20937);
xnor U22372 (N_22372,N_21145,N_20423);
or U22373 (N_22373,N_21239,N_21187);
nand U22374 (N_22374,N_20713,N_21046);
xnor U22375 (N_22375,N_21147,N_20650);
or U22376 (N_22376,N_20859,N_20056);
nor U22377 (N_22377,N_20998,N_20212);
and U22378 (N_22378,N_20435,N_20364);
nand U22379 (N_22379,N_20501,N_20652);
and U22380 (N_22380,N_21068,N_20504);
nand U22381 (N_22381,N_21184,N_20602);
and U22382 (N_22382,N_20135,N_20162);
nor U22383 (N_22383,N_20176,N_20662);
nand U22384 (N_22384,N_20397,N_20226);
or U22385 (N_22385,N_20067,N_20875);
and U22386 (N_22386,N_20272,N_20483);
xor U22387 (N_22387,N_20464,N_20863);
xor U22388 (N_22388,N_20051,N_20581);
nand U22389 (N_22389,N_20333,N_20639);
nand U22390 (N_22390,N_21005,N_20200);
xor U22391 (N_22391,N_20482,N_20919);
and U22392 (N_22392,N_20667,N_20340);
or U22393 (N_22393,N_21194,N_20138);
xnor U22394 (N_22394,N_20873,N_20331);
nand U22395 (N_22395,N_21020,N_20049);
nor U22396 (N_22396,N_20035,N_20193);
and U22397 (N_22397,N_21052,N_20796);
nand U22398 (N_22398,N_20821,N_20152);
nor U22399 (N_22399,N_21181,N_20459);
xnor U22400 (N_22400,N_20219,N_20209);
nor U22401 (N_22401,N_20435,N_20584);
and U22402 (N_22402,N_20885,N_20937);
and U22403 (N_22403,N_20191,N_20396);
nor U22404 (N_22404,N_20611,N_20791);
nand U22405 (N_22405,N_21147,N_20809);
and U22406 (N_22406,N_20076,N_21176);
and U22407 (N_22407,N_20332,N_20616);
xor U22408 (N_22408,N_20546,N_21194);
nand U22409 (N_22409,N_20865,N_21158);
nand U22410 (N_22410,N_20123,N_20815);
nor U22411 (N_22411,N_20791,N_20645);
or U22412 (N_22412,N_20654,N_20255);
xnor U22413 (N_22413,N_20455,N_20188);
xnor U22414 (N_22414,N_20550,N_21093);
and U22415 (N_22415,N_21099,N_20870);
xor U22416 (N_22416,N_20527,N_20615);
xnor U22417 (N_22417,N_20361,N_20015);
and U22418 (N_22418,N_20169,N_20395);
or U22419 (N_22419,N_20792,N_20672);
nand U22420 (N_22420,N_20957,N_20585);
and U22421 (N_22421,N_20368,N_21172);
xor U22422 (N_22422,N_20517,N_20878);
and U22423 (N_22423,N_20996,N_20747);
nor U22424 (N_22424,N_20587,N_20794);
and U22425 (N_22425,N_20945,N_21039);
or U22426 (N_22426,N_21081,N_21111);
xor U22427 (N_22427,N_20062,N_20619);
and U22428 (N_22428,N_20447,N_20839);
or U22429 (N_22429,N_20853,N_20070);
nor U22430 (N_22430,N_20924,N_21175);
nor U22431 (N_22431,N_20077,N_20692);
nor U22432 (N_22432,N_20980,N_20339);
and U22433 (N_22433,N_20617,N_21220);
nor U22434 (N_22434,N_20318,N_21093);
nor U22435 (N_22435,N_20649,N_21225);
nor U22436 (N_22436,N_21219,N_20333);
or U22437 (N_22437,N_20568,N_20385);
and U22438 (N_22438,N_20311,N_20655);
xnor U22439 (N_22439,N_20458,N_21206);
or U22440 (N_22440,N_20555,N_20064);
or U22441 (N_22441,N_20785,N_20454);
nand U22442 (N_22442,N_20479,N_20385);
or U22443 (N_22443,N_20454,N_20233);
xnor U22444 (N_22444,N_20482,N_20233);
nor U22445 (N_22445,N_20590,N_20776);
nor U22446 (N_22446,N_20797,N_20334);
xnor U22447 (N_22447,N_21008,N_20219);
nor U22448 (N_22448,N_21030,N_20826);
and U22449 (N_22449,N_20107,N_20338);
and U22450 (N_22450,N_21148,N_21106);
nor U22451 (N_22451,N_20693,N_20452);
or U22452 (N_22452,N_20277,N_20171);
or U22453 (N_22453,N_20554,N_20951);
or U22454 (N_22454,N_20170,N_21057);
xor U22455 (N_22455,N_20644,N_20461);
nand U22456 (N_22456,N_20395,N_20905);
and U22457 (N_22457,N_20062,N_20823);
nand U22458 (N_22458,N_20912,N_20696);
xnor U22459 (N_22459,N_20510,N_20496);
and U22460 (N_22460,N_20045,N_20978);
xor U22461 (N_22461,N_21151,N_21004);
and U22462 (N_22462,N_21035,N_20250);
xor U22463 (N_22463,N_20249,N_21017);
xnor U22464 (N_22464,N_20768,N_21059);
and U22465 (N_22465,N_20044,N_20644);
or U22466 (N_22466,N_20489,N_20473);
nand U22467 (N_22467,N_20320,N_20103);
xor U22468 (N_22468,N_20314,N_20285);
nand U22469 (N_22469,N_20542,N_20155);
nor U22470 (N_22470,N_20576,N_20601);
nor U22471 (N_22471,N_20055,N_20151);
nand U22472 (N_22472,N_20911,N_20725);
xnor U22473 (N_22473,N_20955,N_21078);
xnor U22474 (N_22474,N_20079,N_20863);
and U22475 (N_22475,N_20585,N_21008);
nand U22476 (N_22476,N_20487,N_20415);
xor U22477 (N_22477,N_20583,N_20031);
or U22478 (N_22478,N_20225,N_20680);
xnor U22479 (N_22479,N_20302,N_20462);
and U22480 (N_22480,N_20997,N_20123);
or U22481 (N_22481,N_20513,N_20944);
xor U22482 (N_22482,N_21021,N_20046);
and U22483 (N_22483,N_20437,N_20746);
or U22484 (N_22484,N_20435,N_20442);
nand U22485 (N_22485,N_20118,N_21236);
nor U22486 (N_22486,N_20928,N_20945);
xnor U22487 (N_22487,N_20970,N_20169);
or U22488 (N_22488,N_21133,N_20605);
and U22489 (N_22489,N_20729,N_21056);
nor U22490 (N_22490,N_20999,N_20209);
nor U22491 (N_22491,N_21105,N_20212);
nor U22492 (N_22492,N_20828,N_20038);
nor U22493 (N_22493,N_20501,N_20270);
nor U22494 (N_22494,N_20116,N_20029);
xnor U22495 (N_22495,N_20499,N_20605);
xnor U22496 (N_22496,N_21164,N_20109);
nand U22497 (N_22497,N_20047,N_20773);
nor U22498 (N_22498,N_20560,N_21166);
nor U22499 (N_22499,N_20619,N_20480);
nand U22500 (N_22500,N_21833,N_21827);
nand U22501 (N_22501,N_21427,N_21678);
or U22502 (N_22502,N_22134,N_21900);
and U22503 (N_22503,N_22248,N_21936);
nor U22504 (N_22504,N_21414,N_22462);
xnor U22505 (N_22505,N_21912,N_22475);
nor U22506 (N_22506,N_21520,N_22394);
nor U22507 (N_22507,N_21880,N_22315);
and U22508 (N_22508,N_21662,N_22142);
and U22509 (N_22509,N_21945,N_22321);
nor U22510 (N_22510,N_21467,N_21637);
nor U22511 (N_22511,N_22211,N_21404);
xnor U22512 (N_22512,N_21633,N_22337);
nand U22513 (N_22513,N_22139,N_21526);
and U22514 (N_22514,N_21680,N_21558);
and U22515 (N_22515,N_21875,N_21596);
xnor U22516 (N_22516,N_21582,N_22207);
nor U22517 (N_22517,N_21436,N_21787);
xnor U22518 (N_22518,N_22178,N_22392);
xor U22519 (N_22519,N_21547,N_22036);
xnor U22520 (N_22520,N_21598,N_21459);
nand U22521 (N_22521,N_21529,N_21472);
or U22522 (N_22522,N_21683,N_22195);
and U22523 (N_22523,N_21870,N_22232);
or U22524 (N_22524,N_22004,N_22084);
and U22525 (N_22525,N_21469,N_22258);
nor U22526 (N_22526,N_21341,N_21280);
xnor U22527 (N_22527,N_21294,N_21758);
and U22528 (N_22528,N_21948,N_21837);
xor U22529 (N_22529,N_22291,N_21482);
nor U22530 (N_22530,N_21279,N_22078);
or U22531 (N_22531,N_21360,N_22125);
xor U22532 (N_22532,N_22229,N_21651);
nand U22533 (N_22533,N_21470,N_21903);
nor U22534 (N_22534,N_21560,N_21854);
nand U22535 (N_22535,N_21431,N_21629);
nor U22536 (N_22536,N_21785,N_22294);
nor U22537 (N_22537,N_21921,N_21869);
nor U22538 (N_22538,N_21579,N_22065);
and U22539 (N_22539,N_21359,N_21725);
nor U22540 (N_22540,N_21707,N_21602);
and U22541 (N_22541,N_21340,N_22069);
or U22542 (N_22542,N_22212,N_21628);
and U22543 (N_22543,N_22374,N_22442);
xor U22544 (N_22544,N_21584,N_22477);
nand U22545 (N_22545,N_21674,N_21899);
or U22546 (N_22546,N_21251,N_21976);
nor U22547 (N_22547,N_22369,N_21834);
nand U22548 (N_22548,N_22100,N_21475);
and U22549 (N_22549,N_22096,N_21874);
nor U22550 (N_22550,N_22062,N_21571);
xor U22551 (N_22551,N_21506,N_21365);
and U22552 (N_22552,N_21298,N_22265);
xnor U22553 (N_22553,N_21375,N_21495);
xnor U22554 (N_22554,N_21743,N_21929);
and U22555 (N_22555,N_22148,N_21855);
nand U22556 (N_22556,N_21413,N_22072);
nor U22557 (N_22557,N_21258,N_22173);
or U22558 (N_22558,N_21738,N_21801);
xnor U22559 (N_22559,N_22323,N_21965);
and U22560 (N_22560,N_21264,N_21873);
and U22561 (N_22561,N_22310,N_21310);
xor U22562 (N_22562,N_21535,N_22433);
or U22563 (N_22563,N_22419,N_21419);
nand U22564 (N_22564,N_21428,N_21452);
xor U22565 (N_22565,N_21887,N_21853);
xor U22566 (N_22566,N_21949,N_21820);
and U22567 (N_22567,N_21543,N_22301);
and U22568 (N_22568,N_21390,N_21980);
or U22569 (N_22569,N_21682,N_21631);
and U22570 (N_22570,N_21661,N_21770);
or U22571 (N_22571,N_22080,N_21957);
nor U22572 (N_22572,N_21252,N_21705);
and U22573 (N_22573,N_21577,N_22144);
nor U22574 (N_22574,N_22160,N_21617);
nand U22575 (N_22575,N_21777,N_21969);
xor U22576 (N_22576,N_21512,N_21805);
or U22577 (N_22577,N_21345,N_21447);
xor U22578 (N_22578,N_21771,N_21395);
and U22579 (N_22579,N_21255,N_21746);
xor U22580 (N_22580,N_22041,N_22040);
or U22581 (N_22581,N_22256,N_22016);
xnor U22582 (N_22582,N_21461,N_22459);
and U22583 (N_22583,N_22060,N_21534);
and U22584 (N_22584,N_22268,N_21963);
and U22585 (N_22585,N_21570,N_22275);
nor U22586 (N_22586,N_22380,N_22428);
and U22587 (N_22587,N_22085,N_21441);
nor U22588 (N_22588,N_21277,N_21305);
nor U22589 (N_22589,N_22124,N_22221);
nor U22590 (N_22590,N_22033,N_21759);
and U22591 (N_22591,N_21859,N_21706);
xor U22592 (N_22592,N_21518,N_21923);
or U22593 (N_22593,N_21293,N_22192);
and U22594 (N_22594,N_22446,N_22222);
and U22595 (N_22595,N_21527,N_21507);
xnor U22596 (N_22596,N_22028,N_21850);
and U22597 (N_22597,N_22172,N_21460);
xor U22598 (N_22598,N_21881,N_22465);
nand U22599 (N_22599,N_21696,N_21438);
or U22600 (N_22600,N_21505,N_21829);
xor U22601 (N_22601,N_21303,N_21807);
nor U22602 (N_22602,N_21615,N_22129);
xnor U22603 (N_22603,N_22279,N_22308);
or U22604 (N_22604,N_22063,N_21799);
or U22605 (N_22605,N_22366,N_22161);
xor U22606 (N_22606,N_21747,N_22481);
nor U22607 (N_22607,N_21319,N_21449);
and U22608 (N_22608,N_21804,N_22295);
xnor U22609 (N_22609,N_21741,N_22316);
xnor U22610 (N_22610,N_22167,N_21721);
nand U22611 (N_22611,N_21626,N_21422);
nand U22612 (N_22612,N_22373,N_21990);
xnor U22613 (N_22613,N_21585,N_21339);
or U22614 (N_22614,N_21781,N_21532);
nand U22615 (N_22615,N_22008,N_21557);
or U22616 (N_22616,N_22297,N_22088);
nor U22617 (N_22617,N_21894,N_21660);
nand U22618 (N_22618,N_21872,N_22480);
or U22619 (N_22619,N_21714,N_21717);
nand U22620 (N_22620,N_22147,N_21645);
nor U22621 (N_22621,N_21440,N_21830);
nand U22622 (N_22622,N_21583,N_22093);
nand U22623 (N_22623,N_21614,N_21627);
nor U22624 (N_22624,N_21407,N_22181);
nor U22625 (N_22625,N_22320,N_21884);
and U22626 (N_22626,N_21425,N_21409);
or U22627 (N_22627,N_21730,N_21367);
xor U22628 (N_22628,N_22292,N_22162);
or U22629 (N_22629,N_21593,N_21966);
xnor U22630 (N_22630,N_21374,N_22424);
xnor U22631 (N_22631,N_21704,N_22024);
nand U22632 (N_22632,N_22006,N_21347);
xor U22633 (N_22633,N_22461,N_22479);
or U22634 (N_22634,N_22344,N_22356);
nor U22635 (N_22635,N_21792,N_21918);
or U22636 (N_22636,N_22404,N_22204);
and U22637 (N_22637,N_21960,N_22146);
xor U22638 (N_22638,N_22498,N_21858);
and U22639 (N_22639,N_21666,N_22044);
nor U22640 (N_22640,N_21754,N_22496);
nand U22641 (N_22641,N_21474,N_21625);
nor U22642 (N_22642,N_21445,N_21938);
and U22643 (N_22643,N_22061,N_21573);
nand U22644 (N_22644,N_21384,N_21906);
nor U22645 (N_22645,N_21896,N_21700);
nand U22646 (N_22646,N_21928,N_22108);
and U22647 (N_22647,N_21810,N_21975);
xor U22648 (N_22648,N_21575,N_21784);
nand U22649 (N_22649,N_22383,N_21321);
nor U22650 (N_22650,N_21403,N_21471);
and U22651 (N_22651,N_22197,N_22255);
nor U22652 (N_22652,N_21304,N_22090);
nand U22653 (N_22653,N_21916,N_22311);
or U22654 (N_22654,N_22478,N_22187);
xor U22655 (N_22655,N_21988,N_22071);
nor U22656 (N_22656,N_21720,N_22246);
nand U22657 (N_22657,N_21517,N_22439);
nand U22658 (N_22658,N_22225,N_21699);
nor U22659 (N_22659,N_21697,N_21656);
or U22660 (N_22660,N_22059,N_22290);
xnor U22661 (N_22661,N_22249,N_22326);
and U22662 (N_22662,N_22052,N_21268);
nand U22663 (N_22663,N_22352,N_22113);
nand U22664 (N_22664,N_22303,N_21417);
and U22665 (N_22665,N_21346,N_22425);
or U22666 (N_22666,N_21795,N_21609);
and U22667 (N_22667,N_21406,N_21983);
nor U22668 (N_22668,N_22163,N_21544);
and U22669 (N_22669,N_22398,N_21967);
xnor U22670 (N_22670,N_21826,N_21767);
or U22671 (N_22671,N_21397,N_22174);
xor U22672 (N_22672,N_22149,N_21276);
or U22673 (N_22673,N_21954,N_21607);
and U22674 (N_22674,N_21864,N_22220);
and U22675 (N_22675,N_22170,N_21260);
nand U22676 (N_22676,N_21994,N_22407);
nor U22677 (N_22677,N_22165,N_22103);
xnor U22678 (N_22678,N_22324,N_21254);
nand U22679 (N_22679,N_21600,N_22436);
and U22680 (N_22680,N_21857,N_21357);
xnor U22681 (N_22681,N_21572,N_21788);
nand U22682 (N_22682,N_21786,N_21311);
nand U22683 (N_22683,N_22132,N_21524);
and U22684 (N_22684,N_21989,N_21592);
xnor U22685 (N_22685,N_21288,N_22367);
xnor U22686 (N_22686,N_21794,N_22241);
xnor U22687 (N_22687,N_21437,N_21984);
or U22688 (N_22688,N_22388,N_21726);
nand U22689 (N_22689,N_21300,N_22081);
xor U22690 (N_22690,N_22397,N_22011);
nor U22691 (N_22691,N_21344,N_21904);
xor U22692 (N_22692,N_21935,N_22046);
nand U22693 (N_22693,N_21639,N_21388);
nor U22694 (N_22694,N_21530,N_21578);
nand U22695 (N_22695,N_22200,N_22395);
nand U22696 (N_22696,N_21692,N_21401);
and U22697 (N_22697,N_22141,N_22066);
nor U22698 (N_22698,N_21362,N_21420);
nand U22699 (N_22699,N_21798,N_22348);
and U22700 (N_22700,N_22346,N_21329);
nand U22701 (N_22701,N_21987,N_21353);
xnor U22702 (N_22702,N_21456,N_22376);
xor U22703 (N_22703,N_22417,N_21971);
xor U22704 (N_22704,N_22128,N_21643);
xnor U22705 (N_22705,N_21942,N_21677);
and U22706 (N_22706,N_21836,N_21316);
xor U22707 (N_22707,N_21632,N_21919);
and U22708 (N_22708,N_22406,N_22032);
xnor U22709 (N_22709,N_21454,N_22372);
or U22710 (N_22710,N_22464,N_21882);
or U22711 (N_22711,N_22411,N_22472);
nand U22712 (N_22712,N_21977,N_22150);
nor U22713 (N_22713,N_21500,N_22420);
or U22714 (N_22714,N_22314,N_21650);
xnor U22715 (N_22715,N_21670,N_22219);
or U22716 (N_22716,N_21369,N_22159);
or U22717 (N_22717,N_21749,N_21542);
and U22718 (N_22718,N_21430,N_22284);
nor U22719 (N_22719,N_22133,N_21755);
xor U22720 (N_22720,N_21930,N_21587);
nor U22721 (N_22721,N_22138,N_21299);
and U22722 (N_22722,N_21986,N_21734);
xnor U22723 (N_22723,N_21306,N_21267);
or U22724 (N_22724,N_21493,N_21462);
nor U22725 (N_22725,N_21657,N_21368);
nand U22726 (N_22726,N_21478,N_22083);
nor U22727 (N_22727,N_21548,N_22179);
or U22728 (N_22728,N_21563,N_22231);
xnor U22729 (N_22729,N_21667,N_21604);
and U22730 (N_22730,N_21519,N_21338);
or U22731 (N_22731,N_21846,N_21839);
nand U22732 (N_22732,N_21812,N_21658);
nand U22733 (N_22733,N_21335,N_22338);
nand U22734 (N_22734,N_21780,N_22243);
xor U22735 (N_22735,N_22019,N_22396);
and U22736 (N_22736,N_21392,N_21433);
or U22737 (N_22737,N_22370,N_21317);
nand U22738 (N_22738,N_21774,N_22131);
nor U22739 (N_22739,N_22115,N_22387);
nand U22740 (N_22740,N_22037,N_21791);
nand U22741 (N_22741,N_21416,N_22274);
and U22742 (N_22742,N_21742,N_21652);
xnor U22743 (N_22743,N_21671,N_22022);
and U22744 (N_22744,N_21708,N_21415);
nand U22745 (N_22745,N_21642,N_21382);
xnor U22746 (N_22746,N_21800,N_21504);
nor U22747 (N_22747,N_21315,N_21497);
xor U22748 (N_22748,N_21995,N_21946);
nand U22749 (N_22749,N_21985,N_22110);
and U22750 (N_22750,N_22023,N_22136);
or U22751 (N_22751,N_22363,N_21509);
nand U22752 (N_22752,N_21937,N_22408);
and U22753 (N_22753,N_22017,N_21793);
nand U22754 (N_22754,N_21411,N_21432);
nand U22755 (N_22755,N_22015,N_22042);
and U22756 (N_22756,N_22191,N_22299);
and U22757 (N_22757,N_22273,N_21510);
xnor U22758 (N_22758,N_21485,N_21398);
nor U22759 (N_22759,N_22127,N_21453);
nor U22760 (N_22760,N_21728,N_22242);
nand U22761 (N_22761,N_21528,N_21418);
nor U22762 (N_22762,N_22313,N_22064);
nor U22763 (N_22763,N_21503,N_22168);
and U22764 (N_22764,N_21426,N_21622);
and U22765 (N_22765,N_22267,N_22206);
nand U22766 (N_22766,N_22432,N_21867);
nor U22767 (N_22767,N_22491,N_21851);
and U22768 (N_22768,N_21443,N_21897);
or U22769 (N_22769,N_22359,N_21483);
and U22770 (N_22770,N_22051,N_21997);
nand U22771 (N_22771,N_22050,N_21769);
nor U22772 (N_22772,N_21342,N_21908);
nand U22773 (N_22773,N_22067,N_22247);
nand U22774 (N_22774,N_21763,N_21623);
and U22775 (N_22775,N_22322,N_21324);
and U22776 (N_22776,N_21647,N_22087);
xor U22777 (N_22777,N_21779,N_21446);
nor U22778 (N_22778,N_21514,N_21688);
and U22779 (N_22779,N_22045,N_21386);
or U22780 (N_22780,N_21408,N_21941);
xnor U22781 (N_22781,N_21323,N_21606);
xnor U22782 (N_22782,N_21297,N_22345);
nor U22783 (N_22783,N_22000,N_22486);
nand U22784 (N_22784,N_21996,N_21400);
or U22785 (N_22785,N_22405,N_21326);
nand U22786 (N_22786,N_21821,N_22106);
xor U22787 (N_22787,N_22300,N_21380);
and U22788 (N_22788,N_22351,N_22448);
nor U22789 (N_22789,N_22287,N_21654);
xnor U22790 (N_22790,N_21924,N_22029);
nor U22791 (N_22791,N_21545,N_21523);
or U22792 (N_22792,N_21366,N_21940);
and U22793 (N_22793,N_21263,N_22403);
nor U22794 (N_22794,N_21845,N_22460);
xor U22795 (N_22795,N_21283,N_22030);
nand U22796 (N_22796,N_22250,N_22457);
xnor U22797 (N_22797,N_22007,N_21405);
and U22798 (N_22798,N_22305,N_21442);
nand U22799 (N_22799,N_21605,N_22018);
nor U22800 (N_22800,N_21838,N_22289);
and U22801 (N_22801,N_21958,N_22259);
nand U22802 (N_22802,N_21723,N_21611);
xor U22803 (N_22803,N_22332,N_22009);
nor U22804 (N_22804,N_22116,N_21256);
xnor U22805 (N_22805,N_21668,N_21665);
or U22806 (N_22806,N_22330,N_21491);
or U22807 (N_22807,N_21358,N_21731);
nor U22808 (N_22808,N_22122,N_21973);
or U22809 (N_22809,N_22254,N_21393);
xnor U22810 (N_22810,N_21396,N_21271);
xor U22811 (N_22811,N_22449,N_21648);
and U22812 (N_22812,N_22013,N_21385);
or U22813 (N_22813,N_22329,N_21831);
nand U22814 (N_22814,N_21819,N_22183);
nor U22815 (N_22815,N_21886,N_21888);
and U22816 (N_22816,N_21693,N_21895);
nand U22817 (N_22817,N_22264,N_21939);
nand U22818 (N_22818,N_21953,N_21722);
or U22819 (N_22819,N_21712,N_22005);
and U22820 (N_22820,N_22270,N_22353);
and U22821 (N_22821,N_21710,N_22010);
xor U22822 (N_22822,N_21451,N_21270);
nor U22823 (N_22823,N_22261,N_22123);
nand U22824 (N_22824,N_21439,N_21612);
or U22825 (N_22825,N_21312,N_22214);
and U22826 (N_22826,N_21580,N_21285);
and U22827 (N_22827,N_21318,N_22328);
and U22828 (N_22828,N_21709,N_21489);
or U22829 (N_22829,N_21686,N_21687);
nand U22830 (N_22830,N_21814,N_22390);
nand U22831 (N_22831,N_21331,N_21259);
or U22832 (N_22832,N_22452,N_21508);
or U22833 (N_22833,N_22077,N_21282);
nand U22834 (N_22834,N_21594,N_22362);
xor U22835 (N_22835,N_21348,N_22269);
xnor U22836 (N_22836,N_22271,N_21624);
and U22837 (N_22837,N_21554,N_21364);
nor U22838 (N_22838,N_21295,N_21822);
and U22839 (N_22839,N_22166,N_21477);
or U22840 (N_22840,N_21640,N_22263);
xor U22841 (N_22841,N_22153,N_21841);
or U22842 (N_22842,N_21434,N_22215);
nor U22843 (N_22843,N_21840,N_21765);
nor U22844 (N_22844,N_22152,N_22276);
nor U22845 (N_22845,N_22319,N_22175);
nor U22846 (N_22846,N_21343,N_21681);
nor U22847 (N_22847,N_22379,N_22234);
nand U22848 (N_22848,N_22119,N_22176);
and U22849 (N_22849,N_21595,N_21421);
nor U22850 (N_22850,N_22483,N_22120);
nand U22851 (N_22851,N_21552,N_22440);
nand U22852 (N_22852,N_21291,N_22143);
or U22853 (N_22853,N_22347,N_22213);
nor U22854 (N_22854,N_22094,N_22495);
or U22855 (N_22855,N_21292,N_21811);
and U22856 (N_22856,N_21531,N_22341);
xnor U22857 (N_22857,N_21956,N_22137);
nand U22858 (N_22858,N_22182,N_22098);
xor U22859 (N_22859,N_21757,N_21603);
nand U22860 (N_22860,N_21328,N_22429);
and U22861 (N_22861,N_22236,N_21702);
or U22862 (N_22862,N_21599,N_21735);
nand U22863 (N_22863,N_22145,N_22184);
or U22864 (N_22864,N_21378,N_21823);
xnor U22865 (N_22865,N_22021,N_21372);
nand U22866 (N_22866,N_21391,N_21745);
and U22867 (N_22867,N_22169,N_21574);
xor U22868 (N_22868,N_21275,N_22157);
nor U22869 (N_22869,N_22058,N_22199);
or U22870 (N_22870,N_21974,N_21308);
nor U22871 (N_22871,N_21736,N_22389);
or U22872 (N_22872,N_21465,N_21852);
xor U22873 (N_22873,N_22431,N_21562);
nand U22874 (N_22874,N_21525,N_22434);
or U22875 (N_22875,N_22245,N_21835);
and U22876 (N_22876,N_21925,N_21515);
xor U22877 (N_22877,N_21790,N_22055);
or U22878 (N_22878,N_21649,N_21978);
nand U22879 (N_22879,N_21302,N_21842);
and U22880 (N_22880,N_22112,N_21636);
nand U22881 (N_22881,N_22109,N_21737);
and U22882 (N_22882,N_21663,N_21951);
nor U22883 (N_22883,N_22031,N_22227);
and U22884 (N_22884,N_21968,N_22224);
nor U22885 (N_22885,N_21484,N_22076);
nor U22886 (N_22886,N_21909,N_22410);
and U22887 (N_22887,N_22277,N_21991);
or U22888 (N_22888,N_22386,N_22223);
xnor U22889 (N_22889,N_21476,N_21890);
xnor U22890 (N_22890,N_21466,N_22283);
xnor U22891 (N_22891,N_22208,N_21892);
or U22892 (N_22892,N_21361,N_22490);
xor U22893 (N_22893,N_21250,N_22360);
and U22894 (N_22894,N_21756,N_21553);
or U22895 (N_22895,N_22118,N_21589);
nor U22896 (N_22896,N_22412,N_21729);
nor U22897 (N_22897,N_21379,N_21901);
or U22898 (N_22898,N_21499,N_22296);
or U22899 (N_22899,N_21676,N_22272);
or U22900 (N_22900,N_21926,N_22444);
and U22901 (N_22901,N_21349,N_21286);
xnor U22902 (N_22902,N_21262,N_22203);
and U22903 (N_22903,N_22468,N_21539);
nor U22904 (N_22904,N_22201,N_22469);
nand U22905 (N_22905,N_22447,N_21773);
nor U22906 (N_22906,N_21257,N_22474);
nand U22907 (N_22907,N_21455,N_22102);
nand U22908 (N_22908,N_22415,N_21337);
nand U22909 (N_22909,N_22317,N_21824);
xor U22910 (N_22910,N_22185,N_21536);
nor U22911 (N_22911,N_21982,N_21435);
or U22912 (N_22912,N_22154,N_21473);
or U22913 (N_22913,N_22092,N_21776);
and U22914 (N_22914,N_21289,N_22075);
nor U22915 (N_22915,N_21907,N_22193);
or U22916 (N_22916,N_21885,N_21943);
or U22917 (N_22917,N_22318,N_21815);
nor U22918 (N_22918,N_22228,N_22099);
and U22919 (N_22919,N_21744,N_22401);
nor U22920 (N_22920,N_21817,N_21389);
or U22921 (N_22921,N_22047,N_21694);
nand U22922 (N_22922,N_22416,N_22057);
xor U22923 (N_22923,N_22377,N_21635);
and U22924 (N_22924,N_21818,N_21399);
xor U22925 (N_22925,N_21444,N_22111);
nor U22926 (N_22926,N_21915,N_21457);
nand U22927 (N_22927,N_22455,N_22335);
and U22928 (N_22928,N_22325,N_22014);
xnor U22929 (N_22929,N_21301,N_21775);
nand U22930 (N_22930,N_21540,N_22070);
xor U22931 (N_22931,N_22336,N_22209);
or U22932 (N_22932,N_21568,N_22230);
or U22933 (N_22933,N_21423,N_22140);
or U22934 (N_22934,N_21480,N_21541);
or U22935 (N_22935,N_22155,N_22393);
or U22936 (N_22936,N_21732,N_21352);
or U22937 (N_22937,N_22251,N_22487);
nor U22938 (N_22938,N_21555,N_21613);
nand U22939 (N_22939,N_22437,N_21998);
and U22940 (N_22940,N_21796,N_21927);
nand U22941 (N_22941,N_22012,N_21549);
and U22942 (N_22942,N_21876,N_22257);
xor U22943 (N_22943,N_21511,N_22034);
nand U22944 (N_22944,N_21487,N_22171);
or U22945 (N_22945,N_22027,N_22384);
or U22946 (N_22946,N_22089,N_21608);
and U22947 (N_22947,N_22282,N_21336);
or U22948 (N_22948,N_22422,N_21586);
and U22949 (N_22949,N_21327,N_21313);
and U22950 (N_22950,N_22216,N_22492);
or U22951 (N_22951,N_21354,N_21813);
nor U22952 (N_22952,N_21659,N_22233);
nor U22953 (N_22953,N_21685,N_22402);
nand U22954 (N_22954,N_22499,N_21959);
or U22955 (N_22955,N_22409,N_22244);
nand U22956 (N_22956,N_22126,N_22020);
and U22957 (N_22957,N_21768,N_22309);
xor U22958 (N_22958,N_21934,N_21646);
or U22959 (N_22959,N_21695,N_21806);
xor U22960 (N_22960,N_21972,N_22476);
or U22961 (N_22961,N_21521,N_22235);
nor U22962 (N_22962,N_22331,N_22095);
xor U22963 (N_22963,N_22107,N_21877);
or U22964 (N_22964,N_22488,N_21905);
and U22965 (N_22965,N_22026,N_22497);
and U22966 (N_22966,N_21641,N_21290);
and U22967 (N_22967,N_22454,N_21891);
nand U22968 (N_22968,N_22189,N_21424);
xnor U22969 (N_22969,N_22278,N_22086);
and U22970 (N_22970,N_21498,N_22049);
xnor U22971 (N_22971,N_21762,N_22156);
nand U22972 (N_22972,N_21581,N_22188);
xnor U22973 (N_22973,N_22082,N_21701);
nor U22974 (N_22974,N_22262,N_21481);
and U22975 (N_22975,N_22482,N_22039);
nand U22976 (N_22976,N_22371,N_21868);
and U22977 (N_22977,N_21448,N_21932);
or U22978 (N_22978,N_21350,N_21740);
xnor U22979 (N_22979,N_22288,N_21488);
and U22980 (N_22980,N_21760,N_22470);
nor U22981 (N_22981,N_22135,N_21621);
or U22982 (N_22982,N_21588,N_21559);
nand U22983 (N_22983,N_21856,N_21591);
nand U22984 (N_22984,N_22427,N_22456);
nor U22985 (N_22985,N_21669,N_21567);
nand U22986 (N_22986,N_22053,N_21653);
nand U22987 (N_22987,N_22035,N_22217);
and U22988 (N_22988,N_21383,N_21278);
or U22989 (N_22989,N_22164,N_21450);
nor U22990 (N_22990,N_22068,N_22056);
nor U22991 (N_22991,N_22304,N_21576);
xor U22992 (N_22992,N_22493,N_21330);
xor U22993 (N_22993,N_21314,N_21828);
nor U22994 (N_22994,N_22378,N_22025);
nand U22995 (N_22995,N_21753,N_22177);
xnor U22996 (N_22996,N_22400,N_22312);
xnor U22997 (N_22997,N_22002,N_21590);
and U22998 (N_22998,N_22450,N_22186);
and U22999 (N_22999,N_22361,N_21803);
nor U23000 (N_23000,N_22121,N_22463);
and U23001 (N_23001,N_22458,N_21878);
nor U23002 (N_23002,N_21797,N_22001);
nor U23003 (N_23003,N_21351,N_21961);
nand U23004 (N_23004,N_21274,N_21501);
and U23005 (N_23005,N_21325,N_21843);
nor U23006 (N_23006,N_21718,N_22358);
nor U23007 (N_23007,N_21860,N_21955);
and U23008 (N_23008,N_21866,N_21281);
and U23009 (N_23009,N_21463,N_22302);
nor U23010 (N_23010,N_22130,N_21296);
xor U23011 (N_23011,N_22343,N_22158);
and U23012 (N_23012,N_21844,N_21848);
nor U23013 (N_23013,N_21703,N_21751);
nand U23014 (N_23014,N_22391,N_21922);
xnor U23015 (N_23015,N_22421,N_21307);
xor U23016 (N_23016,N_21533,N_21716);
and U23017 (N_23017,N_21944,N_22043);
and U23018 (N_23018,N_21468,N_21715);
nand U23019 (N_23019,N_21287,N_22489);
xor U23020 (N_23020,N_21556,N_22307);
xnor U23021 (N_23021,N_21561,N_21802);
nor U23022 (N_23022,N_21889,N_21458);
nor U23023 (N_23023,N_22333,N_22473);
nand U23024 (N_23024,N_21565,N_21752);
or U23025 (N_23025,N_21516,N_21479);
and U23026 (N_23026,N_22365,N_21638);
or U23027 (N_23027,N_21616,N_21816);
xnor U23028 (N_23028,N_21284,N_21634);
or U23029 (N_23029,N_22238,N_21377);
and U23030 (N_23030,N_22117,N_22281);
and U23031 (N_23031,N_21861,N_22190);
nand U23032 (N_23032,N_21673,N_21783);
and U23033 (N_23033,N_21748,N_21334);
xnor U23034 (N_23034,N_22237,N_22441);
or U23035 (N_23035,N_21950,N_22354);
and U23036 (N_23036,N_22382,N_22298);
and U23037 (N_23037,N_21464,N_22423);
or U23038 (N_23038,N_21410,N_21981);
xor U23039 (N_23039,N_22467,N_22430);
nand U23040 (N_23040,N_22466,N_21486);
nand U23041 (N_23041,N_22438,N_22260);
nand U23042 (N_23042,N_21322,N_22342);
nor U23043 (N_23043,N_21566,N_21979);
and U23044 (N_23044,N_22114,N_21914);
nor U23045 (N_23045,N_22306,N_21713);
nand U23046 (N_23046,N_21569,N_22202);
or U23047 (N_23047,N_21332,N_22205);
nor U23048 (N_23048,N_22239,N_22485);
nor U23049 (N_23049,N_21761,N_21644);
nor U23050 (N_23050,N_21490,N_21766);
nor U23051 (N_23051,N_22375,N_22079);
xnor U23052 (N_23052,N_22426,N_21679);
xor U23053 (N_23053,N_21862,N_21373);
and U23054 (N_23054,N_22471,N_21496);
nor U23055 (N_23055,N_21684,N_21999);
nand U23056 (N_23056,N_21381,N_21402);
xor U23057 (N_23057,N_21778,N_22385);
nor U23058 (N_23058,N_21253,N_21750);
nand U23059 (N_23059,N_22293,N_21739);
xor U23060 (N_23060,N_21733,N_21630);
xor U23061 (N_23061,N_21492,N_21513);
and U23062 (N_23062,N_21610,N_21825);
nor U23063 (N_23063,N_21356,N_21893);
nor U23064 (N_23064,N_21789,N_22445);
nor U23065 (N_23065,N_21265,N_21764);
and U23066 (N_23066,N_21564,N_22003);
xnor U23067 (N_23067,N_22104,N_21370);
xnor U23068 (N_23068,N_22334,N_21675);
nand U23069 (N_23069,N_22285,N_21376);
nand U23070 (N_23070,N_21865,N_21363);
or U23071 (N_23071,N_21269,N_21601);
and U23072 (N_23072,N_21546,N_21920);
nor U23073 (N_23073,N_21772,N_21962);
nand U23074 (N_23074,N_21309,N_21522);
and U23075 (N_23075,N_21964,N_21871);
nor U23076 (N_23076,N_22194,N_21724);
xor U23077 (N_23077,N_21537,N_22494);
nor U23078 (N_23078,N_22252,N_22286);
and U23079 (N_23079,N_22105,N_21947);
xor U23080 (N_23080,N_21931,N_21883);
xnor U23081 (N_23081,N_22226,N_21619);
xnor U23082 (N_23082,N_21933,N_21711);
and U23083 (N_23083,N_22340,N_21911);
and U23084 (N_23084,N_22418,N_21898);
xnor U23085 (N_23085,N_21412,N_21266);
nor U23086 (N_23086,N_22327,N_21698);
and U23087 (N_23087,N_22381,N_22074);
xor U23088 (N_23088,N_21394,N_22101);
nor U23089 (N_23089,N_22357,N_21952);
xnor U23090 (N_23090,N_21689,N_22349);
nand U23091 (N_23091,N_21320,N_22435);
and U23092 (N_23092,N_22091,N_22280);
xnor U23093 (N_23093,N_21387,N_22451);
nor U23094 (N_23094,N_21782,N_21620);
nand U23095 (N_23095,N_21672,N_21261);
nand U23096 (N_23096,N_21618,N_22453);
and U23097 (N_23097,N_21913,N_22368);
and U23098 (N_23098,N_21847,N_21371);
xnor U23099 (N_23099,N_21992,N_21655);
nand U23100 (N_23100,N_21917,N_21719);
or U23101 (N_23101,N_21910,N_21355);
nand U23102 (N_23102,N_22484,N_21664);
or U23103 (N_23103,N_21863,N_22180);
nand U23104 (N_23104,N_22253,N_21809);
xnor U23105 (N_23105,N_22097,N_21597);
nor U23106 (N_23106,N_21690,N_22038);
nand U23107 (N_23107,N_22339,N_22266);
xor U23108 (N_23108,N_22196,N_22198);
nor U23109 (N_23109,N_21494,N_22073);
and U23110 (N_23110,N_21273,N_22364);
or U23111 (N_23111,N_22151,N_21502);
and U23112 (N_23112,N_22443,N_22399);
and U23113 (N_23113,N_21993,N_21272);
or U23114 (N_23114,N_21902,N_22414);
nor U23115 (N_23115,N_21691,N_22218);
or U23116 (N_23116,N_22048,N_22240);
or U23117 (N_23117,N_21808,N_22210);
or U23118 (N_23118,N_21727,N_22355);
nand U23119 (N_23119,N_21550,N_21551);
and U23120 (N_23120,N_21879,N_22054);
or U23121 (N_23121,N_21333,N_21429);
and U23122 (N_23122,N_21970,N_21849);
or U23123 (N_23123,N_22413,N_22350);
nand U23124 (N_23124,N_21832,N_21538);
or U23125 (N_23125,N_22474,N_21636);
and U23126 (N_23126,N_21917,N_21318);
nor U23127 (N_23127,N_22273,N_21442);
nor U23128 (N_23128,N_21264,N_22325);
xnor U23129 (N_23129,N_21736,N_21378);
nor U23130 (N_23130,N_21265,N_21650);
or U23131 (N_23131,N_22358,N_21529);
nor U23132 (N_23132,N_21939,N_21655);
nor U23133 (N_23133,N_22433,N_22415);
xor U23134 (N_23134,N_22400,N_22022);
and U23135 (N_23135,N_22086,N_21893);
nor U23136 (N_23136,N_21256,N_21384);
and U23137 (N_23137,N_21265,N_22006);
xor U23138 (N_23138,N_21744,N_21342);
nand U23139 (N_23139,N_22143,N_22464);
xor U23140 (N_23140,N_21458,N_22082);
nand U23141 (N_23141,N_22242,N_21759);
nand U23142 (N_23142,N_21874,N_21347);
and U23143 (N_23143,N_21910,N_21547);
xnor U23144 (N_23144,N_22119,N_21633);
and U23145 (N_23145,N_21939,N_21862);
nor U23146 (N_23146,N_21345,N_22358);
nor U23147 (N_23147,N_22421,N_22482);
nand U23148 (N_23148,N_22273,N_21942);
or U23149 (N_23149,N_21644,N_21846);
and U23150 (N_23150,N_22036,N_21277);
and U23151 (N_23151,N_21852,N_21416);
or U23152 (N_23152,N_21268,N_21598);
and U23153 (N_23153,N_21544,N_22469);
xnor U23154 (N_23154,N_22220,N_21461);
and U23155 (N_23155,N_21588,N_21857);
xor U23156 (N_23156,N_22294,N_22424);
nand U23157 (N_23157,N_22073,N_22052);
nand U23158 (N_23158,N_21462,N_21647);
or U23159 (N_23159,N_22394,N_22347);
xor U23160 (N_23160,N_21320,N_22443);
nand U23161 (N_23161,N_22436,N_22143);
nand U23162 (N_23162,N_22370,N_21853);
or U23163 (N_23163,N_22271,N_21868);
and U23164 (N_23164,N_22134,N_22199);
or U23165 (N_23165,N_21407,N_22257);
xnor U23166 (N_23166,N_21432,N_22182);
xnor U23167 (N_23167,N_21416,N_21600);
nor U23168 (N_23168,N_21455,N_21458);
nand U23169 (N_23169,N_21308,N_22174);
or U23170 (N_23170,N_22446,N_21969);
nand U23171 (N_23171,N_21639,N_22293);
or U23172 (N_23172,N_21575,N_21735);
and U23173 (N_23173,N_21926,N_21516);
nand U23174 (N_23174,N_22249,N_22037);
nand U23175 (N_23175,N_21867,N_21918);
xor U23176 (N_23176,N_22360,N_21883);
xor U23177 (N_23177,N_21559,N_21855);
xnor U23178 (N_23178,N_22361,N_21920);
xnor U23179 (N_23179,N_22398,N_21433);
nor U23180 (N_23180,N_21865,N_21711);
nor U23181 (N_23181,N_22422,N_22030);
xor U23182 (N_23182,N_21888,N_21395);
xor U23183 (N_23183,N_21680,N_21369);
and U23184 (N_23184,N_21881,N_22217);
or U23185 (N_23185,N_21488,N_21896);
or U23186 (N_23186,N_21524,N_21745);
nor U23187 (N_23187,N_21394,N_21529);
nand U23188 (N_23188,N_22016,N_21779);
nor U23189 (N_23189,N_22224,N_22219);
nor U23190 (N_23190,N_21565,N_21992);
nor U23191 (N_23191,N_22479,N_21928);
or U23192 (N_23192,N_21628,N_22170);
xnor U23193 (N_23193,N_21444,N_21493);
nor U23194 (N_23194,N_21273,N_21546);
xor U23195 (N_23195,N_22415,N_21913);
nor U23196 (N_23196,N_22490,N_22387);
or U23197 (N_23197,N_22349,N_21784);
nand U23198 (N_23198,N_22318,N_22327);
nand U23199 (N_23199,N_22233,N_22180);
and U23200 (N_23200,N_21268,N_21926);
and U23201 (N_23201,N_22329,N_21662);
nor U23202 (N_23202,N_21356,N_21820);
nand U23203 (N_23203,N_22142,N_22269);
or U23204 (N_23204,N_21339,N_21462);
or U23205 (N_23205,N_22165,N_22156);
and U23206 (N_23206,N_21817,N_22446);
nand U23207 (N_23207,N_22047,N_21441);
xor U23208 (N_23208,N_21491,N_22190);
nor U23209 (N_23209,N_21536,N_22422);
or U23210 (N_23210,N_21774,N_21647);
or U23211 (N_23211,N_21441,N_21684);
and U23212 (N_23212,N_22316,N_21941);
and U23213 (N_23213,N_21355,N_21732);
nand U23214 (N_23214,N_21266,N_21964);
xor U23215 (N_23215,N_21855,N_21658);
or U23216 (N_23216,N_21825,N_21576);
or U23217 (N_23217,N_21800,N_21587);
and U23218 (N_23218,N_21938,N_21541);
nor U23219 (N_23219,N_22221,N_22052);
xnor U23220 (N_23220,N_21885,N_21607);
or U23221 (N_23221,N_21316,N_22385);
nand U23222 (N_23222,N_22407,N_21286);
nor U23223 (N_23223,N_21474,N_21866);
or U23224 (N_23224,N_22187,N_22412);
and U23225 (N_23225,N_22013,N_21398);
and U23226 (N_23226,N_21350,N_21704);
and U23227 (N_23227,N_22012,N_22169);
or U23228 (N_23228,N_22135,N_21682);
and U23229 (N_23229,N_22468,N_22320);
nor U23230 (N_23230,N_21639,N_22230);
nor U23231 (N_23231,N_22426,N_21458);
nor U23232 (N_23232,N_22105,N_21540);
nand U23233 (N_23233,N_21983,N_21703);
xor U23234 (N_23234,N_22226,N_22410);
or U23235 (N_23235,N_22473,N_22007);
xnor U23236 (N_23236,N_21693,N_21879);
and U23237 (N_23237,N_22214,N_21841);
and U23238 (N_23238,N_21467,N_21945);
xor U23239 (N_23239,N_22313,N_22211);
and U23240 (N_23240,N_21850,N_21290);
nand U23241 (N_23241,N_21314,N_21498);
or U23242 (N_23242,N_21773,N_21524);
nand U23243 (N_23243,N_22169,N_22216);
nand U23244 (N_23244,N_21616,N_22393);
nand U23245 (N_23245,N_21308,N_21464);
or U23246 (N_23246,N_21900,N_22130);
nor U23247 (N_23247,N_22426,N_21335);
and U23248 (N_23248,N_22482,N_21553);
nor U23249 (N_23249,N_21293,N_21312);
or U23250 (N_23250,N_22172,N_21366);
nor U23251 (N_23251,N_21650,N_21480);
nor U23252 (N_23252,N_21659,N_22228);
nand U23253 (N_23253,N_21879,N_22379);
nand U23254 (N_23254,N_21611,N_21612);
nor U23255 (N_23255,N_21822,N_22179);
nand U23256 (N_23256,N_21303,N_21817);
or U23257 (N_23257,N_21585,N_22312);
nor U23258 (N_23258,N_21327,N_21886);
xnor U23259 (N_23259,N_22439,N_21679);
nor U23260 (N_23260,N_21739,N_22017);
xnor U23261 (N_23261,N_21652,N_21293);
or U23262 (N_23262,N_21430,N_22175);
and U23263 (N_23263,N_21990,N_22070);
or U23264 (N_23264,N_22450,N_21858);
and U23265 (N_23265,N_22367,N_22469);
nor U23266 (N_23266,N_21608,N_22220);
and U23267 (N_23267,N_21416,N_21949);
or U23268 (N_23268,N_21436,N_21283);
nor U23269 (N_23269,N_21968,N_21609);
nand U23270 (N_23270,N_22401,N_21874);
and U23271 (N_23271,N_21476,N_21816);
nor U23272 (N_23272,N_22134,N_21459);
nand U23273 (N_23273,N_22295,N_21953);
and U23274 (N_23274,N_21714,N_22160);
and U23275 (N_23275,N_21415,N_21743);
xor U23276 (N_23276,N_21327,N_21967);
or U23277 (N_23277,N_22144,N_21920);
nor U23278 (N_23278,N_22245,N_21700);
nand U23279 (N_23279,N_21443,N_21637);
or U23280 (N_23280,N_21343,N_21830);
xnor U23281 (N_23281,N_22359,N_21931);
nor U23282 (N_23282,N_22393,N_22314);
and U23283 (N_23283,N_22337,N_21615);
xnor U23284 (N_23284,N_21558,N_21598);
xnor U23285 (N_23285,N_21542,N_22371);
nor U23286 (N_23286,N_21780,N_21543);
nor U23287 (N_23287,N_22304,N_21381);
nand U23288 (N_23288,N_22450,N_22305);
xor U23289 (N_23289,N_22338,N_22109);
nor U23290 (N_23290,N_22465,N_21347);
xor U23291 (N_23291,N_21260,N_22191);
nor U23292 (N_23292,N_21856,N_21717);
and U23293 (N_23293,N_21298,N_22389);
nand U23294 (N_23294,N_21735,N_21573);
and U23295 (N_23295,N_21800,N_22028);
or U23296 (N_23296,N_22227,N_22080);
xor U23297 (N_23297,N_22431,N_22457);
nor U23298 (N_23298,N_22480,N_21902);
xnor U23299 (N_23299,N_21689,N_21501);
nor U23300 (N_23300,N_21907,N_22446);
and U23301 (N_23301,N_22496,N_21404);
and U23302 (N_23302,N_21366,N_21590);
nor U23303 (N_23303,N_21916,N_22197);
and U23304 (N_23304,N_22479,N_22048);
nor U23305 (N_23305,N_22436,N_21511);
xnor U23306 (N_23306,N_22211,N_22251);
and U23307 (N_23307,N_22052,N_21805);
nor U23308 (N_23308,N_22085,N_21733);
nor U23309 (N_23309,N_21825,N_21531);
and U23310 (N_23310,N_21445,N_21907);
or U23311 (N_23311,N_22129,N_22137);
nor U23312 (N_23312,N_21391,N_22094);
or U23313 (N_23313,N_21937,N_21320);
nor U23314 (N_23314,N_21437,N_21622);
nor U23315 (N_23315,N_21626,N_21799);
nor U23316 (N_23316,N_22013,N_21809);
xor U23317 (N_23317,N_22450,N_21722);
and U23318 (N_23318,N_21644,N_21290);
and U23319 (N_23319,N_21279,N_21426);
xnor U23320 (N_23320,N_21750,N_21354);
xor U23321 (N_23321,N_22400,N_21977);
nor U23322 (N_23322,N_22169,N_22337);
nor U23323 (N_23323,N_22163,N_21687);
xnor U23324 (N_23324,N_21442,N_21901);
nand U23325 (N_23325,N_21258,N_21927);
or U23326 (N_23326,N_22154,N_21692);
or U23327 (N_23327,N_21332,N_22321);
and U23328 (N_23328,N_21631,N_21870);
xnor U23329 (N_23329,N_22311,N_22180);
or U23330 (N_23330,N_21508,N_21280);
and U23331 (N_23331,N_21475,N_21272);
nor U23332 (N_23332,N_21980,N_22034);
nand U23333 (N_23333,N_22250,N_21592);
xor U23334 (N_23334,N_21488,N_22077);
and U23335 (N_23335,N_22008,N_21587);
xnor U23336 (N_23336,N_21758,N_22273);
nand U23337 (N_23337,N_21307,N_22459);
or U23338 (N_23338,N_21495,N_22411);
xor U23339 (N_23339,N_22097,N_22204);
nor U23340 (N_23340,N_22080,N_21968);
or U23341 (N_23341,N_21374,N_21586);
nor U23342 (N_23342,N_21570,N_21758);
or U23343 (N_23343,N_21493,N_22311);
xor U23344 (N_23344,N_21765,N_21357);
or U23345 (N_23345,N_22257,N_21355);
nand U23346 (N_23346,N_21701,N_21908);
nor U23347 (N_23347,N_21902,N_21447);
nor U23348 (N_23348,N_21361,N_22171);
and U23349 (N_23349,N_22467,N_21555);
nand U23350 (N_23350,N_21904,N_22105);
nand U23351 (N_23351,N_21650,N_21854);
nor U23352 (N_23352,N_21562,N_22419);
or U23353 (N_23353,N_22400,N_21611);
nand U23354 (N_23354,N_22200,N_22088);
nand U23355 (N_23355,N_22298,N_22123);
xnor U23356 (N_23356,N_22429,N_21282);
or U23357 (N_23357,N_21613,N_22304);
xnor U23358 (N_23358,N_22395,N_21948);
nor U23359 (N_23359,N_22339,N_22096);
or U23360 (N_23360,N_22115,N_22239);
and U23361 (N_23361,N_22374,N_22175);
and U23362 (N_23362,N_22445,N_22095);
or U23363 (N_23363,N_21584,N_21939);
xnor U23364 (N_23364,N_21417,N_21910);
and U23365 (N_23365,N_21581,N_21943);
nand U23366 (N_23366,N_21904,N_21723);
or U23367 (N_23367,N_21805,N_21839);
or U23368 (N_23368,N_22325,N_21886);
or U23369 (N_23369,N_22152,N_22222);
or U23370 (N_23370,N_21948,N_22422);
nand U23371 (N_23371,N_21752,N_21678);
nor U23372 (N_23372,N_21277,N_22238);
and U23373 (N_23373,N_22172,N_21386);
nor U23374 (N_23374,N_21687,N_21495);
or U23375 (N_23375,N_21809,N_22141);
nand U23376 (N_23376,N_22151,N_21426);
nand U23377 (N_23377,N_21855,N_21702);
xnor U23378 (N_23378,N_21713,N_22004);
or U23379 (N_23379,N_22463,N_21739);
or U23380 (N_23380,N_21899,N_21678);
xnor U23381 (N_23381,N_22093,N_21483);
or U23382 (N_23382,N_22257,N_22197);
or U23383 (N_23383,N_22150,N_22260);
and U23384 (N_23384,N_21663,N_21546);
xnor U23385 (N_23385,N_22281,N_22448);
and U23386 (N_23386,N_21572,N_22430);
and U23387 (N_23387,N_22065,N_21636);
nand U23388 (N_23388,N_21741,N_21801);
nor U23389 (N_23389,N_21745,N_21853);
nor U23390 (N_23390,N_21697,N_21281);
nand U23391 (N_23391,N_22426,N_21271);
or U23392 (N_23392,N_22283,N_22480);
xnor U23393 (N_23393,N_21610,N_21439);
nor U23394 (N_23394,N_22499,N_21639);
nand U23395 (N_23395,N_21877,N_21786);
xnor U23396 (N_23396,N_21391,N_21690);
nor U23397 (N_23397,N_22107,N_22268);
nand U23398 (N_23398,N_21629,N_22252);
or U23399 (N_23399,N_22422,N_21522);
or U23400 (N_23400,N_21755,N_21573);
or U23401 (N_23401,N_21309,N_21263);
and U23402 (N_23402,N_21451,N_22300);
or U23403 (N_23403,N_22475,N_22180);
and U23404 (N_23404,N_22212,N_21540);
nand U23405 (N_23405,N_21648,N_21865);
nor U23406 (N_23406,N_21728,N_21660);
nor U23407 (N_23407,N_22249,N_22305);
and U23408 (N_23408,N_22062,N_21974);
or U23409 (N_23409,N_21763,N_22354);
nand U23410 (N_23410,N_21563,N_22148);
and U23411 (N_23411,N_21924,N_21478);
xor U23412 (N_23412,N_21687,N_21951);
or U23413 (N_23413,N_22321,N_22006);
nor U23414 (N_23414,N_22155,N_22486);
or U23415 (N_23415,N_21701,N_21862);
nor U23416 (N_23416,N_21847,N_22205);
and U23417 (N_23417,N_21769,N_21503);
xor U23418 (N_23418,N_21429,N_21297);
nor U23419 (N_23419,N_21435,N_22307);
xor U23420 (N_23420,N_22389,N_21658);
nor U23421 (N_23421,N_22189,N_21591);
nor U23422 (N_23422,N_21951,N_22496);
nand U23423 (N_23423,N_21990,N_21703);
or U23424 (N_23424,N_21775,N_21888);
xnor U23425 (N_23425,N_22204,N_21759);
nor U23426 (N_23426,N_21700,N_22364);
and U23427 (N_23427,N_22197,N_21540);
and U23428 (N_23428,N_22461,N_21910);
and U23429 (N_23429,N_21738,N_22280);
xnor U23430 (N_23430,N_21884,N_21769);
or U23431 (N_23431,N_22089,N_22252);
xnor U23432 (N_23432,N_21537,N_21816);
and U23433 (N_23433,N_22321,N_22032);
nand U23434 (N_23434,N_22152,N_21284);
xor U23435 (N_23435,N_21319,N_21446);
nand U23436 (N_23436,N_21989,N_21998);
and U23437 (N_23437,N_22430,N_21719);
or U23438 (N_23438,N_21310,N_21780);
nand U23439 (N_23439,N_22279,N_21937);
and U23440 (N_23440,N_21888,N_22094);
and U23441 (N_23441,N_21470,N_21423);
xor U23442 (N_23442,N_22495,N_21478);
and U23443 (N_23443,N_22410,N_21518);
nand U23444 (N_23444,N_22405,N_21971);
nand U23445 (N_23445,N_21473,N_22373);
or U23446 (N_23446,N_21696,N_21794);
nor U23447 (N_23447,N_21890,N_21715);
and U23448 (N_23448,N_21720,N_21478);
or U23449 (N_23449,N_21740,N_21523);
or U23450 (N_23450,N_22473,N_21873);
and U23451 (N_23451,N_22036,N_21486);
nand U23452 (N_23452,N_21459,N_21713);
xor U23453 (N_23453,N_21345,N_22415);
and U23454 (N_23454,N_21370,N_22043);
nor U23455 (N_23455,N_21258,N_22356);
nand U23456 (N_23456,N_22038,N_21735);
and U23457 (N_23457,N_21589,N_21795);
nand U23458 (N_23458,N_21498,N_21933);
nand U23459 (N_23459,N_22365,N_21551);
and U23460 (N_23460,N_22093,N_21325);
or U23461 (N_23461,N_21929,N_22238);
or U23462 (N_23462,N_22020,N_21387);
xor U23463 (N_23463,N_22160,N_21541);
nand U23464 (N_23464,N_22068,N_21350);
nand U23465 (N_23465,N_22242,N_21925);
and U23466 (N_23466,N_21808,N_21829);
nand U23467 (N_23467,N_22124,N_21978);
and U23468 (N_23468,N_21423,N_21285);
and U23469 (N_23469,N_21946,N_21253);
nor U23470 (N_23470,N_21921,N_22206);
xnor U23471 (N_23471,N_22314,N_21259);
nand U23472 (N_23472,N_22142,N_21919);
nor U23473 (N_23473,N_22383,N_22109);
xor U23474 (N_23474,N_22218,N_21505);
nand U23475 (N_23475,N_22060,N_21669);
or U23476 (N_23476,N_21885,N_21301);
and U23477 (N_23477,N_21310,N_22287);
nand U23478 (N_23478,N_22308,N_22069);
or U23479 (N_23479,N_21844,N_22127);
and U23480 (N_23480,N_22005,N_21298);
nand U23481 (N_23481,N_22412,N_22334);
or U23482 (N_23482,N_21259,N_21730);
or U23483 (N_23483,N_21645,N_21441);
and U23484 (N_23484,N_21436,N_22305);
nor U23485 (N_23485,N_21642,N_21365);
nor U23486 (N_23486,N_22414,N_22369);
xor U23487 (N_23487,N_22447,N_22456);
nor U23488 (N_23488,N_21341,N_22472);
nand U23489 (N_23489,N_22234,N_21512);
xnor U23490 (N_23490,N_21667,N_21903);
or U23491 (N_23491,N_22191,N_21878);
or U23492 (N_23492,N_22189,N_22073);
nor U23493 (N_23493,N_21360,N_21298);
xnor U23494 (N_23494,N_21376,N_21943);
xor U23495 (N_23495,N_21864,N_22112);
xor U23496 (N_23496,N_22070,N_21581);
xnor U23497 (N_23497,N_21319,N_21785);
or U23498 (N_23498,N_21742,N_21753);
xnor U23499 (N_23499,N_22183,N_22492);
or U23500 (N_23500,N_21295,N_21695);
xor U23501 (N_23501,N_22350,N_22483);
xor U23502 (N_23502,N_21961,N_21615);
nor U23503 (N_23503,N_22309,N_21943);
and U23504 (N_23504,N_21434,N_21617);
or U23505 (N_23505,N_21942,N_22425);
nor U23506 (N_23506,N_22201,N_21904);
and U23507 (N_23507,N_22417,N_22490);
xnor U23508 (N_23508,N_22119,N_22435);
or U23509 (N_23509,N_21714,N_22054);
or U23510 (N_23510,N_21585,N_21787);
nand U23511 (N_23511,N_22499,N_21942);
and U23512 (N_23512,N_22240,N_22344);
and U23513 (N_23513,N_22342,N_22001);
or U23514 (N_23514,N_21895,N_22242);
xnor U23515 (N_23515,N_21554,N_22369);
and U23516 (N_23516,N_22137,N_21306);
xor U23517 (N_23517,N_22054,N_21445);
and U23518 (N_23518,N_22378,N_22189);
or U23519 (N_23519,N_22093,N_21629);
or U23520 (N_23520,N_22493,N_21556);
nor U23521 (N_23521,N_21860,N_21561);
or U23522 (N_23522,N_22052,N_21435);
xor U23523 (N_23523,N_21367,N_21474);
nand U23524 (N_23524,N_21425,N_21387);
and U23525 (N_23525,N_22471,N_21265);
nand U23526 (N_23526,N_22151,N_22474);
nor U23527 (N_23527,N_21476,N_21953);
or U23528 (N_23528,N_22198,N_21890);
or U23529 (N_23529,N_22181,N_22394);
nand U23530 (N_23530,N_21257,N_21746);
or U23531 (N_23531,N_22030,N_22392);
nor U23532 (N_23532,N_21545,N_22136);
xor U23533 (N_23533,N_22186,N_21878);
or U23534 (N_23534,N_21761,N_21366);
xnor U23535 (N_23535,N_21503,N_21538);
xor U23536 (N_23536,N_21888,N_22496);
nand U23537 (N_23537,N_22096,N_21772);
xnor U23538 (N_23538,N_21282,N_21961);
or U23539 (N_23539,N_21774,N_21264);
or U23540 (N_23540,N_22289,N_22036);
nand U23541 (N_23541,N_21745,N_21646);
xor U23542 (N_23542,N_22456,N_21725);
xnor U23543 (N_23543,N_21796,N_22264);
xnor U23544 (N_23544,N_21857,N_22432);
xor U23545 (N_23545,N_21859,N_21490);
or U23546 (N_23546,N_22457,N_21995);
nand U23547 (N_23547,N_22329,N_21366);
nor U23548 (N_23548,N_21805,N_21390);
nand U23549 (N_23549,N_22251,N_21747);
or U23550 (N_23550,N_21332,N_22297);
or U23551 (N_23551,N_21424,N_21304);
and U23552 (N_23552,N_21774,N_22336);
and U23553 (N_23553,N_21700,N_21630);
and U23554 (N_23554,N_22051,N_22409);
and U23555 (N_23555,N_22088,N_22288);
xnor U23556 (N_23556,N_21614,N_22498);
or U23557 (N_23557,N_22006,N_21779);
nand U23558 (N_23558,N_21964,N_22454);
nand U23559 (N_23559,N_22407,N_21996);
xnor U23560 (N_23560,N_22305,N_21819);
xor U23561 (N_23561,N_22161,N_22052);
xor U23562 (N_23562,N_22199,N_21266);
xnor U23563 (N_23563,N_22132,N_22101);
or U23564 (N_23564,N_22002,N_21763);
nor U23565 (N_23565,N_22045,N_21412);
xor U23566 (N_23566,N_21855,N_21354);
xnor U23567 (N_23567,N_21737,N_21819);
or U23568 (N_23568,N_21760,N_22362);
nand U23569 (N_23569,N_21478,N_21745);
nand U23570 (N_23570,N_22012,N_21993);
nand U23571 (N_23571,N_21991,N_21884);
and U23572 (N_23572,N_21353,N_21922);
and U23573 (N_23573,N_21279,N_22229);
and U23574 (N_23574,N_22183,N_22095);
nand U23575 (N_23575,N_21776,N_21942);
nor U23576 (N_23576,N_21807,N_22057);
xnor U23577 (N_23577,N_21567,N_21401);
nand U23578 (N_23578,N_22312,N_21475);
and U23579 (N_23579,N_21850,N_22134);
nor U23580 (N_23580,N_21904,N_21902);
nand U23581 (N_23581,N_22208,N_22460);
nor U23582 (N_23582,N_21787,N_22159);
nor U23583 (N_23583,N_22078,N_22279);
xor U23584 (N_23584,N_22427,N_21320);
xnor U23585 (N_23585,N_21277,N_21270);
nand U23586 (N_23586,N_21925,N_21463);
nor U23587 (N_23587,N_22493,N_21629);
or U23588 (N_23588,N_22451,N_21652);
nor U23589 (N_23589,N_21952,N_22131);
and U23590 (N_23590,N_22020,N_22058);
nor U23591 (N_23591,N_21974,N_22490);
xnor U23592 (N_23592,N_21756,N_22203);
or U23593 (N_23593,N_21461,N_22428);
and U23594 (N_23594,N_22370,N_22080);
nand U23595 (N_23595,N_21802,N_22014);
and U23596 (N_23596,N_22375,N_22349);
nand U23597 (N_23597,N_22248,N_21262);
nand U23598 (N_23598,N_21998,N_21664);
nor U23599 (N_23599,N_21715,N_21951);
nand U23600 (N_23600,N_22299,N_21808);
xor U23601 (N_23601,N_22398,N_21827);
xnor U23602 (N_23602,N_21621,N_22391);
nand U23603 (N_23603,N_21983,N_21622);
or U23604 (N_23604,N_21387,N_21933);
xnor U23605 (N_23605,N_21419,N_22065);
nor U23606 (N_23606,N_22002,N_21552);
xor U23607 (N_23607,N_21660,N_22431);
nor U23608 (N_23608,N_21478,N_21823);
nand U23609 (N_23609,N_21339,N_21482);
and U23610 (N_23610,N_21731,N_21604);
or U23611 (N_23611,N_22498,N_21759);
or U23612 (N_23612,N_21445,N_22330);
or U23613 (N_23613,N_21829,N_21764);
nor U23614 (N_23614,N_21301,N_22274);
nor U23615 (N_23615,N_22192,N_21703);
xnor U23616 (N_23616,N_21296,N_21576);
nand U23617 (N_23617,N_22208,N_21839);
nor U23618 (N_23618,N_21657,N_22034);
nand U23619 (N_23619,N_22115,N_22030);
nor U23620 (N_23620,N_22084,N_21722);
and U23621 (N_23621,N_21382,N_22181);
and U23622 (N_23622,N_21332,N_22361);
xor U23623 (N_23623,N_21415,N_21380);
nor U23624 (N_23624,N_22089,N_21706);
nor U23625 (N_23625,N_21947,N_21386);
nand U23626 (N_23626,N_21536,N_21304);
nand U23627 (N_23627,N_22400,N_21466);
nand U23628 (N_23628,N_21426,N_21847);
or U23629 (N_23629,N_21478,N_21599);
and U23630 (N_23630,N_22205,N_21367);
nor U23631 (N_23631,N_21918,N_21376);
xnor U23632 (N_23632,N_21288,N_22387);
nor U23633 (N_23633,N_22060,N_21836);
and U23634 (N_23634,N_21858,N_22253);
nor U23635 (N_23635,N_21810,N_21438);
or U23636 (N_23636,N_22062,N_21405);
nand U23637 (N_23637,N_21850,N_21987);
and U23638 (N_23638,N_21393,N_21591);
or U23639 (N_23639,N_22115,N_22296);
xnor U23640 (N_23640,N_21533,N_22292);
and U23641 (N_23641,N_22269,N_22027);
xor U23642 (N_23642,N_22133,N_21647);
or U23643 (N_23643,N_21621,N_22176);
nor U23644 (N_23644,N_22479,N_21453);
nand U23645 (N_23645,N_22442,N_21292);
and U23646 (N_23646,N_22060,N_21860);
and U23647 (N_23647,N_21991,N_22051);
xor U23648 (N_23648,N_21737,N_21562);
nand U23649 (N_23649,N_21496,N_22053);
or U23650 (N_23650,N_21375,N_21680);
and U23651 (N_23651,N_21545,N_21612);
or U23652 (N_23652,N_21816,N_22219);
or U23653 (N_23653,N_22247,N_21616);
and U23654 (N_23654,N_21503,N_22018);
nor U23655 (N_23655,N_22310,N_22149);
and U23656 (N_23656,N_22328,N_22440);
xnor U23657 (N_23657,N_22363,N_22382);
or U23658 (N_23658,N_22113,N_21621);
nand U23659 (N_23659,N_22208,N_21599);
xnor U23660 (N_23660,N_21753,N_22048);
nand U23661 (N_23661,N_21447,N_22460);
and U23662 (N_23662,N_22165,N_21869);
and U23663 (N_23663,N_21599,N_21631);
and U23664 (N_23664,N_22191,N_21975);
nor U23665 (N_23665,N_21400,N_22181);
or U23666 (N_23666,N_21485,N_22373);
and U23667 (N_23667,N_22166,N_22285);
and U23668 (N_23668,N_22250,N_21353);
and U23669 (N_23669,N_21747,N_21250);
nor U23670 (N_23670,N_22271,N_21888);
or U23671 (N_23671,N_21620,N_21885);
and U23672 (N_23672,N_22479,N_21469);
nand U23673 (N_23673,N_21443,N_21362);
or U23674 (N_23674,N_21765,N_21792);
or U23675 (N_23675,N_21900,N_21726);
nor U23676 (N_23676,N_22410,N_21926);
or U23677 (N_23677,N_21675,N_21928);
nand U23678 (N_23678,N_22446,N_21366);
nand U23679 (N_23679,N_21750,N_21794);
and U23680 (N_23680,N_21914,N_22422);
nand U23681 (N_23681,N_21482,N_21391);
nand U23682 (N_23682,N_21508,N_21465);
xnor U23683 (N_23683,N_22347,N_22211);
nand U23684 (N_23684,N_22484,N_21990);
or U23685 (N_23685,N_21887,N_21334);
nor U23686 (N_23686,N_21341,N_21595);
nand U23687 (N_23687,N_22270,N_21774);
or U23688 (N_23688,N_21382,N_22098);
nor U23689 (N_23689,N_21524,N_22220);
and U23690 (N_23690,N_21583,N_21809);
nand U23691 (N_23691,N_22355,N_22082);
nand U23692 (N_23692,N_22020,N_21440);
nand U23693 (N_23693,N_21989,N_21446);
xnor U23694 (N_23694,N_21660,N_21535);
and U23695 (N_23695,N_21578,N_22314);
and U23696 (N_23696,N_22329,N_22182);
and U23697 (N_23697,N_22014,N_22058);
xnor U23698 (N_23698,N_21520,N_21540);
and U23699 (N_23699,N_21520,N_21391);
nor U23700 (N_23700,N_21583,N_21768);
and U23701 (N_23701,N_22090,N_21273);
or U23702 (N_23702,N_22161,N_22414);
nor U23703 (N_23703,N_21360,N_21594);
or U23704 (N_23704,N_22159,N_21285);
and U23705 (N_23705,N_21831,N_22063);
nand U23706 (N_23706,N_21372,N_21927);
or U23707 (N_23707,N_21665,N_21848);
xor U23708 (N_23708,N_22109,N_21482);
or U23709 (N_23709,N_22454,N_22115);
or U23710 (N_23710,N_21772,N_22041);
xor U23711 (N_23711,N_21994,N_22005);
and U23712 (N_23712,N_22285,N_21473);
or U23713 (N_23713,N_21971,N_21597);
nor U23714 (N_23714,N_22472,N_21459);
xnor U23715 (N_23715,N_22123,N_22232);
nand U23716 (N_23716,N_21749,N_21608);
xor U23717 (N_23717,N_21806,N_22023);
nor U23718 (N_23718,N_21325,N_21547);
nor U23719 (N_23719,N_21672,N_22016);
and U23720 (N_23720,N_21350,N_21283);
or U23721 (N_23721,N_22126,N_21794);
or U23722 (N_23722,N_22375,N_21988);
nand U23723 (N_23723,N_22166,N_21746);
and U23724 (N_23724,N_21587,N_22462);
nand U23725 (N_23725,N_22488,N_21486);
or U23726 (N_23726,N_22473,N_21376);
and U23727 (N_23727,N_21398,N_22011);
or U23728 (N_23728,N_22377,N_21307);
or U23729 (N_23729,N_21301,N_21700);
and U23730 (N_23730,N_21797,N_21891);
and U23731 (N_23731,N_22185,N_21791);
xor U23732 (N_23732,N_21964,N_22416);
xnor U23733 (N_23733,N_21693,N_22419);
nor U23734 (N_23734,N_22120,N_22099);
xnor U23735 (N_23735,N_21289,N_22187);
nand U23736 (N_23736,N_21388,N_21462);
or U23737 (N_23737,N_22358,N_21740);
nand U23738 (N_23738,N_22310,N_21921);
nand U23739 (N_23739,N_21470,N_21981);
or U23740 (N_23740,N_22381,N_21416);
and U23741 (N_23741,N_21635,N_21561);
nand U23742 (N_23742,N_21449,N_21474);
or U23743 (N_23743,N_21797,N_22073);
xnor U23744 (N_23744,N_21316,N_21782);
and U23745 (N_23745,N_21368,N_22369);
xor U23746 (N_23746,N_21614,N_22196);
and U23747 (N_23747,N_21687,N_21737);
nor U23748 (N_23748,N_21785,N_21440);
nor U23749 (N_23749,N_21473,N_22387);
xnor U23750 (N_23750,N_23123,N_22899);
and U23751 (N_23751,N_23241,N_23047);
nand U23752 (N_23752,N_23185,N_23398);
xnor U23753 (N_23753,N_23636,N_23386);
and U23754 (N_23754,N_23472,N_22933);
and U23755 (N_23755,N_22562,N_23626);
and U23756 (N_23756,N_23066,N_23593);
nand U23757 (N_23757,N_22703,N_23006);
xnor U23758 (N_23758,N_22743,N_22865);
and U23759 (N_23759,N_23045,N_22552);
nand U23760 (N_23760,N_22953,N_23606);
nor U23761 (N_23761,N_23265,N_23556);
or U23762 (N_23762,N_23608,N_22840);
nor U23763 (N_23763,N_23745,N_22558);
nand U23764 (N_23764,N_23748,N_23229);
and U23765 (N_23765,N_23187,N_23087);
or U23766 (N_23766,N_22504,N_23350);
nand U23767 (N_23767,N_22734,N_22700);
nor U23768 (N_23768,N_23330,N_22878);
xor U23769 (N_23769,N_22883,N_22637);
or U23770 (N_23770,N_22560,N_22891);
or U23771 (N_23771,N_23296,N_23436);
nor U23772 (N_23772,N_22785,N_22863);
xnor U23773 (N_23773,N_22604,N_23509);
and U23774 (N_23774,N_23297,N_23527);
or U23775 (N_23775,N_22776,N_22751);
xnor U23776 (N_23776,N_22991,N_23740);
xnor U23777 (N_23777,N_23613,N_23703);
nor U23778 (N_23778,N_22744,N_22737);
nor U23779 (N_23779,N_23152,N_22910);
nand U23780 (N_23780,N_23447,N_22733);
nand U23781 (N_23781,N_22729,N_23724);
nor U23782 (N_23782,N_23052,N_22642);
nor U23783 (N_23783,N_22831,N_23396);
or U23784 (N_23784,N_23545,N_23498);
and U23785 (N_23785,N_23487,N_22522);
nand U23786 (N_23786,N_22648,N_23294);
nor U23787 (N_23787,N_22887,N_23729);
or U23788 (N_23788,N_22923,N_23739);
or U23789 (N_23789,N_23523,N_22971);
and U23790 (N_23790,N_23643,N_22727);
nand U23791 (N_23791,N_23146,N_23315);
nand U23792 (N_23792,N_22872,N_23291);
and U23793 (N_23793,N_23081,N_22828);
or U23794 (N_23794,N_23638,N_23639);
and U23795 (N_23795,N_23283,N_22985);
nand U23796 (N_23796,N_22508,N_22928);
and U23797 (N_23797,N_22740,N_22809);
nor U23798 (N_23798,N_22806,N_22871);
or U23799 (N_23799,N_23749,N_23064);
or U23800 (N_23800,N_22870,N_23238);
and U23801 (N_23801,N_23010,N_23595);
nor U23802 (N_23802,N_22681,N_23685);
or U23803 (N_23803,N_23226,N_22800);
or U23804 (N_23804,N_22981,N_22708);
nand U23805 (N_23805,N_23099,N_22797);
and U23806 (N_23806,N_23602,N_22969);
nand U23807 (N_23807,N_22722,N_23687);
and U23808 (N_23808,N_22533,N_23132);
xor U23809 (N_23809,N_23631,N_23412);
nand U23810 (N_23810,N_23597,N_23014);
xnor U23811 (N_23811,N_22812,N_22753);
nand U23812 (N_23812,N_22696,N_22687);
nor U23813 (N_23813,N_22919,N_23374);
nor U23814 (N_23814,N_23660,N_22520);
and U23815 (N_23815,N_22750,N_22741);
nor U23816 (N_23816,N_23600,N_23103);
or U23817 (N_23817,N_23661,N_23275);
nand U23818 (N_23818,N_23526,N_23303);
xnor U23819 (N_23819,N_23278,N_23366);
or U23820 (N_23820,N_23407,N_22548);
nand U23821 (N_23821,N_22852,N_23359);
nand U23822 (N_23822,N_22745,N_22967);
and U23823 (N_23823,N_23255,N_22627);
and U23824 (N_23824,N_23665,N_23369);
nand U23825 (N_23825,N_23502,N_23723);
nor U23826 (N_23826,N_23156,N_23461);
or U23827 (N_23827,N_23092,N_23449);
nor U23828 (N_23828,N_23174,N_22665);
xor U23829 (N_23829,N_23290,N_23694);
xor U23830 (N_23830,N_23355,N_22921);
xnor U23831 (N_23831,N_23673,N_23354);
nor U23832 (N_23832,N_23462,N_23022);
xor U23833 (N_23833,N_23057,N_23628);
xnor U23834 (N_23834,N_23540,N_23188);
or U23835 (N_23835,N_23438,N_23334);
nand U23836 (N_23836,N_23564,N_23281);
xnor U23837 (N_23837,N_22922,N_23307);
or U23838 (N_23838,N_22541,N_23395);
xor U23839 (N_23839,N_22645,N_23051);
xor U23840 (N_23840,N_23002,N_23108);
or U23841 (N_23841,N_23582,N_22643);
nand U23842 (N_23842,N_22688,N_23482);
or U23843 (N_23843,N_23738,N_23417);
nor U23844 (N_23844,N_22918,N_22599);
and U23845 (N_23845,N_22616,N_23216);
nor U23846 (N_23846,N_23094,N_23253);
and U23847 (N_23847,N_22752,N_23085);
and U23848 (N_23848,N_23424,N_22653);
and U23849 (N_23849,N_22996,N_23031);
or U23850 (N_23850,N_23312,N_23543);
or U23851 (N_23851,N_22995,N_22843);
or U23852 (N_23852,N_23339,N_22868);
xnor U23853 (N_23853,N_23023,N_22578);
and U23854 (N_23854,N_23515,N_23504);
nand U23855 (N_23855,N_23073,N_22769);
nor U23856 (N_23856,N_23041,N_22658);
and U23857 (N_23857,N_23194,N_22987);
nor U23858 (N_23858,N_23557,N_22821);
xnor U23859 (N_23859,N_23465,N_22673);
or U23860 (N_23860,N_23599,N_23488);
xnor U23861 (N_23861,N_22655,N_23384);
and U23862 (N_23862,N_23508,N_23389);
nor U23863 (N_23863,N_23393,N_22901);
or U23864 (N_23864,N_23568,N_23243);
xnor U23865 (N_23865,N_23655,N_23474);
nor U23866 (N_23866,N_22770,N_23642);
and U23867 (N_23867,N_22803,N_23548);
nor U23868 (N_23868,N_23443,N_23627);
and U23869 (N_23869,N_22715,N_22986);
xnor U23870 (N_23870,N_23321,N_22720);
nor U23871 (N_23871,N_23712,N_22997);
nor U23872 (N_23872,N_22774,N_22900);
or U23873 (N_23873,N_23381,N_23165);
nand U23874 (N_23874,N_22537,N_23418);
or U23875 (N_23875,N_23121,N_22517);
and U23876 (N_23876,N_22783,N_23088);
or U23877 (N_23877,N_23616,N_23117);
and U23878 (N_23878,N_23214,N_23679);
or U23879 (N_23879,N_23039,N_23507);
nand U23880 (N_23880,N_23533,N_23125);
nand U23881 (N_23881,N_23313,N_23432);
or U23882 (N_23882,N_23489,N_23383);
nand U23883 (N_23883,N_23005,N_23090);
or U23884 (N_23884,N_22962,N_23563);
and U23885 (N_23885,N_23082,N_22609);
or U23886 (N_23886,N_23570,N_22553);
and U23887 (N_23887,N_22906,N_22713);
nor U23888 (N_23888,N_23172,N_23717);
nor U23889 (N_23889,N_22570,N_23483);
xor U23890 (N_23890,N_23222,N_23206);
xor U23891 (N_23891,N_22973,N_23295);
or U23892 (N_23892,N_23336,N_23182);
xnor U23893 (N_23893,N_23040,N_23578);
or U23894 (N_23894,N_22755,N_23445);
nor U23895 (N_23895,N_22880,N_23305);
or U23896 (N_23896,N_23421,N_22853);
or U23897 (N_23897,N_23442,N_22521);
nand U23898 (N_23898,N_22584,N_23078);
nand U23899 (N_23899,N_22633,N_23205);
and U23900 (N_23900,N_22746,N_23370);
nor U23901 (N_23901,N_23378,N_22980);
xor U23902 (N_23902,N_23588,N_23145);
nor U23903 (N_23903,N_22857,N_22822);
and U23904 (N_23904,N_23013,N_22707);
nor U23905 (N_23905,N_23246,N_23621);
xor U23906 (N_23906,N_23495,N_22913);
or U23907 (N_23907,N_23230,N_23168);
xnor U23908 (N_23908,N_23478,N_22657);
xor U23909 (N_23909,N_22825,N_22567);
or U23910 (N_23910,N_23310,N_23618);
xnor U23911 (N_23911,N_22598,N_22575);
nand U23912 (N_23912,N_23697,N_23292);
nor U23913 (N_23913,N_23276,N_23725);
or U23914 (N_23914,N_22539,N_23457);
and U23915 (N_23915,N_23430,N_22896);
nand U23916 (N_23916,N_22866,N_22808);
xor U23917 (N_23917,N_23537,N_23151);
and U23918 (N_23918,N_23178,N_22931);
and U23919 (N_23919,N_23084,N_23361);
nand U23920 (N_23920,N_23195,N_23624);
xnor U23921 (N_23921,N_23542,N_22649);
and U23922 (N_23922,N_22704,N_22591);
xnor U23923 (N_23923,N_23100,N_22735);
xor U23924 (N_23924,N_22585,N_22577);
or U23925 (N_23925,N_23586,N_23245);
and U23926 (N_23926,N_23607,N_22869);
nand U23927 (N_23927,N_23452,N_22613);
nor U23928 (N_23928,N_23467,N_22778);
and U23929 (N_23929,N_23219,N_23539);
or U23930 (N_23930,N_23401,N_23653);
or U23931 (N_23931,N_23622,N_23217);
or U23932 (N_23932,N_22723,N_23630);
nor U23933 (N_23933,N_22698,N_23562);
or U23934 (N_23934,N_22763,N_22544);
or U23935 (N_23935,N_22731,N_23218);
nor U23936 (N_23936,N_22932,N_23373);
and U23937 (N_23937,N_23109,N_23302);
nor U23938 (N_23938,N_22747,N_22719);
xnor U23939 (N_23939,N_22782,N_23404);
xnor U23940 (N_23940,N_23228,N_23377);
or U23941 (N_23941,N_22624,N_23162);
nand U23942 (N_23942,N_23201,N_23416);
xor U23943 (N_23943,N_22659,N_22728);
nor U23944 (N_23944,N_23577,N_22571);
nand U23945 (N_23945,N_22824,N_22671);
nand U23946 (N_23946,N_22989,N_23332);
nor U23947 (N_23947,N_22529,N_22938);
nand U23948 (N_23948,N_23391,N_23667);
nand U23949 (N_23949,N_23362,N_23728);
or U23950 (N_23950,N_23718,N_22817);
xnor U23951 (N_23951,N_23583,N_23063);
nand U23952 (N_23952,N_23306,N_23352);
nor U23953 (N_23953,N_22949,N_22937);
nor U23954 (N_23954,N_23551,N_22582);
or U23955 (N_23955,N_23514,N_22787);
nand U23956 (N_23956,N_23707,N_23609);
nand U23957 (N_23957,N_22668,N_23670);
nor U23958 (N_23958,N_22676,N_23122);
xor U23959 (N_23959,N_23301,N_22507);
and U23960 (N_23960,N_22966,N_22693);
or U23961 (N_23961,N_22630,N_22513);
nand U23962 (N_23962,N_23086,N_22619);
or U23963 (N_23963,N_23271,N_22855);
or U23964 (N_23964,N_23322,N_23196);
or U23965 (N_23965,N_23525,N_23575);
and U23966 (N_23966,N_23505,N_23049);
xnor U23967 (N_23967,N_22897,N_22826);
nor U23968 (N_23968,N_23065,N_22602);
nand U23969 (N_23969,N_22773,N_23554);
nor U23970 (N_23970,N_23069,N_23299);
and U23971 (N_23971,N_23026,N_22695);
xnor U23972 (N_23972,N_23696,N_22816);
and U23973 (N_23973,N_23469,N_22646);
or U23974 (N_23974,N_23688,N_22972);
or U23975 (N_23975,N_23160,N_22959);
or U23976 (N_23976,N_23349,N_23364);
nand U23977 (N_23977,N_23284,N_22586);
or U23978 (N_23978,N_22535,N_22902);
xor U23979 (N_23979,N_22511,N_23426);
or U23980 (N_23980,N_23024,N_23617);
or U23981 (N_23981,N_22982,N_23372);
xnor U23982 (N_23982,N_22538,N_23220);
nand U23983 (N_23983,N_22569,N_22672);
and U23984 (N_23984,N_23662,N_23632);
or U23985 (N_23985,N_23096,N_23183);
xor U23986 (N_23986,N_22764,N_23468);
nor U23987 (N_23987,N_23181,N_22968);
nor U23988 (N_23988,N_22682,N_23419);
nor U23989 (N_23989,N_22509,N_23249);
nand U23990 (N_23990,N_22791,N_22705);
or U23991 (N_23991,N_22994,N_23272);
nor U23992 (N_23992,N_23475,N_23722);
nand U23993 (N_23993,N_22777,N_23644);
nand U23994 (N_23994,N_23314,N_23437);
and U23995 (N_23995,N_22784,N_23133);
or U23996 (N_23996,N_22819,N_22850);
nor U23997 (N_23997,N_22915,N_23671);
or U23998 (N_23998,N_22556,N_22675);
nor U23999 (N_23999,N_23298,N_23387);
and U24000 (N_24000,N_23119,N_22805);
and U24001 (N_24001,N_22641,N_23036);
xnor U24002 (N_24002,N_23319,N_23730);
nor U24003 (N_24003,N_22654,N_22683);
and U24004 (N_24004,N_22796,N_22835);
nand U24005 (N_24005,N_23277,N_22839);
nor U24006 (N_24006,N_23252,N_23280);
nand U24007 (N_24007,N_22628,N_22532);
nand U24008 (N_24008,N_23080,N_23675);
nand U24009 (N_24009,N_23309,N_23136);
nand U24010 (N_24010,N_22608,N_23546);
and U24011 (N_24011,N_22829,N_23158);
or U24012 (N_24012,N_23128,N_23536);
and U24013 (N_24013,N_23360,N_22946);
or U24014 (N_24014,N_23154,N_22974);
or U24015 (N_24015,N_22815,N_22905);
nand U24016 (N_24016,N_23008,N_22951);
nor U24017 (N_24017,N_23333,N_22717);
or U24018 (N_24018,N_22559,N_23325);
nor U24019 (N_24019,N_23204,N_22786);
xor U24020 (N_24020,N_22543,N_23706);
nor U24021 (N_24021,N_22677,N_22638);
and U24022 (N_24022,N_22780,N_23138);
and U24023 (N_24023,N_22589,N_23403);
nand U24024 (N_24024,N_22534,N_23590);
or U24025 (N_24025,N_22847,N_23254);
nand U24026 (N_24026,N_23484,N_22531);
xor U24027 (N_24027,N_22592,N_22622);
xor U24028 (N_24028,N_23463,N_23464);
nor U24029 (N_24029,N_22944,N_22849);
nor U24030 (N_24030,N_22941,N_22930);
nor U24031 (N_24031,N_22739,N_23409);
nor U24032 (N_24032,N_23511,N_23074);
or U24033 (N_24033,N_23574,N_22551);
nand U24034 (N_24034,N_23363,N_22632);
or U24035 (N_24035,N_23439,N_22948);
nor U24036 (N_24036,N_23112,N_23144);
and U24037 (N_24037,N_22975,N_23388);
and U24038 (N_24038,N_22712,N_23155);
xor U24039 (N_24039,N_22998,N_23657);
nor U24040 (N_24040,N_23589,N_22841);
xor U24041 (N_24041,N_23209,N_22542);
nor U24042 (N_24042,N_22939,N_22935);
or U24043 (N_24043,N_23062,N_22781);
nor U24044 (N_24044,N_22793,N_23191);
nor U24045 (N_24045,N_22832,N_22754);
nor U24046 (N_24046,N_22927,N_22779);
nor U24047 (N_24047,N_23000,N_22801);
or U24048 (N_24048,N_23676,N_23528);
and U24049 (N_24049,N_23098,N_23202);
nand U24050 (N_24050,N_22629,N_23732);
and U24051 (N_24051,N_22958,N_22512);
or U24052 (N_24052,N_22768,N_23203);
xnor U24053 (N_24053,N_22718,N_23343);
and U24054 (N_24054,N_23260,N_23454);
nand U24055 (N_24055,N_23274,N_23658);
and U24056 (N_24056,N_23500,N_22684);
and U24057 (N_24057,N_22549,N_23479);
xor U24058 (N_24058,N_23293,N_23455);
and U24059 (N_24059,N_22983,N_23397);
nand U24060 (N_24060,N_22579,N_23674);
and U24061 (N_24061,N_23017,N_23259);
and U24062 (N_24062,N_23025,N_22590);
and U24063 (N_24063,N_22775,N_22886);
nand U24064 (N_24064,N_23571,N_23164);
xor U24065 (N_24065,N_22561,N_23341);
xnor U24066 (N_24066,N_23612,N_23604);
or U24067 (N_24067,N_22732,N_22639);
or U24068 (N_24068,N_22725,N_23170);
or U24069 (N_24069,N_22757,N_23089);
or U24070 (N_24070,N_23032,N_22851);
nor U24071 (N_24071,N_22963,N_23423);
or U24072 (N_24072,N_22957,N_23046);
xor U24073 (N_24073,N_23077,N_23058);
nor U24074 (N_24074,N_22595,N_23385);
nor U24075 (N_24075,N_23736,N_22860);
nand U24076 (N_24076,N_22756,N_23251);
or U24077 (N_24077,N_23646,N_23329);
and U24078 (N_24078,N_23601,N_23692);
or U24079 (N_24079,N_22514,N_23742);
xnor U24080 (N_24080,N_23375,N_23235);
or U24081 (N_24081,N_22563,N_22837);
nor U24082 (N_24082,N_23726,N_23038);
nand U24083 (N_24083,N_23494,N_22518);
nand U24084 (N_24084,N_23471,N_22554);
and U24085 (N_24085,N_23506,N_22909);
nor U24086 (N_24086,N_23264,N_23027);
or U24087 (N_24087,N_22701,N_22929);
or U24088 (N_24088,N_22914,N_23139);
nand U24089 (N_24089,N_23737,N_23415);
nor U24090 (N_24090,N_22947,N_22856);
or U24091 (N_24091,N_23450,N_23001);
and U24092 (N_24092,N_22614,N_23141);
nand U24093 (N_24093,N_23143,N_23328);
or U24094 (N_24094,N_23097,N_23250);
nand U24095 (N_24095,N_23576,N_23734);
nand U24096 (N_24096,N_22664,N_22845);
xor U24097 (N_24097,N_23231,N_22692);
and U24098 (N_24098,N_23242,N_23079);
nor U24099 (N_24099,N_22873,N_23282);
and U24100 (N_24100,N_22594,N_23560);
xnor U24101 (N_24101,N_23104,N_23520);
and U24102 (N_24102,N_23267,N_23054);
xnor U24103 (N_24103,N_23076,N_23611);
nand U24104 (N_24104,N_23060,N_22706);
and U24105 (N_24105,N_22761,N_23503);
and U24106 (N_24106,N_23470,N_23053);
nor U24107 (N_24107,N_23048,N_22954);
xor U24108 (N_24108,N_23716,N_23650);
nand U24109 (N_24109,N_23435,N_23648);
and U24110 (N_24110,N_22674,N_22650);
nand U24111 (N_24111,N_22526,N_22506);
xnor U24112 (N_24112,N_23709,N_23213);
and U24113 (N_24113,N_22842,N_22876);
or U24114 (N_24114,N_23111,N_23248);
nand U24115 (N_24115,N_22620,N_23743);
nor U24116 (N_24116,N_22945,N_23579);
xor U24117 (N_24117,N_23448,N_22820);
xnor U24118 (N_24118,N_22601,N_23193);
nor U24119 (N_24119,N_22862,N_23440);
or U24120 (N_24120,N_22993,N_23207);
xor U24121 (N_24121,N_23425,N_22912);
xnor U24122 (N_24122,N_22540,N_23596);
nand U24123 (N_24123,N_23331,N_22568);
nor U24124 (N_24124,N_23522,N_22724);
and U24125 (N_24125,N_23020,N_23428);
nand U24126 (N_24126,N_22834,N_22612);
nor U24127 (N_24127,N_23592,N_22956);
and U24128 (N_24128,N_22818,N_22636);
xor U24129 (N_24129,N_23101,N_22859);
nor U24130 (N_24130,N_22790,N_23654);
nand U24131 (N_24131,N_23550,N_22502);
or U24132 (N_24132,N_22730,N_23163);
xnor U24133 (N_24133,N_23664,N_23684);
and U24134 (N_24134,N_22924,N_23167);
nor U24135 (N_24135,N_23486,N_22836);
nand U24136 (N_24136,N_23695,N_22999);
and U24137 (N_24137,N_23413,N_22942);
xnor U24138 (N_24138,N_23270,N_23029);
and U24139 (N_24139,N_23652,N_22789);
nor U24140 (N_24140,N_22895,N_22679);
nand U24141 (N_24141,N_23547,N_23367);
xor U24142 (N_24142,N_23656,N_23702);
and U24143 (N_24143,N_22597,N_23427);
nor U24144 (N_24144,N_22530,N_22893);
and U24145 (N_24145,N_22680,N_23279);
xor U24146 (N_24146,N_23698,N_23683);
and U24147 (N_24147,N_23499,N_23115);
or U24148 (N_24148,N_23316,N_22892);
nand U24149 (N_24149,N_22736,N_23033);
or U24150 (N_24150,N_23126,N_23700);
nor U24151 (N_24151,N_22702,N_22884);
nand U24152 (N_24152,N_22709,N_22660);
nand U24153 (N_24153,N_22647,N_22917);
and U24154 (N_24154,N_23149,N_23338);
and U24155 (N_24155,N_23300,N_23190);
nor U24156 (N_24156,N_23519,N_23256);
xnor U24157 (N_24157,N_23422,N_23147);
nor U24158 (N_24158,N_23171,N_22670);
nor U24159 (N_24159,N_22574,N_23093);
or U24160 (N_24160,N_23068,N_23380);
or U24161 (N_24161,N_22978,N_22802);
or U24162 (N_24162,N_23681,N_23446);
or U24163 (N_24163,N_23261,N_23019);
and U24164 (N_24164,N_23635,N_23699);
xnor U24165 (N_24165,N_23567,N_22605);
nor U24166 (N_24166,N_22908,N_22813);
nor U24167 (N_24167,N_23659,N_23311);
xor U24168 (N_24168,N_22867,N_23414);
xor U24169 (N_24169,N_23565,N_23647);
nand U24170 (N_24170,N_22686,N_22588);
nor U24171 (N_24171,N_23573,N_23521);
xor U24172 (N_24172,N_22742,N_23347);
nor U24173 (N_24173,N_23686,N_23641);
or U24174 (N_24174,N_22903,N_22992);
xor U24175 (N_24175,N_22600,N_22984);
and U24176 (N_24176,N_22714,N_23444);
nor U24177 (N_24177,N_22603,N_23150);
xnor U24178 (N_24178,N_23197,N_23598);
or U24179 (N_24179,N_22581,N_23127);
and U24180 (N_24180,N_22823,N_23645);
nand U24181 (N_24181,N_23224,N_23434);
nand U24182 (N_24182,N_22691,N_22694);
or U24183 (N_24183,N_22640,N_22916);
nor U24184 (N_24184,N_23043,N_23492);
or U24185 (N_24185,N_23666,N_23215);
or U24186 (N_24186,N_23225,N_23747);
or U24187 (N_24187,N_22799,N_22699);
and U24188 (N_24188,N_23406,N_22661);
or U24189 (N_24189,N_22749,N_22519);
or U24190 (N_24190,N_23234,N_23371);
and U24191 (N_24191,N_23176,N_23180);
and U24192 (N_24192,N_22758,N_23585);
nand U24193 (N_24193,N_23067,N_23581);
nand U24194 (N_24194,N_23561,N_23114);
or U24195 (N_24195,N_23353,N_23107);
and U24196 (N_24196,N_23584,N_22669);
and U24197 (N_24197,N_22721,N_22848);
nor U24198 (N_24198,N_23134,N_23429);
nand U24199 (N_24199,N_23677,N_22936);
nor U24200 (N_24200,N_22576,N_23634);
nor U24201 (N_24201,N_23346,N_23131);
nor U24202 (N_24202,N_23266,N_22689);
and U24203 (N_24203,N_23368,N_23317);
xnor U24204 (N_24204,N_23529,N_23211);
nand U24205 (N_24205,N_22716,N_23012);
or U24206 (N_24206,N_23189,N_22523);
nor U24207 (N_24207,N_22557,N_23669);
nor U24208 (N_24208,N_23223,N_23257);
nand U24209 (N_24209,N_23701,N_22934);
nand U24210 (N_24210,N_22573,N_23552);
xor U24211 (N_24211,N_23285,N_23420);
and U24212 (N_24212,N_23708,N_22711);
xnor U24213 (N_24213,N_23594,N_23620);
or U24214 (N_24214,N_23623,N_23693);
xnor U24215 (N_24215,N_22587,N_23348);
xor U24216 (N_24216,N_23566,N_23477);
nand U24217 (N_24217,N_23318,N_22875);
nor U24218 (N_24218,N_23135,N_22830);
xor U24219 (N_24219,N_23018,N_23232);
nand U24220 (N_24220,N_23210,N_23061);
or U24221 (N_24221,N_23240,N_23177);
nor U24222 (N_24222,N_23516,N_22528);
and U24223 (N_24223,N_23198,N_22798);
nand U24224 (N_24224,N_22955,N_22771);
nor U24225 (N_24225,N_23715,N_23351);
and U24226 (N_24226,N_23344,N_23569);
or U24227 (N_24227,N_23733,N_22960);
or U24228 (N_24228,N_22885,N_22772);
nand U24229 (N_24229,N_22844,N_22990);
or U24230 (N_24230,N_23510,N_23541);
nand U24231 (N_24231,N_22583,N_22545);
nor U24232 (N_24232,N_23605,N_23714);
and U24233 (N_24233,N_22760,N_23221);
or U24234 (N_24234,N_23460,N_22748);
xor U24235 (N_24235,N_22536,N_23534);
or U24236 (N_24236,N_23345,N_22861);
nand U24237 (N_24237,N_22524,N_23524);
or U24238 (N_24238,N_22596,N_23559);
or U24239 (N_24239,N_23083,N_23239);
nand U24240 (N_24240,N_23179,N_22710);
and U24241 (N_24241,N_23056,N_23184);
and U24242 (N_24242,N_22898,N_23320);
and U24243 (N_24243,N_23095,N_23672);
nor U24244 (N_24244,N_22838,N_22976);
nand U24245 (N_24245,N_23441,N_22881);
nor U24246 (N_24246,N_22516,N_23075);
nor U24247 (N_24247,N_23070,N_22810);
nor U24248 (N_24248,N_22610,N_23433);
or U24249 (N_24249,N_23485,N_23304);
xnor U24250 (N_24250,N_23480,N_23587);
nor U24251 (N_24251,N_23335,N_23402);
xnor U24252 (N_24252,N_23553,N_23493);
xor U24253 (N_24253,N_22907,N_23705);
xor U24254 (N_24254,N_22697,N_22634);
or U24255 (N_24255,N_22505,N_23142);
nor U24256 (N_24256,N_22846,N_23610);
or U24257 (N_24257,N_23663,N_23327);
nand U24258 (N_24258,N_22970,N_22765);
nand U24259 (N_24259,N_23431,N_23517);
nor U24260 (N_24260,N_22617,N_23091);
nand U24261 (N_24261,N_22833,N_23161);
and U24262 (N_24262,N_23518,N_23640);
nand U24263 (N_24263,N_23451,N_23153);
and U24264 (N_24264,N_23130,N_23365);
nor U24265 (N_24265,N_23410,N_23116);
nor U24266 (N_24266,N_22988,N_22940);
and U24267 (N_24267,N_23473,N_22827);
xor U24268 (N_24268,N_23459,N_23035);
xnor U24269 (N_24269,N_23105,N_23501);
nand U24270 (N_24270,N_23113,N_23649);
nor U24271 (N_24271,N_23691,N_23028);
nor U24272 (N_24272,N_23651,N_23615);
nand U24273 (N_24273,N_22926,N_23496);
and U24274 (N_24274,N_22550,N_23258);
nor U24275 (N_24275,N_23558,N_23140);
and U24276 (N_24276,N_22501,N_23244);
nand U24277 (N_24277,N_22767,N_22566);
nand U24278 (N_24278,N_22515,N_23356);
xnor U24279 (N_24279,N_22625,N_22920);
and U24280 (N_24280,N_23050,N_23491);
nor U24281 (N_24281,N_23236,N_22623);
nand U24282 (N_24282,N_22555,N_23288);
xnor U24283 (N_24283,N_23721,N_22925);
and U24284 (N_24284,N_23110,N_22965);
nand U24285 (N_24285,N_23357,N_23591);
nand U24286 (N_24286,N_22814,N_23411);
nor U24287 (N_24287,N_23358,N_23572);
nor U24288 (N_24288,N_23619,N_23735);
nand U24289 (N_24289,N_23269,N_22977);
and U24290 (N_24290,N_23323,N_23030);
nand U24291 (N_24291,N_23009,N_23129);
and U24292 (N_24292,N_22804,N_23490);
and U24293 (N_24293,N_23247,N_22527);
and U24294 (N_24294,N_23173,N_22615);
nand U24295 (N_24295,N_23466,N_22890);
nor U24296 (N_24296,N_23399,N_23166);
nand U24297 (N_24297,N_22979,N_23476);
and U24298 (N_24298,N_23453,N_22795);
nor U24299 (N_24299,N_23458,N_22807);
xnor U24300 (N_24300,N_22882,N_23021);
and U24301 (N_24301,N_23746,N_23118);
and U24302 (N_24302,N_23233,N_22667);
xor U24303 (N_24303,N_22621,N_22606);
nand U24304 (N_24304,N_22662,N_23400);
xnor U24305 (N_24305,N_23633,N_22666);
nand U24306 (N_24306,N_22792,N_23682);
or U24307 (N_24307,N_23208,N_23741);
nor U24308 (N_24308,N_23011,N_22874);
nor U24309 (N_24309,N_23004,N_22911);
or U24310 (N_24310,N_23042,N_22626);
nor U24311 (N_24311,N_22759,N_23262);
xor U24312 (N_24312,N_22690,N_22685);
nand U24313 (N_24313,N_23392,N_23382);
nor U24314 (N_24314,N_23614,N_23102);
xor U24315 (N_24315,N_23273,N_23263);
nor U24316 (N_24316,N_23308,N_23544);
nand U24317 (N_24317,N_22565,N_22766);
nand U24318 (N_24318,N_22788,N_23071);
and U24319 (N_24319,N_23007,N_23186);
nor U24320 (N_24320,N_23037,N_23497);
nand U24321 (N_24321,N_23148,N_22877);
nor U24322 (N_24322,N_23212,N_23159);
nor U24323 (N_24323,N_22510,N_23512);
nor U24324 (N_24324,N_22964,N_23390);
nor U24325 (N_24325,N_23394,N_23538);
xnor U24326 (N_24326,N_23200,N_23072);
nor U24327 (N_24327,N_23287,N_23324);
nor U24328 (N_24328,N_23016,N_23408);
and U24329 (N_24329,N_23603,N_23379);
xnor U24330 (N_24330,N_23456,N_23192);
or U24331 (N_24331,N_23059,N_22678);
xnor U24332 (N_24332,N_23531,N_22631);
nand U24333 (N_24333,N_22635,N_23268);
xnor U24334 (N_24334,N_22738,N_22950);
and U24335 (N_24335,N_22726,N_23711);
or U24336 (N_24336,N_22864,N_22547);
nor U24337 (N_24337,N_23003,N_23680);
xor U24338 (N_24338,N_22961,N_22564);
nand U24339 (N_24339,N_22952,N_23015);
nor U24340 (N_24340,N_23106,N_23689);
or U24341 (N_24341,N_23513,N_22663);
nor U24342 (N_24342,N_23481,N_22794);
xnor U24343 (N_24343,N_23405,N_22525);
nand U24344 (N_24344,N_23580,N_22888);
nor U24345 (N_24345,N_23668,N_22879);
or U24346 (N_24346,N_23549,N_23530);
nand U24347 (N_24347,N_23227,N_22854);
xor U24348 (N_24348,N_23199,N_22889);
and U24349 (N_24349,N_22580,N_22644);
xor U24350 (N_24350,N_22894,N_22762);
xnor U24351 (N_24351,N_23710,N_22811);
xnor U24352 (N_24352,N_23286,N_23175);
nor U24353 (N_24353,N_23044,N_23704);
nand U24354 (N_24354,N_23720,N_22651);
and U24355 (N_24355,N_23731,N_22656);
xnor U24356 (N_24356,N_22904,N_23137);
nand U24357 (N_24357,N_22500,N_23678);
nor U24358 (N_24358,N_22572,N_22618);
nand U24359 (N_24359,N_23629,N_23326);
nor U24360 (N_24360,N_23342,N_23337);
xnor U24361 (N_24361,N_23625,N_23055);
or U24362 (N_24362,N_22503,N_23535);
nand U24363 (N_24363,N_22593,N_23157);
nor U24364 (N_24364,N_22611,N_23124);
and U24365 (N_24365,N_23169,N_23690);
nand U24366 (N_24366,N_23555,N_23719);
and U24367 (N_24367,N_22546,N_22607);
nor U24368 (N_24368,N_23713,N_22652);
xnor U24369 (N_24369,N_23289,N_23637);
or U24370 (N_24370,N_22858,N_23376);
nor U24371 (N_24371,N_23532,N_23237);
nand U24372 (N_24372,N_23034,N_23340);
or U24373 (N_24373,N_22943,N_23727);
and U24374 (N_24374,N_23120,N_23744);
nor U24375 (N_24375,N_23606,N_23291);
nand U24376 (N_24376,N_23031,N_23447);
nor U24377 (N_24377,N_22865,N_22801);
or U24378 (N_24378,N_22877,N_22634);
and U24379 (N_24379,N_22536,N_23314);
and U24380 (N_24380,N_23266,N_23024);
nand U24381 (N_24381,N_23217,N_23201);
nand U24382 (N_24382,N_22673,N_23225);
and U24383 (N_24383,N_22587,N_23720);
or U24384 (N_24384,N_22577,N_22859);
nand U24385 (N_24385,N_23616,N_22840);
nor U24386 (N_24386,N_23066,N_22773);
nand U24387 (N_24387,N_23716,N_23747);
xnor U24388 (N_24388,N_23388,N_22751);
nor U24389 (N_24389,N_22941,N_23351);
or U24390 (N_24390,N_22973,N_23027);
nor U24391 (N_24391,N_22649,N_23655);
nand U24392 (N_24392,N_23567,N_23297);
nor U24393 (N_24393,N_23585,N_23133);
nand U24394 (N_24394,N_22628,N_23029);
or U24395 (N_24395,N_23072,N_23288);
nor U24396 (N_24396,N_23172,N_22842);
and U24397 (N_24397,N_23323,N_22739);
xor U24398 (N_24398,N_22904,N_23298);
nor U24399 (N_24399,N_22670,N_23376);
nand U24400 (N_24400,N_22798,N_23578);
xor U24401 (N_24401,N_23319,N_22548);
and U24402 (N_24402,N_23667,N_22754);
nor U24403 (N_24403,N_23111,N_23232);
or U24404 (N_24404,N_23538,N_22956);
and U24405 (N_24405,N_23459,N_22639);
and U24406 (N_24406,N_22738,N_23743);
nand U24407 (N_24407,N_22804,N_23002);
or U24408 (N_24408,N_23203,N_22502);
nand U24409 (N_24409,N_22610,N_23607);
xnor U24410 (N_24410,N_23190,N_23492);
xor U24411 (N_24411,N_22971,N_23528);
or U24412 (N_24412,N_23200,N_23339);
nand U24413 (N_24413,N_23528,N_23510);
xor U24414 (N_24414,N_22872,N_23615);
or U24415 (N_24415,N_23194,N_23012);
and U24416 (N_24416,N_22557,N_23327);
nand U24417 (N_24417,N_23091,N_23617);
nor U24418 (N_24418,N_22568,N_23388);
or U24419 (N_24419,N_23732,N_23625);
nand U24420 (N_24420,N_23101,N_23673);
or U24421 (N_24421,N_22756,N_22508);
and U24422 (N_24422,N_22739,N_22548);
nand U24423 (N_24423,N_23144,N_23146);
or U24424 (N_24424,N_23546,N_22813);
nor U24425 (N_24425,N_23009,N_23504);
nand U24426 (N_24426,N_23534,N_23089);
nand U24427 (N_24427,N_22979,N_23634);
nand U24428 (N_24428,N_22908,N_23516);
nand U24429 (N_24429,N_22782,N_22714);
xnor U24430 (N_24430,N_22531,N_22771);
nor U24431 (N_24431,N_23179,N_23209);
or U24432 (N_24432,N_23278,N_23429);
nor U24433 (N_24433,N_23662,N_23392);
nand U24434 (N_24434,N_23636,N_23058);
nor U24435 (N_24435,N_23022,N_23529);
nor U24436 (N_24436,N_22821,N_23646);
or U24437 (N_24437,N_23573,N_23223);
nand U24438 (N_24438,N_22859,N_23594);
xor U24439 (N_24439,N_22928,N_23686);
nand U24440 (N_24440,N_23300,N_23221);
and U24441 (N_24441,N_22632,N_23056);
nand U24442 (N_24442,N_22950,N_23520);
and U24443 (N_24443,N_23147,N_23690);
nor U24444 (N_24444,N_22840,N_23491);
and U24445 (N_24445,N_22736,N_22896);
and U24446 (N_24446,N_23027,N_22843);
nand U24447 (N_24447,N_23093,N_23190);
nand U24448 (N_24448,N_22570,N_23721);
nand U24449 (N_24449,N_23018,N_23245);
nand U24450 (N_24450,N_23638,N_23352);
and U24451 (N_24451,N_23008,N_22684);
nand U24452 (N_24452,N_22938,N_22857);
or U24453 (N_24453,N_23281,N_22950);
nand U24454 (N_24454,N_23341,N_23229);
xnor U24455 (N_24455,N_23074,N_23732);
nor U24456 (N_24456,N_22675,N_23009);
or U24457 (N_24457,N_22780,N_22888);
nor U24458 (N_24458,N_23652,N_22673);
xnor U24459 (N_24459,N_23523,N_22840);
nand U24460 (N_24460,N_22950,N_23058);
xor U24461 (N_24461,N_23227,N_23537);
nand U24462 (N_24462,N_22664,N_23477);
xnor U24463 (N_24463,N_23258,N_23337);
nor U24464 (N_24464,N_23745,N_23428);
or U24465 (N_24465,N_23294,N_23096);
or U24466 (N_24466,N_23063,N_23436);
and U24467 (N_24467,N_22689,N_22557);
or U24468 (N_24468,N_23476,N_22610);
xnor U24469 (N_24469,N_23358,N_23580);
nor U24470 (N_24470,N_23719,N_23578);
xor U24471 (N_24471,N_23274,N_23241);
nand U24472 (N_24472,N_23613,N_22854);
and U24473 (N_24473,N_23504,N_23172);
or U24474 (N_24474,N_23450,N_22914);
nand U24475 (N_24475,N_23306,N_23617);
and U24476 (N_24476,N_23686,N_23015);
or U24477 (N_24477,N_23562,N_23249);
or U24478 (N_24478,N_23199,N_22516);
and U24479 (N_24479,N_22601,N_23738);
nor U24480 (N_24480,N_22539,N_22714);
and U24481 (N_24481,N_22595,N_22778);
nand U24482 (N_24482,N_23413,N_23644);
nand U24483 (N_24483,N_23502,N_23732);
and U24484 (N_24484,N_23021,N_23242);
nand U24485 (N_24485,N_23379,N_22762);
xnor U24486 (N_24486,N_23414,N_22738);
and U24487 (N_24487,N_22860,N_22883);
nor U24488 (N_24488,N_22720,N_23494);
nand U24489 (N_24489,N_23573,N_22557);
nor U24490 (N_24490,N_22711,N_22748);
nor U24491 (N_24491,N_23144,N_22592);
xnor U24492 (N_24492,N_23104,N_22817);
and U24493 (N_24493,N_22508,N_22624);
nand U24494 (N_24494,N_23509,N_23165);
and U24495 (N_24495,N_22704,N_23099);
or U24496 (N_24496,N_23105,N_23285);
or U24497 (N_24497,N_22957,N_23369);
or U24498 (N_24498,N_23149,N_23548);
and U24499 (N_24499,N_22920,N_22903);
nand U24500 (N_24500,N_23731,N_23237);
xnor U24501 (N_24501,N_23383,N_23559);
or U24502 (N_24502,N_23176,N_23670);
xnor U24503 (N_24503,N_23251,N_22691);
nand U24504 (N_24504,N_23274,N_23724);
or U24505 (N_24505,N_23308,N_23274);
nand U24506 (N_24506,N_23687,N_23196);
nor U24507 (N_24507,N_22777,N_23213);
xnor U24508 (N_24508,N_22833,N_22724);
nor U24509 (N_24509,N_22900,N_23288);
nor U24510 (N_24510,N_22693,N_23452);
or U24511 (N_24511,N_22604,N_23599);
and U24512 (N_24512,N_23494,N_23362);
nor U24513 (N_24513,N_23022,N_22754);
xor U24514 (N_24514,N_22849,N_22517);
xor U24515 (N_24515,N_22511,N_23714);
xnor U24516 (N_24516,N_22699,N_23106);
nand U24517 (N_24517,N_22503,N_23602);
and U24518 (N_24518,N_22690,N_23228);
nand U24519 (N_24519,N_22639,N_23678);
and U24520 (N_24520,N_22754,N_23445);
or U24521 (N_24521,N_22988,N_23289);
xor U24522 (N_24522,N_23510,N_23383);
and U24523 (N_24523,N_22629,N_23103);
xnor U24524 (N_24524,N_23104,N_23708);
nand U24525 (N_24525,N_23456,N_23699);
and U24526 (N_24526,N_23376,N_23203);
and U24527 (N_24527,N_22560,N_23720);
or U24528 (N_24528,N_23392,N_23537);
nand U24529 (N_24529,N_23138,N_23071);
and U24530 (N_24530,N_22502,N_23647);
xor U24531 (N_24531,N_23103,N_23729);
xnor U24532 (N_24532,N_22716,N_22710);
and U24533 (N_24533,N_23224,N_22814);
nand U24534 (N_24534,N_22823,N_22846);
or U24535 (N_24535,N_22600,N_23220);
nand U24536 (N_24536,N_23550,N_22971);
nand U24537 (N_24537,N_22914,N_23364);
or U24538 (N_24538,N_23556,N_23539);
nand U24539 (N_24539,N_23063,N_23585);
nor U24540 (N_24540,N_22527,N_23723);
xor U24541 (N_24541,N_23177,N_23465);
and U24542 (N_24542,N_23369,N_22620);
xor U24543 (N_24543,N_22501,N_23340);
and U24544 (N_24544,N_23399,N_22781);
nand U24545 (N_24545,N_22640,N_23280);
nor U24546 (N_24546,N_22906,N_23133);
xnor U24547 (N_24547,N_23686,N_23718);
nand U24548 (N_24548,N_22803,N_23516);
and U24549 (N_24549,N_22882,N_23668);
xor U24550 (N_24550,N_23540,N_23227);
nand U24551 (N_24551,N_23696,N_23356);
nand U24552 (N_24552,N_23460,N_23717);
and U24553 (N_24553,N_23652,N_23649);
nand U24554 (N_24554,N_22680,N_23081);
or U24555 (N_24555,N_23232,N_22862);
xor U24556 (N_24556,N_23715,N_23564);
nand U24557 (N_24557,N_22946,N_23017);
xnor U24558 (N_24558,N_22804,N_23071);
nor U24559 (N_24559,N_23551,N_23196);
and U24560 (N_24560,N_23351,N_22726);
nor U24561 (N_24561,N_23181,N_22642);
xor U24562 (N_24562,N_23683,N_23329);
or U24563 (N_24563,N_23088,N_23277);
nor U24564 (N_24564,N_23650,N_22665);
or U24565 (N_24565,N_22504,N_22796);
xnor U24566 (N_24566,N_23028,N_23091);
or U24567 (N_24567,N_23134,N_23582);
or U24568 (N_24568,N_22659,N_23027);
and U24569 (N_24569,N_23042,N_22845);
or U24570 (N_24570,N_23641,N_22675);
nor U24571 (N_24571,N_23113,N_22789);
or U24572 (N_24572,N_23553,N_23263);
nor U24573 (N_24573,N_23593,N_22925);
and U24574 (N_24574,N_23704,N_22969);
nand U24575 (N_24575,N_22686,N_23388);
or U24576 (N_24576,N_23724,N_23208);
nand U24577 (N_24577,N_23740,N_22880);
nor U24578 (N_24578,N_22790,N_23649);
and U24579 (N_24579,N_23101,N_22848);
nor U24580 (N_24580,N_23441,N_23564);
and U24581 (N_24581,N_22855,N_22602);
and U24582 (N_24582,N_23418,N_23576);
nor U24583 (N_24583,N_23611,N_23741);
or U24584 (N_24584,N_23741,N_22827);
and U24585 (N_24585,N_23636,N_22971);
xor U24586 (N_24586,N_22557,N_23514);
and U24587 (N_24587,N_22965,N_23668);
nand U24588 (N_24588,N_23629,N_22702);
nand U24589 (N_24589,N_23114,N_23572);
or U24590 (N_24590,N_23206,N_22861);
or U24591 (N_24591,N_23097,N_22797);
xor U24592 (N_24592,N_23032,N_22521);
xnor U24593 (N_24593,N_23664,N_23532);
xor U24594 (N_24594,N_22783,N_22635);
or U24595 (N_24595,N_23487,N_23074);
nor U24596 (N_24596,N_23360,N_23600);
or U24597 (N_24597,N_22651,N_22860);
or U24598 (N_24598,N_22854,N_23301);
nor U24599 (N_24599,N_23184,N_23736);
nor U24600 (N_24600,N_23202,N_22878);
nand U24601 (N_24601,N_22539,N_23007);
xnor U24602 (N_24602,N_23673,N_22810);
nand U24603 (N_24603,N_22774,N_23633);
nand U24604 (N_24604,N_22915,N_23010);
or U24605 (N_24605,N_22569,N_23043);
xor U24606 (N_24606,N_22925,N_23008);
or U24607 (N_24607,N_23634,N_23446);
or U24608 (N_24608,N_22886,N_23198);
and U24609 (N_24609,N_23223,N_22907);
nand U24610 (N_24610,N_23402,N_23107);
or U24611 (N_24611,N_23528,N_23414);
nand U24612 (N_24612,N_22733,N_22964);
and U24613 (N_24613,N_22716,N_22505);
and U24614 (N_24614,N_22532,N_22640);
and U24615 (N_24615,N_23622,N_22846);
nor U24616 (N_24616,N_23020,N_23628);
nand U24617 (N_24617,N_22589,N_22874);
xnor U24618 (N_24618,N_22812,N_23043);
nor U24619 (N_24619,N_23302,N_23351);
nand U24620 (N_24620,N_23082,N_23257);
or U24621 (N_24621,N_23552,N_23468);
or U24622 (N_24622,N_22870,N_23320);
xnor U24623 (N_24623,N_22584,N_23234);
nor U24624 (N_24624,N_23178,N_23439);
xnor U24625 (N_24625,N_22818,N_22862);
xnor U24626 (N_24626,N_23397,N_22703);
or U24627 (N_24627,N_22845,N_23537);
or U24628 (N_24628,N_22699,N_22557);
nand U24629 (N_24629,N_23542,N_23143);
nor U24630 (N_24630,N_22895,N_22561);
xnor U24631 (N_24631,N_22531,N_23648);
or U24632 (N_24632,N_23516,N_23535);
and U24633 (N_24633,N_22596,N_22754);
nor U24634 (N_24634,N_23718,N_22836);
and U24635 (N_24635,N_23518,N_22803);
nand U24636 (N_24636,N_22898,N_22872);
nand U24637 (N_24637,N_22709,N_22903);
xnor U24638 (N_24638,N_22755,N_23667);
xor U24639 (N_24639,N_23558,N_22902);
and U24640 (N_24640,N_23397,N_23520);
nand U24641 (N_24641,N_22670,N_23322);
nor U24642 (N_24642,N_23022,N_23137);
and U24643 (N_24643,N_23261,N_22671);
xnor U24644 (N_24644,N_22561,N_23085);
nand U24645 (N_24645,N_23396,N_22910);
and U24646 (N_24646,N_23557,N_23682);
nand U24647 (N_24647,N_23666,N_22916);
or U24648 (N_24648,N_23703,N_22508);
nand U24649 (N_24649,N_23187,N_22710);
and U24650 (N_24650,N_23355,N_22729);
xnor U24651 (N_24651,N_22551,N_23180);
xnor U24652 (N_24652,N_23667,N_22800);
and U24653 (N_24653,N_23011,N_23632);
or U24654 (N_24654,N_22800,N_22733);
nor U24655 (N_24655,N_23682,N_23664);
and U24656 (N_24656,N_22989,N_23252);
nor U24657 (N_24657,N_23114,N_22950);
xnor U24658 (N_24658,N_22571,N_23511);
xor U24659 (N_24659,N_22926,N_23137);
nand U24660 (N_24660,N_23071,N_22521);
or U24661 (N_24661,N_22638,N_22943);
xnor U24662 (N_24662,N_22629,N_23271);
or U24663 (N_24663,N_22983,N_23159);
nand U24664 (N_24664,N_23721,N_23095);
nand U24665 (N_24665,N_23412,N_23098);
xor U24666 (N_24666,N_23064,N_22715);
or U24667 (N_24667,N_22927,N_23230);
nand U24668 (N_24668,N_22740,N_23199);
nand U24669 (N_24669,N_22529,N_23641);
nand U24670 (N_24670,N_23149,N_23692);
and U24671 (N_24671,N_23086,N_23338);
nor U24672 (N_24672,N_23580,N_22688);
xnor U24673 (N_24673,N_22589,N_22801);
nor U24674 (N_24674,N_23400,N_22887);
nand U24675 (N_24675,N_23696,N_22681);
nand U24676 (N_24676,N_23514,N_23149);
nor U24677 (N_24677,N_23074,N_23572);
and U24678 (N_24678,N_23669,N_22938);
nor U24679 (N_24679,N_23392,N_23486);
xor U24680 (N_24680,N_23542,N_23073);
xor U24681 (N_24681,N_22660,N_22793);
nor U24682 (N_24682,N_23392,N_23247);
or U24683 (N_24683,N_23063,N_23126);
nand U24684 (N_24684,N_23662,N_22841);
and U24685 (N_24685,N_23031,N_23371);
and U24686 (N_24686,N_23046,N_22852);
nand U24687 (N_24687,N_23719,N_22926);
or U24688 (N_24688,N_23424,N_23106);
nor U24689 (N_24689,N_22979,N_23674);
nor U24690 (N_24690,N_22898,N_22604);
xor U24691 (N_24691,N_23182,N_22875);
nor U24692 (N_24692,N_22621,N_23353);
or U24693 (N_24693,N_23485,N_22890);
nand U24694 (N_24694,N_23675,N_23453);
nor U24695 (N_24695,N_22746,N_22725);
nor U24696 (N_24696,N_23667,N_23417);
xnor U24697 (N_24697,N_22601,N_22815);
and U24698 (N_24698,N_23409,N_23696);
nor U24699 (N_24699,N_22726,N_23542);
xor U24700 (N_24700,N_23580,N_23067);
or U24701 (N_24701,N_22763,N_23607);
or U24702 (N_24702,N_23161,N_23281);
nor U24703 (N_24703,N_22847,N_23024);
or U24704 (N_24704,N_23327,N_22932);
or U24705 (N_24705,N_22596,N_22961);
and U24706 (N_24706,N_23723,N_23508);
and U24707 (N_24707,N_22731,N_23453);
nand U24708 (N_24708,N_23321,N_23014);
nor U24709 (N_24709,N_22816,N_22507);
xor U24710 (N_24710,N_23163,N_23590);
and U24711 (N_24711,N_23218,N_23022);
and U24712 (N_24712,N_23109,N_23639);
xnor U24713 (N_24713,N_23454,N_22702);
nor U24714 (N_24714,N_22712,N_22595);
and U24715 (N_24715,N_22904,N_23420);
nand U24716 (N_24716,N_23487,N_23301);
xnor U24717 (N_24717,N_23364,N_22993);
or U24718 (N_24718,N_22757,N_22989);
or U24719 (N_24719,N_23493,N_22692);
nor U24720 (N_24720,N_23665,N_22883);
nand U24721 (N_24721,N_23594,N_23727);
and U24722 (N_24722,N_23031,N_23117);
nand U24723 (N_24723,N_23406,N_23375);
and U24724 (N_24724,N_23424,N_23201);
nand U24725 (N_24725,N_22805,N_22907);
and U24726 (N_24726,N_23460,N_23382);
xor U24727 (N_24727,N_23506,N_23165);
nor U24728 (N_24728,N_22500,N_22721);
xnor U24729 (N_24729,N_23221,N_22890);
nand U24730 (N_24730,N_23459,N_22946);
and U24731 (N_24731,N_22515,N_23705);
and U24732 (N_24732,N_23584,N_22854);
nor U24733 (N_24733,N_22905,N_22699);
or U24734 (N_24734,N_23579,N_23337);
xor U24735 (N_24735,N_23278,N_23386);
and U24736 (N_24736,N_23334,N_22549);
nor U24737 (N_24737,N_23300,N_22599);
nand U24738 (N_24738,N_23739,N_23495);
and U24739 (N_24739,N_22572,N_22523);
xnor U24740 (N_24740,N_23429,N_23625);
and U24741 (N_24741,N_23246,N_23557);
and U24742 (N_24742,N_22696,N_22963);
xor U24743 (N_24743,N_23362,N_23533);
nor U24744 (N_24744,N_22903,N_22590);
and U24745 (N_24745,N_23730,N_22852);
or U24746 (N_24746,N_23383,N_23387);
and U24747 (N_24747,N_23038,N_22554);
xor U24748 (N_24748,N_23049,N_22812);
nand U24749 (N_24749,N_22778,N_22673);
or U24750 (N_24750,N_22656,N_23524);
nand U24751 (N_24751,N_23661,N_22615);
xor U24752 (N_24752,N_23430,N_23025);
nand U24753 (N_24753,N_23149,N_22563);
nor U24754 (N_24754,N_23018,N_22538);
nand U24755 (N_24755,N_23050,N_23396);
xnor U24756 (N_24756,N_23036,N_23001);
nor U24757 (N_24757,N_23517,N_22908);
or U24758 (N_24758,N_22951,N_22636);
nand U24759 (N_24759,N_23626,N_23634);
and U24760 (N_24760,N_22938,N_22771);
or U24761 (N_24761,N_22654,N_23041);
and U24762 (N_24762,N_23174,N_22744);
xnor U24763 (N_24763,N_23721,N_23134);
or U24764 (N_24764,N_22713,N_23003);
or U24765 (N_24765,N_23275,N_23679);
xnor U24766 (N_24766,N_22732,N_23103);
nand U24767 (N_24767,N_22595,N_23669);
nor U24768 (N_24768,N_22721,N_23235);
xor U24769 (N_24769,N_23072,N_23173);
nand U24770 (N_24770,N_23033,N_23165);
nand U24771 (N_24771,N_23097,N_23739);
nand U24772 (N_24772,N_22735,N_23189);
or U24773 (N_24773,N_22885,N_23387);
nand U24774 (N_24774,N_23689,N_23486);
or U24775 (N_24775,N_22839,N_23635);
or U24776 (N_24776,N_22718,N_22982);
nand U24777 (N_24777,N_23300,N_23142);
or U24778 (N_24778,N_22815,N_23689);
or U24779 (N_24779,N_23050,N_22848);
or U24780 (N_24780,N_22788,N_22545);
nand U24781 (N_24781,N_23157,N_23589);
nor U24782 (N_24782,N_23522,N_23392);
nor U24783 (N_24783,N_22649,N_22732);
xor U24784 (N_24784,N_22633,N_22753);
nor U24785 (N_24785,N_22716,N_23278);
nor U24786 (N_24786,N_22906,N_23045);
or U24787 (N_24787,N_23041,N_22646);
and U24788 (N_24788,N_22545,N_23058);
xnor U24789 (N_24789,N_22588,N_23371);
or U24790 (N_24790,N_23280,N_22794);
nand U24791 (N_24791,N_23658,N_23232);
nand U24792 (N_24792,N_23056,N_23725);
and U24793 (N_24793,N_23399,N_22699);
and U24794 (N_24794,N_23227,N_22580);
nand U24795 (N_24795,N_23214,N_23611);
xor U24796 (N_24796,N_22937,N_23020);
nor U24797 (N_24797,N_22851,N_23128);
nor U24798 (N_24798,N_22525,N_23013);
xnor U24799 (N_24799,N_23448,N_22548);
nor U24800 (N_24800,N_22688,N_23589);
xnor U24801 (N_24801,N_23303,N_23579);
nor U24802 (N_24802,N_23636,N_23293);
nand U24803 (N_24803,N_23176,N_22949);
and U24804 (N_24804,N_23445,N_23616);
nand U24805 (N_24805,N_22513,N_22524);
xor U24806 (N_24806,N_22680,N_22730);
or U24807 (N_24807,N_23164,N_22877);
or U24808 (N_24808,N_23253,N_23470);
and U24809 (N_24809,N_22582,N_23226);
or U24810 (N_24810,N_23271,N_23440);
xnor U24811 (N_24811,N_22788,N_23133);
and U24812 (N_24812,N_23601,N_23000);
and U24813 (N_24813,N_22546,N_23098);
and U24814 (N_24814,N_23417,N_22701);
nor U24815 (N_24815,N_23184,N_22709);
and U24816 (N_24816,N_23329,N_23673);
or U24817 (N_24817,N_23081,N_23304);
xnor U24818 (N_24818,N_22668,N_23747);
xnor U24819 (N_24819,N_23264,N_22993);
nor U24820 (N_24820,N_23699,N_23170);
or U24821 (N_24821,N_22534,N_23215);
nor U24822 (N_24822,N_23182,N_23292);
and U24823 (N_24823,N_23100,N_22876);
and U24824 (N_24824,N_22997,N_23148);
or U24825 (N_24825,N_22890,N_23330);
or U24826 (N_24826,N_23406,N_22816);
and U24827 (N_24827,N_23386,N_23721);
and U24828 (N_24828,N_23233,N_23127);
nor U24829 (N_24829,N_23613,N_23269);
nor U24830 (N_24830,N_22560,N_23744);
xnor U24831 (N_24831,N_22812,N_23468);
xor U24832 (N_24832,N_22705,N_22919);
nor U24833 (N_24833,N_23541,N_22978);
xor U24834 (N_24834,N_23115,N_23683);
xnor U24835 (N_24835,N_22907,N_23257);
or U24836 (N_24836,N_22979,N_23425);
and U24837 (N_24837,N_23047,N_23466);
and U24838 (N_24838,N_23528,N_23029);
and U24839 (N_24839,N_23237,N_23357);
and U24840 (N_24840,N_23104,N_23712);
and U24841 (N_24841,N_23274,N_22915);
and U24842 (N_24842,N_23472,N_22520);
or U24843 (N_24843,N_23629,N_23448);
xor U24844 (N_24844,N_22545,N_23691);
xnor U24845 (N_24845,N_22582,N_23383);
or U24846 (N_24846,N_23740,N_23450);
xnor U24847 (N_24847,N_22584,N_22539);
and U24848 (N_24848,N_23279,N_23215);
or U24849 (N_24849,N_23355,N_22506);
and U24850 (N_24850,N_23383,N_22937);
nand U24851 (N_24851,N_22995,N_23544);
and U24852 (N_24852,N_23006,N_22993);
and U24853 (N_24853,N_23065,N_23119);
or U24854 (N_24854,N_23334,N_23284);
xnor U24855 (N_24855,N_23628,N_23166);
nand U24856 (N_24856,N_22657,N_22874);
nand U24857 (N_24857,N_22575,N_22748);
xor U24858 (N_24858,N_23382,N_23666);
nor U24859 (N_24859,N_23545,N_23547);
or U24860 (N_24860,N_23271,N_23579);
nor U24861 (N_24861,N_23702,N_22531);
nand U24862 (N_24862,N_22848,N_23664);
nor U24863 (N_24863,N_23183,N_23651);
xnor U24864 (N_24864,N_23191,N_23154);
and U24865 (N_24865,N_22828,N_22672);
nor U24866 (N_24866,N_22652,N_22836);
nor U24867 (N_24867,N_22964,N_22744);
nor U24868 (N_24868,N_23405,N_22801);
or U24869 (N_24869,N_23140,N_23484);
and U24870 (N_24870,N_23108,N_22873);
and U24871 (N_24871,N_23015,N_23630);
nor U24872 (N_24872,N_22861,N_22571);
nor U24873 (N_24873,N_22550,N_22528);
nor U24874 (N_24874,N_23381,N_22653);
xnor U24875 (N_24875,N_22530,N_22677);
and U24876 (N_24876,N_22705,N_22921);
and U24877 (N_24877,N_22619,N_23220);
or U24878 (N_24878,N_23013,N_23745);
or U24879 (N_24879,N_22520,N_22549);
and U24880 (N_24880,N_23164,N_22961);
nand U24881 (N_24881,N_23627,N_23461);
nand U24882 (N_24882,N_23603,N_23589);
nand U24883 (N_24883,N_23692,N_23669);
and U24884 (N_24884,N_22688,N_23028);
xnor U24885 (N_24885,N_23265,N_23002);
nand U24886 (N_24886,N_23331,N_23155);
and U24887 (N_24887,N_22520,N_22692);
nor U24888 (N_24888,N_23548,N_23692);
xor U24889 (N_24889,N_22534,N_23575);
xor U24890 (N_24890,N_23247,N_23263);
or U24891 (N_24891,N_23411,N_23704);
xor U24892 (N_24892,N_23174,N_22661);
or U24893 (N_24893,N_23571,N_23454);
and U24894 (N_24894,N_23449,N_23648);
xnor U24895 (N_24895,N_22637,N_23579);
nor U24896 (N_24896,N_23702,N_22881);
nor U24897 (N_24897,N_22714,N_23153);
nand U24898 (N_24898,N_23104,N_23022);
xor U24899 (N_24899,N_22798,N_22741);
xnor U24900 (N_24900,N_23068,N_23237);
nand U24901 (N_24901,N_23021,N_23340);
xor U24902 (N_24902,N_23092,N_22857);
or U24903 (N_24903,N_22752,N_23150);
and U24904 (N_24904,N_22953,N_23294);
nor U24905 (N_24905,N_22999,N_23342);
nor U24906 (N_24906,N_23186,N_23098);
or U24907 (N_24907,N_22921,N_23732);
or U24908 (N_24908,N_23247,N_23736);
or U24909 (N_24909,N_22539,N_23160);
nand U24910 (N_24910,N_23459,N_22670);
or U24911 (N_24911,N_22792,N_22784);
xor U24912 (N_24912,N_22715,N_22950);
xnor U24913 (N_24913,N_23228,N_23693);
and U24914 (N_24914,N_23259,N_23473);
and U24915 (N_24915,N_23112,N_22657);
or U24916 (N_24916,N_23529,N_22834);
or U24917 (N_24917,N_23533,N_22825);
nor U24918 (N_24918,N_23643,N_23258);
nand U24919 (N_24919,N_22790,N_23399);
or U24920 (N_24920,N_23402,N_23074);
or U24921 (N_24921,N_22592,N_23474);
nand U24922 (N_24922,N_22519,N_22753);
or U24923 (N_24923,N_23262,N_23599);
nor U24924 (N_24924,N_22694,N_23333);
and U24925 (N_24925,N_23107,N_23434);
nand U24926 (N_24926,N_22869,N_22917);
and U24927 (N_24927,N_23439,N_23115);
and U24928 (N_24928,N_23171,N_23559);
nand U24929 (N_24929,N_23070,N_23469);
nand U24930 (N_24930,N_22677,N_23097);
or U24931 (N_24931,N_22583,N_23030);
nand U24932 (N_24932,N_23279,N_23101);
and U24933 (N_24933,N_23030,N_22690);
nand U24934 (N_24934,N_23005,N_22522);
nor U24935 (N_24935,N_23005,N_22880);
nor U24936 (N_24936,N_23062,N_22760);
xnor U24937 (N_24937,N_23380,N_22912);
xnor U24938 (N_24938,N_23175,N_23224);
and U24939 (N_24939,N_22599,N_22851);
xnor U24940 (N_24940,N_23339,N_22615);
nor U24941 (N_24941,N_23011,N_22945);
nand U24942 (N_24942,N_22796,N_23707);
nor U24943 (N_24943,N_22649,N_23211);
and U24944 (N_24944,N_23099,N_22834);
xnor U24945 (N_24945,N_22972,N_23643);
and U24946 (N_24946,N_23009,N_22995);
and U24947 (N_24947,N_23121,N_22884);
nand U24948 (N_24948,N_23596,N_23152);
xnor U24949 (N_24949,N_22726,N_23701);
and U24950 (N_24950,N_22599,N_23451);
and U24951 (N_24951,N_23439,N_22523);
or U24952 (N_24952,N_23358,N_22892);
or U24953 (N_24953,N_22781,N_23180);
or U24954 (N_24954,N_23668,N_22676);
or U24955 (N_24955,N_22857,N_23267);
nand U24956 (N_24956,N_23646,N_23247);
or U24957 (N_24957,N_23431,N_22953);
or U24958 (N_24958,N_22528,N_23518);
nor U24959 (N_24959,N_23531,N_23026);
nand U24960 (N_24960,N_23119,N_22926);
nand U24961 (N_24961,N_23510,N_23360);
or U24962 (N_24962,N_22850,N_22943);
and U24963 (N_24963,N_22778,N_22626);
nor U24964 (N_24964,N_23208,N_23006);
or U24965 (N_24965,N_22940,N_22771);
or U24966 (N_24966,N_23736,N_23376);
nor U24967 (N_24967,N_23408,N_23413);
xor U24968 (N_24968,N_23080,N_23440);
or U24969 (N_24969,N_23228,N_23376);
xor U24970 (N_24970,N_23508,N_23394);
xnor U24971 (N_24971,N_22738,N_23353);
nand U24972 (N_24972,N_23521,N_23429);
xnor U24973 (N_24973,N_23546,N_22829);
nand U24974 (N_24974,N_23188,N_23008);
nor U24975 (N_24975,N_23179,N_23332);
or U24976 (N_24976,N_22720,N_23484);
nor U24977 (N_24977,N_22648,N_23469);
or U24978 (N_24978,N_22935,N_23160);
xnor U24979 (N_24979,N_23162,N_23160);
or U24980 (N_24980,N_23634,N_23699);
or U24981 (N_24981,N_23557,N_22912);
or U24982 (N_24982,N_22918,N_23058);
xnor U24983 (N_24983,N_22571,N_23215);
or U24984 (N_24984,N_22516,N_22566);
nand U24985 (N_24985,N_23396,N_23185);
and U24986 (N_24986,N_23579,N_22750);
xnor U24987 (N_24987,N_23507,N_23073);
xor U24988 (N_24988,N_22645,N_23028);
or U24989 (N_24989,N_22964,N_23641);
nor U24990 (N_24990,N_23180,N_23468);
nor U24991 (N_24991,N_22575,N_22735);
xor U24992 (N_24992,N_23113,N_22673);
and U24993 (N_24993,N_23516,N_22564);
and U24994 (N_24994,N_23477,N_23016);
or U24995 (N_24995,N_23307,N_22833);
or U24996 (N_24996,N_23516,N_23039);
nand U24997 (N_24997,N_23604,N_23629);
nand U24998 (N_24998,N_23162,N_23738);
nor U24999 (N_24999,N_22935,N_23139);
or UO_0 (O_0,N_24581,N_24220);
and UO_1 (O_1,N_24590,N_23835);
or UO_2 (O_2,N_24108,N_23776);
nor UO_3 (O_3,N_24053,N_24875);
nand UO_4 (O_4,N_24396,N_24461);
and UO_5 (O_5,N_24724,N_24386);
xor UO_6 (O_6,N_24735,N_24229);
nor UO_7 (O_7,N_24283,N_24671);
or UO_8 (O_8,N_23912,N_24315);
or UO_9 (O_9,N_24987,N_23850);
xor UO_10 (O_10,N_24597,N_24619);
xnor UO_11 (O_11,N_23809,N_24127);
xor UO_12 (O_12,N_24453,N_24202);
xnor UO_13 (O_13,N_23784,N_24926);
xor UO_14 (O_14,N_24029,N_24321);
nor UO_15 (O_15,N_24246,N_24663);
xnor UO_16 (O_16,N_24553,N_24344);
nand UO_17 (O_17,N_23894,N_24016);
nand UO_18 (O_18,N_24943,N_23998);
nand UO_19 (O_19,N_23919,N_24244);
nand UO_20 (O_20,N_23960,N_24984);
and UO_21 (O_21,N_23796,N_24572);
or UO_22 (O_22,N_24469,N_23848);
nor UO_23 (O_23,N_24203,N_24301);
xor UO_24 (O_24,N_24523,N_23888);
nand UO_25 (O_25,N_24275,N_24534);
nor UO_26 (O_26,N_24475,N_24181);
and UO_27 (O_27,N_24041,N_23989);
nor UO_28 (O_28,N_24698,N_24187);
and UO_29 (O_29,N_24725,N_24907);
or UO_30 (O_30,N_24516,N_24669);
xnor UO_31 (O_31,N_24082,N_24675);
xnor UO_32 (O_32,N_24562,N_24682);
nor UO_33 (O_33,N_24707,N_24252);
xnor UO_34 (O_34,N_24214,N_24556);
or UO_35 (O_35,N_24720,N_24611);
nor UO_36 (O_36,N_24394,N_24487);
xor UO_37 (O_37,N_24170,N_24945);
nor UO_38 (O_38,N_24882,N_23855);
nand UO_39 (O_39,N_24741,N_23985);
nand UO_40 (O_40,N_24440,N_24470);
nor UO_41 (O_41,N_24021,N_24304);
or UO_42 (O_42,N_24319,N_24891);
xnor UO_43 (O_43,N_24134,N_24294);
and UO_44 (O_44,N_24690,N_23970);
or UO_45 (O_45,N_24790,N_24858);
xnor UO_46 (O_46,N_24555,N_23916);
and UO_47 (O_47,N_24763,N_24503);
xor UO_48 (O_48,N_24227,N_23754);
or UO_49 (O_49,N_23948,N_24019);
or UO_50 (O_50,N_24439,N_23910);
xor UO_51 (O_51,N_24193,N_23820);
or UO_52 (O_52,N_24755,N_24706);
nor UO_53 (O_53,N_23996,N_24840);
nor UO_54 (O_54,N_24867,N_23983);
nand UO_55 (O_55,N_24494,N_24471);
nor UO_56 (O_56,N_24102,N_24434);
xnor UO_57 (O_57,N_24645,N_24111);
and UO_58 (O_58,N_24346,N_24748);
nor UO_59 (O_59,N_23863,N_24038);
nor UO_60 (O_60,N_24432,N_24083);
nor UO_61 (O_61,N_24767,N_23911);
xor UO_62 (O_62,N_24226,N_23845);
xor UO_63 (O_63,N_24750,N_24316);
xnor UO_64 (O_64,N_23858,N_24222);
xnor UO_65 (O_65,N_24390,N_24240);
or UO_66 (O_66,N_23772,N_23937);
nand UO_67 (O_67,N_24531,N_24906);
xor UO_68 (O_68,N_24908,N_24343);
nor UO_69 (O_69,N_24352,N_24405);
or UO_70 (O_70,N_23774,N_23752);
nand UO_71 (O_71,N_24383,N_23775);
nand UO_72 (O_72,N_24493,N_24295);
nand UO_73 (O_73,N_24955,N_24794);
nor UO_74 (O_74,N_24802,N_23968);
nor UO_75 (O_75,N_24349,N_24191);
or UO_76 (O_76,N_23897,N_23898);
nand UO_77 (O_77,N_24586,N_24048);
nor UO_78 (O_78,N_23841,N_24095);
xnor UO_79 (O_79,N_23759,N_24753);
and UO_80 (O_80,N_23887,N_24098);
nand UO_81 (O_81,N_24093,N_24065);
nand UO_82 (O_82,N_23956,N_24124);
nor UO_83 (O_83,N_24743,N_23892);
and UO_84 (O_84,N_24365,N_24771);
or UO_85 (O_85,N_23944,N_24683);
and UO_86 (O_86,N_24911,N_24002);
or UO_87 (O_87,N_24737,N_23750);
nor UO_88 (O_88,N_24459,N_23905);
or UO_89 (O_89,N_24460,N_24190);
and UO_90 (O_90,N_24335,N_24501);
and UO_91 (O_91,N_24185,N_24915);
nor UO_92 (O_92,N_24178,N_24551);
nand UO_93 (O_93,N_24277,N_23864);
and UO_94 (O_94,N_24885,N_24371);
xnor UO_95 (O_95,N_24435,N_24017);
nand UO_96 (O_96,N_24670,N_23756);
or UO_97 (O_97,N_24705,N_24600);
nand UO_98 (O_98,N_24922,N_23765);
xor UO_99 (O_99,N_24580,N_24001);
nor UO_100 (O_100,N_23795,N_24476);
nor UO_101 (O_101,N_24243,N_23908);
and UO_102 (O_102,N_24860,N_24280);
nor UO_103 (O_103,N_24901,N_24883);
and UO_104 (O_104,N_24554,N_24601);
nand UO_105 (O_105,N_24101,N_23943);
and UO_106 (O_106,N_23813,N_23881);
nor UO_107 (O_107,N_24798,N_24629);
and UO_108 (O_108,N_24261,N_24426);
or UO_109 (O_109,N_24161,N_24954);
or UO_110 (O_110,N_24122,N_24746);
and UO_111 (O_111,N_24828,N_24379);
and UO_112 (O_112,N_24895,N_24980);
nand UO_113 (O_113,N_24579,N_24135);
nand UO_114 (O_114,N_24338,N_24512);
xnor UO_115 (O_115,N_24188,N_24960);
or UO_116 (O_116,N_24307,N_24993);
or UO_117 (O_117,N_24722,N_24931);
and UO_118 (O_118,N_24511,N_24859);
xor UO_119 (O_119,N_24543,N_24966);
nand UO_120 (O_120,N_24995,N_24286);
or UO_121 (O_121,N_24637,N_23758);
or UO_122 (O_122,N_24873,N_23836);
and UO_123 (O_123,N_24267,N_24620);
or UO_124 (O_124,N_24458,N_24529);
nor UO_125 (O_125,N_24868,N_23868);
nor UO_126 (O_126,N_23933,N_24429);
nand UO_127 (O_127,N_24231,N_24423);
nand UO_128 (O_128,N_24800,N_24538);
or UO_129 (O_129,N_24367,N_24042);
xor UO_130 (O_130,N_24912,N_24414);
nand UO_131 (O_131,N_24677,N_24944);
nand UO_132 (O_132,N_24018,N_23926);
or UO_133 (O_133,N_23965,N_24078);
and UO_134 (O_134,N_24342,N_24696);
xnor UO_135 (O_135,N_24413,N_23900);
xnor UO_136 (O_136,N_23871,N_24605);
and UO_137 (O_137,N_23769,N_24213);
nand UO_138 (O_138,N_24140,N_24415);
and UO_139 (O_139,N_24025,N_24160);
or UO_140 (O_140,N_23992,N_24096);
xnor UO_141 (O_141,N_24730,N_24035);
and UO_142 (O_142,N_24479,N_23969);
and UO_143 (O_143,N_24333,N_24902);
xor UO_144 (O_144,N_24350,N_24905);
and UO_145 (O_145,N_24330,N_24633);
and UO_146 (O_146,N_24667,N_23798);
or UO_147 (O_147,N_24255,N_23870);
nand UO_148 (O_148,N_24162,N_24010);
nor UO_149 (O_149,N_24810,N_23928);
or UO_150 (O_150,N_24211,N_24951);
xnor UO_151 (O_151,N_24574,N_24589);
xnor UO_152 (O_152,N_24146,N_24805);
nor UO_153 (O_153,N_24120,N_23904);
nand UO_154 (O_154,N_24417,N_24376);
nor UO_155 (O_155,N_24686,N_24988);
nand UO_156 (O_156,N_24657,N_24583);
and UO_157 (O_157,N_24540,N_24732);
or UO_158 (O_158,N_24985,N_24389);
or UO_159 (O_159,N_24477,N_24994);
nor UO_160 (O_160,N_24353,N_24929);
xnor UO_161 (O_161,N_24497,N_24269);
or UO_162 (O_162,N_23935,N_24786);
nor UO_163 (O_163,N_24892,N_23982);
and UO_164 (O_164,N_24197,N_24808);
nor UO_165 (O_165,N_24351,N_24692);
nor UO_166 (O_166,N_24688,N_24979);
xnor UO_167 (O_167,N_24004,N_24697);
nand UO_168 (O_168,N_24143,N_24391);
xor UO_169 (O_169,N_23815,N_23915);
and UO_170 (O_170,N_23846,N_23947);
and UO_171 (O_171,N_24466,N_24846);
and UO_172 (O_172,N_24525,N_23893);
or UO_173 (O_173,N_24648,N_23976);
xor UO_174 (O_174,N_24145,N_24762);
and UO_175 (O_175,N_24627,N_23924);
nand UO_176 (O_176,N_24395,N_23847);
or UO_177 (O_177,N_24625,N_24862);
xor UO_178 (O_178,N_24151,N_24207);
and UO_179 (O_179,N_24409,N_23839);
or UO_180 (O_180,N_24842,N_24863);
or UO_181 (O_181,N_24115,N_24630);
and UO_182 (O_182,N_24714,N_23791);
nor UO_183 (O_183,N_24660,N_23907);
nor UO_184 (O_184,N_24799,N_24643);
xor UO_185 (O_185,N_23901,N_24681);
xor UO_186 (O_186,N_23945,N_24431);
nor UO_187 (O_187,N_24199,N_23869);
nand UO_188 (O_188,N_24463,N_23966);
xor UO_189 (O_189,N_24997,N_24265);
nor UO_190 (O_190,N_24871,N_24087);
and UO_191 (O_191,N_23961,N_24264);
nand UO_192 (O_192,N_24530,N_24289);
and UO_193 (O_193,N_24050,N_24173);
or UO_194 (O_194,N_24180,N_23762);
xor UO_195 (O_195,N_23806,N_24587);
or UO_196 (O_196,N_24266,N_24573);
or UO_197 (O_197,N_24034,N_23934);
xnor UO_198 (O_198,N_24056,N_24872);
nand UO_199 (O_199,N_24628,N_23891);
or UO_200 (O_200,N_24839,N_24372);
xor UO_201 (O_201,N_24152,N_23941);
and UO_202 (O_202,N_24772,N_24704);
nand UO_203 (O_203,N_24793,N_24869);
or UO_204 (O_204,N_24399,N_24826);
or UO_205 (O_205,N_24816,N_24595);
nor UO_206 (O_206,N_24804,N_24285);
or UO_207 (O_207,N_24259,N_24088);
or UO_208 (O_208,N_24938,N_24451);
nor UO_209 (O_209,N_24662,N_24974);
nor UO_210 (O_210,N_24847,N_24789);
or UO_211 (O_211,N_24069,N_23753);
nor UO_212 (O_212,N_23826,N_24299);
and UO_213 (O_213,N_24615,N_24402);
nor UO_214 (O_214,N_24225,N_24401);
nand UO_215 (O_215,N_24761,N_24518);
and UO_216 (O_216,N_24559,N_23854);
xor UO_217 (O_217,N_24206,N_24565);
nor UO_218 (O_218,N_24989,N_23882);
and UO_219 (O_219,N_24110,N_23792);
and UO_220 (O_220,N_24811,N_24485);
nor UO_221 (O_221,N_24421,N_24099);
and UO_222 (O_222,N_24712,N_23914);
xnor UO_223 (O_223,N_24976,N_24358);
or UO_224 (O_224,N_24654,N_24602);
nor UO_225 (O_225,N_24544,N_24052);
and UO_226 (O_226,N_24936,N_23957);
nand UO_227 (O_227,N_24599,N_24448);
or UO_228 (O_228,N_24273,N_24526);
nand UO_229 (O_229,N_24000,N_24205);
nor UO_230 (O_230,N_23991,N_24355);
and UO_231 (O_231,N_24136,N_24903);
nand UO_232 (O_232,N_23838,N_24950);
nand UO_233 (O_233,N_24673,N_23940);
or UO_234 (O_234,N_23866,N_24764);
or UO_235 (O_235,N_24070,N_24201);
or UO_236 (O_236,N_24801,N_24830);
xnor UO_237 (O_237,N_24123,N_24570);
and UO_238 (O_238,N_24369,N_24506);
or UO_239 (O_239,N_23840,N_24332);
nand UO_240 (O_240,N_24884,N_24022);
or UO_241 (O_241,N_24303,N_24887);
nand UO_242 (O_242,N_24480,N_23949);
nand UO_243 (O_243,N_23874,N_24779);
or UO_244 (O_244,N_24024,N_24566);
or UO_245 (O_245,N_23797,N_24658);
nor UO_246 (O_246,N_24596,N_24496);
nor UO_247 (O_247,N_24807,N_23860);
xnor UO_248 (O_248,N_24484,N_24392);
nand UO_249 (O_249,N_24086,N_24129);
nor UO_250 (O_250,N_23981,N_24064);
xor UO_251 (O_251,N_24591,N_24293);
and UO_252 (O_252,N_23959,N_24612);
nand UO_253 (O_253,N_24011,N_24900);
xnor UO_254 (O_254,N_23853,N_24442);
and UO_255 (O_255,N_24788,N_24715);
or UO_256 (O_256,N_23946,N_24861);
xnor UO_257 (O_257,N_24169,N_24505);
nor UO_258 (O_258,N_24744,N_24624);
nand UO_259 (O_259,N_24614,N_24569);
xnor UO_260 (O_260,N_23865,N_24568);
nor UO_261 (O_261,N_24292,N_24040);
xnor UO_262 (O_262,N_24059,N_24416);
nand UO_263 (O_263,N_24138,N_24878);
nor UO_264 (O_264,N_24502,N_24796);
nor UO_265 (O_265,N_24783,N_24106);
or UO_266 (O_266,N_23827,N_24456);
and UO_267 (O_267,N_24068,N_24340);
xor UO_268 (O_268,N_24306,N_23942);
nand UO_269 (O_269,N_24661,N_24242);
or UO_270 (O_270,N_23984,N_24928);
or UO_271 (O_271,N_24679,N_24258);
nand UO_272 (O_272,N_24850,N_23780);
nand UO_273 (O_273,N_24282,N_23975);
xnor UO_274 (O_274,N_24621,N_24921);
xnor UO_275 (O_275,N_24917,N_24067);
or UO_276 (O_276,N_24787,N_24713);
and UO_277 (O_277,N_24952,N_24418);
xnor UO_278 (O_278,N_24100,N_24881);
and UO_279 (O_279,N_23917,N_23902);
nor UO_280 (O_280,N_24888,N_24403);
nor UO_281 (O_281,N_24118,N_24279);
or UO_282 (O_282,N_24009,N_24632);
or UO_283 (O_283,N_24532,N_24927);
or UO_284 (O_284,N_24689,N_24184);
nand UO_285 (O_285,N_23921,N_24128);
xnor UO_286 (O_286,N_24665,N_23972);
or UO_287 (O_287,N_24825,N_23955);
nor UO_288 (O_288,N_24150,N_24381);
xor UO_289 (O_289,N_24091,N_24158);
and UO_290 (O_290,N_24548,N_24736);
and UO_291 (O_291,N_24345,N_24462);
or UO_292 (O_292,N_23997,N_24608);
and UO_293 (O_293,N_23883,N_24163);
nor UO_294 (O_294,N_24819,N_24754);
nand UO_295 (O_295,N_24969,N_24121);
xnor UO_296 (O_296,N_24939,N_24849);
nand UO_297 (O_297,N_24147,N_23849);
and UO_298 (O_298,N_24020,N_24514);
nand UO_299 (O_299,N_24238,N_24896);
nor UO_300 (O_300,N_23755,N_23830);
or UO_301 (O_301,N_24323,N_23990);
nor UO_302 (O_302,N_23785,N_24576);
nand UO_303 (O_303,N_24433,N_24412);
xor UO_304 (O_304,N_24420,N_24879);
nor UO_305 (O_305,N_24045,N_24820);
xor UO_306 (O_306,N_23950,N_24320);
nor UO_307 (O_307,N_24864,N_24959);
nand UO_308 (O_308,N_24428,N_24194);
or UO_309 (O_309,N_24622,N_23811);
and UO_310 (O_310,N_24427,N_24649);
xor UO_311 (O_311,N_24057,N_24215);
nand UO_312 (O_312,N_23890,N_24302);
nor UO_313 (O_313,N_24674,N_24618);
or UO_314 (O_314,N_24444,N_24899);
xnor UO_315 (O_315,N_24836,N_24835);
xnor UO_316 (O_316,N_23922,N_24613);
xor UO_317 (O_317,N_24972,N_24560);
nor UO_318 (O_318,N_24012,N_24854);
and UO_319 (O_319,N_24026,N_24103);
and UO_320 (O_320,N_24313,N_24827);
or UO_321 (O_321,N_24924,N_24256);
and UO_322 (O_322,N_24005,N_24079);
nor UO_323 (O_323,N_24198,N_24141);
nand UO_324 (O_324,N_24874,N_24233);
or UO_325 (O_325,N_23777,N_24920);
or UO_326 (O_326,N_24982,N_24992);
and UO_327 (O_327,N_24521,N_24008);
or UO_328 (O_328,N_24584,N_24308);
and UO_329 (O_329,N_24015,N_24217);
and UO_330 (O_330,N_23903,N_24054);
nor UO_331 (O_331,N_24894,N_24708);
or UO_332 (O_332,N_24216,N_24710);
nand UO_333 (O_333,N_24189,N_24116);
xor UO_334 (O_334,N_23843,N_24653);
or UO_335 (O_335,N_24691,N_24953);
xnor UO_336 (O_336,N_24311,N_24112);
or UO_337 (O_337,N_24155,N_24314);
or UO_338 (O_338,N_24288,N_24564);
nand UO_339 (O_339,N_24780,N_24765);
nor UO_340 (O_340,N_24609,N_23927);
or UO_341 (O_341,N_24739,N_24652);
nor UO_342 (O_342,N_24478,N_24200);
or UO_343 (O_343,N_24999,N_24575);
or UO_344 (O_344,N_24366,N_24368);
or UO_345 (O_345,N_24131,N_24774);
nor UO_346 (O_346,N_24133,N_24577);
and UO_347 (O_347,N_24228,N_24236);
nand UO_348 (O_348,N_24550,N_23931);
nand UO_349 (O_349,N_24886,N_24348);
nand UO_350 (O_350,N_24373,N_24235);
nor UO_351 (O_351,N_24925,N_24781);
xor UO_352 (O_352,N_24676,N_24910);
xnor UO_353 (O_353,N_23779,N_23763);
nor UO_354 (O_354,N_24137,N_24322);
nor UO_355 (O_355,N_24492,N_24515);
nor UO_356 (O_356,N_24659,N_24341);
nand UO_357 (O_357,N_24183,N_24062);
nor UO_358 (O_358,N_23793,N_23973);
or UO_359 (O_359,N_24766,N_24378);
or UO_360 (O_360,N_24784,N_23923);
xor UO_361 (O_361,N_23925,N_24468);
xnor UO_362 (O_362,N_24327,N_24937);
nor UO_363 (O_363,N_23978,N_24474);
xor UO_364 (O_364,N_24071,N_24646);
xor UO_365 (O_365,N_24196,N_24347);
and UO_366 (O_366,N_23958,N_24388);
nand UO_367 (O_367,N_24125,N_24339);
nand UO_368 (O_368,N_24186,N_24318);
xor UO_369 (O_369,N_24734,N_23884);
xnor UO_370 (O_370,N_24664,N_24549);
or UO_371 (O_371,N_24809,N_24935);
nor UO_372 (O_372,N_24370,N_24909);
or UO_373 (O_373,N_24080,N_24606);
and UO_374 (O_374,N_23929,N_24791);
nor UO_375 (O_375,N_24006,N_24360);
nor UO_376 (O_376,N_24387,N_24723);
nor UO_377 (O_377,N_24507,N_23909);
or UO_378 (O_378,N_24305,N_23880);
and UO_379 (O_379,N_24221,N_23856);
and UO_380 (O_380,N_24411,N_24234);
or UO_381 (O_381,N_24962,N_24876);
and UO_382 (O_382,N_23987,N_23862);
xor UO_383 (O_383,N_24375,N_24357);
or UO_384 (O_384,N_24964,N_24384);
nor UO_385 (O_385,N_24159,N_24751);
xor UO_386 (O_386,N_23993,N_24956);
xnor UO_387 (O_387,N_24144,N_24393);
and UO_388 (O_388,N_24167,N_24239);
nor UO_389 (O_389,N_24212,N_24241);
nor UO_390 (O_390,N_24776,N_24117);
xnor UO_391 (O_391,N_24483,N_24445);
nand UO_392 (O_392,N_24536,N_24806);
and UO_393 (O_393,N_24527,N_24272);
nand UO_394 (O_394,N_24329,N_24044);
or UO_395 (O_395,N_24558,N_24449);
nor UO_396 (O_396,N_24934,N_24407);
xnor UO_397 (O_397,N_23768,N_24014);
nand UO_398 (O_398,N_24635,N_24795);
or UO_399 (O_399,N_24870,N_24422);
xor UO_400 (O_400,N_24647,N_24097);
and UO_401 (O_401,N_24594,N_24524);
and UO_402 (O_402,N_24182,N_24711);
xnor UO_403 (O_403,N_24636,N_24967);
or UO_404 (O_404,N_24957,N_24821);
xnor UO_405 (O_405,N_23788,N_23913);
xnor UO_406 (O_406,N_24380,N_24727);
nand UO_407 (O_407,N_24274,N_24824);
xor UO_408 (O_408,N_23807,N_24153);
or UO_409 (O_409,N_24400,N_24398);
nand UO_410 (O_410,N_23879,N_23767);
or UO_411 (O_411,N_24678,N_24814);
nor UO_412 (O_412,N_23770,N_23810);
nand UO_413 (O_413,N_24728,N_24604);
or UO_414 (O_414,N_24312,N_24760);
or UO_415 (O_415,N_23787,N_24996);
xor UO_416 (O_416,N_23971,N_24965);
xor UO_417 (O_417,N_23936,N_24176);
nor UO_418 (O_418,N_24437,N_23802);
and UO_419 (O_419,N_24317,N_23930);
nor UO_420 (O_420,N_23764,N_23781);
xor UO_421 (O_421,N_23805,N_24651);
and UO_422 (O_422,N_24165,N_24049);
xor UO_423 (O_423,N_24641,N_24537);
nand UO_424 (O_424,N_23979,N_24813);
nor UO_425 (O_425,N_24857,N_24094);
or UO_426 (O_426,N_24192,N_24567);
and UO_427 (O_427,N_23873,N_23877);
nor UO_428 (O_428,N_24687,N_24616);
nor UO_429 (O_429,N_24585,N_23821);
nand UO_430 (O_430,N_24509,N_24918);
xor UO_431 (O_431,N_24785,N_24610);
xor UO_432 (O_432,N_24223,N_24547);
nor UO_433 (O_433,N_24948,N_24076);
nor UO_434 (O_434,N_23828,N_24893);
xor UO_435 (O_435,N_23896,N_24592);
or UO_436 (O_436,N_24464,N_23932);
or UO_437 (O_437,N_24204,N_24336);
and UO_438 (O_438,N_24709,N_24060);
nand UO_439 (O_439,N_24946,N_24702);
and UO_440 (O_440,N_23844,N_24047);
or UO_441 (O_441,N_23872,N_24061);
nor UO_442 (O_442,N_23977,N_23967);
nor UO_443 (O_443,N_24263,N_24623);
or UO_444 (O_444,N_24541,N_24446);
and UO_445 (O_445,N_24114,N_24703);
and UO_446 (O_446,N_24844,N_24406);
or UO_447 (O_447,N_24013,N_24377);
or UO_448 (O_448,N_24598,N_24084);
or UO_449 (O_449,N_24631,N_24561);
and UO_450 (O_450,N_24656,N_24300);
nor UO_451 (O_451,N_23804,N_24495);
xnor UO_452 (O_452,N_24769,N_23801);
nor UO_453 (O_453,N_23875,N_24270);
xor UO_454 (O_454,N_23808,N_24841);
nor UO_455 (O_455,N_23818,N_24374);
nand UO_456 (O_456,N_24963,N_24650);
and UO_457 (O_457,N_24833,N_24104);
nor UO_458 (O_458,N_24454,N_23766);
or UO_459 (O_459,N_24699,N_24626);
xor UO_460 (O_460,N_24970,N_24749);
nand UO_461 (O_461,N_24975,N_24362);
xnor UO_462 (O_462,N_24171,N_24856);
xnor UO_463 (O_463,N_24430,N_24499);
or UO_464 (O_464,N_24419,N_23895);
nor UO_465 (O_465,N_24981,N_24037);
xnor UO_466 (O_466,N_24919,N_24668);
or UO_467 (O_467,N_24890,N_23812);
and UO_468 (O_468,N_23790,N_24172);
nor UO_469 (O_469,N_23771,N_24074);
nor UO_470 (O_470,N_24382,N_24473);
and UO_471 (O_471,N_23823,N_24498);
xor UO_472 (O_472,N_24866,N_23899);
or UO_473 (O_473,N_24157,N_24467);
nand UO_474 (O_474,N_24324,N_24331);
and UO_475 (O_475,N_24156,N_23952);
or UO_476 (O_476,N_24166,N_23906);
nor UO_477 (O_477,N_24582,N_24768);
nor UO_478 (O_478,N_24260,N_23786);
xor UO_479 (O_479,N_24639,N_24533);
xnor UO_480 (O_480,N_24109,N_24508);
or UO_481 (O_481,N_24481,N_24218);
nor UO_482 (O_482,N_24593,N_24491);
or UO_483 (O_483,N_24224,N_24356);
and UO_484 (O_484,N_24758,N_24897);
nor UO_485 (O_485,N_24528,N_23876);
and UO_486 (O_486,N_24364,N_24672);
nor UO_487 (O_487,N_24880,N_24923);
nor UO_488 (O_488,N_24113,N_23834);
nand UO_489 (O_489,N_24230,N_24043);
nor UO_490 (O_490,N_24803,N_24254);
nor UO_491 (O_491,N_24797,N_24535);
and UO_492 (O_492,N_23859,N_23939);
xnor UO_493 (O_493,N_23886,N_23800);
xor UO_494 (O_494,N_24142,N_24644);
and UO_495 (O_495,N_23938,N_23878);
or UO_496 (O_496,N_24865,N_24326);
or UO_497 (O_497,N_24334,N_24425);
or UO_498 (O_498,N_23988,N_24291);
nor UO_499 (O_499,N_24742,N_24852);
nor UO_500 (O_500,N_24695,N_24055);
or UO_501 (O_501,N_23783,N_24132);
nand UO_502 (O_502,N_24253,N_24759);
nand UO_503 (O_503,N_24666,N_24085);
or UO_504 (O_504,N_24490,N_24913);
xnor UO_505 (O_505,N_24232,N_24757);
and UO_506 (O_506,N_24838,N_24031);
nor UO_507 (O_507,N_24361,N_24328);
and UO_508 (O_508,N_24843,N_23964);
xnor UO_509 (O_509,N_24046,N_24770);
xor UO_510 (O_510,N_23920,N_24916);
xnor UO_511 (O_511,N_23974,N_24310);
xnor UO_512 (O_512,N_24978,N_24904);
nor UO_513 (O_513,N_24832,N_24773);
xnor UO_514 (O_514,N_23842,N_24853);
and UO_515 (O_515,N_23953,N_24410);
nor UO_516 (O_516,N_24063,N_24778);
or UO_517 (O_517,N_24877,N_24139);
nand UO_518 (O_518,N_24486,N_24268);
or UO_519 (O_519,N_24717,N_24397);
or UO_520 (O_520,N_24424,N_24296);
nor UO_521 (O_521,N_24195,N_24251);
and UO_522 (O_522,N_24914,N_24539);
nor UO_523 (O_523,N_24489,N_24028);
nand UO_524 (O_524,N_24731,N_24278);
nor UO_525 (O_525,N_23773,N_23819);
nand UO_526 (O_526,N_24845,N_24066);
nand UO_527 (O_527,N_24090,N_24947);
and UO_528 (O_528,N_24039,N_24716);
or UO_529 (O_529,N_24510,N_23799);
or UO_530 (O_530,N_24089,N_23918);
and UO_531 (O_531,N_24700,N_24822);
nand UO_532 (O_532,N_24107,N_24968);
and UO_533 (O_533,N_23803,N_23829);
nand UO_534 (O_534,N_24298,N_24655);
and UO_535 (O_535,N_24823,N_24262);
or UO_536 (O_536,N_24745,N_24949);
xor UO_537 (O_537,N_23951,N_24848);
or UO_538 (O_538,N_24775,N_24325);
and UO_539 (O_539,N_24023,N_24247);
xor UO_540 (O_540,N_24290,N_24179);
xor UO_541 (O_541,N_23889,N_23760);
and UO_542 (O_542,N_24718,N_24105);
or UO_543 (O_543,N_23857,N_24812);
nor UO_544 (O_544,N_23817,N_24961);
xnor UO_545 (O_545,N_23962,N_24007);
nor UO_546 (O_546,N_24752,N_23824);
and UO_547 (O_547,N_24032,N_23831);
xnor UO_548 (O_548,N_24003,N_23751);
xnor UO_549 (O_549,N_24815,N_24973);
xnor UO_550 (O_550,N_24058,N_24245);
or UO_551 (O_551,N_24685,N_24175);
and UO_552 (O_552,N_24942,N_24237);
nand UO_553 (O_553,N_23822,N_24287);
or UO_554 (O_554,N_24488,N_24617);
nand UO_555 (O_555,N_23814,N_23995);
and UO_556 (O_556,N_24588,N_24557);
nor UO_557 (O_557,N_24309,N_23816);
nor UO_558 (O_558,N_24354,N_24036);
and UO_559 (O_559,N_24051,N_23794);
and UO_560 (O_560,N_24634,N_24740);
and UO_561 (O_561,N_24208,N_24075);
or UO_562 (O_562,N_23994,N_24404);
xor UO_563 (O_563,N_24033,N_24831);
and UO_564 (O_564,N_24990,N_24281);
nor UO_565 (O_565,N_24542,N_24834);
and UO_566 (O_566,N_24472,N_24276);
and UO_567 (O_567,N_24729,N_23999);
or UO_568 (O_568,N_24563,N_23778);
and UO_569 (O_569,N_24148,N_24738);
nor UO_570 (O_570,N_24337,N_24719);
nor UO_571 (O_571,N_24504,N_24126);
xnor UO_572 (O_572,N_24998,N_24248);
and UO_573 (O_573,N_24500,N_23761);
nand UO_574 (O_574,N_24219,N_24694);
xor UO_575 (O_575,N_23837,N_24271);
nand UO_576 (O_576,N_24027,N_24701);
nand UO_577 (O_577,N_24482,N_24941);
nand UO_578 (O_578,N_24257,N_24436);
xor UO_579 (O_579,N_24450,N_24408);
nand UO_580 (O_580,N_24385,N_24081);
nor UO_581 (O_581,N_24520,N_24452);
nand UO_582 (O_582,N_24930,N_24513);
nor UO_583 (O_583,N_24855,N_24817);
nand UO_584 (O_584,N_24940,N_23986);
and UO_585 (O_585,N_24363,N_24607);
xor UO_586 (O_586,N_24933,N_24829);
and UO_587 (O_587,N_24932,N_24721);
xnor UO_588 (O_588,N_24837,N_24792);
nor UO_589 (O_589,N_24986,N_24571);
xor UO_590 (O_590,N_24851,N_24603);
xnor UO_591 (O_591,N_24818,N_24777);
or UO_592 (O_592,N_23782,N_24073);
xor UO_593 (O_593,N_24578,N_24072);
and UO_594 (O_594,N_24210,N_24522);
nor UO_595 (O_595,N_24457,N_24640);
and UO_596 (O_596,N_23789,N_23833);
nand UO_597 (O_597,N_24164,N_24438);
and UO_598 (O_598,N_23867,N_24177);
nor UO_599 (O_599,N_24154,N_24638);
nor UO_600 (O_600,N_24545,N_24756);
nor UO_601 (O_601,N_24174,N_23963);
xnor UO_602 (O_602,N_24130,N_24250);
or UO_603 (O_603,N_24726,N_24782);
and UO_604 (O_604,N_24284,N_24359);
xnor UO_605 (O_605,N_23885,N_24983);
xor UO_606 (O_606,N_24747,N_24168);
nor UO_607 (O_607,N_24733,N_24077);
or UO_608 (O_608,N_23861,N_24447);
nand UO_609 (O_609,N_24898,N_24552);
and UO_610 (O_610,N_23832,N_23852);
nor UO_611 (O_611,N_24519,N_24680);
and UO_612 (O_612,N_24209,N_24297);
xnor UO_613 (O_613,N_24465,N_23851);
xnor UO_614 (O_614,N_23954,N_23980);
or UO_615 (O_615,N_24684,N_24149);
xor UO_616 (O_616,N_24958,N_24119);
nand UO_617 (O_617,N_24455,N_24441);
and UO_618 (O_618,N_24546,N_24030);
and UO_619 (O_619,N_24517,N_23757);
nand UO_620 (O_620,N_24971,N_24642);
nand UO_621 (O_621,N_24092,N_24443);
xnor UO_622 (O_622,N_23825,N_24249);
nand UO_623 (O_623,N_24977,N_24991);
nor UO_624 (O_624,N_24889,N_24693);
nor UO_625 (O_625,N_24977,N_24219);
nor UO_626 (O_626,N_24276,N_24194);
and UO_627 (O_627,N_23976,N_24205);
xor UO_628 (O_628,N_24413,N_24074);
or UO_629 (O_629,N_24012,N_24019);
nor UO_630 (O_630,N_24899,N_24605);
xor UO_631 (O_631,N_24914,N_24503);
xor UO_632 (O_632,N_24638,N_24003);
or UO_633 (O_633,N_24665,N_24709);
nor UO_634 (O_634,N_24197,N_24636);
and UO_635 (O_635,N_24914,N_24302);
or UO_636 (O_636,N_24312,N_24823);
and UO_637 (O_637,N_24176,N_23847);
and UO_638 (O_638,N_24095,N_23972);
nor UO_639 (O_639,N_24113,N_24432);
nor UO_640 (O_640,N_23835,N_24195);
nor UO_641 (O_641,N_24305,N_24011);
or UO_642 (O_642,N_24571,N_23777);
or UO_643 (O_643,N_24307,N_24539);
nor UO_644 (O_644,N_24102,N_23902);
or UO_645 (O_645,N_24294,N_24127);
xnor UO_646 (O_646,N_24929,N_24149);
and UO_647 (O_647,N_24426,N_23889);
and UO_648 (O_648,N_23783,N_24581);
or UO_649 (O_649,N_24275,N_24771);
nand UO_650 (O_650,N_24688,N_24818);
or UO_651 (O_651,N_24874,N_24057);
xor UO_652 (O_652,N_24446,N_24883);
and UO_653 (O_653,N_24374,N_24640);
nor UO_654 (O_654,N_24297,N_23813);
nor UO_655 (O_655,N_24233,N_24577);
nand UO_656 (O_656,N_24825,N_24602);
nand UO_657 (O_657,N_24052,N_24726);
or UO_658 (O_658,N_24037,N_24463);
and UO_659 (O_659,N_24502,N_24379);
and UO_660 (O_660,N_23882,N_24199);
nor UO_661 (O_661,N_24261,N_24021);
and UO_662 (O_662,N_24814,N_24670);
and UO_663 (O_663,N_24863,N_23787);
or UO_664 (O_664,N_24276,N_24637);
nor UO_665 (O_665,N_23835,N_23980);
and UO_666 (O_666,N_24386,N_24882);
nor UO_667 (O_667,N_23787,N_24459);
nand UO_668 (O_668,N_24383,N_24256);
and UO_669 (O_669,N_23905,N_24443);
nor UO_670 (O_670,N_24621,N_24686);
xor UO_671 (O_671,N_24802,N_24873);
or UO_672 (O_672,N_23796,N_24215);
xor UO_673 (O_673,N_24856,N_24121);
xor UO_674 (O_674,N_24212,N_24149);
nand UO_675 (O_675,N_24309,N_24357);
xor UO_676 (O_676,N_24939,N_23790);
nor UO_677 (O_677,N_24527,N_24332);
xor UO_678 (O_678,N_24294,N_24378);
nor UO_679 (O_679,N_24836,N_24971);
or UO_680 (O_680,N_24228,N_24687);
or UO_681 (O_681,N_23984,N_24121);
and UO_682 (O_682,N_24617,N_23981);
and UO_683 (O_683,N_23795,N_24507);
xnor UO_684 (O_684,N_24827,N_24360);
nand UO_685 (O_685,N_24930,N_24582);
nand UO_686 (O_686,N_24081,N_23919);
xor UO_687 (O_687,N_24902,N_24193);
nor UO_688 (O_688,N_23866,N_24134);
xnor UO_689 (O_689,N_23981,N_23755);
nor UO_690 (O_690,N_23794,N_24483);
and UO_691 (O_691,N_24046,N_24303);
nor UO_692 (O_692,N_24442,N_24226);
and UO_693 (O_693,N_24859,N_24470);
nor UO_694 (O_694,N_24427,N_24678);
or UO_695 (O_695,N_24561,N_24266);
and UO_696 (O_696,N_24605,N_24327);
or UO_697 (O_697,N_24681,N_24989);
or UO_698 (O_698,N_23866,N_24515);
or UO_699 (O_699,N_24990,N_24063);
nand UO_700 (O_700,N_24084,N_24099);
nor UO_701 (O_701,N_24479,N_23928);
and UO_702 (O_702,N_24609,N_24055);
xor UO_703 (O_703,N_23886,N_24917);
nor UO_704 (O_704,N_24241,N_23984);
xor UO_705 (O_705,N_24112,N_24751);
xnor UO_706 (O_706,N_24885,N_24625);
nor UO_707 (O_707,N_24021,N_24563);
or UO_708 (O_708,N_24675,N_24628);
and UO_709 (O_709,N_24962,N_24030);
or UO_710 (O_710,N_23848,N_23867);
nand UO_711 (O_711,N_24833,N_24054);
nand UO_712 (O_712,N_24375,N_24898);
and UO_713 (O_713,N_24284,N_24595);
or UO_714 (O_714,N_24161,N_24525);
or UO_715 (O_715,N_23853,N_24753);
nor UO_716 (O_716,N_24098,N_24845);
or UO_717 (O_717,N_24991,N_24387);
or UO_718 (O_718,N_24518,N_23786);
xnor UO_719 (O_719,N_24069,N_24098);
or UO_720 (O_720,N_24976,N_23847);
nor UO_721 (O_721,N_24056,N_24236);
and UO_722 (O_722,N_24042,N_24085);
and UO_723 (O_723,N_24826,N_24248);
or UO_724 (O_724,N_24395,N_23871);
nand UO_725 (O_725,N_24309,N_24340);
nand UO_726 (O_726,N_24414,N_24141);
or UO_727 (O_727,N_24951,N_24138);
nor UO_728 (O_728,N_24835,N_23915);
nor UO_729 (O_729,N_24767,N_24808);
or UO_730 (O_730,N_24259,N_24176);
nand UO_731 (O_731,N_24358,N_23986);
or UO_732 (O_732,N_24415,N_24724);
and UO_733 (O_733,N_24402,N_24094);
nand UO_734 (O_734,N_23762,N_24471);
xor UO_735 (O_735,N_24466,N_23802);
xor UO_736 (O_736,N_24871,N_24103);
nand UO_737 (O_737,N_24208,N_24685);
and UO_738 (O_738,N_24279,N_24850);
or UO_739 (O_739,N_24193,N_24637);
nor UO_740 (O_740,N_24700,N_24134);
nand UO_741 (O_741,N_24754,N_24818);
nand UO_742 (O_742,N_24432,N_23780);
nand UO_743 (O_743,N_23782,N_23912);
xor UO_744 (O_744,N_24385,N_24105);
or UO_745 (O_745,N_24826,N_24535);
or UO_746 (O_746,N_24333,N_24074);
nand UO_747 (O_747,N_24404,N_24551);
or UO_748 (O_748,N_23784,N_24214);
or UO_749 (O_749,N_24656,N_24827);
xnor UO_750 (O_750,N_24535,N_24381);
nand UO_751 (O_751,N_24613,N_23811);
nor UO_752 (O_752,N_24876,N_24911);
nand UO_753 (O_753,N_24758,N_24318);
and UO_754 (O_754,N_24019,N_23853);
xor UO_755 (O_755,N_24959,N_23815);
and UO_756 (O_756,N_24168,N_24401);
xor UO_757 (O_757,N_24130,N_24035);
nor UO_758 (O_758,N_24313,N_24242);
and UO_759 (O_759,N_24683,N_24676);
nor UO_760 (O_760,N_24089,N_24387);
nor UO_761 (O_761,N_24419,N_24685);
and UO_762 (O_762,N_24179,N_24905);
or UO_763 (O_763,N_24443,N_24743);
nor UO_764 (O_764,N_24305,N_24277);
xor UO_765 (O_765,N_24811,N_24673);
and UO_766 (O_766,N_24435,N_24483);
or UO_767 (O_767,N_23881,N_24145);
xnor UO_768 (O_768,N_24798,N_24352);
nand UO_769 (O_769,N_24309,N_24183);
xnor UO_770 (O_770,N_24855,N_24020);
or UO_771 (O_771,N_24070,N_24223);
xor UO_772 (O_772,N_24484,N_24846);
xor UO_773 (O_773,N_24673,N_24039);
and UO_774 (O_774,N_23943,N_24994);
xor UO_775 (O_775,N_24992,N_24728);
xnor UO_776 (O_776,N_23872,N_24014);
xor UO_777 (O_777,N_24582,N_24879);
and UO_778 (O_778,N_23968,N_23952);
or UO_779 (O_779,N_24846,N_24639);
xnor UO_780 (O_780,N_24190,N_24896);
or UO_781 (O_781,N_24907,N_24042);
nand UO_782 (O_782,N_24125,N_24375);
nand UO_783 (O_783,N_24315,N_24032);
xnor UO_784 (O_784,N_24459,N_24870);
nor UO_785 (O_785,N_23755,N_24949);
nand UO_786 (O_786,N_24582,N_24297);
and UO_787 (O_787,N_24784,N_24811);
nor UO_788 (O_788,N_24404,N_24677);
or UO_789 (O_789,N_23881,N_23989);
or UO_790 (O_790,N_24575,N_24881);
nand UO_791 (O_791,N_24188,N_24410);
xnor UO_792 (O_792,N_24140,N_23774);
or UO_793 (O_793,N_24458,N_24672);
nand UO_794 (O_794,N_24383,N_24088);
nor UO_795 (O_795,N_23754,N_24413);
nand UO_796 (O_796,N_23794,N_23865);
nor UO_797 (O_797,N_24247,N_24055);
nand UO_798 (O_798,N_23878,N_24072);
xor UO_799 (O_799,N_24473,N_24115);
nand UO_800 (O_800,N_24748,N_24751);
nand UO_801 (O_801,N_24567,N_24651);
nand UO_802 (O_802,N_24034,N_24507);
xor UO_803 (O_803,N_24725,N_24384);
nor UO_804 (O_804,N_24100,N_24487);
and UO_805 (O_805,N_24058,N_24939);
nor UO_806 (O_806,N_24644,N_24859);
nand UO_807 (O_807,N_23761,N_24077);
or UO_808 (O_808,N_24697,N_24404);
and UO_809 (O_809,N_23911,N_23882);
xnor UO_810 (O_810,N_23934,N_24438);
nor UO_811 (O_811,N_24015,N_24485);
and UO_812 (O_812,N_24846,N_24365);
or UO_813 (O_813,N_24871,N_24244);
nand UO_814 (O_814,N_23994,N_24942);
or UO_815 (O_815,N_24174,N_24503);
or UO_816 (O_816,N_24129,N_24751);
xnor UO_817 (O_817,N_24875,N_23866);
nor UO_818 (O_818,N_24229,N_24782);
nand UO_819 (O_819,N_24308,N_24540);
or UO_820 (O_820,N_23929,N_24541);
nand UO_821 (O_821,N_24233,N_24083);
nor UO_822 (O_822,N_24301,N_24480);
or UO_823 (O_823,N_23819,N_24003);
xor UO_824 (O_824,N_24709,N_24103);
xor UO_825 (O_825,N_24779,N_24716);
xor UO_826 (O_826,N_24605,N_24297);
nor UO_827 (O_827,N_23892,N_24546);
and UO_828 (O_828,N_24782,N_23822);
nand UO_829 (O_829,N_24222,N_24827);
nand UO_830 (O_830,N_24492,N_24877);
and UO_831 (O_831,N_24004,N_24749);
and UO_832 (O_832,N_24410,N_24711);
or UO_833 (O_833,N_24962,N_24199);
or UO_834 (O_834,N_24212,N_24780);
and UO_835 (O_835,N_23789,N_24507);
or UO_836 (O_836,N_24522,N_24733);
and UO_837 (O_837,N_24528,N_24727);
nor UO_838 (O_838,N_24190,N_24595);
nand UO_839 (O_839,N_24646,N_23944);
nor UO_840 (O_840,N_24894,N_24505);
nand UO_841 (O_841,N_24291,N_24469);
and UO_842 (O_842,N_23878,N_24367);
or UO_843 (O_843,N_23920,N_24151);
or UO_844 (O_844,N_24242,N_24452);
nor UO_845 (O_845,N_24875,N_24017);
or UO_846 (O_846,N_24506,N_24631);
nand UO_847 (O_847,N_24357,N_24243);
and UO_848 (O_848,N_24056,N_24081);
or UO_849 (O_849,N_23894,N_24374);
and UO_850 (O_850,N_24457,N_24091);
nor UO_851 (O_851,N_24433,N_24233);
nor UO_852 (O_852,N_24389,N_24032);
or UO_853 (O_853,N_24177,N_24096);
and UO_854 (O_854,N_24366,N_24084);
xnor UO_855 (O_855,N_24458,N_24709);
xnor UO_856 (O_856,N_24092,N_24781);
nand UO_857 (O_857,N_24459,N_24942);
xnor UO_858 (O_858,N_23836,N_23957);
or UO_859 (O_859,N_23886,N_23996);
xnor UO_860 (O_860,N_24753,N_24613);
nand UO_861 (O_861,N_24822,N_24929);
nor UO_862 (O_862,N_24507,N_23942);
nor UO_863 (O_863,N_24157,N_23882);
or UO_864 (O_864,N_24731,N_23998);
and UO_865 (O_865,N_23804,N_24928);
and UO_866 (O_866,N_23819,N_24556);
and UO_867 (O_867,N_23850,N_24109);
nand UO_868 (O_868,N_24466,N_24110);
xor UO_869 (O_869,N_24949,N_23811);
xnor UO_870 (O_870,N_24441,N_24088);
nor UO_871 (O_871,N_24316,N_24487);
nor UO_872 (O_872,N_24526,N_24894);
nand UO_873 (O_873,N_24964,N_24649);
or UO_874 (O_874,N_24136,N_24118);
or UO_875 (O_875,N_24289,N_24177);
nand UO_876 (O_876,N_24996,N_24847);
xor UO_877 (O_877,N_24185,N_23828);
and UO_878 (O_878,N_24754,N_23955);
nor UO_879 (O_879,N_23862,N_24661);
xnor UO_880 (O_880,N_24321,N_24509);
or UO_881 (O_881,N_23860,N_24891);
nand UO_882 (O_882,N_24969,N_24783);
and UO_883 (O_883,N_24403,N_24511);
or UO_884 (O_884,N_23811,N_24790);
nand UO_885 (O_885,N_24854,N_24857);
or UO_886 (O_886,N_24421,N_24899);
and UO_887 (O_887,N_23769,N_24540);
nor UO_888 (O_888,N_24779,N_23751);
or UO_889 (O_889,N_24821,N_24265);
nand UO_890 (O_890,N_23880,N_24416);
or UO_891 (O_891,N_24934,N_24916);
and UO_892 (O_892,N_24880,N_24175);
nor UO_893 (O_893,N_23830,N_24283);
nor UO_894 (O_894,N_24366,N_24056);
nor UO_895 (O_895,N_24842,N_24512);
nand UO_896 (O_896,N_23799,N_24343);
or UO_897 (O_897,N_24407,N_24644);
or UO_898 (O_898,N_24867,N_24260);
or UO_899 (O_899,N_24985,N_24255);
xor UO_900 (O_900,N_24725,N_23879);
xnor UO_901 (O_901,N_24435,N_24314);
nor UO_902 (O_902,N_24813,N_24069);
or UO_903 (O_903,N_24021,N_24935);
nand UO_904 (O_904,N_23874,N_24321);
nand UO_905 (O_905,N_24699,N_24061);
xnor UO_906 (O_906,N_24621,N_24462);
nor UO_907 (O_907,N_24586,N_24148);
xor UO_908 (O_908,N_24369,N_24234);
nand UO_909 (O_909,N_24940,N_24235);
or UO_910 (O_910,N_24252,N_24492);
and UO_911 (O_911,N_24693,N_24391);
xor UO_912 (O_912,N_23767,N_24879);
or UO_913 (O_913,N_24900,N_23887);
and UO_914 (O_914,N_23893,N_24629);
nand UO_915 (O_915,N_24811,N_24678);
or UO_916 (O_916,N_24320,N_24575);
and UO_917 (O_917,N_24995,N_24839);
or UO_918 (O_918,N_24471,N_24613);
or UO_919 (O_919,N_24841,N_24489);
or UO_920 (O_920,N_24458,N_24870);
or UO_921 (O_921,N_24103,N_24166);
nor UO_922 (O_922,N_24683,N_24611);
xor UO_923 (O_923,N_24283,N_24790);
nand UO_924 (O_924,N_23792,N_24208);
nor UO_925 (O_925,N_24632,N_24059);
or UO_926 (O_926,N_24786,N_24547);
nand UO_927 (O_927,N_24503,N_24212);
or UO_928 (O_928,N_24545,N_24281);
or UO_929 (O_929,N_24363,N_24151);
xnor UO_930 (O_930,N_24098,N_24738);
and UO_931 (O_931,N_23953,N_24782);
nand UO_932 (O_932,N_24236,N_24582);
nor UO_933 (O_933,N_24533,N_24372);
nand UO_934 (O_934,N_23949,N_24831);
xor UO_935 (O_935,N_24494,N_24747);
or UO_936 (O_936,N_24413,N_24940);
or UO_937 (O_937,N_24758,N_24463);
xor UO_938 (O_938,N_23967,N_24629);
nor UO_939 (O_939,N_24767,N_24919);
xor UO_940 (O_940,N_24993,N_23913);
xnor UO_941 (O_941,N_24927,N_24826);
nand UO_942 (O_942,N_24034,N_24050);
nor UO_943 (O_943,N_23955,N_24112);
or UO_944 (O_944,N_24254,N_24621);
nand UO_945 (O_945,N_24797,N_24802);
nand UO_946 (O_946,N_24806,N_23801);
nand UO_947 (O_947,N_24785,N_24181);
and UO_948 (O_948,N_24276,N_24079);
nand UO_949 (O_949,N_24557,N_24158);
and UO_950 (O_950,N_24822,N_24907);
xor UO_951 (O_951,N_23789,N_24458);
nor UO_952 (O_952,N_24944,N_24013);
nor UO_953 (O_953,N_24915,N_23750);
and UO_954 (O_954,N_24144,N_24844);
or UO_955 (O_955,N_24131,N_23858);
xor UO_956 (O_956,N_24400,N_24122);
nor UO_957 (O_957,N_24903,N_24783);
and UO_958 (O_958,N_24650,N_24858);
nand UO_959 (O_959,N_24735,N_24959);
and UO_960 (O_960,N_24096,N_23861);
nand UO_961 (O_961,N_24591,N_24960);
and UO_962 (O_962,N_24749,N_24591);
nand UO_963 (O_963,N_23802,N_24634);
nor UO_964 (O_964,N_24070,N_24616);
and UO_965 (O_965,N_24699,N_24986);
nand UO_966 (O_966,N_24672,N_24144);
xnor UO_967 (O_967,N_24282,N_24163);
nor UO_968 (O_968,N_24733,N_24258);
nand UO_969 (O_969,N_23988,N_24284);
and UO_970 (O_970,N_24322,N_24121);
xnor UO_971 (O_971,N_24161,N_24224);
and UO_972 (O_972,N_24438,N_24122);
nand UO_973 (O_973,N_24064,N_24966);
or UO_974 (O_974,N_24049,N_24866);
nand UO_975 (O_975,N_24397,N_24815);
nor UO_976 (O_976,N_24201,N_24241);
or UO_977 (O_977,N_24591,N_24376);
and UO_978 (O_978,N_23851,N_24065);
nand UO_979 (O_979,N_24141,N_23897);
nand UO_980 (O_980,N_23984,N_24924);
nor UO_981 (O_981,N_24105,N_24108);
or UO_982 (O_982,N_23779,N_24555);
xor UO_983 (O_983,N_24463,N_24124);
or UO_984 (O_984,N_24931,N_24908);
xor UO_985 (O_985,N_24673,N_24991);
or UO_986 (O_986,N_23923,N_24720);
or UO_987 (O_987,N_24757,N_24124);
xnor UO_988 (O_988,N_23911,N_24397);
and UO_989 (O_989,N_24637,N_24873);
nand UO_990 (O_990,N_24604,N_24748);
and UO_991 (O_991,N_24941,N_24200);
nand UO_992 (O_992,N_24255,N_23835);
or UO_993 (O_993,N_24581,N_24858);
nor UO_994 (O_994,N_23863,N_24766);
nand UO_995 (O_995,N_24106,N_24939);
nand UO_996 (O_996,N_24507,N_24573);
and UO_997 (O_997,N_24596,N_24046);
nor UO_998 (O_998,N_24753,N_24728);
or UO_999 (O_999,N_23841,N_24754);
xor UO_1000 (O_1000,N_24865,N_23916);
and UO_1001 (O_1001,N_24102,N_24226);
and UO_1002 (O_1002,N_24135,N_24650);
or UO_1003 (O_1003,N_23891,N_24467);
xnor UO_1004 (O_1004,N_24499,N_24045);
and UO_1005 (O_1005,N_24623,N_24796);
and UO_1006 (O_1006,N_24936,N_24345);
nor UO_1007 (O_1007,N_24536,N_24108);
nor UO_1008 (O_1008,N_24255,N_24214);
nand UO_1009 (O_1009,N_24736,N_24887);
nand UO_1010 (O_1010,N_24022,N_23967);
or UO_1011 (O_1011,N_24490,N_24544);
nor UO_1012 (O_1012,N_24647,N_24160);
or UO_1013 (O_1013,N_24256,N_24773);
nand UO_1014 (O_1014,N_23934,N_24311);
and UO_1015 (O_1015,N_24969,N_24603);
or UO_1016 (O_1016,N_24995,N_24972);
nor UO_1017 (O_1017,N_24768,N_24882);
xor UO_1018 (O_1018,N_23831,N_24186);
and UO_1019 (O_1019,N_24213,N_24597);
nor UO_1020 (O_1020,N_24742,N_24759);
nor UO_1021 (O_1021,N_24832,N_24525);
nand UO_1022 (O_1022,N_24193,N_24231);
nand UO_1023 (O_1023,N_24013,N_24623);
nor UO_1024 (O_1024,N_24838,N_24082);
nand UO_1025 (O_1025,N_24865,N_24417);
nand UO_1026 (O_1026,N_24636,N_24565);
xor UO_1027 (O_1027,N_23750,N_24793);
nand UO_1028 (O_1028,N_24272,N_24549);
nand UO_1029 (O_1029,N_23752,N_24190);
or UO_1030 (O_1030,N_24324,N_24528);
and UO_1031 (O_1031,N_24319,N_24413);
xor UO_1032 (O_1032,N_24702,N_23963);
xnor UO_1033 (O_1033,N_23752,N_23816);
and UO_1034 (O_1034,N_23945,N_24970);
nand UO_1035 (O_1035,N_24454,N_24409);
nand UO_1036 (O_1036,N_24536,N_24175);
and UO_1037 (O_1037,N_24714,N_24690);
or UO_1038 (O_1038,N_24216,N_23750);
xnor UO_1039 (O_1039,N_24897,N_23769);
and UO_1040 (O_1040,N_24741,N_24499);
or UO_1041 (O_1041,N_24279,N_23911);
and UO_1042 (O_1042,N_24981,N_24428);
nand UO_1043 (O_1043,N_23964,N_24848);
nand UO_1044 (O_1044,N_24468,N_24800);
xnor UO_1045 (O_1045,N_24625,N_24337);
nor UO_1046 (O_1046,N_23760,N_24138);
nor UO_1047 (O_1047,N_24027,N_24356);
and UO_1048 (O_1048,N_24735,N_24009);
xor UO_1049 (O_1049,N_24379,N_24883);
and UO_1050 (O_1050,N_24383,N_24684);
nand UO_1051 (O_1051,N_24507,N_23904);
xor UO_1052 (O_1052,N_24926,N_24694);
xnor UO_1053 (O_1053,N_24005,N_24604);
nor UO_1054 (O_1054,N_23959,N_24008);
and UO_1055 (O_1055,N_24377,N_24516);
xnor UO_1056 (O_1056,N_24581,N_24131);
and UO_1057 (O_1057,N_24859,N_24398);
or UO_1058 (O_1058,N_24084,N_24386);
and UO_1059 (O_1059,N_23930,N_24799);
or UO_1060 (O_1060,N_23984,N_24176);
or UO_1061 (O_1061,N_24575,N_24075);
xnor UO_1062 (O_1062,N_23833,N_24496);
xor UO_1063 (O_1063,N_24489,N_24413);
nand UO_1064 (O_1064,N_24510,N_24907);
nand UO_1065 (O_1065,N_24411,N_23759);
and UO_1066 (O_1066,N_24834,N_24892);
nor UO_1067 (O_1067,N_24731,N_23865);
and UO_1068 (O_1068,N_24021,N_24662);
nand UO_1069 (O_1069,N_24328,N_24215);
or UO_1070 (O_1070,N_24077,N_24872);
xor UO_1071 (O_1071,N_24274,N_24396);
nand UO_1072 (O_1072,N_24183,N_24133);
and UO_1073 (O_1073,N_23868,N_24193);
and UO_1074 (O_1074,N_24473,N_23945);
nor UO_1075 (O_1075,N_24032,N_24373);
nand UO_1076 (O_1076,N_24122,N_23959);
nand UO_1077 (O_1077,N_24817,N_24165);
or UO_1078 (O_1078,N_24318,N_24062);
nor UO_1079 (O_1079,N_24226,N_24283);
and UO_1080 (O_1080,N_24494,N_24385);
nor UO_1081 (O_1081,N_23815,N_24909);
nor UO_1082 (O_1082,N_24651,N_24347);
or UO_1083 (O_1083,N_24011,N_24045);
xor UO_1084 (O_1084,N_24600,N_23897);
or UO_1085 (O_1085,N_24864,N_24709);
nor UO_1086 (O_1086,N_24789,N_24705);
nand UO_1087 (O_1087,N_24263,N_24726);
or UO_1088 (O_1088,N_24638,N_23985);
and UO_1089 (O_1089,N_24892,N_24179);
and UO_1090 (O_1090,N_23977,N_24958);
nor UO_1091 (O_1091,N_24805,N_23981);
xor UO_1092 (O_1092,N_24042,N_24378);
nand UO_1093 (O_1093,N_23762,N_24290);
and UO_1094 (O_1094,N_24720,N_24187);
nor UO_1095 (O_1095,N_24847,N_24539);
nand UO_1096 (O_1096,N_24598,N_23965);
xnor UO_1097 (O_1097,N_24260,N_24383);
or UO_1098 (O_1098,N_24058,N_24194);
and UO_1099 (O_1099,N_23851,N_24554);
nor UO_1100 (O_1100,N_24634,N_24926);
xnor UO_1101 (O_1101,N_24687,N_24297);
nand UO_1102 (O_1102,N_24369,N_23773);
nor UO_1103 (O_1103,N_24830,N_24779);
xor UO_1104 (O_1104,N_23930,N_24406);
or UO_1105 (O_1105,N_24685,N_24503);
nor UO_1106 (O_1106,N_24936,N_24570);
nand UO_1107 (O_1107,N_24170,N_24308);
xor UO_1108 (O_1108,N_24437,N_24606);
nor UO_1109 (O_1109,N_24354,N_24968);
or UO_1110 (O_1110,N_24933,N_24589);
or UO_1111 (O_1111,N_24131,N_23911);
or UO_1112 (O_1112,N_23824,N_24184);
nor UO_1113 (O_1113,N_24095,N_24181);
or UO_1114 (O_1114,N_24286,N_24038);
nand UO_1115 (O_1115,N_23983,N_24249);
xnor UO_1116 (O_1116,N_24682,N_23861);
and UO_1117 (O_1117,N_24497,N_24046);
or UO_1118 (O_1118,N_24183,N_24474);
nor UO_1119 (O_1119,N_24862,N_24288);
or UO_1120 (O_1120,N_24872,N_24292);
or UO_1121 (O_1121,N_24000,N_24116);
xor UO_1122 (O_1122,N_24912,N_24658);
nor UO_1123 (O_1123,N_24625,N_23972);
xnor UO_1124 (O_1124,N_23857,N_24548);
and UO_1125 (O_1125,N_24882,N_24092);
or UO_1126 (O_1126,N_24552,N_24116);
and UO_1127 (O_1127,N_24258,N_24099);
xnor UO_1128 (O_1128,N_23851,N_24231);
nand UO_1129 (O_1129,N_24220,N_24223);
nor UO_1130 (O_1130,N_23857,N_24265);
and UO_1131 (O_1131,N_24378,N_23909);
nor UO_1132 (O_1132,N_24228,N_24119);
and UO_1133 (O_1133,N_24337,N_24364);
nor UO_1134 (O_1134,N_24243,N_23750);
nor UO_1135 (O_1135,N_23828,N_24330);
or UO_1136 (O_1136,N_24951,N_24583);
nor UO_1137 (O_1137,N_24189,N_24772);
or UO_1138 (O_1138,N_24556,N_24147);
nor UO_1139 (O_1139,N_24990,N_24375);
and UO_1140 (O_1140,N_24146,N_24038);
or UO_1141 (O_1141,N_24274,N_23780);
nand UO_1142 (O_1142,N_24989,N_24640);
nor UO_1143 (O_1143,N_24888,N_23887);
nor UO_1144 (O_1144,N_24190,N_24015);
nand UO_1145 (O_1145,N_24874,N_24916);
or UO_1146 (O_1146,N_24677,N_24894);
nand UO_1147 (O_1147,N_24318,N_24032);
nor UO_1148 (O_1148,N_24514,N_24942);
nand UO_1149 (O_1149,N_23981,N_24635);
and UO_1150 (O_1150,N_24009,N_23954);
nor UO_1151 (O_1151,N_24496,N_23768);
nand UO_1152 (O_1152,N_23840,N_24828);
or UO_1153 (O_1153,N_24466,N_24619);
and UO_1154 (O_1154,N_24143,N_24078);
or UO_1155 (O_1155,N_23986,N_23827);
nor UO_1156 (O_1156,N_24930,N_24086);
and UO_1157 (O_1157,N_24791,N_24893);
or UO_1158 (O_1158,N_23959,N_24723);
and UO_1159 (O_1159,N_23780,N_24176);
and UO_1160 (O_1160,N_24437,N_24494);
or UO_1161 (O_1161,N_24953,N_23834);
and UO_1162 (O_1162,N_24374,N_23921);
nor UO_1163 (O_1163,N_23965,N_24252);
or UO_1164 (O_1164,N_23880,N_23776);
or UO_1165 (O_1165,N_24557,N_24471);
nor UO_1166 (O_1166,N_24922,N_24242);
xnor UO_1167 (O_1167,N_24226,N_24815);
nor UO_1168 (O_1168,N_24708,N_24648);
nand UO_1169 (O_1169,N_24625,N_24770);
nor UO_1170 (O_1170,N_23780,N_24345);
nor UO_1171 (O_1171,N_24421,N_24288);
nand UO_1172 (O_1172,N_24184,N_24633);
xnor UO_1173 (O_1173,N_24670,N_23849);
and UO_1174 (O_1174,N_24167,N_24915);
or UO_1175 (O_1175,N_24512,N_24272);
or UO_1176 (O_1176,N_23817,N_23888);
or UO_1177 (O_1177,N_23818,N_24392);
or UO_1178 (O_1178,N_23835,N_23759);
nor UO_1179 (O_1179,N_24350,N_23827);
nand UO_1180 (O_1180,N_24861,N_24467);
xnor UO_1181 (O_1181,N_24766,N_24468);
nor UO_1182 (O_1182,N_24509,N_23791);
and UO_1183 (O_1183,N_23759,N_24144);
and UO_1184 (O_1184,N_24898,N_24584);
xor UO_1185 (O_1185,N_24242,N_24983);
or UO_1186 (O_1186,N_24905,N_24655);
nand UO_1187 (O_1187,N_23870,N_24777);
or UO_1188 (O_1188,N_23854,N_24173);
nand UO_1189 (O_1189,N_24489,N_24464);
or UO_1190 (O_1190,N_23875,N_24795);
and UO_1191 (O_1191,N_24495,N_24746);
xor UO_1192 (O_1192,N_24305,N_24706);
xnor UO_1193 (O_1193,N_23789,N_23939);
or UO_1194 (O_1194,N_24828,N_24424);
nand UO_1195 (O_1195,N_24644,N_24200);
nand UO_1196 (O_1196,N_24108,N_24077);
nand UO_1197 (O_1197,N_23961,N_23972);
or UO_1198 (O_1198,N_24855,N_24943);
nor UO_1199 (O_1199,N_23860,N_23954);
xor UO_1200 (O_1200,N_24073,N_23913);
or UO_1201 (O_1201,N_23783,N_24232);
nor UO_1202 (O_1202,N_24227,N_24807);
nand UO_1203 (O_1203,N_24304,N_23863);
nor UO_1204 (O_1204,N_24607,N_24285);
and UO_1205 (O_1205,N_23983,N_23895);
or UO_1206 (O_1206,N_23810,N_24543);
and UO_1207 (O_1207,N_24395,N_24602);
nand UO_1208 (O_1208,N_23761,N_24890);
and UO_1209 (O_1209,N_24542,N_23820);
and UO_1210 (O_1210,N_24722,N_24712);
xnor UO_1211 (O_1211,N_24983,N_24163);
or UO_1212 (O_1212,N_24084,N_23991);
xnor UO_1213 (O_1213,N_24125,N_24967);
xor UO_1214 (O_1214,N_23822,N_24708);
xnor UO_1215 (O_1215,N_24347,N_23894);
nand UO_1216 (O_1216,N_24983,N_23985);
nor UO_1217 (O_1217,N_23891,N_23781);
xnor UO_1218 (O_1218,N_24940,N_24310);
nand UO_1219 (O_1219,N_24264,N_24482);
and UO_1220 (O_1220,N_24907,N_24980);
xor UO_1221 (O_1221,N_24088,N_24912);
and UO_1222 (O_1222,N_24718,N_24474);
nand UO_1223 (O_1223,N_24915,N_23821);
nor UO_1224 (O_1224,N_24107,N_23856);
or UO_1225 (O_1225,N_24099,N_24102);
or UO_1226 (O_1226,N_24314,N_24375);
and UO_1227 (O_1227,N_24085,N_24003);
xor UO_1228 (O_1228,N_24722,N_24140);
nor UO_1229 (O_1229,N_24000,N_23752);
or UO_1230 (O_1230,N_24650,N_24911);
nor UO_1231 (O_1231,N_23959,N_24168);
and UO_1232 (O_1232,N_24907,N_24261);
nor UO_1233 (O_1233,N_23864,N_24072);
or UO_1234 (O_1234,N_24545,N_23896);
nor UO_1235 (O_1235,N_24358,N_24873);
or UO_1236 (O_1236,N_24429,N_24898);
nor UO_1237 (O_1237,N_24679,N_23985);
nor UO_1238 (O_1238,N_23893,N_24234);
and UO_1239 (O_1239,N_24618,N_24179);
nor UO_1240 (O_1240,N_23891,N_23923);
nand UO_1241 (O_1241,N_24561,N_24623);
or UO_1242 (O_1242,N_24085,N_24435);
xor UO_1243 (O_1243,N_24592,N_24116);
and UO_1244 (O_1244,N_24801,N_24332);
and UO_1245 (O_1245,N_23765,N_24244);
nor UO_1246 (O_1246,N_24559,N_23995);
and UO_1247 (O_1247,N_24885,N_24623);
xnor UO_1248 (O_1248,N_23797,N_24309);
nand UO_1249 (O_1249,N_23988,N_23752);
nor UO_1250 (O_1250,N_23858,N_24336);
or UO_1251 (O_1251,N_23978,N_24486);
nand UO_1252 (O_1252,N_23765,N_23793);
and UO_1253 (O_1253,N_24098,N_24704);
or UO_1254 (O_1254,N_23987,N_23888);
nand UO_1255 (O_1255,N_23920,N_24498);
nor UO_1256 (O_1256,N_24964,N_23838);
nor UO_1257 (O_1257,N_24782,N_24103);
or UO_1258 (O_1258,N_24611,N_24224);
xnor UO_1259 (O_1259,N_24692,N_24879);
nor UO_1260 (O_1260,N_24615,N_23913);
nor UO_1261 (O_1261,N_24204,N_24069);
nand UO_1262 (O_1262,N_24335,N_24673);
nor UO_1263 (O_1263,N_24896,N_24500);
or UO_1264 (O_1264,N_23811,N_23857);
and UO_1265 (O_1265,N_24164,N_24435);
and UO_1266 (O_1266,N_24843,N_24618);
nand UO_1267 (O_1267,N_24934,N_24623);
xnor UO_1268 (O_1268,N_24650,N_24235);
nor UO_1269 (O_1269,N_24261,N_24729);
nor UO_1270 (O_1270,N_24354,N_24430);
and UO_1271 (O_1271,N_24404,N_23922);
xor UO_1272 (O_1272,N_24502,N_24077);
xnor UO_1273 (O_1273,N_24774,N_24506);
nor UO_1274 (O_1274,N_24064,N_24950);
and UO_1275 (O_1275,N_23899,N_23822);
or UO_1276 (O_1276,N_24053,N_24695);
and UO_1277 (O_1277,N_24393,N_24081);
nand UO_1278 (O_1278,N_24058,N_23953);
and UO_1279 (O_1279,N_24760,N_23974);
nor UO_1280 (O_1280,N_24426,N_24742);
and UO_1281 (O_1281,N_24558,N_24023);
nor UO_1282 (O_1282,N_24936,N_24003);
nor UO_1283 (O_1283,N_23992,N_24923);
nor UO_1284 (O_1284,N_24894,N_24758);
xor UO_1285 (O_1285,N_24837,N_24338);
xor UO_1286 (O_1286,N_24605,N_24353);
xnor UO_1287 (O_1287,N_24408,N_24723);
and UO_1288 (O_1288,N_24296,N_24638);
nand UO_1289 (O_1289,N_24548,N_24470);
or UO_1290 (O_1290,N_24141,N_24063);
and UO_1291 (O_1291,N_23830,N_24260);
or UO_1292 (O_1292,N_24668,N_23992);
nand UO_1293 (O_1293,N_24015,N_24018);
nand UO_1294 (O_1294,N_23997,N_24807);
nand UO_1295 (O_1295,N_24750,N_24602);
nor UO_1296 (O_1296,N_24834,N_24748);
xor UO_1297 (O_1297,N_24742,N_24311);
nor UO_1298 (O_1298,N_23874,N_24597);
nand UO_1299 (O_1299,N_23944,N_24874);
nand UO_1300 (O_1300,N_23868,N_24706);
nor UO_1301 (O_1301,N_24367,N_24108);
nand UO_1302 (O_1302,N_24379,N_24726);
and UO_1303 (O_1303,N_24335,N_24315);
nor UO_1304 (O_1304,N_24735,N_24188);
xor UO_1305 (O_1305,N_24062,N_24262);
nand UO_1306 (O_1306,N_24392,N_24657);
nand UO_1307 (O_1307,N_24582,N_24632);
or UO_1308 (O_1308,N_24821,N_24945);
and UO_1309 (O_1309,N_24515,N_24856);
nand UO_1310 (O_1310,N_24829,N_24022);
nor UO_1311 (O_1311,N_24516,N_24173);
nor UO_1312 (O_1312,N_23873,N_24095);
nor UO_1313 (O_1313,N_24182,N_24187);
xor UO_1314 (O_1314,N_24828,N_23998);
xnor UO_1315 (O_1315,N_24978,N_24295);
nand UO_1316 (O_1316,N_24256,N_24927);
nand UO_1317 (O_1317,N_24507,N_24467);
xnor UO_1318 (O_1318,N_24532,N_24337);
nand UO_1319 (O_1319,N_23751,N_24937);
or UO_1320 (O_1320,N_24089,N_24158);
or UO_1321 (O_1321,N_24387,N_24926);
and UO_1322 (O_1322,N_24371,N_24352);
nand UO_1323 (O_1323,N_24184,N_23825);
xor UO_1324 (O_1324,N_24590,N_24844);
nand UO_1325 (O_1325,N_24182,N_24222);
and UO_1326 (O_1326,N_23903,N_24950);
nand UO_1327 (O_1327,N_24607,N_24520);
or UO_1328 (O_1328,N_24996,N_24537);
xor UO_1329 (O_1329,N_24030,N_24604);
nor UO_1330 (O_1330,N_24446,N_24833);
xnor UO_1331 (O_1331,N_24529,N_23800);
nand UO_1332 (O_1332,N_24708,N_24988);
nand UO_1333 (O_1333,N_24418,N_24627);
nor UO_1334 (O_1334,N_23969,N_23776);
and UO_1335 (O_1335,N_24617,N_23921);
nor UO_1336 (O_1336,N_24388,N_23764);
and UO_1337 (O_1337,N_24975,N_24953);
nand UO_1338 (O_1338,N_24840,N_24925);
or UO_1339 (O_1339,N_24280,N_23993);
nor UO_1340 (O_1340,N_23828,N_24158);
and UO_1341 (O_1341,N_24338,N_24286);
xor UO_1342 (O_1342,N_24270,N_24661);
xnor UO_1343 (O_1343,N_24656,N_24369);
xor UO_1344 (O_1344,N_24270,N_24435);
nor UO_1345 (O_1345,N_23976,N_24258);
nand UO_1346 (O_1346,N_24672,N_24234);
and UO_1347 (O_1347,N_24347,N_24507);
nand UO_1348 (O_1348,N_24768,N_24933);
or UO_1349 (O_1349,N_24517,N_24259);
nor UO_1350 (O_1350,N_23833,N_23933);
nor UO_1351 (O_1351,N_24394,N_24876);
nor UO_1352 (O_1352,N_24661,N_24772);
or UO_1353 (O_1353,N_24213,N_23924);
nand UO_1354 (O_1354,N_24785,N_23805);
nand UO_1355 (O_1355,N_23860,N_24829);
nand UO_1356 (O_1356,N_24995,N_24627);
and UO_1357 (O_1357,N_24756,N_23769);
xnor UO_1358 (O_1358,N_23922,N_24744);
nand UO_1359 (O_1359,N_24778,N_24372);
and UO_1360 (O_1360,N_24856,N_23929);
xnor UO_1361 (O_1361,N_24033,N_23876);
and UO_1362 (O_1362,N_24801,N_24164);
nor UO_1363 (O_1363,N_23976,N_24707);
and UO_1364 (O_1364,N_24247,N_24582);
xnor UO_1365 (O_1365,N_24378,N_24616);
or UO_1366 (O_1366,N_23898,N_24592);
and UO_1367 (O_1367,N_24548,N_24838);
xnor UO_1368 (O_1368,N_23752,N_24173);
nor UO_1369 (O_1369,N_24980,N_24793);
or UO_1370 (O_1370,N_24402,N_24720);
and UO_1371 (O_1371,N_23968,N_24857);
nand UO_1372 (O_1372,N_24189,N_24529);
nand UO_1373 (O_1373,N_24483,N_23957);
nand UO_1374 (O_1374,N_23842,N_24877);
xnor UO_1375 (O_1375,N_24296,N_23799);
or UO_1376 (O_1376,N_24300,N_23771);
or UO_1377 (O_1377,N_24718,N_24866);
xnor UO_1378 (O_1378,N_24702,N_23869);
nor UO_1379 (O_1379,N_23834,N_24838);
or UO_1380 (O_1380,N_24328,N_24330);
xnor UO_1381 (O_1381,N_24096,N_23825);
nand UO_1382 (O_1382,N_24671,N_24743);
nand UO_1383 (O_1383,N_24357,N_24845);
nor UO_1384 (O_1384,N_24599,N_24102);
or UO_1385 (O_1385,N_24017,N_23761);
or UO_1386 (O_1386,N_24053,N_23865);
nor UO_1387 (O_1387,N_23855,N_24298);
nor UO_1388 (O_1388,N_24292,N_23818);
nand UO_1389 (O_1389,N_24943,N_24701);
xnor UO_1390 (O_1390,N_23778,N_24313);
nor UO_1391 (O_1391,N_23973,N_23870);
nand UO_1392 (O_1392,N_23990,N_24178);
nor UO_1393 (O_1393,N_24030,N_24542);
nor UO_1394 (O_1394,N_24948,N_24925);
and UO_1395 (O_1395,N_24140,N_24748);
nand UO_1396 (O_1396,N_24536,N_24231);
xnor UO_1397 (O_1397,N_24685,N_23915);
nor UO_1398 (O_1398,N_24716,N_24486);
or UO_1399 (O_1399,N_24711,N_24026);
or UO_1400 (O_1400,N_24802,N_24023);
nor UO_1401 (O_1401,N_24737,N_24438);
nor UO_1402 (O_1402,N_24973,N_24430);
or UO_1403 (O_1403,N_24004,N_24855);
xnor UO_1404 (O_1404,N_24289,N_23789);
nand UO_1405 (O_1405,N_23923,N_24563);
or UO_1406 (O_1406,N_24318,N_24182);
xnor UO_1407 (O_1407,N_24430,N_24392);
or UO_1408 (O_1408,N_24402,N_24633);
or UO_1409 (O_1409,N_24846,N_24513);
nand UO_1410 (O_1410,N_24002,N_24053);
nor UO_1411 (O_1411,N_24342,N_24248);
and UO_1412 (O_1412,N_23844,N_23878);
or UO_1413 (O_1413,N_23839,N_24256);
xnor UO_1414 (O_1414,N_24643,N_24018);
xor UO_1415 (O_1415,N_24621,N_23820);
nor UO_1416 (O_1416,N_24582,N_24890);
nor UO_1417 (O_1417,N_24020,N_24516);
or UO_1418 (O_1418,N_24564,N_24275);
xor UO_1419 (O_1419,N_24578,N_24591);
and UO_1420 (O_1420,N_24555,N_24791);
and UO_1421 (O_1421,N_24201,N_24136);
nand UO_1422 (O_1422,N_24021,N_24146);
nand UO_1423 (O_1423,N_24042,N_24767);
nor UO_1424 (O_1424,N_24158,N_24673);
nor UO_1425 (O_1425,N_24579,N_24868);
nand UO_1426 (O_1426,N_24358,N_23919);
or UO_1427 (O_1427,N_24141,N_24424);
xor UO_1428 (O_1428,N_24068,N_24634);
nand UO_1429 (O_1429,N_23931,N_24765);
nand UO_1430 (O_1430,N_24161,N_24209);
nand UO_1431 (O_1431,N_24781,N_24695);
nand UO_1432 (O_1432,N_24452,N_24934);
xor UO_1433 (O_1433,N_24091,N_23830);
and UO_1434 (O_1434,N_23848,N_24304);
nand UO_1435 (O_1435,N_24066,N_24424);
or UO_1436 (O_1436,N_24470,N_24077);
or UO_1437 (O_1437,N_24107,N_24506);
nor UO_1438 (O_1438,N_23976,N_24942);
nand UO_1439 (O_1439,N_24176,N_23832);
nand UO_1440 (O_1440,N_24923,N_24611);
or UO_1441 (O_1441,N_23970,N_24394);
xnor UO_1442 (O_1442,N_24742,N_24443);
and UO_1443 (O_1443,N_24670,N_24266);
nor UO_1444 (O_1444,N_24085,N_24247);
or UO_1445 (O_1445,N_24145,N_24100);
nor UO_1446 (O_1446,N_24773,N_24954);
or UO_1447 (O_1447,N_24760,N_23850);
and UO_1448 (O_1448,N_23915,N_24287);
nor UO_1449 (O_1449,N_23872,N_24984);
nor UO_1450 (O_1450,N_24587,N_24801);
or UO_1451 (O_1451,N_24584,N_23774);
and UO_1452 (O_1452,N_24474,N_24283);
nand UO_1453 (O_1453,N_24650,N_24515);
nand UO_1454 (O_1454,N_24120,N_24279);
xnor UO_1455 (O_1455,N_23995,N_24036);
nand UO_1456 (O_1456,N_24722,N_24041);
and UO_1457 (O_1457,N_24758,N_23937);
and UO_1458 (O_1458,N_24244,N_24388);
nor UO_1459 (O_1459,N_23830,N_24994);
or UO_1460 (O_1460,N_24428,N_24020);
xor UO_1461 (O_1461,N_24466,N_24923);
nand UO_1462 (O_1462,N_24859,N_23758);
and UO_1463 (O_1463,N_24331,N_24762);
nand UO_1464 (O_1464,N_24387,N_24481);
xnor UO_1465 (O_1465,N_24056,N_24825);
nand UO_1466 (O_1466,N_24048,N_23930);
or UO_1467 (O_1467,N_24267,N_24500);
nand UO_1468 (O_1468,N_24127,N_24320);
nor UO_1469 (O_1469,N_24723,N_24757);
and UO_1470 (O_1470,N_24466,N_24482);
nand UO_1471 (O_1471,N_24071,N_23832);
nand UO_1472 (O_1472,N_24647,N_24009);
nand UO_1473 (O_1473,N_24565,N_24669);
nor UO_1474 (O_1474,N_24732,N_24515);
nor UO_1475 (O_1475,N_24587,N_24983);
and UO_1476 (O_1476,N_24155,N_24742);
or UO_1477 (O_1477,N_24060,N_23967);
or UO_1478 (O_1478,N_24155,N_23800);
nor UO_1479 (O_1479,N_24692,N_24579);
nand UO_1480 (O_1480,N_24737,N_24351);
or UO_1481 (O_1481,N_23799,N_24391);
or UO_1482 (O_1482,N_24144,N_24686);
nand UO_1483 (O_1483,N_24336,N_24649);
nand UO_1484 (O_1484,N_24156,N_24217);
or UO_1485 (O_1485,N_24501,N_24462);
xnor UO_1486 (O_1486,N_24570,N_24089);
nor UO_1487 (O_1487,N_23988,N_23798);
and UO_1488 (O_1488,N_23972,N_24035);
nand UO_1489 (O_1489,N_23803,N_24332);
nor UO_1490 (O_1490,N_24143,N_24801);
and UO_1491 (O_1491,N_24479,N_24592);
and UO_1492 (O_1492,N_24667,N_24795);
or UO_1493 (O_1493,N_24665,N_24855);
or UO_1494 (O_1494,N_24109,N_24959);
xnor UO_1495 (O_1495,N_24311,N_24561);
xnor UO_1496 (O_1496,N_24312,N_24976);
nand UO_1497 (O_1497,N_23909,N_24255);
xor UO_1498 (O_1498,N_24865,N_24653);
xor UO_1499 (O_1499,N_24290,N_24374);
nand UO_1500 (O_1500,N_24531,N_23882);
or UO_1501 (O_1501,N_24526,N_24121);
nand UO_1502 (O_1502,N_23778,N_24929);
xnor UO_1503 (O_1503,N_24951,N_24750);
nor UO_1504 (O_1504,N_23901,N_24152);
and UO_1505 (O_1505,N_23904,N_23948);
nand UO_1506 (O_1506,N_24032,N_23964);
and UO_1507 (O_1507,N_24634,N_24390);
or UO_1508 (O_1508,N_24582,N_24851);
or UO_1509 (O_1509,N_24893,N_24057);
xnor UO_1510 (O_1510,N_24789,N_24877);
or UO_1511 (O_1511,N_23975,N_24876);
or UO_1512 (O_1512,N_24306,N_24634);
nand UO_1513 (O_1513,N_24245,N_24519);
or UO_1514 (O_1514,N_24639,N_24488);
xnor UO_1515 (O_1515,N_24330,N_24429);
or UO_1516 (O_1516,N_24912,N_24561);
xnor UO_1517 (O_1517,N_23952,N_24023);
xnor UO_1518 (O_1518,N_24655,N_24210);
or UO_1519 (O_1519,N_24876,N_24727);
nand UO_1520 (O_1520,N_24451,N_24922);
or UO_1521 (O_1521,N_24930,N_24700);
or UO_1522 (O_1522,N_24713,N_24089);
xnor UO_1523 (O_1523,N_24160,N_24345);
nor UO_1524 (O_1524,N_24701,N_24343);
and UO_1525 (O_1525,N_23760,N_24211);
xor UO_1526 (O_1526,N_24916,N_23819);
or UO_1527 (O_1527,N_24409,N_24301);
nand UO_1528 (O_1528,N_24545,N_24208);
or UO_1529 (O_1529,N_24651,N_24424);
and UO_1530 (O_1530,N_24813,N_24512);
and UO_1531 (O_1531,N_24689,N_24508);
xor UO_1532 (O_1532,N_24845,N_24361);
xor UO_1533 (O_1533,N_24230,N_23800);
nand UO_1534 (O_1534,N_24974,N_24511);
and UO_1535 (O_1535,N_24491,N_24242);
nand UO_1536 (O_1536,N_24744,N_24291);
and UO_1537 (O_1537,N_24057,N_24477);
nor UO_1538 (O_1538,N_24441,N_24198);
nor UO_1539 (O_1539,N_24151,N_24534);
xor UO_1540 (O_1540,N_23878,N_24450);
xnor UO_1541 (O_1541,N_24705,N_24363);
and UO_1542 (O_1542,N_23945,N_24424);
nor UO_1543 (O_1543,N_24705,N_24813);
and UO_1544 (O_1544,N_24727,N_23865);
nand UO_1545 (O_1545,N_23832,N_24871);
and UO_1546 (O_1546,N_24777,N_24085);
and UO_1547 (O_1547,N_24180,N_24455);
or UO_1548 (O_1548,N_24791,N_24627);
nor UO_1549 (O_1549,N_24724,N_24360);
or UO_1550 (O_1550,N_24976,N_24065);
xnor UO_1551 (O_1551,N_24992,N_24232);
xnor UO_1552 (O_1552,N_24077,N_24647);
nand UO_1553 (O_1553,N_24549,N_24607);
nand UO_1554 (O_1554,N_23992,N_24538);
and UO_1555 (O_1555,N_24184,N_24402);
xor UO_1556 (O_1556,N_24670,N_24517);
xor UO_1557 (O_1557,N_24887,N_23787);
and UO_1558 (O_1558,N_23869,N_24068);
xnor UO_1559 (O_1559,N_24533,N_23892);
or UO_1560 (O_1560,N_24512,N_24649);
nand UO_1561 (O_1561,N_24529,N_23942);
or UO_1562 (O_1562,N_24434,N_23875);
nand UO_1563 (O_1563,N_23925,N_24697);
xnor UO_1564 (O_1564,N_23986,N_23810);
or UO_1565 (O_1565,N_24867,N_24681);
nand UO_1566 (O_1566,N_24515,N_24314);
nand UO_1567 (O_1567,N_24466,N_23902);
nor UO_1568 (O_1568,N_24587,N_23783);
nand UO_1569 (O_1569,N_24158,N_24602);
and UO_1570 (O_1570,N_24747,N_24930);
xnor UO_1571 (O_1571,N_24110,N_24153);
nor UO_1572 (O_1572,N_23905,N_23985);
xor UO_1573 (O_1573,N_24904,N_24837);
or UO_1574 (O_1574,N_24257,N_24107);
or UO_1575 (O_1575,N_24178,N_24555);
nor UO_1576 (O_1576,N_23983,N_24979);
or UO_1577 (O_1577,N_24408,N_24464);
and UO_1578 (O_1578,N_24543,N_24488);
nor UO_1579 (O_1579,N_24427,N_24651);
nand UO_1580 (O_1580,N_24403,N_24106);
and UO_1581 (O_1581,N_24366,N_24669);
xor UO_1582 (O_1582,N_24849,N_24155);
and UO_1583 (O_1583,N_23954,N_24736);
nor UO_1584 (O_1584,N_23848,N_23890);
nand UO_1585 (O_1585,N_24118,N_24562);
nand UO_1586 (O_1586,N_24859,N_24273);
xnor UO_1587 (O_1587,N_24193,N_23857);
xor UO_1588 (O_1588,N_24077,N_24849);
xor UO_1589 (O_1589,N_24040,N_24818);
and UO_1590 (O_1590,N_24296,N_24254);
and UO_1591 (O_1591,N_24704,N_23898);
xnor UO_1592 (O_1592,N_24573,N_24367);
xor UO_1593 (O_1593,N_24568,N_23810);
xnor UO_1594 (O_1594,N_23988,N_24197);
nor UO_1595 (O_1595,N_24225,N_24534);
or UO_1596 (O_1596,N_23951,N_24941);
and UO_1597 (O_1597,N_24238,N_24506);
xor UO_1598 (O_1598,N_24958,N_24716);
or UO_1599 (O_1599,N_23917,N_24582);
or UO_1600 (O_1600,N_24808,N_24069);
nor UO_1601 (O_1601,N_24074,N_24231);
nand UO_1602 (O_1602,N_24326,N_23861);
xor UO_1603 (O_1603,N_24871,N_24150);
and UO_1604 (O_1604,N_23785,N_24165);
xnor UO_1605 (O_1605,N_23829,N_23824);
xor UO_1606 (O_1606,N_24243,N_24483);
xor UO_1607 (O_1607,N_24129,N_24493);
or UO_1608 (O_1608,N_24205,N_24268);
nor UO_1609 (O_1609,N_24917,N_23871);
nand UO_1610 (O_1610,N_23839,N_24347);
nor UO_1611 (O_1611,N_24507,N_24082);
and UO_1612 (O_1612,N_24960,N_24048);
nand UO_1613 (O_1613,N_24290,N_23895);
xnor UO_1614 (O_1614,N_23781,N_24862);
or UO_1615 (O_1615,N_24883,N_24718);
and UO_1616 (O_1616,N_24848,N_24376);
nor UO_1617 (O_1617,N_24099,N_24501);
nand UO_1618 (O_1618,N_24661,N_24558);
or UO_1619 (O_1619,N_24243,N_24220);
xnor UO_1620 (O_1620,N_24306,N_24950);
nand UO_1621 (O_1621,N_24880,N_24426);
nor UO_1622 (O_1622,N_24300,N_23772);
nor UO_1623 (O_1623,N_23952,N_23970);
or UO_1624 (O_1624,N_24835,N_24855);
or UO_1625 (O_1625,N_23953,N_23830);
nand UO_1626 (O_1626,N_23985,N_24086);
nor UO_1627 (O_1627,N_24309,N_23826);
xor UO_1628 (O_1628,N_24063,N_24426);
nor UO_1629 (O_1629,N_24119,N_24280);
and UO_1630 (O_1630,N_24261,N_23837);
nand UO_1631 (O_1631,N_24288,N_24849);
nor UO_1632 (O_1632,N_24162,N_24845);
nand UO_1633 (O_1633,N_24111,N_24062);
xnor UO_1634 (O_1634,N_24227,N_24382);
xnor UO_1635 (O_1635,N_23767,N_24076);
and UO_1636 (O_1636,N_24686,N_24036);
or UO_1637 (O_1637,N_24607,N_24465);
nand UO_1638 (O_1638,N_24940,N_24047);
nor UO_1639 (O_1639,N_24006,N_23825);
xor UO_1640 (O_1640,N_24689,N_23830);
and UO_1641 (O_1641,N_23822,N_23863);
and UO_1642 (O_1642,N_24148,N_24707);
and UO_1643 (O_1643,N_24149,N_24399);
or UO_1644 (O_1644,N_23862,N_24395);
nor UO_1645 (O_1645,N_23894,N_24332);
nor UO_1646 (O_1646,N_24489,N_24479);
nor UO_1647 (O_1647,N_24817,N_23965);
or UO_1648 (O_1648,N_24014,N_24187);
and UO_1649 (O_1649,N_24934,N_24523);
or UO_1650 (O_1650,N_24863,N_24875);
nor UO_1651 (O_1651,N_24981,N_24274);
nand UO_1652 (O_1652,N_24039,N_24097);
nor UO_1653 (O_1653,N_24489,N_23988);
or UO_1654 (O_1654,N_23941,N_24636);
or UO_1655 (O_1655,N_24409,N_24235);
nor UO_1656 (O_1656,N_24842,N_24356);
xnor UO_1657 (O_1657,N_23955,N_23963);
xor UO_1658 (O_1658,N_24737,N_24902);
or UO_1659 (O_1659,N_24498,N_24892);
and UO_1660 (O_1660,N_24923,N_24950);
and UO_1661 (O_1661,N_24426,N_24623);
or UO_1662 (O_1662,N_24288,N_24258);
or UO_1663 (O_1663,N_24917,N_24343);
xnor UO_1664 (O_1664,N_24083,N_24029);
and UO_1665 (O_1665,N_23802,N_24548);
xnor UO_1666 (O_1666,N_24968,N_24327);
nor UO_1667 (O_1667,N_24476,N_23753);
xnor UO_1668 (O_1668,N_24522,N_24349);
nand UO_1669 (O_1669,N_24472,N_24596);
nor UO_1670 (O_1670,N_24166,N_24970);
nand UO_1671 (O_1671,N_24372,N_24515);
nand UO_1672 (O_1672,N_24632,N_24670);
nor UO_1673 (O_1673,N_24421,N_24382);
xor UO_1674 (O_1674,N_23905,N_24001);
and UO_1675 (O_1675,N_23762,N_24597);
nor UO_1676 (O_1676,N_23963,N_24746);
nand UO_1677 (O_1677,N_23905,N_24926);
or UO_1678 (O_1678,N_24116,N_24838);
nor UO_1679 (O_1679,N_24440,N_24626);
nor UO_1680 (O_1680,N_24190,N_24971);
nand UO_1681 (O_1681,N_24546,N_24325);
and UO_1682 (O_1682,N_24215,N_23848);
xnor UO_1683 (O_1683,N_24980,N_24606);
xor UO_1684 (O_1684,N_24007,N_23863);
xnor UO_1685 (O_1685,N_24311,N_24868);
nor UO_1686 (O_1686,N_24181,N_24736);
nor UO_1687 (O_1687,N_24855,N_23974);
or UO_1688 (O_1688,N_24314,N_24254);
and UO_1689 (O_1689,N_24323,N_24981);
xnor UO_1690 (O_1690,N_24785,N_23941);
and UO_1691 (O_1691,N_23782,N_23789);
nand UO_1692 (O_1692,N_24749,N_24595);
xnor UO_1693 (O_1693,N_23943,N_24638);
xnor UO_1694 (O_1694,N_24488,N_24853);
xor UO_1695 (O_1695,N_24606,N_24605);
and UO_1696 (O_1696,N_23766,N_24825);
nand UO_1697 (O_1697,N_24649,N_24063);
nor UO_1698 (O_1698,N_24107,N_23891);
and UO_1699 (O_1699,N_24375,N_23908);
and UO_1700 (O_1700,N_24027,N_24203);
and UO_1701 (O_1701,N_24490,N_24737);
nor UO_1702 (O_1702,N_24379,N_24328);
xor UO_1703 (O_1703,N_23966,N_24876);
and UO_1704 (O_1704,N_23886,N_23788);
nand UO_1705 (O_1705,N_23758,N_24816);
nor UO_1706 (O_1706,N_24834,N_24886);
or UO_1707 (O_1707,N_24138,N_24050);
or UO_1708 (O_1708,N_24825,N_24677);
or UO_1709 (O_1709,N_24861,N_23795);
nor UO_1710 (O_1710,N_24100,N_24211);
nor UO_1711 (O_1711,N_24232,N_23992);
or UO_1712 (O_1712,N_24659,N_24066);
and UO_1713 (O_1713,N_24752,N_23787);
or UO_1714 (O_1714,N_24144,N_24243);
xnor UO_1715 (O_1715,N_24189,N_23851);
nor UO_1716 (O_1716,N_24343,N_24329);
nor UO_1717 (O_1717,N_24115,N_24153);
xnor UO_1718 (O_1718,N_24765,N_24187);
nor UO_1719 (O_1719,N_24911,N_24381);
nand UO_1720 (O_1720,N_24360,N_23766);
and UO_1721 (O_1721,N_24465,N_24825);
and UO_1722 (O_1722,N_24417,N_24854);
nor UO_1723 (O_1723,N_23968,N_24910);
or UO_1724 (O_1724,N_24144,N_24335);
and UO_1725 (O_1725,N_24177,N_24076);
nor UO_1726 (O_1726,N_24068,N_24476);
nor UO_1727 (O_1727,N_24219,N_24731);
nor UO_1728 (O_1728,N_24904,N_24823);
or UO_1729 (O_1729,N_23949,N_24214);
or UO_1730 (O_1730,N_24084,N_24380);
nand UO_1731 (O_1731,N_24754,N_24013);
nor UO_1732 (O_1732,N_24259,N_24263);
nor UO_1733 (O_1733,N_24156,N_24505);
and UO_1734 (O_1734,N_23772,N_24327);
nor UO_1735 (O_1735,N_24449,N_24761);
nor UO_1736 (O_1736,N_23770,N_24750);
nand UO_1737 (O_1737,N_24656,N_24238);
nor UO_1738 (O_1738,N_24305,N_24511);
nand UO_1739 (O_1739,N_24990,N_24641);
xor UO_1740 (O_1740,N_24556,N_23833);
nand UO_1741 (O_1741,N_24421,N_24076);
nor UO_1742 (O_1742,N_24616,N_24472);
and UO_1743 (O_1743,N_24697,N_24163);
xor UO_1744 (O_1744,N_23783,N_23844);
or UO_1745 (O_1745,N_24211,N_24568);
xor UO_1746 (O_1746,N_24552,N_24548);
and UO_1747 (O_1747,N_24331,N_23763);
nand UO_1748 (O_1748,N_24699,N_24665);
nand UO_1749 (O_1749,N_24974,N_24782);
or UO_1750 (O_1750,N_24911,N_24027);
nand UO_1751 (O_1751,N_23882,N_24104);
and UO_1752 (O_1752,N_24212,N_23897);
and UO_1753 (O_1753,N_23826,N_24478);
nor UO_1754 (O_1754,N_23975,N_24788);
nor UO_1755 (O_1755,N_24759,N_24782);
and UO_1756 (O_1756,N_24353,N_24455);
nor UO_1757 (O_1757,N_24459,N_23857);
or UO_1758 (O_1758,N_24206,N_24522);
xor UO_1759 (O_1759,N_23988,N_24282);
xor UO_1760 (O_1760,N_23909,N_24743);
nor UO_1761 (O_1761,N_24971,N_24233);
nand UO_1762 (O_1762,N_24720,N_23818);
and UO_1763 (O_1763,N_23769,N_24075);
or UO_1764 (O_1764,N_23875,N_24369);
or UO_1765 (O_1765,N_24794,N_24178);
xor UO_1766 (O_1766,N_23753,N_24010);
or UO_1767 (O_1767,N_24873,N_24233);
and UO_1768 (O_1768,N_24890,N_24577);
xnor UO_1769 (O_1769,N_24412,N_24602);
nor UO_1770 (O_1770,N_23877,N_24689);
xnor UO_1771 (O_1771,N_24598,N_24388);
nor UO_1772 (O_1772,N_24073,N_24633);
xnor UO_1773 (O_1773,N_23987,N_24561);
xnor UO_1774 (O_1774,N_24902,N_23908);
xor UO_1775 (O_1775,N_24426,N_24406);
and UO_1776 (O_1776,N_24163,N_24687);
xor UO_1777 (O_1777,N_24107,N_24537);
and UO_1778 (O_1778,N_24345,N_24527);
nor UO_1779 (O_1779,N_24321,N_24060);
nand UO_1780 (O_1780,N_24423,N_24561);
or UO_1781 (O_1781,N_24353,N_24088);
and UO_1782 (O_1782,N_24665,N_23750);
xor UO_1783 (O_1783,N_24739,N_24938);
nand UO_1784 (O_1784,N_24731,N_24860);
nor UO_1785 (O_1785,N_24389,N_24904);
nor UO_1786 (O_1786,N_24030,N_24640);
nor UO_1787 (O_1787,N_23876,N_24743);
and UO_1788 (O_1788,N_23947,N_24512);
xnor UO_1789 (O_1789,N_24838,N_24773);
and UO_1790 (O_1790,N_24815,N_24295);
or UO_1791 (O_1791,N_24820,N_24159);
nor UO_1792 (O_1792,N_24537,N_23843);
and UO_1793 (O_1793,N_24660,N_24974);
and UO_1794 (O_1794,N_24813,N_24771);
or UO_1795 (O_1795,N_24425,N_24149);
and UO_1796 (O_1796,N_24125,N_24680);
xor UO_1797 (O_1797,N_24665,N_23824);
or UO_1798 (O_1798,N_23756,N_23797);
nor UO_1799 (O_1799,N_24382,N_24635);
or UO_1800 (O_1800,N_24900,N_24853);
and UO_1801 (O_1801,N_24562,N_24693);
nor UO_1802 (O_1802,N_24996,N_24878);
nand UO_1803 (O_1803,N_24079,N_24559);
xnor UO_1804 (O_1804,N_24127,N_24663);
nand UO_1805 (O_1805,N_24474,N_24968);
xnor UO_1806 (O_1806,N_24768,N_24133);
nor UO_1807 (O_1807,N_24850,N_24656);
nor UO_1808 (O_1808,N_24459,N_23884);
or UO_1809 (O_1809,N_23861,N_24050);
nor UO_1810 (O_1810,N_24248,N_23754);
xor UO_1811 (O_1811,N_24738,N_24627);
nand UO_1812 (O_1812,N_24412,N_24291);
nand UO_1813 (O_1813,N_24383,N_24615);
nor UO_1814 (O_1814,N_24696,N_24890);
or UO_1815 (O_1815,N_24961,N_24138);
or UO_1816 (O_1816,N_24573,N_23909);
xor UO_1817 (O_1817,N_23842,N_23844);
xnor UO_1818 (O_1818,N_24651,N_24255);
nor UO_1819 (O_1819,N_24001,N_23906);
or UO_1820 (O_1820,N_24312,N_24464);
and UO_1821 (O_1821,N_24090,N_23957);
and UO_1822 (O_1822,N_24466,N_23876);
and UO_1823 (O_1823,N_24734,N_24562);
or UO_1824 (O_1824,N_24820,N_24847);
or UO_1825 (O_1825,N_24720,N_24809);
xor UO_1826 (O_1826,N_23802,N_24563);
nor UO_1827 (O_1827,N_24664,N_24846);
xor UO_1828 (O_1828,N_24185,N_24780);
xnor UO_1829 (O_1829,N_24635,N_24084);
xor UO_1830 (O_1830,N_24020,N_23909);
nand UO_1831 (O_1831,N_24869,N_24248);
or UO_1832 (O_1832,N_24596,N_24598);
or UO_1833 (O_1833,N_24615,N_24626);
xor UO_1834 (O_1834,N_24334,N_24492);
nand UO_1835 (O_1835,N_24267,N_24873);
nor UO_1836 (O_1836,N_23876,N_24814);
and UO_1837 (O_1837,N_24551,N_24791);
nor UO_1838 (O_1838,N_24219,N_23752);
xnor UO_1839 (O_1839,N_24067,N_24940);
xnor UO_1840 (O_1840,N_24361,N_24945);
and UO_1841 (O_1841,N_24260,N_24588);
nand UO_1842 (O_1842,N_24641,N_24163);
and UO_1843 (O_1843,N_24169,N_24817);
and UO_1844 (O_1844,N_24387,N_23961);
and UO_1845 (O_1845,N_24239,N_23924);
and UO_1846 (O_1846,N_24788,N_24374);
and UO_1847 (O_1847,N_24839,N_23750);
nor UO_1848 (O_1848,N_24560,N_24337);
or UO_1849 (O_1849,N_24170,N_24621);
or UO_1850 (O_1850,N_24863,N_24328);
nand UO_1851 (O_1851,N_23882,N_24759);
or UO_1852 (O_1852,N_24212,N_24933);
nor UO_1853 (O_1853,N_24211,N_24856);
nor UO_1854 (O_1854,N_24299,N_24818);
nand UO_1855 (O_1855,N_24336,N_24345);
or UO_1856 (O_1856,N_23923,N_24301);
xor UO_1857 (O_1857,N_24863,N_23864);
nand UO_1858 (O_1858,N_24878,N_24865);
and UO_1859 (O_1859,N_23903,N_24691);
xor UO_1860 (O_1860,N_24324,N_24998);
and UO_1861 (O_1861,N_24108,N_24995);
and UO_1862 (O_1862,N_24543,N_24280);
nor UO_1863 (O_1863,N_24478,N_24438);
nand UO_1864 (O_1864,N_24562,N_23835);
and UO_1865 (O_1865,N_24236,N_24516);
nand UO_1866 (O_1866,N_24093,N_23821);
or UO_1867 (O_1867,N_24847,N_24732);
or UO_1868 (O_1868,N_24257,N_24202);
or UO_1869 (O_1869,N_23951,N_24015);
and UO_1870 (O_1870,N_24221,N_24113);
or UO_1871 (O_1871,N_24114,N_24334);
xor UO_1872 (O_1872,N_24318,N_23824);
nor UO_1873 (O_1873,N_23789,N_24490);
nand UO_1874 (O_1874,N_24182,N_23909);
and UO_1875 (O_1875,N_24687,N_24989);
and UO_1876 (O_1876,N_24787,N_24363);
and UO_1877 (O_1877,N_23815,N_24423);
xnor UO_1878 (O_1878,N_23834,N_24112);
nand UO_1879 (O_1879,N_24700,N_24915);
xnor UO_1880 (O_1880,N_24453,N_23788);
xor UO_1881 (O_1881,N_23931,N_24669);
nor UO_1882 (O_1882,N_23780,N_24237);
xnor UO_1883 (O_1883,N_24747,N_24639);
xnor UO_1884 (O_1884,N_24107,N_24340);
nand UO_1885 (O_1885,N_24908,N_24865);
xnor UO_1886 (O_1886,N_23805,N_24040);
and UO_1887 (O_1887,N_24867,N_24779);
or UO_1888 (O_1888,N_24109,N_24413);
or UO_1889 (O_1889,N_24429,N_24741);
nor UO_1890 (O_1890,N_24401,N_24141);
nand UO_1891 (O_1891,N_24294,N_24824);
and UO_1892 (O_1892,N_23837,N_24807);
and UO_1893 (O_1893,N_24605,N_23988);
nor UO_1894 (O_1894,N_24893,N_24843);
or UO_1895 (O_1895,N_24687,N_24405);
nor UO_1896 (O_1896,N_24648,N_24227);
nor UO_1897 (O_1897,N_24184,N_24368);
and UO_1898 (O_1898,N_24774,N_24146);
nand UO_1899 (O_1899,N_24405,N_24748);
nor UO_1900 (O_1900,N_24054,N_23871);
and UO_1901 (O_1901,N_23813,N_24445);
nor UO_1902 (O_1902,N_24820,N_24854);
nand UO_1903 (O_1903,N_23999,N_24678);
nand UO_1904 (O_1904,N_24521,N_24142);
nand UO_1905 (O_1905,N_23963,N_24907);
and UO_1906 (O_1906,N_24664,N_24567);
or UO_1907 (O_1907,N_24882,N_24998);
and UO_1908 (O_1908,N_24867,N_24375);
and UO_1909 (O_1909,N_24505,N_24174);
nand UO_1910 (O_1910,N_24997,N_24886);
nor UO_1911 (O_1911,N_24285,N_24660);
nor UO_1912 (O_1912,N_24804,N_24950);
nand UO_1913 (O_1913,N_24630,N_23751);
nor UO_1914 (O_1914,N_24684,N_23979);
nand UO_1915 (O_1915,N_23933,N_24605);
xnor UO_1916 (O_1916,N_24182,N_24812);
or UO_1917 (O_1917,N_24620,N_23937);
or UO_1918 (O_1918,N_24779,N_24216);
nand UO_1919 (O_1919,N_24871,N_23986);
or UO_1920 (O_1920,N_24115,N_23755);
and UO_1921 (O_1921,N_23785,N_24657);
xor UO_1922 (O_1922,N_24909,N_23905);
nand UO_1923 (O_1923,N_24461,N_24082);
or UO_1924 (O_1924,N_24456,N_23777);
xnor UO_1925 (O_1925,N_24538,N_24365);
and UO_1926 (O_1926,N_24833,N_24947);
nor UO_1927 (O_1927,N_23794,N_24964);
nor UO_1928 (O_1928,N_23785,N_24958);
nand UO_1929 (O_1929,N_24388,N_24035);
nand UO_1930 (O_1930,N_24144,N_24509);
nor UO_1931 (O_1931,N_24988,N_24725);
nor UO_1932 (O_1932,N_23817,N_24414);
xor UO_1933 (O_1933,N_24191,N_24202);
and UO_1934 (O_1934,N_23821,N_24104);
nor UO_1935 (O_1935,N_24894,N_24996);
nand UO_1936 (O_1936,N_24261,N_23912);
or UO_1937 (O_1937,N_24375,N_24470);
and UO_1938 (O_1938,N_24264,N_24884);
nand UO_1939 (O_1939,N_24937,N_24474);
nor UO_1940 (O_1940,N_24895,N_24755);
and UO_1941 (O_1941,N_24594,N_24138);
and UO_1942 (O_1942,N_23905,N_24540);
or UO_1943 (O_1943,N_24201,N_24577);
and UO_1944 (O_1944,N_23858,N_24133);
or UO_1945 (O_1945,N_23838,N_24895);
nand UO_1946 (O_1946,N_24074,N_24125);
xnor UO_1947 (O_1947,N_24744,N_24434);
nor UO_1948 (O_1948,N_24874,N_24487);
and UO_1949 (O_1949,N_23924,N_23889);
nor UO_1950 (O_1950,N_24072,N_24524);
nor UO_1951 (O_1951,N_24767,N_24476);
or UO_1952 (O_1952,N_24627,N_24258);
nand UO_1953 (O_1953,N_24289,N_24964);
nand UO_1954 (O_1954,N_23956,N_24724);
xnor UO_1955 (O_1955,N_24815,N_24624);
and UO_1956 (O_1956,N_24740,N_24040);
nand UO_1957 (O_1957,N_24079,N_24694);
or UO_1958 (O_1958,N_24808,N_23953);
or UO_1959 (O_1959,N_24596,N_24933);
or UO_1960 (O_1960,N_24481,N_24271);
nand UO_1961 (O_1961,N_24938,N_23770);
and UO_1962 (O_1962,N_24337,N_24887);
and UO_1963 (O_1963,N_24926,N_24178);
xnor UO_1964 (O_1964,N_24906,N_23802);
xor UO_1965 (O_1965,N_23955,N_24827);
nor UO_1966 (O_1966,N_24920,N_24560);
nor UO_1967 (O_1967,N_24526,N_23947);
and UO_1968 (O_1968,N_24766,N_24364);
nand UO_1969 (O_1969,N_24152,N_23781);
xnor UO_1970 (O_1970,N_23886,N_24759);
nand UO_1971 (O_1971,N_23787,N_24761);
nand UO_1972 (O_1972,N_23948,N_24707);
or UO_1973 (O_1973,N_23776,N_24618);
nor UO_1974 (O_1974,N_24468,N_24198);
or UO_1975 (O_1975,N_24704,N_23918);
and UO_1976 (O_1976,N_24926,N_24102);
and UO_1977 (O_1977,N_24525,N_24729);
and UO_1978 (O_1978,N_24363,N_24131);
and UO_1979 (O_1979,N_24927,N_24123);
xor UO_1980 (O_1980,N_24783,N_24218);
xnor UO_1981 (O_1981,N_24982,N_24706);
xor UO_1982 (O_1982,N_24398,N_23868);
and UO_1983 (O_1983,N_24485,N_23946);
or UO_1984 (O_1984,N_24270,N_23901);
or UO_1985 (O_1985,N_24194,N_23896);
nand UO_1986 (O_1986,N_24035,N_24674);
xor UO_1987 (O_1987,N_24345,N_24656);
nand UO_1988 (O_1988,N_24025,N_24878);
nor UO_1989 (O_1989,N_24658,N_23994);
or UO_1990 (O_1990,N_24925,N_24445);
nand UO_1991 (O_1991,N_24977,N_24063);
or UO_1992 (O_1992,N_24941,N_24914);
and UO_1993 (O_1993,N_24781,N_24621);
nand UO_1994 (O_1994,N_24014,N_24740);
xnor UO_1995 (O_1995,N_24190,N_24433);
and UO_1996 (O_1996,N_24982,N_24151);
nor UO_1997 (O_1997,N_24352,N_24809);
xor UO_1998 (O_1998,N_24715,N_24152);
xor UO_1999 (O_1999,N_24871,N_24574);
nor UO_2000 (O_2000,N_24106,N_24919);
nand UO_2001 (O_2001,N_23902,N_23783);
nand UO_2002 (O_2002,N_23790,N_24651);
nand UO_2003 (O_2003,N_24907,N_23797);
or UO_2004 (O_2004,N_24456,N_23927);
or UO_2005 (O_2005,N_23789,N_24073);
or UO_2006 (O_2006,N_24790,N_23893);
nand UO_2007 (O_2007,N_24885,N_24897);
and UO_2008 (O_2008,N_24837,N_24396);
nand UO_2009 (O_2009,N_24464,N_24577);
or UO_2010 (O_2010,N_23828,N_24529);
nand UO_2011 (O_2011,N_24248,N_24250);
nand UO_2012 (O_2012,N_23877,N_24189);
and UO_2013 (O_2013,N_24558,N_23924);
xnor UO_2014 (O_2014,N_24122,N_24171);
nand UO_2015 (O_2015,N_24186,N_24884);
nand UO_2016 (O_2016,N_24888,N_23864);
and UO_2017 (O_2017,N_24733,N_24656);
and UO_2018 (O_2018,N_24573,N_24036);
xnor UO_2019 (O_2019,N_24030,N_24194);
or UO_2020 (O_2020,N_24224,N_24065);
nand UO_2021 (O_2021,N_24480,N_24609);
nand UO_2022 (O_2022,N_24356,N_24688);
or UO_2023 (O_2023,N_23864,N_24590);
and UO_2024 (O_2024,N_24006,N_24546);
and UO_2025 (O_2025,N_24745,N_24368);
nand UO_2026 (O_2026,N_24706,N_24877);
nor UO_2027 (O_2027,N_24369,N_24216);
nor UO_2028 (O_2028,N_24121,N_24390);
nor UO_2029 (O_2029,N_23875,N_24870);
nand UO_2030 (O_2030,N_23876,N_23800);
or UO_2031 (O_2031,N_23794,N_24435);
nor UO_2032 (O_2032,N_24352,N_24872);
nand UO_2033 (O_2033,N_24981,N_24157);
nor UO_2034 (O_2034,N_24197,N_23778);
nand UO_2035 (O_2035,N_24121,N_24844);
nand UO_2036 (O_2036,N_24931,N_24427);
nand UO_2037 (O_2037,N_24775,N_24686);
or UO_2038 (O_2038,N_24185,N_24191);
and UO_2039 (O_2039,N_24537,N_24162);
or UO_2040 (O_2040,N_24075,N_24450);
xor UO_2041 (O_2041,N_24623,N_24923);
nor UO_2042 (O_2042,N_24555,N_24629);
or UO_2043 (O_2043,N_24774,N_24703);
nor UO_2044 (O_2044,N_24331,N_24139);
xor UO_2045 (O_2045,N_24782,N_24080);
and UO_2046 (O_2046,N_23882,N_24934);
or UO_2047 (O_2047,N_24480,N_24667);
or UO_2048 (O_2048,N_24856,N_24471);
nor UO_2049 (O_2049,N_24776,N_23845);
or UO_2050 (O_2050,N_24895,N_24330);
and UO_2051 (O_2051,N_24628,N_24057);
and UO_2052 (O_2052,N_24502,N_24926);
or UO_2053 (O_2053,N_23892,N_23793);
nand UO_2054 (O_2054,N_24818,N_24177);
or UO_2055 (O_2055,N_24716,N_24641);
xnor UO_2056 (O_2056,N_24400,N_24360);
xor UO_2057 (O_2057,N_23834,N_24492);
and UO_2058 (O_2058,N_24595,N_24468);
or UO_2059 (O_2059,N_24458,N_23774);
xor UO_2060 (O_2060,N_24805,N_24043);
nor UO_2061 (O_2061,N_24495,N_24165);
nor UO_2062 (O_2062,N_24493,N_24976);
and UO_2063 (O_2063,N_24517,N_24375);
or UO_2064 (O_2064,N_24118,N_24614);
and UO_2065 (O_2065,N_24976,N_24960);
xor UO_2066 (O_2066,N_24083,N_24161);
or UO_2067 (O_2067,N_24091,N_23857);
and UO_2068 (O_2068,N_24095,N_24214);
and UO_2069 (O_2069,N_23951,N_23893);
and UO_2070 (O_2070,N_23908,N_24105);
xor UO_2071 (O_2071,N_24418,N_23890);
nand UO_2072 (O_2072,N_24156,N_24047);
and UO_2073 (O_2073,N_24548,N_24914);
nand UO_2074 (O_2074,N_24405,N_23923);
and UO_2075 (O_2075,N_24420,N_23955);
or UO_2076 (O_2076,N_24706,N_24957);
nand UO_2077 (O_2077,N_24734,N_23856);
xnor UO_2078 (O_2078,N_24566,N_24404);
and UO_2079 (O_2079,N_24356,N_24472);
nor UO_2080 (O_2080,N_24481,N_24334);
and UO_2081 (O_2081,N_24300,N_23760);
nand UO_2082 (O_2082,N_24501,N_23952);
nor UO_2083 (O_2083,N_24493,N_24039);
nor UO_2084 (O_2084,N_24242,N_24998);
xor UO_2085 (O_2085,N_24188,N_23859);
or UO_2086 (O_2086,N_24481,N_24734);
or UO_2087 (O_2087,N_24851,N_24232);
xor UO_2088 (O_2088,N_24606,N_24381);
nor UO_2089 (O_2089,N_23838,N_24903);
nor UO_2090 (O_2090,N_24996,N_23920);
xnor UO_2091 (O_2091,N_24655,N_24237);
nor UO_2092 (O_2092,N_23758,N_24998);
and UO_2093 (O_2093,N_24524,N_24423);
or UO_2094 (O_2094,N_24599,N_23900);
or UO_2095 (O_2095,N_24952,N_23880);
nor UO_2096 (O_2096,N_24661,N_24854);
nor UO_2097 (O_2097,N_24362,N_24189);
or UO_2098 (O_2098,N_24457,N_24186);
nand UO_2099 (O_2099,N_24562,N_24324);
and UO_2100 (O_2100,N_24652,N_23917);
nand UO_2101 (O_2101,N_23911,N_24577);
nand UO_2102 (O_2102,N_24705,N_24226);
xnor UO_2103 (O_2103,N_24414,N_24699);
or UO_2104 (O_2104,N_24050,N_24798);
xnor UO_2105 (O_2105,N_24185,N_24726);
xor UO_2106 (O_2106,N_24297,N_24042);
and UO_2107 (O_2107,N_23839,N_24143);
and UO_2108 (O_2108,N_24182,N_23857);
nor UO_2109 (O_2109,N_24846,N_23965);
nand UO_2110 (O_2110,N_24801,N_24017);
nor UO_2111 (O_2111,N_24274,N_24889);
or UO_2112 (O_2112,N_23986,N_24534);
xnor UO_2113 (O_2113,N_24281,N_24590);
or UO_2114 (O_2114,N_24512,N_24712);
or UO_2115 (O_2115,N_24013,N_24299);
or UO_2116 (O_2116,N_24047,N_24197);
xnor UO_2117 (O_2117,N_24986,N_23762);
or UO_2118 (O_2118,N_24305,N_24594);
nor UO_2119 (O_2119,N_24324,N_24589);
or UO_2120 (O_2120,N_24078,N_23750);
nand UO_2121 (O_2121,N_24515,N_24545);
nor UO_2122 (O_2122,N_24704,N_24726);
or UO_2123 (O_2123,N_24984,N_24084);
nand UO_2124 (O_2124,N_24002,N_24928);
and UO_2125 (O_2125,N_23992,N_24744);
or UO_2126 (O_2126,N_24150,N_24519);
nand UO_2127 (O_2127,N_23917,N_24542);
xor UO_2128 (O_2128,N_24542,N_24649);
nor UO_2129 (O_2129,N_23815,N_24460);
nand UO_2130 (O_2130,N_24666,N_23819);
and UO_2131 (O_2131,N_24250,N_24548);
nor UO_2132 (O_2132,N_24725,N_24822);
nand UO_2133 (O_2133,N_23770,N_23831);
nor UO_2134 (O_2134,N_24025,N_24430);
xnor UO_2135 (O_2135,N_24787,N_24018);
nor UO_2136 (O_2136,N_24920,N_23940);
xor UO_2137 (O_2137,N_24034,N_24138);
or UO_2138 (O_2138,N_24210,N_24581);
xor UO_2139 (O_2139,N_24552,N_24370);
xor UO_2140 (O_2140,N_24499,N_24039);
or UO_2141 (O_2141,N_24122,N_23947);
and UO_2142 (O_2142,N_24481,N_24461);
and UO_2143 (O_2143,N_23834,N_24714);
xnor UO_2144 (O_2144,N_24463,N_24017);
xnor UO_2145 (O_2145,N_24609,N_24523);
or UO_2146 (O_2146,N_24333,N_24340);
or UO_2147 (O_2147,N_24346,N_24132);
and UO_2148 (O_2148,N_24384,N_23796);
xnor UO_2149 (O_2149,N_24980,N_24451);
nor UO_2150 (O_2150,N_24337,N_24771);
and UO_2151 (O_2151,N_24036,N_24675);
or UO_2152 (O_2152,N_23971,N_24913);
nand UO_2153 (O_2153,N_23765,N_24707);
or UO_2154 (O_2154,N_24316,N_24591);
nand UO_2155 (O_2155,N_23821,N_24231);
nand UO_2156 (O_2156,N_24206,N_24105);
nor UO_2157 (O_2157,N_23809,N_24740);
nand UO_2158 (O_2158,N_24665,N_23765);
nand UO_2159 (O_2159,N_24305,N_24450);
nor UO_2160 (O_2160,N_24850,N_24945);
or UO_2161 (O_2161,N_24855,N_24586);
nor UO_2162 (O_2162,N_24201,N_24418);
or UO_2163 (O_2163,N_24630,N_24728);
nor UO_2164 (O_2164,N_24492,N_24880);
or UO_2165 (O_2165,N_23985,N_24777);
and UO_2166 (O_2166,N_23901,N_23812);
and UO_2167 (O_2167,N_24441,N_23812);
nor UO_2168 (O_2168,N_23921,N_24438);
and UO_2169 (O_2169,N_24440,N_24712);
nor UO_2170 (O_2170,N_24690,N_24126);
nor UO_2171 (O_2171,N_24573,N_24630);
nor UO_2172 (O_2172,N_24057,N_24032);
nand UO_2173 (O_2173,N_24794,N_24795);
or UO_2174 (O_2174,N_23873,N_24292);
nand UO_2175 (O_2175,N_24749,N_24203);
and UO_2176 (O_2176,N_24735,N_24773);
and UO_2177 (O_2177,N_24021,N_23930);
and UO_2178 (O_2178,N_24870,N_24320);
and UO_2179 (O_2179,N_24028,N_24035);
xnor UO_2180 (O_2180,N_24444,N_24096);
nand UO_2181 (O_2181,N_24833,N_24782);
nand UO_2182 (O_2182,N_24316,N_24925);
nand UO_2183 (O_2183,N_24838,N_24137);
and UO_2184 (O_2184,N_24120,N_24386);
or UO_2185 (O_2185,N_24317,N_24690);
nor UO_2186 (O_2186,N_24989,N_24619);
nor UO_2187 (O_2187,N_23774,N_24211);
and UO_2188 (O_2188,N_24934,N_24175);
or UO_2189 (O_2189,N_23775,N_24196);
xor UO_2190 (O_2190,N_24316,N_24843);
and UO_2191 (O_2191,N_23820,N_23960);
or UO_2192 (O_2192,N_24331,N_24736);
and UO_2193 (O_2193,N_24712,N_24114);
and UO_2194 (O_2194,N_24084,N_24787);
and UO_2195 (O_2195,N_23948,N_24885);
and UO_2196 (O_2196,N_24314,N_24241);
and UO_2197 (O_2197,N_24697,N_24653);
and UO_2198 (O_2198,N_23863,N_24156);
xnor UO_2199 (O_2199,N_23984,N_24986);
xor UO_2200 (O_2200,N_23925,N_23881);
or UO_2201 (O_2201,N_24157,N_24299);
xor UO_2202 (O_2202,N_24402,N_24618);
xnor UO_2203 (O_2203,N_24460,N_24174);
nor UO_2204 (O_2204,N_24544,N_24968);
nor UO_2205 (O_2205,N_24946,N_24536);
and UO_2206 (O_2206,N_24265,N_23854);
nand UO_2207 (O_2207,N_24828,N_24139);
or UO_2208 (O_2208,N_24178,N_23857);
or UO_2209 (O_2209,N_24929,N_24652);
nor UO_2210 (O_2210,N_23811,N_24549);
and UO_2211 (O_2211,N_24120,N_23975);
and UO_2212 (O_2212,N_24397,N_24462);
xnor UO_2213 (O_2213,N_24459,N_24360);
nand UO_2214 (O_2214,N_24762,N_24347);
nor UO_2215 (O_2215,N_24095,N_24176);
nor UO_2216 (O_2216,N_24195,N_24318);
nor UO_2217 (O_2217,N_24390,N_23779);
and UO_2218 (O_2218,N_24775,N_24819);
xnor UO_2219 (O_2219,N_24087,N_24877);
nor UO_2220 (O_2220,N_23832,N_23867);
or UO_2221 (O_2221,N_24018,N_24516);
xor UO_2222 (O_2222,N_24347,N_24493);
and UO_2223 (O_2223,N_24361,N_24458);
xnor UO_2224 (O_2224,N_24365,N_24631);
or UO_2225 (O_2225,N_24893,N_24427);
or UO_2226 (O_2226,N_24263,N_23979);
and UO_2227 (O_2227,N_24562,N_24876);
nor UO_2228 (O_2228,N_24768,N_23792);
nand UO_2229 (O_2229,N_24210,N_24715);
and UO_2230 (O_2230,N_24784,N_24928);
and UO_2231 (O_2231,N_24380,N_24850);
or UO_2232 (O_2232,N_24805,N_24314);
xor UO_2233 (O_2233,N_24385,N_24891);
and UO_2234 (O_2234,N_24545,N_23823);
nor UO_2235 (O_2235,N_24865,N_24821);
and UO_2236 (O_2236,N_24540,N_24264);
and UO_2237 (O_2237,N_24428,N_24174);
nand UO_2238 (O_2238,N_24434,N_24789);
nand UO_2239 (O_2239,N_23951,N_23878);
and UO_2240 (O_2240,N_24766,N_24217);
or UO_2241 (O_2241,N_24817,N_24373);
nor UO_2242 (O_2242,N_24248,N_24476);
nor UO_2243 (O_2243,N_23891,N_24654);
nor UO_2244 (O_2244,N_24486,N_24183);
nand UO_2245 (O_2245,N_23976,N_24547);
nand UO_2246 (O_2246,N_24690,N_24988);
and UO_2247 (O_2247,N_24489,N_24980);
or UO_2248 (O_2248,N_24855,N_24068);
nand UO_2249 (O_2249,N_24098,N_24587);
nor UO_2250 (O_2250,N_24275,N_23995);
xor UO_2251 (O_2251,N_24629,N_23991);
nand UO_2252 (O_2252,N_24404,N_24074);
and UO_2253 (O_2253,N_24192,N_24734);
and UO_2254 (O_2254,N_24192,N_24281);
xor UO_2255 (O_2255,N_24208,N_24613);
or UO_2256 (O_2256,N_24198,N_24877);
and UO_2257 (O_2257,N_24601,N_23774);
nor UO_2258 (O_2258,N_24803,N_23843);
xnor UO_2259 (O_2259,N_24744,N_23854);
or UO_2260 (O_2260,N_24333,N_24645);
nand UO_2261 (O_2261,N_24019,N_24672);
nor UO_2262 (O_2262,N_24463,N_24751);
or UO_2263 (O_2263,N_23916,N_24780);
or UO_2264 (O_2264,N_23851,N_24145);
xor UO_2265 (O_2265,N_24115,N_24191);
or UO_2266 (O_2266,N_24995,N_24030);
xnor UO_2267 (O_2267,N_23957,N_24700);
nor UO_2268 (O_2268,N_24382,N_23764);
and UO_2269 (O_2269,N_24468,N_23905);
and UO_2270 (O_2270,N_24006,N_24422);
or UO_2271 (O_2271,N_23825,N_24097);
and UO_2272 (O_2272,N_23907,N_24320);
nand UO_2273 (O_2273,N_24760,N_24765);
or UO_2274 (O_2274,N_24290,N_23885);
or UO_2275 (O_2275,N_24456,N_24622);
or UO_2276 (O_2276,N_24320,N_23752);
nor UO_2277 (O_2277,N_24918,N_24142);
nand UO_2278 (O_2278,N_24721,N_23848);
nor UO_2279 (O_2279,N_24363,N_24531);
nand UO_2280 (O_2280,N_24252,N_24072);
xor UO_2281 (O_2281,N_24688,N_24953);
nand UO_2282 (O_2282,N_24153,N_23811);
and UO_2283 (O_2283,N_23980,N_23888);
or UO_2284 (O_2284,N_24835,N_24893);
xnor UO_2285 (O_2285,N_23864,N_24988);
nand UO_2286 (O_2286,N_24669,N_24473);
and UO_2287 (O_2287,N_24791,N_24682);
and UO_2288 (O_2288,N_24845,N_24045);
xnor UO_2289 (O_2289,N_24081,N_23907);
or UO_2290 (O_2290,N_24947,N_24779);
nand UO_2291 (O_2291,N_24075,N_24033);
and UO_2292 (O_2292,N_24954,N_24222);
nand UO_2293 (O_2293,N_23912,N_24535);
xnor UO_2294 (O_2294,N_24107,N_24525);
nor UO_2295 (O_2295,N_24203,N_23791);
and UO_2296 (O_2296,N_24515,N_23841);
nand UO_2297 (O_2297,N_24955,N_24979);
or UO_2298 (O_2298,N_24055,N_24500);
nand UO_2299 (O_2299,N_24495,N_24548);
xnor UO_2300 (O_2300,N_23936,N_24468);
xor UO_2301 (O_2301,N_24670,N_24910);
nand UO_2302 (O_2302,N_23862,N_24799);
nand UO_2303 (O_2303,N_23784,N_23792);
and UO_2304 (O_2304,N_23757,N_23929);
nor UO_2305 (O_2305,N_24588,N_24900);
nand UO_2306 (O_2306,N_24857,N_24755);
nor UO_2307 (O_2307,N_24556,N_24859);
nor UO_2308 (O_2308,N_24033,N_24438);
and UO_2309 (O_2309,N_24165,N_23822);
nor UO_2310 (O_2310,N_24345,N_24202);
xnor UO_2311 (O_2311,N_24192,N_23835);
xor UO_2312 (O_2312,N_24270,N_24220);
nand UO_2313 (O_2313,N_24358,N_24468);
nor UO_2314 (O_2314,N_23784,N_24105);
xor UO_2315 (O_2315,N_24604,N_24834);
nand UO_2316 (O_2316,N_24983,N_24233);
xnor UO_2317 (O_2317,N_24726,N_24288);
nand UO_2318 (O_2318,N_24626,N_23907);
nor UO_2319 (O_2319,N_24912,N_24689);
nor UO_2320 (O_2320,N_24149,N_24125);
xnor UO_2321 (O_2321,N_24589,N_24254);
nor UO_2322 (O_2322,N_24471,N_23947);
and UO_2323 (O_2323,N_24666,N_23877);
or UO_2324 (O_2324,N_24517,N_24721);
xnor UO_2325 (O_2325,N_24518,N_24702);
nor UO_2326 (O_2326,N_24940,N_23751);
xnor UO_2327 (O_2327,N_24692,N_24188);
nand UO_2328 (O_2328,N_24875,N_24042);
xnor UO_2329 (O_2329,N_24994,N_24671);
and UO_2330 (O_2330,N_24066,N_23877);
xor UO_2331 (O_2331,N_24733,N_24616);
xor UO_2332 (O_2332,N_24240,N_24920);
nor UO_2333 (O_2333,N_24895,N_24099);
and UO_2334 (O_2334,N_24249,N_24706);
xor UO_2335 (O_2335,N_24057,N_24275);
nand UO_2336 (O_2336,N_23906,N_24702);
nor UO_2337 (O_2337,N_23945,N_24066);
or UO_2338 (O_2338,N_24705,N_24005);
nor UO_2339 (O_2339,N_23866,N_23768);
or UO_2340 (O_2340,N_24998,N_23876);
or UO_2341 (O_2341,N_24530,N_24536);
or UO_2342 (O_2342,N_24808,N_24789);
nor UO_2343 (O_2343,N_24687,N_24385);
or UO_2344 (O_2344,N_24065,N_23850);
xor UO_2345 (O_2345,N_24815,N_24758);
nand UO_2346 (O_2346,N_24536,N_24619);
nand UO_2347 (O_2347,N_23779,N_24798);
nor UO_2348 (O_2348,N_24948,N_23908);
nor UO_2349 (O_2349,N_24099,N_24816);
nand UO_2350 (O_2350,N_24052,N_23807);
nor UO_2351 (O_2351,N_23932,N_24748);
or UO_2352 (O_2352,N_24413,N_24905);
nand UO_2353 (O_2353,N_24479,N_24115);
xor UO_2354 (O_2354,N_24624,N_23949);
and UO_2355 (O_2355,N_24203,N_23862);
and UO_2356 (O_2356,N_24585,N_23931);
or UO_2357 (O_2357,N_24811,N_24682);
nand UO_2358 (O_2358,N_24915,N_23947);
and UO_2359 (O_2359,N_24183,N_24825);
and UO_2360 (O_2360,N_24092,N_24906);
nand UO_2361 (O_2361,N_23784,N_24335);
xnor UO_2362 (O_2362,N_24566,N_24351);
nor UO_2363 (O_2363,N_24608,N_24339);
and UO_2364 (O_2364,N_24644,N_24761);
or UO_2365 (O_2365,N_24133,N_24847);
nor UO_2366 (O_2366,N_24582,N_24091);
and UO_2367 (O_2367,N_24154,N_24447);
nand UO_2368 (O_2368,N_24556,N_23809);
or UO_2369 (O_2369,N_24516,N_24415);
xor UO_2370 (O_2370,N_24685,N_24626);
or UO_2371 (O_2371,N_23941,N_24756);
nand UO_2372 (O_2372,N_24036,N_23764);
and UO_2373 (O_2373,N_24314,N_24223);
nand UO_2374 (O_2374,N_24050,N_24070);
or UO_2375 (O_2375,N_23867,N_24158);
xor UO_2376 (O_2376,N_24400,N_24795);
nand UO_2377 (O_2377,N_24361,N_23815);
nor UO_2378 (O_2378,N_23801,N_24235);
and UO_2379 (O_2379,N_24129,N_24289);
nor UO_2380 (O_2380,N_24598,N_24407);
xor UO_2381 (O_2381,N_23980,N_24371);
nor UO_2382 (O_2382,N_24697,N_23990);
xor UO_2383 (O_2383,N_24826,N_24066);
nand UO_2384 (O_2384,N_23847,N_24989);
or UO_2385 (O_2385,N_23948,N_24307);
nand UO_2386 (O_2386,N_24020,N_24406);
xor UO_2387 (O_2387,N_24423,N_24472);
and UO_2388 (O_2388,N_24191,N_24581);
nand UO_2389 (O_2389,N_23947,N_24536);
or UO_2390 (O_2390,N_24952,N_24609);
or UO_2391 (O_2391,N_24007,N_24589);
nor UO_2392 (O_2392,N_24909,N_24713);
nand UO_2393 (O_2393,N_24274,N_24763);
nand UO_2394 (O_2394,N_24915,N_24787);
or UO_2395 (O_2395,N_24863,N_24652);
nand UO_2396 (O_2396,N_23993,N_24296);
nor UO_2397 (O_2397,N_24695,N_24434);
or UO_2398 (O_2398,N_24087,N_24335);
and UO_2399 (O_2399,N_24256,N_24377);
and UO_2400 (O_2400,N_24736,N_24150);
nand UO_2401 (O_2401,N_24197,N_23795);
and UO_2402 (O_2402,N_24865,N_24161);
nor UO_2403 (O_2403,N_24826,N_23840);
or UO_2404 (O_2404,N_24210,N_24378);
xnor UO_2405 (O_2405,N_23764,N_24246);
nand UO_2406 (O_2406,N_24309,N_24064);
xnor UO_2407 (O_2407,N_24626,N_24390);
xor UO_2408 (O_2408,N_24061,N_24979);
nand UO_2409 (O_2409,N_23948,N_23856);
or UO_2410 (O_2410,N_24185,N_24540);
nor UO_2411 (O_2411,N_23831,N_24522);
or UO_2412 (O_2412,N_24273,N_23979);
and UO_2413 (O_2413,N_24141,N_24806);
nor UO_2414 (O_2414,N_24904,N_24666);
nor UO_2415 (O_2415,N_23911,N_23819);
xnor UO_2416 (O_2416,N_24826,N_24407);
xnor UO_2417 (O_2417,N_24816,N_24007);
and UO_2418 (O_2418,N_24074,N_24814);
and UO_2419 (O_2419,N_23771,N_24787);
and UO_2420 (O_2420,N_24598,N_23926);
nand UO_2421 (O_2421,N_24686,N_23997);
and UO_2422 (O_2422,N_23898,N_23999);
and UO_2423 (O_2423,N_24198,N_23926);
and UO_2424 (O_2424,N_24369,N_24105);
and UO_2425 (O_2425,N_24943,N_24938);
nor UO_2426 (O_2426,N_24610,N_24810);
and UO_2427 (O_2427,N_24248,N_23942);
nor UO_2428 (O_2428,N_23919,N_24183);
nor UO_2429 (O_2429,N_24924,N_24723);
and UO_2430 (O_2430,N_24118,N_23781);
nor UO_2431 (O_2431,N_24844,N_23909);
or UO_2432 (O_2432,N_24256,N_24413);
or UO_2433 (O_2433,N_24653,N_24498);
nand UO_2434 (O_2434,N_24975,N_24887);
and UO_2435 (O_2435,N_24259,N_24326);
nor UO_2436 (O_2436,N_24647,N_24125);
or UO_2437 (O_2437,N_24588,N_24421);
and UO_2438 (O_2438,N_24121,N_23862);
and UO_2439 (O_2439,N_23772,N_24394);
or UO_2440 (O_2440,N_24927,N_24966);
nor UO_2441 (O_2441,N_23758,N_24720);
nor UO_2442 (O_2442,N_24962,N_23806);
xnor UO_2443 (O_2443,N_24370,N_24275);
xnor UO_2444 (O_2444,N_24223,N_24354);
and UO_2445 (O_2445,N_24275,N_24148);
nor UO_2446 (O_2446,N_24232,N_24294);
nand UO_2447 (O_2447,N_24080,N_24012);
and UO_2448 (O_2448,N_23783,N_23969);
and UO_2449 (O_2449,N_24165,N_24245);
nand UO_2450 (O_2450,N_24480,N_24424);
nor UO_2451 (O_2451,N_24704,N_24517);
and UO_2452 (O_2452,N_23955,N_24663);
xnor UO_2453 (O_2453,N_24918,N_24340);
or UO_2454 (O_2454,N_24030,N_23837);
nand UO_2455 (O_2455,N_24096,N_24689);
nand UO_2456 (O_2456,N_24281,N_24939);
xor UO_2457 (O_2457,N_24122,N_24204);
nor UO_2458 (O_2458,N_24523,N_23873);
xnor UO_2459 (O_2459,N_24042,N_24851);
nand UO_2460 (O_2460,N_24335,N_24793);
nor UO_2461 (O_2461,N_24020,N_24945);
or UO_2462 (O_2462,N_24044,N_24322);
and UO_2463 (O_2463,N_24286,N_24787);
nor UO_2464 (O_2464,N_24956,N_24073);
or UO_2465 (O_2465,N_24406,N_24015);
and UO_2466 (O_2466,N_24972,N_24269);
nor UO_2467 (O_2467,N_24334,N_24777);
nand UO_2468 (O_2468,N_24822,N_24858);
and UO_2469 (O_2469,N_23991,N_24390);
and UO_2470 (O_2470,N_24140,N_24982);
and UO_2471 (O_2471,N_24253,N_24488);
nand UO_2472 (O_2472,N_23790,N_24263);
and UO_2473 (O_2473,N_23986,N_24512);
nand UO_2474 (O_2474,N_24220,N_24336);
and UO_2475 (O_2475,N_24133,N_24631);
nand UO_2476 (O_2476,N_24691,N_24633);
nand UO_2477 (O_2477,N_24327,N_24833);
xnor UO_2478 (O_2478,N_24914,N_24970);
nand UO_2479 (O_2479,N_24975,N_24659);
nand UO_2480 (O_2480,N_24319,N_23767);
xnor UO_2481 (O_2481,N_23933,N_24853);
nand UO_2482 (O_2482,N_24213,N_24932);
xor UO_2483 (O_2483,N_24360,N_24782);
or UO_2484 (O_2484,N_24768,N_24654);
or UO_2485 (O_2485,N_24070,N_23977);
xor UO_2486 (O_2486,N_24842,N_23796);
or UO_2487 (O_2487,N_24534,N_24202);
nand UO_2488 (O_2488,N_24349,N_24411);
xnor UO_2489 (O_2489,N_24266,N_24380);
nor UO_2490 (O_2490,N_24516,N_23986);
xnor UO_2491 (O_2491,N_23804,N_24900);
or UO_2492 (O_2492,N_23993,N_24964);
nor UO_2493 (O_2493,N_24176,N_24092);
xnor UO_2494 (O_2494,N_24255,N_24228);
nor UO_2495 (O_2495,N_24000,N_24135);
nor UO_2496 (O_2496,N_23881,N_24744);
nor UO_2497 (O_2497,N_24569,N_24582);
or UO_2498 (O_2498,N_24233,N_24461);
and UO_2499 (O_2499,N_24748,N_24765);
or UO_2500 (O_2500,N_24677,N_24824);
nand UO_2501 (O_2501,N_23974,N_24824);
xor UO_2502 (O_2502,N_24580,N_23924);
and UO_2503 (O_2503,N_24827,N_24183);
xor UO_2504 (O_2504,N_23825,N_23977);
nor UO_2505 (O_2505,N_24406,N_24526);
nand UO_2506 (O_2506,N_24705,N_24681);
nor UO_2507 (O_2507,N_24533,N_24543);
xor UO_2508 (O_2508,N_24832,N_24815);
and UO_2509 (O_2509,N_23991,N_23870);
nor UO_2510 (O_2510,N_24539,N_23990);
and UO_2511 (O_2511,N_24401,N_24266);
or UO_2512 (O_2512,N_24004,N_24451);
xor UO_2513 (O_2513,N_24372,N_24674);
or UO_2514 (O_2514,N_24453,N_24530);
and UO_2515 (O_2515,N_24276,N_24564);
and UO_2516 (O_2516,N_24434,N_23850);
nand UO_2517 (O_2517,N_24182,N_24924);
or UO_2518 (O_2518,N_24068,N_24059);
xor UO_2519 (O_2519,N_24282,N_24732);
nand UO_2520 (O_2520,N_24722,N_24571);
or UO_2521 (O_2521,N_24752,N_24073);
and UO_2522 (O_2522,N_24761,N_24950);
or UO_2523 (O_2523,N_24384,N_24672);
nand UO_2524 (O_2524,N_23873,N_24842);
or UO_2525 (O_2525,N_24418,N_24934);
nand UO_2526 (O_2526,N_24727,N_23814);
nor UO_2527 (O_2527,N_24978,N_24639);
nand UO_2528 (O_2528,N_24413,N_24182);
and UO_2529 (O_2529,N_23882,N_24991);
nand UO_2530 (O_2530,N_24252,N_24861);
and UO_2531 (O_2531,N_24814,N_24385);
and UO_2532 (O_2532,N_23813,N_24668);
nor UO_2533 (O_2533,N_24590,N_24309);
and UO_2534 (O_2534,N_24419,N_23993);
nor UO_2535 (O_2535,N_24065,N_24412);
nand UO_2536 (O_2536,N_24663,N_24096);
or UO_2537 (O_2537,N_24609,N_24835);
nand UO_2538 (O_2538,N_24480,N_24571);
nand UO_2539 (O_2539,N_24668,N_23810);
nor UO_2540 (O_2540,N_24630,N_24930);
or UO_2541 (O_2541,N_23795,N_23981);
xnor UO_2542 (O_2542,N_24433,N_24694);
or UO_2543 (O_2543,N_24914,N_24500);
or UO_2544 (O_2544,N_24649,N_24619);
nor UO_2545 (O_2545,N_24621,N_24822);
and UO_2546 (O_2546,N_24219,N_24659);
xor UO_2547 (O_2547,N_24062,N_24624);
nor UO_2548 (O_2548,N_24480,N_24566);
nor UO_2549 (O_2549,N_23970,N_24379);
nand UO_2550 (O_2550,N_24950,N_24080);
or UO_2551 (O_2551,N_24261,N_24996);
xor UO_2552 (O_2552,N_24868,N_24468);
or UO_2553 (O_2553,N_24679,N_24238);
xor UO_2554 (O_2554,N_23845,N_24414);
nor UO_2555 (O_2555,N_24743,N_24467);
xor UO_2556 (O_2556,N_24438,N_24535);
nor UO_2557 (O_2557,N_24739,N_24033);
xnor UO_2558 (O_2558,N_24358,N_24793);
nand UO_2559 (O_2559,N_24932,N_24983);
nor UO_2560 (O_2560,N_24255,N_24755);
or UO_2561 (O_2561,N_24304,N_23885);
and UO_2562 (O_2562,N_24205,N_23931);
and UO_2563 (O_2563,N_24646,N_24576);
or UO_2564 (O_2564,N_24974,N_23935);
nor UO_2565 (O_2565,N_24276,N_24727);
xor UO_2566 (O_2566,N_24406,N_24790);
nor UO_2567 (O_2567,N_24141,N_24758);
and UO_2568 (O_2568,N_23859,N_24844);
xnor UO_2569 (O_2569,N_24810,N_23953);
or UO_2570 (O_2570,N_24804,N_24875);
and UO_2571 (O_2571,N_24109,N_24157);
and UO_2572 (O_2572,N_23755,N_23945);
or UO_2573 (O_2573,N_24175,N_24310);
and UO_2574 (O_2574,N_24719,N_24014);
nand UO_2575 (O_2575,N_24146,N_24172);
and UO_2576 (O_2576,N_24030,N_24905);
nor UO_2577 (O_2577,N_23980,N_24606);
and UO_2578 (O_2578,N_23947,N_23986);
xnor UO_2579 (O_2579,N_23834,N_24003);
nand UO_2580 (O_2580,N_24794,N_23963);
nor UO_2581 (O_2581,N_24784,N_24373);
nand UO_2582 (O_2582,N_24104,N_24851);
nor UO_2583 (O_2583,N_24045,N_23917);
xor UO_2584 (O_2584,N_24412,N_24933);
and UO_2585 (O_2585,N_24820,N_23935);
or UO_2586 (O_2586,N_24540,N_23856);
nand UO_2587 (O_2587,N_23808,N_24955);
nand UO_2588 (O_2588,N_24502,N_24444);
and UO_2589 (O_2589,N_23829,N_24742);
nor UO_2590 (O_2590,N_24364,N_24004);
xnor UO_2591 (O_2591,N_24134,N_23945);
or UO_2592 (O_2592,N_24988,N_24616);
nor UO_2593 (O_2593,N_24023,N_24695);
nand UO_2594 (O_2594,N_23957,N_24600);
nand UO_2595 (O_2595,N_23868,N_24514);
nand UO_2596 (O_2596,N_24531,N_24960);
nor UO_2597 (O_2597,N_24609,N_24501);
or UO_2598 (O_2598,N_24729,N_24361);
or UO_2599 (O_2599,N_24817,N_24185);
nor UO_2600 (O_2600,N_24243,N_24119);
nand UO_2601 (O_2601,N_24952,N_24706);
and UO_2602 (O_2602,N_23896,N_24165);
nor UO_2603 (O_2603,N_24138,N_24770);
and UO_2604 (O_2604,N_23846,N_24445);
nand UO_2605 (O_2605,N_24921,N_24276);
or UO_2606 (O_2606,N_24180,N_24507);
nor UO_2607 (O_2607,N_24914,N_24913);
and UO_2608 (O_2608,N_24778,N_24426);
and UO_2609 (O_2609,N_23798,N_24399);
nor UO_2610 (O_2610,N_23780,N_24057);
and UO_2611 (O_2611,N_24764,N_24237);
and UO_2612 (O_2612,N_24552,N_24925);
xor UO_2613 (O_2613,N_24533,N_24879);
nand UO_2614 (O_2614,N_23823,N_23970);
or UO_2615 (O_2615,N_24392,N_23899);
or UO_2616 (O_2616,N_24492,N_23801);
and UO_2617 (O_2617,N_24180,N_23948);
nor UO_2618 (O_2618,N_24327,N_23766);
xor UO_2619 (O_2619,N_24632,N_24267);
or UO_2620 (O_2620,N_24002,N_23865);
and UO_2621 (O_2621,N_24290,N_24017);
nand UO_2622 (O_2622,N_24641,N_24612);
nand UO_2623 (O_2623,N_24784,N_23885);
nand UO_2624 (O_2624,N_24898,N_24810);
nand UO_2625 (O_2625,N_24359,N_24879);
nor UO_2626 (O_2626,N_24064,N_24807);
and UO_2627 (O_2627,N_23767,N_24877);
nand UO_2628 (O_2628,N_24153,N_24046);
xnor UO_2629 (O_2629,N_24299,N_24745);
or UO_2630 (O_2630,N_24458,N_23969);
nand UO_2631 (O_2631,N_23932,N_24146);
or UO_2632 (O_2632,N_24115,N_24228);
or UO_2633 (O_2633,N_24089,N_24938);
and UO_2634 (O_2634,N_24426,N_24582);
xor UO_2635 (O_2635,N_23868,N_23954);
xor UO_2636 (O_2636,N_24042,N_24587);
or UO_2637 (O_2637,N_24541,N_24749);
or UO_2638 (O_2638,N_24770,N_24340);
nand UO_2639 (O_2639,N_24061,N_24586);
or UO_2640 (O_2640,N_24508,N_24024);
or UO_2641 (O_2641,N_24649,N_23981);
nor UO_2642 (O_2642,N_24977,N_24548);
xnor UO_2643 (O_2643,N_24956,N_24294);
and UO_2644 (O_2644,N_24040,N_24899);
xnor UO_2645 (O_2645,N_24271,N_24717);
nand UO_2646 (O_2646,N_24519,N_24010);
xnor UO_2647 (O_2647,N_24715,N_24386);
or UO_2648 (O_2648,N_24147,N_23916);
and UO_2649 (O_2649,N_24517,N_24269);
nor UO_2650 (O_2650,N_24667,N_24790);
or UO_2651 (O_2651,N_24237,N_24528);
or UO_2652 (O_2652,N_24612,N_24607);
and UO_2653 (O_2653,N_23783,N_24326);
nand UO_2654 (O_2654,N_24051,N_24322);
and UO_2655 (O_2655,N_24869,N_24752);
or UO_2656 (O_2656,N_24009,N_24175);
or UO_2657 (O_2657,N_24800,N_24194);
and UO_2658 (O_2658,N_24657,N_24920);
or UO_2659 (O_2659,N_24098,N_23777);
or UO_2660 (O_2660,N_23959,N_24056);
and UO_2661 (O_2661,N_23890,N_24245);
and UO_2662 (O_2662,N_24231,N_24105);
or UO_2663 (O_2663,N_24141,N_24178);
and UO_2664 (O_2664,N_24713,N_24006);
nor UO_2665 (O_2665,N_24373,N_24435);
or UO_2666 (O_2666,N_24832,N_24378);
nor UO_2667 (O_2667,N_24463,N_23938);
xor UO_2668 (O_2668,N_23884,N_24371);
nor UO_2669 (O_2669,N_24015,N_24853);
and UO_2670 (O_2670,N_24397,N_23797);
nand UO_2671 (O_2671,N_24220,N_23866);
or UO_2672 (O_2672,N_24111,N_23997);
and UO_2673 (O_2673,N_24896,N_23913);
and UO_2674 (O_2674,N_24208,N_23770);
xor UO_2675 (O_2675,N_24955,N_23780);
xor UO_2676 (O_2676,N_24198,N_24711);
nand UO_2677 (O_2677,N_24545,N_24470);
xnor UO_2678 (O_2678,N_24331,N_23782);
and UO_2679 (O_2679,N_24272,N_23853);
and UO_2680 (O_2680,N_23952,N_24129);
nor UO_2681 (O_2681,N_24819,N_23779);
nand UO_2682 (O_2682,N_24099,N_23773);
and UO_2683 (O_2683,N_24417,N_24598);
nand UO_2684 (O_2684,N_23803,N_24629);
xor UO_2685 (O_2685,N_24144,N_24580);
nor UO_2686 (O_2686,N_24588,N_24901);
xor UO_2687 (O_2687,N_24071,N_24550);
or UO_2688 (O_2688,N_24202,N_24268);
xnor UO_2689 (O_2689,N_24059,N_24883);
xor UO_2690 (O_2690,N_24724,N_24529);
xor UO_2691 (O_2691,N_24238,N_24863);
xnor UO_2692 (O_2692,N_24575,N_23763);
and UO_2693 (O_2693,N_24382,N_24984);
xnor UO_2694 (O_2694,N_24023,N_24806);
xnor UO_2695 (O_2695,N_24431,N_24904);
or UO_2696 (O_2696,N_24038,N_23989);
and UO_2697 (O_2697,N_24481,N_24666);
and UO_2698 (O_2698,N_24482,N_24656);
nor UO_2699 (O_2699,N_23828,N_24344);
or UO_2700 (O_2700,N_24769,N_23787);
xor UO_2701 (O_2701,N_24971,N_24351);
nor UO_2702 (O_2702,N_24704,N_24930);
or UO_2703 (O_2703,N_23942,N_24032);
or UO_2704 (O_2704,N_23750,N_24580);
xnor UO_2705 (O_2705,N_23774,N_24959);
nand UO_2706 (O_2706,N_24314,N_24301);
or UO_2707 (O_2707,N_24322,N_23837);
xnor UO_2708 (O_2708,N_24089,N_23772);
or UO_2709 (O_2709,N_24323,N_23763);
or UO_2710 (O_2710,N_23803,N_24027);
nor UO_2711 (O_2711,N_24328,N_24707);
nand UO_2712 (O_2712,N_24063,N_24180);
xnor UO_2713 (O_2713,N_24334,N_24799);
or UO_2714 (O_2714,N_24742,N_24904);
xnor UO_2715 (O_2715,N_24136,N_24876);
nand UO_2716 (O_2716,N_24346,N_24452);
nor UO_2717 (O_2717,N_24830,N_23847);
nor UO_2718 (O_2718,N_24501,N_24836);
and UO_2719 (O_2719,N_24791,N_24237);
nand UO_2720 (O_2720,N_24716,N_24656);
nor UO_2721 (O_2721,N_24164,N_24434);
xor UO_2722 (O_2722,N_24638,N_23859);
nand UO_2723 (O_2723,N_24099,N_24668);
xnor UO_2724 (O_2724,N_24472,N_23897);
and UO_2725 (O_2725,N_24510,N_24685);
and UO_2726 (O_2726,N_23927,N_24738);
nor UO_2727 (O_2727,N_24607,N_24534);
and UO_2728 (O_2728,N_24555,N_24463);
or UO_2729 (O_2729,N_24959,N_23944);
and UO_2730 (O_2730,N_24438,N_24503);
or UO_2731 (O_2731,N_24252,N_24956);
or UO_2732 (O_2732,N_24723,N_24494);
or UO_2733 (O_2733,N_23860,N_24611);
or UO_2734 (O_2734,N_24077,N_24822);
xor UO_2735 (O_2735,N_24473,N_24559);
or UO_2736 (O_2736,N_24246,N_24358);
nand UO_2737 (O_2737,N_24268,N_23947);
nand UO_2738 (O_2738,N_24695,N_24502);
nor UO_2739 (O_2739,N_24479,N_24428);
xor UO_2740 (O_2740,N_23913,N_24699);
or UO_2741 (O_2741,N_24764,N_24055);
nand UO_2742 (O_2742,N_23996,N_23948);
nor UO_2743 (O_2743,N_24122,N_23782);
or UO_2744 (O_2744,N_24952,N_23995);
or UO_2745 (O_2745,N_24837,N_24791);
nor UO_2746 (O_2746,N_24184,N_24182);
xnor UO_2747 (O_2747,N_24137,N_23846);
nand UO_2748 (O_2748,N_24455,N_23954);
xor UO_2749 (O_2749,N_24757,N_23908);
or UO_2750 (O_2750,N_24218,N_24052);
or UO_2751 (O_2751,N_23788,N_23858);
and UO_2752 (O_2752,N_23768,N_24084);
nand UO_2753 (O_2753,N_24659,N_24200);
nor UO_2754 (O_2754,N_24734,N_24603);
xor UO_2755 (O_2755,N_24045,N_24910);
and UO_2756 (O_2756,N_24592,N_24145);
or UO_2757 (O_2757,N_24491,N_24136);
xnor UO_2758 (O_2758,N_24615,N_23906);
nor UO_2759 (O_2759,N_24372,N_23953);
nand UO_2760 (O_2760,N_24494,N_23882);
xor UO_2761 (O_2761,N_24885,N_23958);
and UO_2762 (O_2762,N_24680,N_24246);
and UO_2763 (O_2763,N_24944,N_24925);
or UO_2764 (O_2764,N_24458,N_24536);
and UO_2765 (O_2765,N_24467,N_24701);
or UO_2766 (O_2766,N_24854,N_24842);
or UO_2767 (O_2767,N_24068,N_24363);
and UO_2768 (O_2768,N_24995,N_24923);
nor UO_2769 (O_2769,N_24925,N_23913);
and UO_2770 (O_2770,N_24420,N_23838);
nand UO_2771 (O_2771,N_24662,N_24598);
nor UO_2772 (O_2772,N_24797,N_24662);
and UO_2773 (O_2773,N_24587,N_24033);
and UO_2774 (O_2774,N_24922,N_24823);
xor UO_2775 (O_2775,N_24968,N_24244);
and UO_2776 (O_2776,N_24429,N_24887);
nor UO_2777 (O_2777,N_24902,N_23894);
xnor UO_2778 (O_2778,N_24582,N_24243);
or UO_2779 (O_2779,N_24062,N_24597);
or UO_2780 (O_2780,N_24802,N_24397);
xor UO_2781 (O_2781,N_24226,N_24831);
nand UO_2782 (O_2782,N_24700,N_24221);
or UO_2783 (O_2783,N_24725,N_24308);
nor UO_2784 (O_2784,N_23899,N_24854);
or UO_2785 (O_2785,N_24720,N_24591);
or UO_2786 (O_2786,N_23900,N_24324);
nor UO_2787 (O_2787,N_24190,N_24294);
and UO_2788 (O_2788,N_24605,N_24289);
nor UO_2789 (O_2789,N_24283,N_24653);
nand UO_2790 (O_2790,N_23802,N_24524);
nand UO_2791 (O_2791,N_24828,N_23894);
nand UO_2792 (O_2792,N_24397,N_24557);
and UO_2793 (O_2793,N_23755,N_24543);
nand UO_2794 (O_2794,N_24265,N_24376);
and UO_2795 (O_2795,N_24220,N_24487);
and UO_2796 (O_2796,N_24752,N_24541);
xnor UO_2797 (O_2797,N_24500,N_24879);
nor UO_2798 (O_2798,N_24999,N_24432);
nand UO_2799 (O_2799,N_23757,N_24579);
or UO_2800 (O_2800,N_24660,N_23794);
or UO_2801 (O_2801,N_24339,N_23857);
xnor UO_2802 (O_2802,N_24265,N_24427);
or UO_2803 (O_2803,N_24991,N_24047);
or UO_2804 (O_2804,N_24150,N_24589);
nand UO_2805 (O_2805,N_24158,N_24250);
nand UO_2806 (O_2806,N_24773,N_24498);
nor UO_2807 (O_2807,N_23905,N_23968);
nor UO_2808 (O_2808,N_24712,N_24730);
nor UO_2809 (O_2809,N_24581,N_24955);
xnor UO_2810 (O_2810,N_24770,N_23884);
nand UO_2811 (O_2811,N_23908,N_24230);
xnor UO_2812 (O_2812,N_24998,N_24539);
xnor UO_2813 (O_2813,N_23816,N_24681);
and UO_2814 (O_2814,N_24093,N_24149);
or UO_2815 (O_2815,N_23835,N_24855);
and UO_2816 (O_2816,N_24970,N_24261);
and UO_2817 (O_2817,N_24601,N_24194);
xnor UO_2818 (O_2818,N_24894,N_24167);
nor UO_2819 (O_2819,N_24721,N_24045);
nor UO_2820 (O_2820,N_24150,N_24467);
or UO_2821 (O_2821,N_24932,N_24711);
and UO_2822 (O_2822,N_24820,N_24014);
nand UO_2823 (O_2823,N_23883,N_24872);
or UO_2824 (O_2824,N_24286,N_24179);
or UO_2825 (O_2825,N_24871,N_24629);
nand UO_2826 (O_2826,N_24222,N_24735);
xor UO_2827 (O_2827,N_24962,N_24457);
xor UO_2828 (O_2828,N_24805,N_23905);
and UO_2829 (O_2829,N_24985,N_24080);
nor UO_2830 (O_2830,N_24778,N_23997);
or UO_2831 (O_2831,N_24883,N_24563);
and UO_2832 (O_2832,N_24876,N_24084);
nor UO_2833 (O_2833,N_23824,N_24006);
nor UO_2834 (O_2834,N_24005,N_24678);
and UO_2835 (O_2835,N_24761,N_24589);
xnor UO_2836 (O_2836,N_24047,N_24976);
or UO_2837 (O_2837,N_24166,N_24361);
and UO_2838 (O_2838,N_23751,N_24893);
nand UO_2839 (O_2839,N_24063,N_24070);
or UO_2840 (O_2840,N_23934,N_23926);
nand UO_2841 (O_2841,N_24655,N_24704);
nor UO_2842 (O_2842,N_24913,N_24967);
nand UO_2843 (O_2843,N_24200,N_24120);
and UO_2844 (O_2844,N_24012,N_24830);
xor UO_2845 (O_2845,N_23917,N_24244);
or UO_2846 (O_2846,N_23912,N_24856);
xor UO_2847 (O_2847,N_24270,N_24340);
xnor UO_2848 (O_2848,N_24517,N_24176);
and UO_2849 (O_2849,N_24650,N_23791);
or UO_2850 (O_2850,N_24240,N_23962);
nor UO_2851 (O_2851,N_24087,N_24414);
xor UO_2852 (O_2852,N_24255,N_24442);
nor UO_2853 (O_2853,N_23932,N_24690);
xnor UO_2854 (O_2854,N_24014,N_24446);
xor UO_2855 (O_2855,N_24472,N_23756);
nor UO_2856 (O_2856,N_24648,N_24418);
and UO_2857 (O_2857,N_23844,N_24517);
nand UO_2858 (O_2858,N_24417,N_24152);
and UO_2859 (O_2859,N_24624,N_23785);
or UO_2860 (O_2860,N_24183,N_24966);
xor UO_2861 (O_2861,N_24867,N_24510);
or UO_2862 (O_2862,N_24722,N_24736);
xor UO_2863 (O_2863,N_24739,N_24501);
nor UO_2864 (O_2864,N_24795,N_24090);
nand UO_2865 (O_2865,N_24320,N_24901);
and UO_2866 (O_2866,N_24669,N_23817);
nand UO_2867 (O_2867,N_24632,N_24574);
xnor UO_2868 (O_2868,N_24152,N_24467);
or UO_2869 (O_2869,N_24699,N_24820);
or UO_2870 (O_2870,N_23905,N_23849);
xor UO_2871 (O_2871,N_24055,N_23759);
nor UO_2872 (O_2872,N_24421,N_24169);
and UO_2873 (O_2873,N_24933,N_24734);
nor UO_2874 (O_2874,N_24466,N_24136);
nand UO_2875 (O_2875,N_24468,N_24765);
nor UO_2876 (O_2876,N_24076,N_23952);
nand UO_2877 (O_2877,N_24303,N_24609);
and UO_2878 (O_2878,N_24406,N_24435);
xnor UO_2879 (O_2879,N_24892,N_24483);
or UO_2880 (O_2880,N_24915,N_24636);
nor UO_2881 (O_2881,N_24507,N_24172);
or UO_2882 (O_2882,N_24342,N_23976);
or UO_2883 (O_2883,N_24346,N_24683);
nor UO_2884 (O_2884,N_23783,N_24252);
xor UO_2885 (O_2885,N_24120,N_24203);
or UO_2886 (O_2886,N_24126,N_23837);
nand UO_2887 (O_2887,N_23939,N_24245);
or UO_2888 (O_2888,N_23841,N_23812);
xnor UO_2889 (O_2889,N_24211,N_24304);
or UO_2890 (O_2890,N_23966,N_24943);
nor UO_2891 (O_2891,N_24220,N_23884);
and UO_2892 (O_2892,N_24125,N_24201);
or UO_2893 (O_2893,N_23836,N_24929);
nand UO_2894 (O_2894,N_23788,N_24255);
xnor UO_2895 (O_2895,N_24864,N_24884);
nand UO_2896 (O_2896,N_24946,N_23925);
nand UO_2897 (O_2897,N_24561,N_24788);
nor UO_2898 (O_2898,N_24435,N_24083);
and UO_2899 (O_2899,N_23816,N_24004);
and UO_2900 (O_2900,N_24673,N_24450);
nand UO_2901 (O_2901,N_24295,N_24603);
and UO_2902 (O_2902,N_24079,N_24751);
nand UO_2903 (O_2903,N_24881,N_24607);
or UO_2904 (O_2904,N_24565,N_24652);
or UO_2905 (O_2905,N_24318,N_23758);
nand UO_2906 (O_2906,N_24058,N_23811);
and UO_2907 (O_2907,N_24364,N_23960);
nand UO_2908 (O_2908,N_24802,N_24767);
nor UO_2909 (O_2909,N_24651,N_24342);
nor UO_2910 (O_2910,N_23939,N_24244);
nor UO_2911 (O_2911,N_23844,N_24797);
nor UO_2912 (O_2912,N_24210,N_24941);
or UO_2913 (O_2913,N_24446,N_24642);
and UO_2914 (O_2914,N_23842,N_24540);
or UO_2915 (O_2915,N_24239,N_24977);
xor UO_2916 (O_2916,N_24523,N_24217);
xnor UO_2917 (O_2917,N_24434,N_23990);
nand UO_2918 (O_2918,N_24790,N_24997);
or UO_2919 (O_2919,N_24968,N_24825);
or UO_2920 (O_2920,N_24617,N_23801);
nor UO_2921 (O_2921,N_24486,N_23773);
nand UO_2922 (O_2922,N_24191,N_23982);
and UO_2923 (O_2923,N_24804,N_24818);
nand UO_2924 (O_2924,N_24773,N_24334);
nor UO_2925 (O_2925,N_24369,N_24201);
and UO_2926 (O_2926,N_24583,N_24367);
and UO_2927 (O_2927,N_24461,N_24059);
or UO_2928 (O_2928,N_23812,N_24852);
xnor UO_2929 (O_2929,N_24851,N_24827);
or UO_2930 (O_2930,N_24675,N_24157);
and UO_2931 (O_2931,N_23930,N_23880);
nor UO_2932 (O_2932,N_24290,N_24669);
nor UO_2933 (O_2933,N_24125,N_24809);
or UO_2934 (O_2934,N_24424,N_24530);
nand UO_2935 (O_2935,N_23819,N_23804);
and UO_2936 (O_2936,N_23755,N_24615);
and UO_2937 (O_2937,N_24309,N_24587);
xor UO_2938 (O_2938,N_24284,N_24287);
nand UO_2939 (O_2939,N_24451,N_24763);
xor UO_2940 (O_2940,N_24267,N_24579);
and UO_2941 (O_2941,N_24439,N_24288);
and UO_2942 (O_2942,N_24619,N_23787);
and UO_2943 (O_2943,N_23947,N_24067);
or UO_2944 (O_2944,N_24485,N_23954);
and UO_2945 (O_2945,N_23804,N_23792);
xor UO_2946 (O_2946,N_24043,N_24771);
nand UO_2947 (O_2947,N_24312,N_24095);
and UO_2948 (O_2948,N_24979,N_23781);
and UO_2949 (O_2949,N_23946,N_24982);
xnor UO_2950 (O_2950,N_24195,N_24248);
and UO_2951 (O_2951,N_24494,N_24530);
xor UO_2952 (O_2952,N_24519,N_24863);
nor UO_2953 (O_2953,N_24096,N_24873);
nor UO_2954 (O_2954,N_24383,N_23973);
nand UO_2955 (O_2955,N_24586,N_23781);
or UO_2956 (O_2956,N_24272,N_24093);
or UO_2957 (O_2957,N_24815,N_24305);
nor UO_2958 (O_2958,N_24613,N_23908);
nor UO_2959 (O_2959,N_24589,N_24121);
nor UO_2960 (O_2960,N_23972,N_23989);
nor UO_2961 (O_2961,N_24118,N_24106);
nand UO_2962 (O_2962,N_23806,N_24153);
nand UO_2963 (O_2963,N_24793,N_24671);
nor UO_2964 (O_2964,N_24158,N_24805);
or UO_2965 (O_2965,N_24487,N_24631);
and UO_2966 (O_2966,N_24919,N_24250);
xor UO_2967 (O_2967,N_23917,N_24866);
xor UO_2968 (O_2968,N_24569,N_24219);
or UO_2969 (O_2969,N_24899,N_24773);
xor UO_2970 (O_2970,N_23838,N_23855);
or UO_2971 (O_2971,N_23826,N_24832);
nor UO_2972 (O_2972,N_24037,N_23971);
and UO_2973 (O_2973,N_23876,N_24204);
xor UO_2974 (O_2974,N_23960,N_24991);
nand UO_2975 (O_2975,N_23760,N_24165);
nor UO_2976 (O_2976,N_24588,N_24881);
or UO_2977 (O_2977,N_23788,N_24139);
or UO_2978 (O_2978,N_23802,N_24424);
or UO_2979 (O_2979,N_23839,N_24646);
nand UO_2980 (O_2980,N_24660,N_24515);
and UO_2981 (O_2981,N_24566,N_24357);
nand UO_2982 (O_2982,N_24169,N_24024);
and UO_2983 (O_2983,N_24581,N_24409);
nor UO_2984 (O_2984,N_24277,N_24851);
nand UO_2985 (O_2985,N_24456,N_24151);
nand UO_2986 (O_2986,N_24140,N_24635);
nor UO_2987 (O_2987,N_24142,N_24310);
or UO_2988 (O_2988,N_24557,N_24258);
and UO_2989 (O_2989,N_24402,N_24244);
xor UO_2990 (O_2990,N_24111,N_24879);
nand UO_2991 (O_2991,N_24219,N_24387);
xor UO_2992 (O_2992,N_23895,N_24269);
nand UO_2993 (O_2993,N_24965,N_24239);
xnor UO_2994 (O_2994,N_24409,N_24578);
nand UO_2995 (O_2995,N_23809,N_24619);
and UO_2996 (O_2996,N_24152,N_23874);
or UO_2997 (O_2997,N_23834,N_24406);
and UO_2998 (O_2998,N_24197,N_23883);
or UO_2999 (O_2999,N_24348,N_24951);
endmodule