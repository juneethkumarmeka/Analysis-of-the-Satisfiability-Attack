module basic_2000_20000_2500_5_levels_5xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
xor U0 (N_0,In_278,In_1957);
or U1 (N_1,In_929,In_96);
or U2 (N_2,In_1781,In_995);
or U3 (N_3,In_1908,In_639);
or U4 (N_4,In_773,In_1652);
nor U5 (N_5,In_1940,In_1367);
nor U6 (N_6,In_1846,In_1920);
nor U7 (N_7,In_1290,In_1450);
and U8 (N_8,In_990,In_1611);
nor U9 (N_9,In_835,In_1637);
nand U10 (N_10,In_312,In_1058);
nor U11 (N_11,In_1913,In_1771);
nor U12 (N_12,In_1980,In_1901);
and U13 (N_13,In_1778,In_13);
nand U14 (N_14,In_1448,In_1514);
xnor U15 (N_15,In_1363,In_1090);
or U16 (N_16,In_1995,In_1910);
nand U17 (N_17,In_980,In_94);
nor U18 (N_18,In_214,In_146);
nor U19 (N_19,In_1257,In_451);
xnor U20 (N_20,In_1074,In_1244);
nand U21 (N_21,In_612,In_91);
nand U22 (N_22,In_514,In_252);
or U23 (N_23,In_24,In_1342);
nor U24 (N_24,In_966,In_1261);
nand U25 (N_25,In_1805,In_262);
nand U26 (N_26,In_1966,In_836);
or U27 (N_27,In_1681,In_295);
nor U28 (N_28,In_1807,In_1304);
nand U29 (N_29,In_463,In_1275);
nand U30 (N_30,In_618,In_634);
nor U31 (N_31,In_1630,In_501);
nand U32 (N_32,In_1680,In_826);
nor U33 (N_33,In_1856,In_363);
or U34 (N_34,In_1106,In_1126);
nor U35 (N_35,In_83,In_1173);
or U36 (N_36,In_884,In_1129);
nand U37 (N_37,In_1286,In_1458);
or U38 (N_38,In_39,In_103);
and U39 (N_39,In_1171,In_253);
nand U40 (N_40,In_1205,In_1946);
nor U41 (N_41,In_204,In_1839);
or U42 (N_42,In_1315,In_753);
nand U43 (N_43,In_415,In_168);
nor U44 (N_44,In_525,In_965);
nor U45 (N_45,In_563,In_1958);
nor U46 (N_46,In_1260,In_185);
nor U47 (N_47,In_814,In_731);
nor U48 (N_48,In_600,In_849);
and U49 (N_49,In_900,In_382);
xor U50 (N_50,In_971,In_1387);
xnor U51 (N_51,In_1557,In_1595);
nor U52 (N_52,In_1788,In_1499);
or U53 (N_53,In_1293,In_306);
or U54 (N_54,In_1258,In_1016);
or U55 (N_55,In_1024,In_1810);
and U56 (N_56,In_258,In_1408);
or U57 (N_57,In_187,In_810);
xnor U58 (N_58,In_341,In_877);
or U59 (N_59,In_65,In_1424);
nand U60 (N_60,In_346,In_249);
and U61 (N_61,In_165,In_603);
xnor U62 (N_62,In_1789,In_1020);
and U63 (N_63,In_1123,In_704);
nand U64 (N_64,In_1761,In_1785);
nor U65 (N_65,In_1110,In_1197);
nor U66 (N_66,In_637,In_284);
or U67 (N_67,In_645,In_1142);
nor U68 (N_68,In_1382,In_661);
xor U69 (N_69,In_1010,In_1442);
xnor U70 (N_70,In_869,In_366);
and U71 (N_71,In_699,In_1501);
nor U72 (N_72,In_1289,In_1555);
or U73 (N_73,In_678,In_1721);
nor U74 (N_74,In_1421,In_120);
nor U75 (N_75,In_1180,In_905);
or U76 (N_76,In_915,In_838);
xnor U77 (N_77,In_851,In_759);
nand U78 (N_78,In_410,In_938);
nor U79 (N_79,In_908,In_1337);
nand U80 (N_80,In_1797,In_1462);
xor U81 (N_81,In_1490,In_1075);
nand U82 (N_82,In_1202,In_62);
nor U83 (N_83,In_744,In_576);
and U84 (N_84,In_1496,In_1842);
and U85 (N_85,In_935,In_1230);
or U86 (N_86,In_356,In_767);
xor U87 (N_87,In_1553,In_104);
or U88 (N_88,In_556,In_1774);
nor U89 (N_89,In_1863,In_504);
and U90 (N_90,In_528,In_872);
nand U91 (N_91,In_1684,In_1606);
and U92 (N_92,In_1441,In_1597);
nand U93 (N_93,In_1883,In_850);
and U94 (N_94,In_1725,In_855);
nand U95 (N_95,In_1269,In_1067);
or U96 (N_96,In_1044,In_1766);
xnor U97 (N_97,In_397,In_11);
nand U98 (N_98,In_1219,In_1822);
nor U99 (N_99,In_301,In_469);
xnor U100 (N_100,In_739,In_414);
nor U101 (N_101,In_1537,In_74);
xor U102 (N_102,In_1800,In_196);
nor U103 (N_103,In_257,In_396);
or U104 (N_104,In_1339,In_1377);
or U105 (N_105,In_1517,In_994);
nand U106 (N_106,In_530,In_348);
or U107 (N_107,In_721,In_125);
nand U108 (N_108,In_619,In_1633);
nor U109 (N_109,In_314,In_539);
nor U110 (N_110,In_565,In_1610);
nor U111 (N_111,In_687,In_1368);
or U112 (N_112,In_1519,In_1479);
nand U113 (N_113,In_1878,In_1598);
nand U114 (N_114,In_1876,In_212);
or U115 (N_115,In_495,In_732);
or U116 (N_116,In_1984,In_49);
or U117 (N_117,In_1264,In_734);
nand U118 (N_118,In_1237,In_1941);
nor U119 (N_119,In_1943,In_1407);
nand U120 (N_120,In_351,In_1592);
nor U121 (N_121,In_1146,In_1283);
nand U122 (N_122,In_1979,In_119);
or U123 (N_123,In_142,In_1100);
and U124 (N_124,In_1647,In_1151);
nand U125 (N_125,In_1987,In_1163);
and U126 (N_126,In_1743,In_456);
nor U127 (N_127,In_1410,In_616);
nand U128 (N_128,In_447,In_570);
xnor U129 (N_129,In_1591,In_726);
and U130 (N_130,In_1133,In_1613);
and U131 (N_131,In_335,In_195);
and U132 (N_132,In_520,In_1470);
nor U133 (N_133,In_960,In_73);
nor U134 (N_134,In_1256,In_503);
xnor U135 (N_135,In_1340,In_1777);
xnor U136 (N_136,In_395,In_1086);
and U137 (N_137,In_1709,In_1073);
nor U138 (N_138,In_169,In_985);
or U139 (N_139,In_419,In_1992);
nand U140 (N_140,In_886,In_729);
nor U141 (N_141,In_1472,In_1926);
xor U142 (N_142,In_1053,In_1302);
or U143 (N_143,In_483,In_1981);
nand U144 (N_144,In_1798,In_344);
nor U145 (N_145,In_1738,In_280);
nor U146 (N_146,In_1046,In_1423);
and U147 (N_147,In_776,In_518);
xor U148 (N_148,In_519,In_1989);
xnor U149 (N_149,In_1525,In_631);
or U150 (N_150,In_756,In_1025);
xor U151 (N_151,In_1212,In_774);
nand U152 (N_152,In_244,In_1198);
and U153 (N_153,In_595,In_626);
and U154 (N_154,In_1120,In_19);
or U155 (N_155,In_1536,In_67);
xnor U156 (N_156,In_1348,In_1203);
and U157 (N_157,In_260,In_71);
nor U158 (N_158,In_1760,In_100);
or U159 (N_159,In_1150,In_1651);
nor U160 (N_160,In_928,In_1397);
nand U161 (N_161,In_462,In_878);
nor U162 (N_162,In_1216,In_1844);
nor U163 (N_163,In_1001,In_1460);
nor U164 (N_164,In_1182,In_571);
nand U165 (N_165,In_989,In_76);
or U166 (N_166,In_975,In_1013);
nand U167 (N_167,In_77,In_955);
and U168 (N_168,In_684,In_35);
or U169 (N_169,In_1770,In_1579);
and U170 (N_170,In_353,In_880);
or U171 (N_171,In_1706,In_1454);
nor U172 (N_172,In_1308,In_1051);
or U173 (N_173,In_802,In_246);
and U174 (N_174,In_1921,In_1109);
and U175 (N_175,In_1838,In_1035);
or U176 (N_176,In_1322,In_1378);
nor U177 (N_177,In_1279,In_203);
and U178 (N_178,In_858,In_476);
and U179 (N_179,In_890,In_370);
nand U180 (N_180,In_621,In_513);
nor U181 (N_181,In_1440,In_175);
nand U182 (N_182,In_1922,In_1451);
and U183 (N_183,In_1612,In_1791);
nand U184 (N_184,In_422,In_765);
nor U185 (N_185,In_1799,In_467);
or U186 (N_186,In_671,In_1009);
nand U187 (N_187,In_713,In_733);
xor U188 (N_188,In_566,In_310);
nor U189 (N_189,In_1699,In_1115);
nor U190 (N_190,In_380,In_1281);
xnor U191 (N_191,In_837,In_32);
and U192 (N_192,In_1779,In_1712);
nand U193 (N_193,In_1998,In_882);
nor U194 (N_194,In_1635,In_1070);
nand U195 (N_195,In_807,In_242);
or U196 (N_196,In_763,In_1179);
or U197 (N_197,In_1003,In_443);
nor U198 (N_198,In_285,In_227);
nor U199 (N_199,In_116,In_1232);
and U200 (N_200,In_25,In_1986);
nor U201 (N_201,In_199,In_108);
or U202 (N_202,In_1643,In_264);
and U203 (N_203,In_486,In_1088);
or U204 (N_204,In_736,In_1307);
and U205 (N_205,In_793,In_286);
nand U206 (N_206,In_1875,In_1621);
nor U207 (N_207,In_1185,In_326);
xnor U208 (N_208,In_892,In_682);
or U209 (N_209,In_1616,In_1891);
or U210 (N_210,In_1136,In_1911);
and U211 (N_211,In_232,In_1380);
nor U212 (N_212,In_479,In_1412);
xor U213 (N_213,In_1676,In_1114);
or U214 (N_214,In_215,In_403);
nand U215 (N_215,In_1650,In_1149);
nor U216 (N_216,In_670,In_1990);
nand U217 (N_217,In_381,In_14);
or U218 (N_218,In_1028,In_615);
xor U219 (N_219,In_1014,In_584);
and U220 (N_220,In_1802,In_95);
nor U221 (N_221,In_220,In_330);
nor U222 (N_222,In_1793,In_413);
nor U223 (N_223,In_572,In_794);
nand U224 (N_224,In_948,In_963);
nor U225 (N_225,In_1622,In_847);
nor U226 (N_226,In_1601,In_29);
nand U227 (N_227,In_1632,In_1480);
nor U228 (N_228,In_269,In_1329);
and U229 (N_229,In_811,In_446);
nand U230 (N_230,In_31,In_1434);
or U231 (N_231,In_48,In_1860);
nor U232 (N_232,In_1964,In_460);
or U233 (N_233,In_970,In_685);
nand U234 (N_234,In_548,In_1713);
nor U235 (N_235,In_597,In_1696);
and U236 (N_236,In_1933,In_1562);
nand U237 (N_237,In_1700,In_740);
and U238 (N_238,In_1145,In_1975);
xnor U239 (N_239,In_433,In_797);
nand U240 (N_240,In_452,In_93);
nor U241 (N_241,In_1411,In_1573);
and U242 (N_242,In_1841,In_686);
nor U243 (N_243,In_1165,In_1148);
and U244 (N_244,In_749,In_465);
nor U245 (N_245,In_464,In_585);
nor U246 (N_246,In_511,In_693);
nor U247 (N_247,In_1231,In_1850);
nand U248 (N_248,In_1226,In_1135);
or U249 (N_249,In_221,In_206);
nor U250 (N_250,In_1041,In_1094);
nor U251 (N_251,In_606,In_854);
or U252 (N_252,In_1960,In_752);
and U253 (N_253,In_255,In_668);
nand U254 (N_254,In_1330,In_1017);
nor U255 (N_255,In_912,In_1005);
nor U256 (N_256,In_20,In_1871);
nand U257 (N_257,In_1473,In_47);
nor U258 (N_258,In_1081,In_61);
nor U259 (N_259,In_226,In_1213);
and U260 (N_260,In_643,In_1343);
nand U261 (N_261,In_428,In_1732);
nor U262 (N_262,In_1143,In_833);
and U263 (N_263,In_1574,In_1736);
or U264 (N_264,In_1147,In_1688);
or U265 (N_265,In_1787,In_16);
nand U266 (N_266,In_1042,In_1900);
and U267 (N_267,In_277,In_1641);
nor U268 (N_268,In_1756,In_54);
nor U269 (N_269,In_1168,In_343);
nand U270 (N_270,In_978,In_412);
xnor U271 (N_271,In_1930,In_1973);
and U272 (N_272,In_1566,In_780);
xor U273 (N_273,In_979,In_784);
nor U274 (N_274,In_1455,In_1288);
nand U275 (N_275,In_667,In_426);
and U276 (N_276,In_496,In_1038);
or U277 (N_277,In_12,In_712);
nor U278 (N_278,In_924,In_1855);
or U279 (N_279,In_1371,In_735);
or U280 (N_280,In_1693,In_1008);
nor U281 (N_281,In_649,In_825);
nor U282 (N_282,In_805,In_1045);
and U283 (N_283,In_416,In_288);
and U284 (N_284,In_1814,In_473);
or U285 (N_285,In_1547,In_1703);
nand U286 (N_286,In_491,In_321);
and U287 (N_287,In_136,In_1445);
or U288 (N_288,In_582,In_1324);
nand U289 (N_289,In_1331,In_1730);
or U290 (N_290,In_201,In_1518);
and U291 (N_291,In_1731,In_1456);
xnor U292 (N_292,In_1996,In_228);
or U293 (N_293,In_654,In_522);
or U294 (N_294,In_891,In_41);
nor U295 (N_295,In_1019,In_1162);
and U296 (N_296,In_715,In_1865);
xnor U297 (N_297,In_225,In_1358);
or U298 (N_298,In_1813,In_1832);
nor U299 (N_299,In_1429,In_859);
and U300 (N_300,In_640,In_623);
or U301 (N_301,In_409,In_1649);
nand U302 (N_302,In_1488,In_427);
and U303 (N_303,In_782,In_498);
nand U304 (N_304,In_302,In_230);
nor U305 (N_305,In_786,In_1744);
nand U306 (N_306,In_111,In_137);
and U307 (N_307,In_282,In_1769);
nor U308 (N_308,In_834,In_475);
nand U309 (N_309,In_184,In_1483);
nor U310 (N_310,In_1121,In_390);
and U311 (N_311,In_1816,In_1541);
xor U312 (N_312,In_59,In_231);
and U313 (N_313,In_1386,In_540);
xor U314 (N_314,In_663,In_1064);
and U315 (N_315,In_1117,In_904);
nor U316 (N_316,In_1193,In_1963);
nor U317 (N_317,In_1240,In_1453);
nor U318 (N_318,In_992,In_1665);
or U319 (N_319,In_207,In_916);
nand U320 (N_320,In_482,In_1510);
or U321 (N_321,In_543,In_1134);
or U322 (N_322,In_1549,In_1072);
nor U323 (N_323,In_1837,In_303);
xor U324 (N_324,In_78,In_702);
or U325 (N_325,In_499,In_1494);
xor U326 (N_326,In_1753,In_155);
and U327 (N_327,In_489,In_128);
and U328 (N_328,In_1266,In_1972);
and U329 (N_329,In_160,In_150);
nor U330 (N_330,In_1222,In_399);
nand U331 (N_331,In_1656,In_842);
nor U332 (N_332,In_1638,In_764);
nand U333 (N_333,In_81,In_339);
or U334 (N_334,In_1927,In_1678);
and U335 (N_335,In_1988,In_1464);
xnor U336 (N_336,In_789,In_1722);
xor U337 (N_337,In_554,In_1784);
and U338 (N_338,In_1707,In_1742);
nand U339 (N_339,In_754,In_320);
and U340 (N_340,In_1554,In_445);
and U341 (N_341,In_1446,In_1991);
or U342 (N_342,In_1945,In_1199);
nand U343 (N_343,In_1748,In_1277);
and U344 (N_344,In_383,In_352);
xor U345 (N_345,In_1204,In_1102);
nand U346 (N_346,In_586,In_770);
nor U347 (N_347,In_1211,In_1740);
or U348 (N_348,In_1535,In_964);
nand U349 (N_349,In_1141,In_1297);
and U350 (N_350,In_1345,In_129);
and U351 (N_351,In_673,In_779);
nand U352 (N_352,In_1629,In_1273);
nand U353 (N_353,In_1040,In_1310);
or U354 (N_354,In_1449,In_1127);
nand U355 (N_355,In_1505,In_92);
or U356 (N_356,In_843,In_1426);
and U357 (N_357,In_1419,In_1884);
nand U358 (N_358,In_82,In_102);
nor U359 (N_359,In_646,In_294);
nor U360 (N_360,In_127,In_3);
or U361 (N_361,In_152,In_23);
nand U362 (N_362,In_839,In_1138);
nand U363 (N_363,In_1854,In_149);
and U364 (N_364,In_40,In_1570);
or U365 (N_365,In_1057,In_1191);
nor U366 (N_366,In_977,In_632);
xor U367 (N_367,In_1604,In_987);
nand U368 (N_368,In_930,In_642);
nand U369 (N_369,In_517,In_931);
or U370 (N_370,In_1754,In_299);
and U371 (N_371,In_1619,In_524);
or U372 (N_372,In_1082,In_506);
nand U373 (N_373,In_17,In_154);
nor U374 (N_374,In_722,In_939);
or U375 (N_375,In_112,In_1096);
nand U376 (N_376,In_655,In_1022);
nand U377 (N_377,In_647,In_1895);
or U378 (N_378,In_967,In_243);
and U379 (N_379,In_828,In_188);
or U380 (N_380,In_601,In_1765);
xor U381 (N_381,In_1885,In_98);
xnor U382 (N_382,In_998,In_653);
or U383 (N_383,In_1758,In_1111);
xnor U384 (N_384,In_625,In_1834);
or U385 (N_385,In_1790,In_202);
nand U386 (N_386,In_1430,In_1463);
nor U387 (N_387,In_400,In_1607);
or U388 (N_388,In_665,In_1326);
nor U389 (N_389,In_881,In_99);
and U390 (N_390,In_1873,In_1824);
xnor U391 (N_391,In_472,In_800);
nor U392 (N_392,In_1720,In_575);
nand U393 (N_393,In_455,In_1605);
nand U394 (N_394,In_461,In_1679);
or U395 (N_395,In_1625,In_853);
and U396 (N_396,In_438,In_1899);
nor U397 (N_397,In_307,In_323);
nor U398 (N_398,In_1773,In_1724);
nand U399 (N_399,In_1154,In_769);
nor U400 (N_400,In_388,In_547);
and U401 (N_401,In_1015,In_1903);
nor U402 (N_402,In_1296,In_692);
nand U403 (N_403,In_115,In_1803);
nor U404 (N_404,In_1228,In_509);
and U405 (N_405,In_1229,In_318);
and U406 (N_406,In_1285,In_1209);
nor U407 (N_407,In_1545,In_1527);
and U408 (N_408,In_435,In_313);
xnor U409 (N_409,In_1033,In_1508);
nand U410 (N_410,In_26,In_594);
and U411 (N_411,In_1623,In_1085);
and U412 (N_412,In_1772,In_1819);
and U413 (N_413,In_1939,In_182);
and U414 (N_414,In_1417,In_123);
or U415 (N_415,In_1925,In_1007);
and U416 (N_416,In_669,In_1299);
nand U417 (N_417,In_1055,In_1533);
nand U418 (N_418,In_785,In_660);
xnor U419 (N_419,In_1919,In_1585);
and U420 (N_420,In_981,In_1669);
or U421 (N_421,In_425,In_43);
nand U422 (N_422,In_1952,In_1011);
or U423 (N_423,In_1775,In_1671);
nor U424 (N_424,In_378,In_1474);
nor U425 (N_425,In_896,In_126);
or U426 (N_426,In_85,In_535);
nand U427 (N_427,In_1481,In_695);
nand U428 (N_428,In_561,In_1192);
xnor U429 (N_429,In_1504,In_932);
and U430 (N_430,In_829,In_1924);
and U431 (N_431,In_508,In_1786);
and U432 (N_432,In_902,In_1872);
nand U433 (N_433,In_868,In_1534);
nand U434 (N_434,In_440,In_1947);
nor U435 (N_435,In_490,In_1325);
and U436 (N_436,In_106,In_1608);
nor U437 (N_437,In_1404,In_1780);
nor U438 (N_438,In_1714,In_1);
xnor U439 (N_439,In_1936,In_743);
or U440 (N_440,In_1124,In_1529);
and U441 (N_441,In_976,In_680);
and U442 (N_442,In_1402,In_1139);
nand U443 (N_443,In_1729,In_1880);
and U444 (N_444,In_1660,In_1130);
or U445 (N_445,In_635,In_861);
nand U446 (N_446,In_1233,In_1356);
or U447 (N_447,In_1418,In_459);
or U448 (N_448,In_1664,In_1831);
or U449 (N_449,In_1866,In_1828);
xnor U450 (N_450,In_1931,In_1956);
and U451 (N_451,In_276,In_153);
xnor U452 (N_452,In_292,In_384);
and U453 (N_453,In_862,In_122);
nor U454 (N_454,In_1065,In_1398);
nand U455 (N_455,In_274,In_101);
nand U456 (N_456,In_1376,In_1870);
xor U457 (N_457,In_863,In_747);
nor U458 (N_458,In_1178,In_1321);
nor U459 (N_459,In_534,In_1467);
or U460 (N_460,In_1653,In_454);
nor U461 (N_461,In_1357,In_1689);
nand U462 (N_462,In_1112,In_962);
and U463 (N_463,In_1385,In_953);
nor U464 (N_464,In_1166,In_349);
nor U465 (N_465,In_537,In_57);
or U466 (N_466,In_250,In_1580);
and U467 (N_467,In_1654,In_404);
xor U468 (N_468,In_969,In_694);
xor U469 (N_469,In_6,In_1413);
or U470 (N_470,In_1561,In_373);
nor U471 (N_471,In_1727,In_1750);
or U472 (N_472,In_652,In_430);
nor U473 (N_473,In_1857,In_174);
and U474 (N_474,In_516,In_1836);
nor U475 (N_475,In_417,In_166);
nor U476 (N_476,In_442,In_1347);
and U477 (N_477,In_958,In_1091);
and U478 (N_478,In_988,In_1432);
or U479 (N_479,In_267,In_1311);
and U480 (N_480,In_1144,In_1639);
and U481 (N_481,In_439,In_263);
or U482 (N_482,In_710,In_361);
or U483 (N_483,In_1835,In_617);
and U484 (N_484,In_1023,In_1677);
nand U485 (N_485,In_1801,In_558);
xnor U486 (N_486,In_672,In_1217);
or U487 (N_487,In_1615,In_1224);
or U488 (N_488,In_1351,In_745);
nand U489 (N_489,In_7,In_1888);
and U490 (N_490,In_15,In_1221);
xor U491 (N_491,In_1245,In_1189);
nand U492 (N_492,In_148,In_1004);
and U493 (N_493,In_1466,In_1176);
xnor U494 (N_494,In_218,In_1190);
and U495 (N_495,In_138,In_1476);
nor U496 (N_496,In_1069,In_18);
nor U497 (N_497,In_1047,In_79);
and U498 (N_498,In_972,In_1572);
and U499 (N_499,In_1512,In_1563);
or U500 (N_500,In_792,In_1118);
or U501 (N_501,In_758,In_1080);
nor U502 (N_502,In_944,In_577);
and U503 (N_503,In_474,In_118);
and U504 (N_504,In_1896,In_229);
or U505 (N_505,In_1032,In_1548);
or U506 (N_506,In_1993,In_1886);
nor U507 (N_507,In_529,In_502);
nor U508 (N_508,In_291,In_1728);
or U509 (N_509,In_234,In_1251);
nor U510 (N_510,In_1098,In_650);
or U511 (N_511,In_338,In_1379);
and U512 (N_512,In_936,In_481);
or U513 (N_513,In_1294,In_484);
nor U514 (N_514,In_762,In_1636);
and U515 (N_515,In_358,In_1847);
and U516 (N_516,In_131,In_1783);
or U517 (N_517,In_559,In_984);
xor U518 (N_518,In_588,In_555);
nand U519 (N_519,In_893,In_911);
and U520 (N_520,In_1917,In_816);
nand U521 (N_521,In_385,In_701);
or U522 (N_522,In_870,In_1581);
or U523 (N_523,In_1867,In_304);
nor U524 (N_524,In_1752,In_1609);
nor U525 (N_525,In_107,In_1312);
nand U526 (N_526,In_1543,In_1320);
nand U527 (N_527,In_290,In_1252);
nor U528 (N_528,In_162,In_799);
nor U529 (N_529,In_1640,In_1994);
and U530 (N_530,In_1531,In_485);
or U531 (N_531,In_1845,In_720);
and U532 (N_532,In_121,In_848);
and U533 (N_533,In_1172,In_748);
and U534 (N_534,In_982,In_172);
nand U535 (N_535,In_133,In_1515);
or U536 (N_536,In_1270,In_856);
and U537 (N_537,In_923,In_1043);
or U538 (N_538,In_730,In_1600);
nor U539 (N_539,In_1596,In_1352);
or U540 (N_540,In_1624,In_1161);
and U541 (N_541,In_1459,In_1465);
or U542 (N_542,In_1879,In_697);
or U543 (N_543,In_1428,In_401);
and U544 (N_544,In_1565,In_1056);
or U545 (N_545,In_1420,In_1815);
nor U546 (N_546,In_170,In_1242);
nand U547 (N_547,In_1049,In_251);
xnor U548 (N_548,In_599,In_1532);
or U549 (N_549,In_375,In_376);
nand U550 (N_550,In_493,In_1132);
nand U551 (N_551,In_105,In_1436);
or U552 (N_552,In_841,In_1373);
nand U553 (N_553,In_1661,In_1659);
nor U554 (N_554,In_1327,In_1087);
nand U555 (N_555,In_360,In_830);
or U556 (N_556,In_75,In_1267);
nand U557 (N_557,In_327,In_377);
nor U558 (N_558,In_141,In_832);
nand U559 (N_559,In_674,In_1391);
or U560 (N_560,In_432,In_500);
or U561 (N_561,In_322,In_1904);
and U562 (N_562,In_1923,In_365);
nand U563 (N_563,In_1280,In_198);
and U564 (N_564,In_134,In_1223);
nor U565 (N_565,In_630,In_1158);
xor U566 (N_566,In_217,In_1962);
or U567 (N_567,In_901,In_1687);
nor U568 (N_568,In_1951,In_1715);
and U569 (N_569,In_186,In_1444);
or U570 (N_570,In_706,In_1355);
and U571 (N_571,In_1062,In_159);
nand U572 (N_572,In_783,In_300);
nand U573 (N_573,In_708,In_614);
and U574 (N_574,In_1313,In_275);
nand U575 (N_575,In_1012,In_110);
and U576 (N_576,In_1762,In_1131);
nand U577 (N_577,In_27,In_477);
nor U578 (N_578,In_1157,In_1137);
or U579 (N_579,In_1344,In_1971);
xor U580 (N_580,In_1594,In_1006);
nand U581 (N_581,In_354,In_544);
nand U582 (N_582,In_1809,In_1965);
and U583 (N_583,In_1383,In_1739);
and U584 (N_584,In_596,In_240);
or U585 (N_585,In_191,In_578);
xor U586 (N_586,In_999,In_696);
and U587 (N_587,In_1116,In_1516);
and U588 (N_588,In_505,In_342);
or U589 (N_589,In_568,In_1364);
nand U590 (N_590,In_1843,In_1177);
nor U591 (N_591,In_194,In_1907);
nor U592 (N_592,In_1447,In_1201);
and U593 (N_593,In_768,In_1830);
or U594 (N_594,In_874,In_407);
and U595 (N_595,In_1603,In_183);
and U596 (N_596,In_845,In_564);
nor U597 (N_597,In_1215,In_406);
and U598 (N_598,In_991,In_236);
nor U599 (N_599,In_587,In_1194);
nand U600 (N_600,In_553,In_937);
or U601 (N_601,In_1912,In_46);
nand U602 (N_602,In_1396,In_1833);
nand U603 (N_603,In_959,In_1817);
or U604 (N_604,In_1571,In_641);
or U605 (N_605,In_1452,In_1167);
or U606 (N_606,In_1425,In_355);
nand U607 (N_607,In_1169,In_1427);
or U608 (N_608,In_145,In_798);
or U609 (N_609,In_223,In_512);
or U610 (N_610,In_927,In_1818);
or U611 (N_611,In_398,In_200);
or U612 (N_612,In_1759,In_1066);
or U613 (N_613,In_638,In_63);
nand U614 (N_614,In_405,In_1848);
and U615 (N_615,In_55,In_1674);
nand U616 (N_616,In_362,In_973);
nor U617 (N_617,In_1349,In_56);
xor U618 (N_618,In_457,In_823);
nor U619 (N_619,In_213,In_997);
and U620 (N_620,In_4,In_1593);
nor U621 (N_621,In_1587,In_1977);
or U622 (N_622,In_1372,In_724);
and U623 (N_623,In_261,In_1254);
nor U624 (N_624,In_1303,In_742);
nor U625 (N_625,In_161,In_1546);
nor U626 (N_626,In_171,In_1849);
and U627 (N_627,In_44,In_347);
nand U628 (N_628,In_808,In_1627);
and U629 (N_629,In_393,In_1335);
nor U630 (N_630,In_507,In_1097);
nand U631 (N_631,In_737,In_1523);
and U632 (N_632,In_1967,In_167);
nand U633 (N_633,In_1734,In_1292);
and U634 (N_634,In_1916,In_628);
xor U635 (N_635,In_1862,In_30);
nor U636 (N_636,In_1122,In_1726);
or U637 (N_637,In_1160,In_703);
and U638 (N_638,In_1914,In_1018);
xnor U639 (N_639,In_714,In_345);
nor U640 (N_640,In_775,In_1050);
nor U641 (N_641,In_163,In_1333);
nand U642 (N_642,In_297,In_1489);
or U643 (N_643,In_247,In_392);
or U644 (N_644,In_894,In_315);
nor U645 (N_645,In_899,In_1184);
xor U646 (N_646,In_256,In_1265);
nand U647 (N_647,In_1893,In_1298);
or U648 (N_648,In_36,In_1568);
and U649 (N_649,In_389,In_827);
nor U650 (N_650,In_1366,In_1059);
nor U651 (N_651,In_598,In_1234);
and U652 (N_652,In_718,In_755);
nor U653 (N_653,In_1882,In_238);
nor U654 (N_654,In_950,In_679);
or U655 (N_655,In_1414,In_316);
or U656 (N_656,In_89,In_1897);
or U657 (N_657,In_1235,In_666);
nand U658 (N_658,In_1618,In_177);
nor U659 (N_659,In_391,In_1982);
or U660 (N_660,In_1953,In_1078);
and U661 (N_661,In_907,In_777);
nand U662 (N_662,In_1682,In_1238);
and U663 (N_663,In_560,In_205);
or U664 (N_664,In_1438,In_1084);
or U665 (N_665,In_1881,In_817);
nand U666 (N_666,In_919,In_1586);
nor U667 (N_667,In_132,In_898);
and U668 (N_668,In_593,In_1582);
nand U669 (N_669,In_1186,In_181);
nand U670 (N_670,In_1858,In_846);
nor U671 (N_671,In_1485,In_478);
nor U672 (N_672,In_1301,In_1443);
nand U673 (N_673,In_1175,In_1188);
nor U674 (N_674,In_324,In_648);
nand U675 (N_675,In_1511,In_219);
or U676 (N_676,In_308,In_538);
or U677 (N_677,In_325,In_925);
and U678 (N_678,In_1999,In_532);
nor U679 (N_679,In_1210,In_1673);
nand U680 (N_680,In_144,In_681);
nor U681 (N_681,In_470,In_1314);
xor U682 (N_682,In_1478,In_60);
nor U683 (N_683,In_51,In_949);
or U684 (N_684,In_604,In_716);
or U685 (N_685,In_1026,In_45);
nand U686 (N_686,In_1300,In_368);
nand U687 (N_687,In_1670,In_515);
nor U688 (N_688,In_728,In_1864);
and U689 (N_689,In_1218,In_1524);
or U690 (N_690,In_1718,In_741);
or U691 (N_691,In_411,In_844);
or U692 (N_692,In_38,In_66);
nor U693 (N_693,In_974,In_1334);
nand U694 (N_694,In_279,In_510);
nand U695 (N_695,In_1929,In_266);
nor U696 (N_696,In_951,In_254);
and U697 (N_697,In_609,In_781);
xnor U698 (N_698,In_273,In_1544);
nor U699 (N_699,In_1093,In_436);
or U700 (N_700,In_1976,In_956);
and U701 (N_701,In_1400,In_918);
and U702 (N_702,In_466,In_331);
nand U703 (N_703,In_1105,In_209);
and U704 (N_704,In_1710,In_1542);
and U705 (N_705,In_757,In_497);
or U706 (N_706,In_1390,In_917);
nor U707 (N_707,In_494,In_1031);
nand U708 (N_708,In_1645,In_934);
nand U709 (N_709,In_709,In_1374);
nand U710 (N_710,In_1658,In_1503);
xnor U711 (N_711,In_333,In_942);
and U712 (N_712,In_487,In_1083);
and U713 (N_713,In_1353,In_1642);
nand U714 (N_714,In_156,In_1584);
or U715 (N_715,In_803,In_1751);
nor U716 (N_716,In_579,In_1657);
and U717 (N_717,In_527,In_1905);
nor U718 (N_718,In_272,In_790);
xor U719 (N_719,In_374,In_526);
and U720 (N_720,In_1317,In_189);
nor U721 (N_721,In_1997,In_1246);
and U722 (N_722,In_449,In_1493);
or U723 (N_723,In_1068,In_983);
and U724 (N_724,In_42,In_1890);
and U725 (N_725,In_444,In_1021);
nor U726 (N_726,In_1422,In_173);
nor U727 (N_727,In_1909,In_1968);
xor U728 (N_728,In_1119,In_492);
nor U729 (N_729,In_109,In_1220);
nand U730 (N_730,In_488,In_1389);
or U731 (N_731,In_1705,In_804);
nand U732 (N_732,In_1249,In_387);
nor U733 (N_733,In_1092,In_705);
and U734 (N_734,In_158,In_831);
xnor U735 (N_735,In_541,In_1037);
nor U736 (N_736,In_1107,In_1564);
nor U737 (N_737,In_656,In_866);
and U738 (N_738,In_1634,In_921);
nor U739 (N_739,In_450,In_480);
and U740 (N_740,In_943,In_1795);
nand U741 (N_741,In_309,In_190);
nand U742 (N_742,In_1859,In_1942);
or U743 (N_743,In_1268,In_1915);
nor U744 (N_744,In_659,In_1513);
or U745 (N_745,In_1063,In_84);
nand U746 (N_746,In_429,In_657);
or U747 (N_747,In_1284,In_58);
and U748 (N_748,In_1393,In_806);
nand U749 (N_749,In_1502,In_1077);
or U750 (N_750,In_420,In_1170);
or U751 (N_751,In_1937,In_1354);
and U752 (N_752,In_1764,In_1027);
and U753 (N_753,In_1469,In_1892);
and U754 (N_754,In_1435,In_690);
nor U755 (N_755,In_357,In_542);
or U756 (N_756,In_887,In_562);
nand U757 (N_757,In_1540,In_766);
or U758 (N_758,In_265,In_1583);
nand U759 (N_759,In_1507,In_1401);
xor U760 (N_760,In_1644,In_287);
xor U761 (N_761,In_1255,In_1365);
nor U762 (N_762,In_1851,In_1668);
xnor U763 (N_763,In_1437,In_791);
and U764 (N_764,In_1755,In_421);
or U765 (N_765,In_337,In_867);
and U766 (N_766,In_1576,In_364);
nor U767 (N_767,In_1128,In_523);
nor U768 (N_768,In_1757,In_1248);
and U769 (N_769,In_1617,In_1207);
nor U770 (N_770,In_986,In_1409);
nand U771 (N_771,In_1667,In_531);
and U772 (N_772,In_1359,In_910);
xor U773 (N_773,In_448,In_1874);
or U774 (N_774,In_259,In_1646);
xnor U775 (N_775,In_1306,In_9);
nand U776 (N_776,In_1560,In_1520);
and U777 (N_777,In_332,In_1716);
nand U778 (N_778,In_812,In_72);
or U779 (N_779,In_239,In_1944);
nand U780 (N_780,In_613,In_394);
nor U781 (N_781,In_139,In_130);
and U782 (N_782,In_1558,In_97);
or U783 (N_783,In_1551,In_857);
nor U784 (N_784,In_8,In_1577);
nand U785 (N_785,In_241,In_1108);
nor U786 (N_786,In_1030,In_675);
nor U787 (N_787,In_1431,In_157);
or U788 (N_788,In_873,In_885);
nand U789 (N_789,In_340,In_1969);
or U790 (N_790,In_1717,In_1889);
xnor U791 (N_791,In_1852,In_1701);
or U792 (N_792,In_677,In_1521);
or U793 (N_793,In_1125,In_658);
nand U794 (N_794,In_795,In_1291);
or U795 (N_795,In_1811,In_1243);
xnor U796 (N_796,In_1768,In_1711);
xor U797 (N_797,In_37,In_386);
nand U798 (N_798,In_903,In_10);
nand U799 (N_799,In_1626,In_2);
nor U800 (N_800,In_1155,In_1539);
and U801 (N_801,In_1978,In_1685);
and U802 (N_802,In_1208,In_233);
nand U803 (N_803,In_968,In_441);
or U804 (N_804,In_296,In_1156);
nor U805 (N_805,In_33,In_591);
nand U806 (N_806,In_636,In_1295);
nor U807 (N_807,In_1336,In_633);
nor U808 (N_808,In_70,In_283);
and U809 (N_809,In_914,In_664);
and U810 (N_810,In_222,In_1079);
nand U811 (N_811,In_1938,In_1655);
or U812 (N_812,In_1538,In_210);
nand U813 (N_813,In_453,In_1934);
xnor U814 (N_814,In_458,In_760);
xor U815 (N_815,In_610,In_369);
nand U816 (N_816,In_1792,In_1241);
nor U817 (N_817,In_651,In_1433);
and U818 (N_818,In_581,In_605);
nor U819 (N_819,In_437,In_424);
and U820 (N_820,In_179,In_1095);
or U821 (N_821,In_418,In_1253);
nand U822 (N_822,In_592,In_52);
and U823 (N_823,In_897,In_197);
or U824 (N_824,In_1825,In_1282);
or U825 (N_825,In_871,In_920);
or U826 (N_826,In_809,In_135);
nand U827 (N_827,In_1820,In_622);
nor U828 (N_828,In_1341,In_1492);
and U829 (N_829,In_1868,In_114);
nand U830 (N_830,In_5,In_1898);
nand U831 (N_831,In_1439,In_1974);
nor U832 (N_832,In_926,In_1362);
or U833 (N_833,In_1589,In_237);
xnor U834 (N_834,In_0,In_1227);
nor U835 (N_835,In_788,In_235);
nor U836 (N_836,In_922,In_771);
nor U837 (N_837,In_683,In_1276);
xnor U838 (N_838,In_1704,In_550);
nor U839 (N_839,In_468,In_957);
and U840 (N_840,In_1360,In_143);
nand U841 (N_841,In_545,In_1153);
nand U842 (N_842,In_402,In_1332);
nand U843 (N_843,In_1697,In_1316);
and U844 (N_844,In_1187,In_1475);
nand U845 (N_845,In_1959,In_1196);
or U846 (N_846,In_1763,In_818);
and U847 (N_847,In_569,In_822);
or U848 (N_848,In_1262,In_1113);
and U849 (N_849,In_698,In_1000);
nor U850 (N_850,In_707,In_840);
or U851 (N_851,In_329,In_1468);
xnor U852 (N_852,In_1970,In_113);
or U853 (N_853,In_21,In_1578);
xnor U854 (N_854,In_1477,In_1271);
nor U855 (N_855,In_1602,In_772);
nor U856 (N_856,In_371,In_607);
nor U857 (N_857,In_1278,In_551);
nor U858 (N_858,In_1029,In_372);
nor U859 (N_859,In_1794,In_350);
nor U860 (N_860,In_1686,In_725);
and U861 (N_861,In_1506,In_1247);
nor U862 (N_862,In_379,In_289);
xnor U863 (N_863,In_876,In_750);
or U864 (N_864,In_359,In_1918);
xnor U865 (N_865,In_941,In_408);
or U866 (N_866,In_1200,In_1949);
and U867 (N_867,In_1628,In_1034);
and U868 (N_868,In_1236,In_1804);
nor U869 (N_869,In_140,In_1906);
nand U870 (N_870,In_305,In_1672);
or U871 (N_871,In_1675,In_1698);
nand U872 (N_872,In_1948,In_676);
and U873 (N_873,In_311,In_367);
nand U874 (N_874,In_268,In_1089);
nor U875 (N_875,In_945,In_1274);
or U876 (N_876,In_1735,In_1099);
and U877 (N_877,In_796,In_1403);
or U878 (N_878,In_1381,In_147);
or U879 (N_879,In_1776,In_1509);
nand U880 (N_880,In_1620,In_1782);
or U881 (N_881,In_574,In_691);
and U882 (N_882,In_281,In_946);
nand U883 (N_883,In_883,In_1528);
or U884 (N_884,In_271,In_1747);
nand U885 (N_885,In_913,In_1694);
nand U886 (N_886,In_86,In_549);
nor U887 (N_887,In_1983,In_1599);
nor U888 (N_888,In_761,In_557);
nand U889 (N_889,In_1461,In_1388);
and U890 (N_890,In_1745,In_627);
nand U891 (N_891,In_1484,In_1250);
and U892 (N_892,In_1840,In_1497);
nand U893 (N_893,In_471,In_1950);
nor U894 (N_894,In_711,In_1590);
and U895 (N_895,In_69,In_22);
or U896 (N_896,In_954,In_1806);
xnor U897 (N_897,In_1181,In_1195);
nor U898 (N_898,In_1323,In_820);
and U899 (N_899,In_1575,In_778);
nor U900 (N_900,In_1319,In_1495);
nor U901 (N_901,In_1733,In_624);
nor U902 (N_902,In_552,In_1985);
nand U903 (N_903,In_1159,In_1482);
nand U904 (N_904,In_1861,In_1826);
nor U905 (N_905,In_1174,In_1588);
and U906 (N_906,In_164,In_180);
nand U907 (N_907,In_1395,In_28);
and U908 (N_908,In_889,In_1071);
xnor U909 (N_909,In_431,In_1500);
nand U910 (N_910,In_719,In_1767);
nor U911 (N_911,In_1183,In_1737);
or U912 (N_912,In_1328,In_176);
and U913 (N_913,In_1955,In_117);
nor U914 (N_914,In_1796,In_1808);
and U915 (N_915,In_80,In_1690);
nor U916 (N_916,In_573,In_1206);
nand U917 (N_917,In_865,In_1152);
and U918 (N_918,In_1823,In_1061);
or U919 (N_919,In_1457,In_1104);
and U920 (N_920,In_1526,In_1002);
xnor U921 (N_921,In_589,In_53);
and U922 (N_922,In_1415,In_1902);
xor U923 (N_923,In_1708,In_1530);
and U924 (N_924,In_334,In_90);
and U925 (N_925,In_1954,In_590);
or U926 (N_926,In_1214,In_933);
xor U927 (N_927,In_947,In_813);
nand U928 (N_928,In_1666,In_87);
nor U929 (N_929,In_1853,In_1932);
nor U930 (N_930,In_151,In_1749);
or U931 (N_931,In_1498,In_1103);
and U932 (N_932,In_1350,In_940);
or U933 (N_933,In_1829,In_1662);
xnor U934 (N_934,In_1695,In_909);
nand U935 (N_935,In_689,In_208);
and U936 (N_936,In_1487,In_751);
or U937 (N_937,In_224,In_1225);
nand U938 (N_938,In_434,In_852);
xor U939 (N_939,In_801,In_738);
and U940 (N_940,In_1894,In_1550);
xnor U941 (N_941,In_1259,In_1683);
nand U942 (N_942,In_1052,In_1370);
xnor U943 (N_943,In_895,In_629);
nand U944 (N_944,In_270,In_583);
and U945 (N_945,In_819,In_1060);
or U946 (N_946,In_952,In_211);
xor U947 (N_947,In_1036,In_961);
and U948 (N_948,In_1719,In_1691);
nor U949 (N_949,In_1746,In_298);
nand U950 (N_950,In_1522,In_1239);
or U951 (N_951,In_1392,In_1491);
and U952 (N_952,In_993,In_787);
and U953 (N_953,In_336,In_1663);
nor U954 (N_954,In_1416,In_875);
or U955 (N_955,In_1406,In_1309);
and U956 (N_956,In_1692,In_860);
and U957 (N_957,In_717,In_1164);
nor U958 (N_958,In_1287,In_193);
and U959 (N_959,In_1812,In_1723);
xor U960 (N_960,In_1384,In_906);
and U961 (N_961,In_1648,In_536);
or U962 (N_962,In_815,In_1263);
and U963 (N_963,In_1076,In_1935);
nor U964 (N_964,In_192,In_611);
or U965 (N_965,In_580,In_1338);
or U966 (N_966,In_1827,In_546);
nor U967 (N_967,In_423,In_1399);
or U968 (N_968,In_1559,In_88);
or U969 (N_969,In_1928,In_1887);
nand U970 (N_970,In_293,In_1821);
nand U971 (N_971,In_64,In_1961);
nand U972 (N_972,In_1101,In_727);
xor U973 (N_973,In_1375,In_178);
nor U974 (N_974,In_317,In_1346);
nor U975 (N_975,In_1394,In_644);
nand U976 (N_976,In_1552,In_50);
and U977 (N_977,In_124,In_1405);
nor U978 (N_978,In_1556,In_1140);
nor U979 (N_979,In_746,In_1631);
nand U980 (N_980,In_662,In_328);
or U981 (N_981,In_1305,In_245);
nand U982 (N_982,In_1569,In_216);
nor U983 (N_983,In_1054,In_1877);
xor U984 (N_984,In_533,In_824);
xnor U985 (N_985,In_521,In_1039);
nand U986 (N_986,In_821,In_319);
xnor U987 (N_987,In_879,In_1741);
and U988 (N_988,In_688,In_888);
nor U989 (N_989,In_1048,In_68);
and U990 (N_990,In_608,In_1318);
nand U991 (N_991,In_602,In_567);
or U992 (N_992,In_1614,In_1702);
xnor U993 (N_993,In_996,In_700);
or U994 (N_994,In_1272,In_34);
xnor U995 (N_995,In_1567,In_620);
nand U996 (N_996,In_248,In_723);
nand U997 (N_997,In_1486,In_864);
nor U998 (N_998,In_1869,In_1369);
or U999 (N_999,In_1361,In_1471);
and U1000 (N_1000,In_1204,In_424);
xor U1001 (N_1001,In_1739,In_708);
and U1002 (N_1002,In_829,In_348);
or U1003 (N_1003,In_1201,In_858);
nand U1004 (N_1004,In_284,In_439);
nor U1005 (N_1005,In_1087,In_1886);
and U1006 (N_1006,In_1829,In_1678);
nor U1007 (N_1007,In_576,In_872);
and U1008 (N_1008,In_1788,In_1965);
nor U1009 (N_1009,In_1628,In_1827);
xnor U1010 (N_1010,In_1229,In_476);
nand U1011 (N_1011,In_25,In_969);
xor U1012 (N_1012,In_81,In_743);
or U1013 (N_1013,In_1621,In_535);
nor U1014 (N_1014,In_1421,In_1681);
or U1015 (N_1015,In_1300,In_652);
nor U1016 (N_1016,In_1227,In_37);
nand U1017 (N_1017,In_1419,In_840);
xor U1018 (N_1018,In_1543,In_1689);
or U1019 (N_1019,In_1805,In_531);
or U1020 (N_1020,In_1384,In_1079);
nor U1021 (N_1021,In_1453,In_1737);
nand U1022 (N_1022,In_1935,In_350);
nand U1023 (N_1023,In_78,In_1196);
nor U1024 (N_1024,In_1193,In_782);
nand U1025 (N_1025,In_23,In_1363);
nand U1026 (N_1026,In_246,In_638);
and U1027 (N_1027,In_590,In_206);
and U1028 (N_1028,In_261,In_830);
xor U1029 (N_1029,In_1471,In_972);
nor U1030 (N_1030,In_1678,In_371);
nand U1031 (N_1031,In_129,In_1965);
and U1032 (N_1032,In_239,In_216);
xor U1033 (N_1033,In_1647,In_1071);
xnor U1034 (N_1034,In_410,In_335);
nand U1035 (N_1035,In_102,In_223);
nor U1036 (N_1036,In_1646,In_818);
nand U1037 (N_1037,In_194,In_196);
nor U1038 (N_1038,In_1627,In_1272);
nor U1039 (N_1039,In_258,In_849);
nand U1040 (N_1040,In_1342,In_1333);
xnor U1041 (N_1041,In_1913,In_35);
and U1042 (N_1042,In_1639,In_1348);
and U1043 (N_1043,In_1623,In_69);
and U1044 (N_1044,In_1808,In_1262);
nor U1045 (N_1045,In_948,In_812);
nor U1046 (N_1046,In_1155,In_1334);
or U1047 (N_1047,In_372,In_1790);
and U1048 (N_1048,In_1173,In_1814);
and U1049 (N_1049,In_1068,In_1607);
or U1050 (N_1050,In_337,In_1866);
xnor U1051 (N_1051,In_1397,In_196);
nand U1052 (N_1052,In_1916,In_1586);
nor U1053 (N_1053,In_1295,In_1002);
or U1054 (N_1054,In_840,In_1825);
or U1055 (N_1055,In_815,In_547);
nand U1056 (N_1056,In_56,In_622);
or U1057 (N_1057,In_98,In_705);
xnor U1058 (N_1058,In_20,In_1051);
nand U1059 (N_1059,In_1382,In_528);
xnor U1060 (N_1060,In_109,In_778);
or U1061 (N_1061,In_21,In_1131);
xor U1062 (N_1062,In_1073,In_1163);
and U1063 (N_1063,In_1865,In_1831);
xor U1064 (N_1064,In_895,In_569);
nor U1065 (N_1065,In_720,In_1423);
or U1066 (N_1066,In_221,In_1272);
or U1067 (N_1067,In_381,In_1703);
and U1068 (N_1068,In_622,In_1611);
and U1069 (N_1069,In_406,In_68);
nor U1070 (N_1070,In_120,In_1301);
and U1071 (N_1071,In_1161,In_201);
nand U1072 (N_1072,In_754,In_1686);
or U1073 (N_1073,In_1142,In_856);
xor U1074 (N_1074,In_979,In_1823);
and U1075 (N_1075,In_1483,In_1661);
or U1076 (N_1076,In_1217,In_33);
or U1077 (N_1077,In_1804,In_1595);
or U1078 (N_1078,In_1448,In_1362);
and U1079 (N_1079,In_957,In_1108);
and U1080 (N_1080,In_189,In_1367);
nor U1081 (N_1081,In_96,In_1322);
nor U1082 (N_1082,In_1766,In_306);
nand U1083 (N_1083,In_712,In_1269);
nor U1084 (N_1084,In_1874,In_1090);
xor U1085 (N_1085,In_1621,In_1228);
or U1086 (N_1086,In_345,In_1607);
and U1087 (N_1087,In_1993,In_1802);
nor U1088 (N_1088,In_867,In_1719);
and U1089 (N_1089,In_468,In_541);
nand U1090 (N_1090,In_41,In_155);
or U1091 (N_1091,In_1400,In_1943);
or U1092 (N_1092,In_1733,In_1049);
nand U1093 (N_1093,In_186,In_710);
or U1094 (N_1094,In_1315,In_1410);
nand U1095 (N_1095,In_1798,In_940);
or U1096 (N_1096,In_1323,In_1794);
or U1097 (N_1097,In_1900,In_376);
nand U1098 (N_1098,In_625,In_1647);
nor U1099 (N_1099,In_1781,In_21);
nor U1100 (N_1100,In_25,In_732);
or U1101 (N_1101,In_1085,In_643);
nand U1102 (N_1102,In_1246,In_1769);
nand U1103 (N_1103,In_1138,In_1488);
nand U1104 (N_1104,In_158,In_960);
nor U1105 (N_1105,In_1391,In_607);
xnor U1106 (N_1106,In_765,In_446);
or U1107 (N_1107,In_1109,In_1903);
nor U1108 (N_1108,In_1943,In_1260);
nor U1109 (N_1109,In_1343,In_236);
nor U1110 (N_1110,In_58,In_681);
nand U1111 (N_1111,In_1872,In_1847);
and U1112 (N_1112,In_14,In_1117);
and U1113 (N_1113,In_69,In_1543);
or U1114 (N_1114,In_672,In_172);
and U1115 (N_1115,In_708,In_1583);
or U1116 (N_1116,In_388,In_526);
xor U1117 (N_1117,In_333,In_304);
or U1118 (N_1118,In_1127,In_68);
xnor U1119 (N_1119,In_537,In_543);
nand U1120 (N_1120,In_1228,In_1364);
nand U1121 (N_1121,In_1153,In_773);
nor U1122 (N_1122,In_825,In_349);
nand U1123 (N_1123,In_1139,In_1968);
nor U1124 (N_1124,In_1654,In_736);
nor U1125 (N_1125,In_393,In_1609);
xor U1126 (N_1126,In_547,In_234);
or U1127 (N_1127,In_289,In_646);
nor U1128 (N_1128,In_32,In_700);
or U1129 (N_1129,In_109,In_103);
nand U1130 (N_1130,In_668,In_1423);
or U1131 (N_1131,In_1045,In_1808);
nor U1132 (N_1132,In_736,In_717);
xor U1133 (N_1133,In_1754,In_1941);
or U1134 (N_1134,In_1329,In_527);
nand U1135 (N_1135,In_738,In_1703);
nand U1136 (N_1136,In_950,In_123);
and U1137 (N_1137,In_335,In_319);
nor U1138 (N_1138,In_1119,In_1613);
xnor U1139 (N_1139,In_1994,In_1083);
and U1140 (N_1140,In_878,In_1833);
or U1141 (N_1141,In_1975,In_1935);
xor U1142 (N_1142,In_1390,In_1660);
nand U1143 (N_1143,In_298,In_1029);
and U1144 (N_1144,In_960,In_1422);
and U1145 (N_1145,In_1306,In_1803);
nand U1146 (N_1146,In_511,In_518);
or U1147 (N_1147,In_370,In_705);
nor U1148 (N_1148,In_701,In_608);
xnor U1149 (N_1149,In_954,In_1950);
xnor U1150 (N_1150,In_1808,In_344);
xnor U1151 (N_1151,In_1963,In_1623);
nand U1152 (N_1152,In_1501,In_218);
xnor U1153 (N_1153,In_1837,In_1461);
xor U1154 (N_1154,In_525,In_550);
nand U1155 (N_1155,In_720,In_49);
or U1156 (N_1156,In_723,In_1514);
nand U1157 (N_1157,In_1897,In_1610);
or U1158 (N_1158,In_338,In_498);
and U1159 (N_1159,In_4,In_1001);
nand U1160 (N_1160,In_113,In_178);
nand U1161 (N_1161,In_59,In_1181);
xor U1162 (N_1162,In_983,In_973);
or U1163 (N_1163,In_564,In_1464);
xnor U1164 (N_1164,In_726,In_357);
nand U1165 (N_1165,In_1811,In_1455);
nand U1166 (N_1166,In_364,In_1370);
xor U1167 (N_1167,In_1485,In_637);
nor U1168 (N_1168,In_300,In_329);
or U1169 (N_1169,In_1231,In_1668);
nor U1170 (N_1170,In_1994,In_167);
nor U1171 (N_1171,In_785,In_1433);
nor U1172 (N_1172,In_1951,In_402);
nor U1173 (N_1173,In_425,In_315);
nor U1174 (N_1174,In_100,In_1095);
xnor U1175 (N_1175,In_553,In_962);
nand U1176 (N_1176,In_587,In_792);
nand U1177 (N_1177,In_1672,In_787);
nand U1178 (N_1178,In_347,In_167);
nor U1179 (N_1179,In_1157,In_1830);
and U1180 (N_1180,In_520,In_1673);
and U1181 (N_1181,In_1799,In_828);
xor U1182 (N_1182,In_1976,In_1899);
nand U1183 (N_1183,In_1514,In_761);
and U1184 (N_1184,In_741,In_7);
nor U1185 (N_1185,In_565,In_1445);
nor U1186 (N_1186,In_672,In_1547);
nor U1187 (N_1187,In_34,In_415);
nand U1188 (N_1188,In_1284,In_670);
xor U1189 (N_1189,In_1162,In_333);
nor U1190 (N_1190,In_92,In_1328);
nand U1191 (N_1191,In_867,In_17);
and U1192 (N_1192,In_1875,In_139);
nor U1193 (N_1193,In_1520,In_336);
or U1194 (N_1194,In_815,In_196);
and U1195 (N_1195,In_1840,In_152);
nand U1196 (N_1196,In_726,In_96);
nand U1197 (N_1197,In_183,In_841);
or U1198 (N_1198,In_278,In_1880);
or U1199 (N_1199,In_985,In_703);
or U1200 (N_1200,In_1530,In_120);
or U1201 (N_1201,In_1399,In_705);
nor U1202 (N_1202,In_511,In_186);
nand U1203 (N_1203,In_1564,In_1905);
nor U1204 (N_1204,In_1873,In_1838);
or U1205 (N_1205,In_1905,In_1538);
nor U1206 (N_1206,In_1944,In_889);
nor U1207 (N_1207,In_1224,In_1841);
nand U1208 (N_1208,In_1136,In_1319);
and U1209 (N_1209,In_597,In_1350);
nand U1210 (N_1210,In_1429,In_971);
and U1211 (N_1211,In_221,In_939);
and U1212 (N_1212,In_653,In_1318);
nor U1213 (N_1213,In_1419,In_1510);
or U1214 (N_1214,In_1224,In_850);
xor U1215 (N_1215,In_641,In_339);
or U1216 (N_1216,In_1595,In_68);
or U1217 (N_1217,In_1244,In_1689);
or U1218 (N_1218,In_1632,In_241);
or U1219 (N_1219,In_384,In_488);
nor U1220 (N_1220,In_867,In_671);
nor U1221 (N_1221,In_1656,In_500);
nor U1222 (N_1222,In_852,In_524);
or U1223 (N_1223,In_1274,In_776);
xor U1224 (N_1224,In_1679,In_1004);
xor U1225 (N_1225,In_1867,In_1334);
or U1226 (N_1226,In_1862,In_187);
or U1227 (N_1227,In_1719,In_1041);
and U1228 (N_1228,In_1106,In_1163);
nor U1229 (N_1229,In_1730,In_877);
and U1230 (N_1230,In_596,In_179);
or U1231 (N_1231,In_1331,In_1685);
or U1232 (N_1232,In_892,In_1047);
or U1233 (N_1233,In_813,In_1968);
or U1234 (N_1234,In_1099,In_307);
and U1235 (N_1235,In_925,In_1823);
and U1236 (N_1236,In_1178,In_408);
nor U1237 (N_1237,In_398,In_667);
nor U1238 (N_1238,In_365,In_1786);
nor U1239 (N_1239,In_523,In_157);
nor U1240 (N_1240,In_1306,In_631);
nand U1241 (N_1241,In_1708,In_1221);
nand U1242 (N_1242,In_764,In_1513);
xor U1243 (N_1243,In_1863,In_1185);
and U1244 (N_1244,In_1928,In_701);
xor U1245 (N_1245,In_50,In_1262);
nand U1246 (N_1246,In_380,In_808);
xnor U1247 (N_1247,In_970,In_1943);
and U1248 (N_1248,In_449,In_473);
and U1249 (N_1249,In_1225,In_398);
or U1250 (N_1250,In_606,In_972);
nand U1251 (N_1251,In_408,In_1924);
nand U1252 (N_1252,In_1055,In_330);
or U1253 (N_1253,In_1269,In_1877);
nand U1254 (N_1254,In_647,In_347);
or U1255 (N_1255,In_1094,In_1101);
nand U1256 (N_1256,In_1326,In_1170);
and U1257 (N_1257,In_1051,In_413);
and U1258 (N_1258,In_1275,In_948);
or U1259 (N_1259,In_297,In_172);
nand U1260 (N_1260,In_1934,In_911);
nor U1261 (N_1261,In_1108,In_1545);
and U1262 (N_1262,In_808,In_1828);
and U1263 (N_1263,In_761,In_494);
nand U1264 (N_1264,In_1876,In_790);
or U1265 (N_1265,In_1,In_1516);
nand U1266 (N_1266,In_89,In_463);
nor U1267 (N_1267,In_1739,In_1890);
nand U1268 (N_1268,In_1378,In_164);
or U1269 (N_1269,In_1257,In_1221);
nor U1270 (N_1270,In_1191,In_1094);
and U1271 (N_1271,In_645,In_438);
and U1272 (N_1272,In_646,In_408);
or U1273 (N_1273,In_936,In_1048);
nor U1274 (N_1274,In_1154,In_775);
xnor U1275 (N_1275,In_1382,In_833);
nor U1276 (N_1276,In_593,In_1050);
nor U1277 (N_1277,In_1652,In_1932);
or U1278 (N_1278,In_1154,In_1064);
or U1279 (N_1279,In_636,In_1985);
xnor U1280 (N_1280,In_98,In_1484);
nand U1281 (N_1281,In_926,In_1628);
and U1282 (N_1282,In_1214,In_1656);
nor U1283 (N_1283,In_1019,In_1509);
nor U1284 (N_1284,In_1556,In_235);
nand U1285 (N_1285,In_1200,In_1085);
or U1286 (N_1286,In_290,In_960);
xor U1287 (N_1287,In_425,In_679);
nor U1288 (N_1288,In_478,In_1457);
xnor U1289 (N_1289,In_1411,In_1681);
and U1290 (N_1290,In_1787,In_1684);
and U1291 (N_1291,In_25,In_1135);
and U1292 (N_1292,In_1616,In_1936);
or U1293 (N_1293,In_1113,In_1231);
nor U1294 (N_1294,In_421,In_1708);
nand U1295 (N_1295,In_683,In_318);
xnor U1296 (N_1296,In_1781,In_1242);
and U1297 (N_1297,In_747,In_321);
nor U1298 (N_1298,In_912,In_1916);
nor U1299 (N_1299,In_324,In_558);
nand U1300 (N_1300,In_1915,In_613);
nand U1301 (N_1301,In_1773,In_1212);
nor U1302 (N_1302,In_1187,In_1222);
nand U1303 (N_1303,In_972,In_1197);
and U1304 (N_1304,In_1381,In_1276);
nor U1305 (N_1305,In_52,In_318);
and U1306 (N_1306,In_739,In_1611);
and U1307 (N_1307,In_979,In_1793);
nor U1308 (N_1308,In_1749,In_1492);
and U1309 (N_1309,In_1203,In_332);
and U1310 (N_1310,In_755,In_193);
and U1311 (N_1311,In_1116,In_499);
nor U1312 (N_1312,In_1105,In_1975);
and U1313 (N_1313,In_1990,In_237);
or U1314 (N_1314,In_788,In_1040);
nand U1315 (N_1315,In_1355,In_1799);
nand U1316 (N_1316,In_654,In_557);
or U1317 (N_1317,In_253,In_1586);
or U1318 (N_1318,In_1898,In_408);
nor U1319 (N_1319,In_507,In_592);
nand U1320 (N_1320,In_1049,In_1010);
nand U1321 (N_1321,In_487,In_1028);
nand U1322 (N_1322,In_1236,In_1623);
and U1323 (N_1323,In_1377,In_902);
or U1324 (N_1324,In_443,In_1685);
nand U1325 (N_1325,In_1738,In_774);
nand U1326 (N_1326,In_1843,In_753);
or U1327 (N_1327,In_703,In_1836);
xor U1328 (N_1328,In_1371,In_830);
and U1329 (N_1329,In_818,In_1302);
nand U1330 (N_1330,In_1366,In_1237);
and U1331 (N_1331,In_83,In_685);
and U1332 (N_1332,In_840,In_1946);
nand U1333 (N_1333,In_1097,In_1085);
nor U1334 (N_1334,In_924,In_1067);
or U1335 (N_1335,In_1725,In_755);
or U1336 (N_1336,In_663,In_604);
nand U1337 (N_1337,In_1704,In_166);
nor U1338 (N_1338,In_1120,In_654);
or U1339 (N_1339,In_826,In_1786);
and U1340 (N_1340,In_109,In_968);
and U1341 (N_1341,In_1657,In_156);
nor U1342 (N_1342,In_637,In_1110);
or U1343 (N_1343,In_1295,In_517);
nor U1344 (N_1344,In_978,In_42);
nand U1345 (N_1345,In_480,In_1718);
nor U1346 (N_1346,In_1758,In_1554);
xor U1347 (N_1347,In_1731,In_1558);
nor U1348 (N_1348,In_1214,In_603);
or U1349 (N_1349,In_1895,In_184);
or U1350 (N_1350,In_874,In_746);
nor U1351 (N_1351,In_255,In_1093);
and U1352 (N_1352,In_1280,In_1743);
and U1353 (N_1353,In_1336,In_300);
or U1354 (N_1354,In_597,In_1855);
and U1355 (N_1355,In_129,In_60);
or U1356 (N_1356,In_1673,In_49);
nor U1357 (N_1357,In_769,In_620);
or U1358 (N_1358,In_1314,In_708);
and U1359 (N_1359,In_1629,In_1336);
and U1360 (N_1360,In_477,In_311);
xnor U1361 (N_1361,In_424,In_833);
or U1362 (N_1362,In_1838,In_901);
and U1363 (N_1363,In_1228,In_1355);
xor U1364 (N_1364,In_1416,In_774);
nor U1365 (N_1365,In_1190,In_1153);
xnor U1366 (N_1366,In_279,In_1628);
nor U1367 (N_1367,In_1798,In_911);
or U1368 (N_1368,In_890,In_905);
xnor U1369 (N_1369,In_1631,In_1281);
and U1370 (N_1370,In_1879,In_117);
or U1371 (N_1371,In_1543,In_442);
xor U1372 (N_1372,In_1512,In_299);
or U1373 (N_1373,In_992,In_1109);
nor U1374 (N_1374,In_95,In_1309);
or U1375 (N_1375,In_1493,In_236);
nor U1376 (N_1376,In_316,In_276);
or U1377 (N_1377,In_24,In_1444);
nand U1378 (N_1378,In_1596,In_459);
and U1379 (N_1379,In_460,In_680);
and U1380 (N_1380,In_1840,In_1456);
or U1381 (N_1381,In_127,In_514);
nand U1382 (N_1382,In_1951,In_1381);
nand U1383 (N_1383,In_165,In_672);
nand U1384 (N_1384,In_1109,In_269);
nor U1385 (N_1385,In_870,In_1998);
nor U1386 (N_1386,In_1166,In_1056);
nor U1387 (N_1387,In_1309,In_1438);
nor U1388 (N_1388,In_373,In_1313);
nor U1389 (N_1389,In_1503,In_1840);
xor U1390 (N_1390,In_1720,In_776);
nor U1391 (N_1391,In_1934,In_1423);
nand U1392 (N_1392,In_90,In_272);
or U1393 (N_1393,In_1385,In_1689);
or U1394 (N_1394,In_1329,In_1528);
or U1395 (N_1395,In_131,In_1409);
nand U1396 (N_1396,In_1946,In_880);
nor U1397 (N_1397,In_155,In_1222);
nor U1398 (N_1398,In_1282,In_1864);
or U1399 (N_1399,In_1745,In_139);
nand U1400 (N_1400,In_643,In_414);
or U1401 (N_1401,In_13,In_68);
nor U1402 (N_1402,In_1551,In_1670);
or U1403 (N_1403,In_1325,In_1228);
and U1404 (N_1404,In_626,In_1071);
xor U1405 (N_1405,In_428,In_1015);
xnor U1406 (N_1406,In_1928,In_1729);
nand U1407 (N_1407,In_1358,In_1603);
nor U1408 (N_1408,In_1046,In_1194);
nor U1409 (N_1409,In_1318,In_1815);
or U1410 (N_1410,In_1217,In_83);
nand U1411 (N_1411,In_315,In_589);
and U1412 (N_1412,In_1562,In_547);
or U1413 (N_1413,In_481,In_867);
nand U1414 (N_1414,In_438,In_905);
and U1415 (N_1415,In_921,In_96);
nor U1416 (N_1416,In_1194,In_291);
nand U1417 (N_1417,In_87,In_637);
or U1418 (N_1418,In_425,In_1001);
xnor U1419 (N_1419,In_1987,In_1951);
nor U1420 (N_1420,In_676,In_1039);
nor U1421 (N_1421,In_585,In_46);
and U1422 (N_1422,In_592,In_1462);
xor U1423 (N_1423,In_1346,In_49);
nand U1424 (N_1424,In_584,In_1824);
and U1425 (N_1425,In_881,In_992);
or U1426 (N_1426,In_494,In_1471);
or U1427 (N_1427,In_583,In_70);
nand U1428 (N_1428,In_974,In_466);
xor U1429 (N_1429,In_1940,In_214);
xor U1430 (N_1430,In_1694,In_940);
or U1431 (N_1431,In_1184,In_1185);
nor U1432 (N_1432,In_1473,In_177);
nor U1433 (N_1433,In_1987,In_1400);
nand U1434 (N_1434,In_1718,In_1026);
nor U1435 (N_1435,In_1473,In_233);
nor U1436 (N_1436,In_1985,In_1913);
nand U1437 (N_1437,In_1499,In_464);
and U1438 (N_1438,In_560,In_317);
and U1439 (N_1439,In_628,In_956);
xor U1440 (N_1440,In_343,In_1807);
or U1441 (N_1441,In_1664,In_1869);
and U1442 (N_1442,In_1482,In_321);
and U1443 (N_1443,In_1479,In_1788);
nand U1444 (N_1444,In_1297,In_1803);
nand U1445 (N_1445,In_607,In_1781);
nor U1446 (N_1446,In_246,In_235);
or U1447 (N_1447,In_1865,In_1333);
nand U1448 (N_1448,In_18,In_126);
or U1449 (N_1449,In_1941,In_1649);
nor U1450 (N_1450,In_1662,In_51);
xor U1451 (N_1451,In_1106,In_361);
and U1452 (N_1452,In_1985,In_1880);
nand U1453 (N_1453,In_18,In_469);
xnor U1454 (N_1454,In_839,In_1885);
and U1455 (N_1455,In_1535,In_1915);
nor U1456 (N_1456,In_848,In_151);
and U1457 (N_1457,In_1029,In_1273);
or U1458 (N_1458,In_355,In_1621);
nand U1459 (N_1459,In_1946,In_1649);
and U1460 (N_1460,In_1043,In_276);
or U1461 (N_1461,In_1990,In_437);
nor U1462 (N_1462,In_478,In_938);
or U1463 (N_1463,In_991,In_1431);
nand U1464 (N_1464,In_178,In_1496);
nor U1465 (N_1465,In_176,In_1937);
nand U1466 (N_1466,In_939,In_1950);
and U1467 (N_1467,In_19,In_196);
nor U1468 (N_1468,In_1842,In_823);
or U1469 (N_1469,In_700,In_1045);
and U1470 (N_1470,In_281,In_1475);
nor U1471 (N_1471,In_414,In_519);
or U1472 (N_1472,In_1399,In_276);
or U1473 (N_1473,In_1418,In_862);
nand U1474 (N_1474,In_1173,In_416);
or U1475 (N_1475,In_906,In_1984);
and U1476 (N_1476,In_1665,In_1485);
nand U1477 (N_1477,In_1926,In_1866);
and U1478 (N_1478,In_1656,In_1684);
or U1479 (N_1479,In_1919,In_1423);
nand U1480 (N_1480,In_1665,In_1563);
xor U1481 (N_1481,In_1753,In_300);
and U1482 (N_1482,In_934,In_388);
nand U1483 (N_1483,In_448,In_1244);
or U1484 (N_1484,In_582,In_1771);
nand U1485 (N_1485,In_370,In_916);
nor U1486 (N_1486,In_818,In_1132);
and U1487 (N_1487,In_422,In_190);
nand U1488 (N_1488,In_597,In_357);
or U1489 (N_1489,In_483,In_615);
nor U1490 (N_1490,In_668,In_197);
nor U1491 (N_1491,In_220,In_1452);
nor U1492 (N_1492,In_811,In_124);
nand U1493 (N_1493,In_1282,In_1905);
or U1494 (N_1494,In_980,In_151);
or U1495 (N_1495,In_490,In_1646);
xor U1496 (N_1496,In_409,In_86);
nor U1497 (N_1497,In_1024,In_1195);
or U1498 (N_1498,In_653,In_815);
nand U1499 (N_1499,In_1324,In_1282);
nor U1500 (N_1500,In_349,In_1837);
nand U1501 (N_1501,In_719,In_625);
xor U1502 (N_1502,In_1287,In_371);
xnor U1503 (N_1503,In_870,In_1966);
and U1504 (N_1504,In_217,In_1509);
nor U1505 (N_1505,In_985,In_513);
xor U1506 (N_1506,In_266,In_131);
and U1507 (N_1507,In_1247,In_362);
and U1508 (N_1508,In_1936,In_1339);
nand U1509 (N_1509,In_14,In_369);
and U1510 (N_1510,In_163,In_932);
and U1511 (N_1511,In_648,In_1316);
xor U1512 (N_1512,In_159,In_770);
or U1513 (N_1513,In_763,In_777);
or U1514 (N_1514,In_1643,In_1898);
and U1515 (N_1515,In_1939,In_910);
and U1516 (N_1516,In_375,In_876);
and U1517 (N_1517,In_671,In_207);
or U1518 (N_1518,In_1602,In_924);
nand U1519 (N_1519,In_116,In_976);
nor U1520 (N_1520,In_337,In_1334);
nor U1521 (N_1521,In_1664,In_175);
or U1522 (N_1522,In_785,In_399);
nor U1523 (N_1523,In_1017,In_111);
xor U1524 (N_1524,In_1241,In_1479);
or U1525 (N_1525,In_128,In_1030);
and U1526 (N_1526,In_704,In_146);
nand U1527 (N_1527,In_278,In_1184);
or U1528 (N_1528,In_854,In_608);
and U1529 (N_1529,In_1575,In_1894);
nor U1530 (N_1530,In_371,In_291);
nor U1531 (N_1531,In_907,In_906);
xnor U1532 (N_1532,In_1908,In_1977);
nand U1533 (N_1533,In_660,In_1078);
nor U1534 (N_1534,In_1082,In_1312);
and U1535 (N_1535,In_937,In_1978);
nand U1536 (N_1536,In_1751,In_1960);
or U1537 (N_1537,In_1461,In_1439);
nand U1538 (N_1538,In_84,In_1680);
and U1539 (N_1539,In_393,In_1879);
and U1540 (N_1540,In_1448,In_969);
xor U1541 (N_1541,In_562,In_841);
nor U1542 (N_1542,In_1815,In_1182);
nand U1543 (N_1543,In_1568,In_1523);
and U1544 (N_1544,In_348,In_183);
and U1545 (N_1545,In_1657,In_1771);
nor U1546 (N_1546,In_380,In_1986);
nor U1547 (N_1547,In_244,In_1670);
and U1548 (N_1548,In_1176,In_1769);
nor U1549 (N_1549,In_203,In_63);
or U1550 (N_1550,In_1074,In_1982);
nand U1551 (N_1551,In_160,In_4);
nand U1552 (N_1552,In_788,In_748);
nor U1553 (N_1553,In_1936,In_122);
nand U1554 (N_1554,In_591,In_1919);
or U1555 (N_1555,In_1173,In_962);
nor U1556 (N_1556,In_291,In_632);
nand U1557 (N_1557,In_1868,In_1675);
or U1558 (N_1558,In_691,In_270);
nor U1559 (N_1559,In_1110,In_1858);
and U1560 (N_1560,In_100,In_645);
nor U1561 (N_1561,In_584,In_739);
and U1562 (N_1562,In_543,In_1796);
or U1563 (N_1563,In_683,In_1236);
nand U1564 (N_1564,In_732,In_676);
and U1565 (N_1565,In_1024,In_389);
nor U1566 (N_1566,In_1712,In_991);
and U1567 (N_1567,In_1313,In_1083);
nor U1568 (N_1568,In_1314,In_1987);
or U1569 (N_1569,In_860,In_657);
or U1570 (N_1570,In_1114,In_1497);
and U1571 (N_1571,In_509,In_554);
and U1572 (N_1572,In_1093,In_1458);
and U1573 (N_1573,In_75,In_177);
or U1574 (N_1574,In_365,In_909);
nor U1575 (N_1575,In_496,In_1535);
nand U1576 (N_1576,In_1161,In_477);
and U1577 (N_1577,In_1659,In_558);
nor U1578 (N_1578,In_1141,In_1426);
and U1579 (N_1579,In_697,In_409);
nor U1580 (N_1580,In_1444,In_378);
and U1581 (N_1581,In_186,In_625);
and U1582 (N_1582,In_1031,In_592);
nand U1583 (N_1583,In_1014,In_1594);
or U1584 (N_1584,In_1768,In_980);
nand U1585 (N_1585,In_1029,In_759);
or U1586 (N_1586,In_345,In_703);
nor U1587 (N_1587,In_1939,In_956);
nor U1588 (N_1588,In_1181,In_1193);
nand U1589 (N_1589,In_536,In_1479);
nand U1590 (N_1590,In_1698,In_763);
and U1591 (N_1591,In_83,In_1412);
or U1592 (N_1592,In_1295,In_874);
nor U1593 (N_1593,In_1689,In_777);
nor U1594 (N_1594,In_634,In_1780);
xnor U1595 (N_1595,In_154,In_1841);
nor U1596 (N_1596,In_1376,In_1244);
nand U1597 (N_1597,In_910,In_1272);
nand U1598 (N_1598,In_1268,In_938);
or U1599 (N_1599,In_102,In_1082);
nand U1600 (N_1600,In_1548,In_913);
nor U1601 (N_1601,In_1783,In_25);
and U1602 (N_1602,In_262,In_1715);
or U1603 (N_1603,In_490,In_221);
nand U1604 (N_1604,In_1919,In_22);
and U1605 (N_1605,In_732,In_777);
and U1606 (N_1606,In_202,In_1805);
and U1607 (N_1607,In_1665,In_1620);
nand U1608 (N_1608,In_1590,In_1750);
and U1609 (N_1609,In_1837,In_1583);
or U1610 (N_1610,In_1397,In_670);
nor U1611 (N_1611,In_1208,In_379);
nor U1612 (N_1612,In_1271,In_1199);
nand U1613 (N_1613,In_78,In_1386);
and U1614 (N_1614,In_270,In_334);
nand U1615 (N_1615,In_467,In_1323);
nand U1616 (N_1616,In_1040,In_1652);
nand U1617 (N_1617,In_425,In_509);
and U1618 (N_1618,In_1585,In_682);
and U1619 (N_1619,In_1700,In_584);
or U1620 (N_1620,In_188,In_638);
xnor U1621 (N_1621,In_1476,In_1696);
and U1622 (N_1622,In_977,In_476);
and U1623 (N_1623,In_1473,In_1720);
or U1624 (N_1624,In_1729,In_1526);
or U1625 (N_1625,In_25,In_303);
and U1626 (N_1626,In_1051,In_1131);
nor U1627 (N_1627,In_535,In_1265);
or U1628 (N_1628,In_1258,In_811);
nand U1629 (N_1629,In_72,In_1090);
xor U1630 (N_1630,In_1776,In_381);
nor U1631 (N_1631,In_1171,In_862);
nor U1632 (N_1632,In_448,In_754);
and U1633 (N_1633,In_179,In_1346);
nor U1634 (N_1634,In_1505,In_1414);
or U1635 (N_1635,In_156,In_1656);
nor U1636 (N_1636,In_1492,In_172);
nand U1637 (N_1637,In_1904,In_1139);
or U1638 (N_1638,In_38,In_1522);
xor U1639 (N_1639,In_427,In_1303);
and U1640 (N_1640,In_1024,In_329);
nor U1641 (N_1641,In_412,In_140);
nor U1642 (N_1642,In_1061,In_1758);
and U1643 (N_1643,In_1874,In_685);
nor U1644 (N_1644,In_1898,In_1743);
nor U1645 (N_1645,In_1903,In_1444);
nand U1646 (N_1646,In_513,In_1223);
nor U1647 (N_1647,In_1043,In_1784);
nand U1648 (N_1648,In_1108,In_65);
nand U1649 (N_1649,In_1259,In_1218);
and U1650 (N_1650,In_532,In_965);
nor U1651 (N_1651,In_462,In_1488);
or U1652 (N_1652,In_1605,In_752);
or U1653 (N_1653,In_1383,In_1454);
or U1654 (N_1654,In_1039,In_1291);
or U1655 (N_1655,In_1717,In_109);
nand U1656 (N_1656,In_1818,In_1708);
or U1657 (N_1657,In_1493,In_694);
and U1658 (N_1658,In_1196,In_292);
nor U1659 (N_1659,In_27,In_1772);
and U1660 (N_1660,In_877,In_1989);
xor U1661 (N_1661,In_1052,In_1198);
nor U1662 (N_1662,In_175,In_1344);
nor U1663 (N_1663,In_950,In_1229);
nor U1664 (N_1664,In_314,In_1654);
xor U1665 (N_1665,In_107,In_465);
and U1666 (N_1666,In_1082,In_1234);
or U1667 (N_1667,In_1136,In_348);
nand U1668 (N_1668,In_1582,In_617);
and U1669 (N_1669,In_483,In_608);
nor U1670 (N_1670,In_306,In_1713);
nand U1671 (N_1671,In_1582,In_1449);
or U1672 (N_1672,In_1633,In_1592);
nand U1673 (N_1673,In_762,In_1584);
nor U1674 (N_1674,In_1124,In_1584);
or U1675 (N_1675,In_153,In_1685);
xor U1676 (N_1676,In_1502,In_1110);
or U1677 (N_1677,In_906,In_873);
or U1678 (N_1678,In_1474,In_858);
nor U1679 (N_1679,In_56,In_430);
or U1680 (N_1680,In_268,In_448);
nor U1681 (N_1681,In_145,In_63);
nor U1682 (N_1682,In_598,In_1735);
nand U1683 (N_1683,In_1108,In_896);
or U1684 (N_1684,In_489,In_369);
nor U1685 (N_1685,In_718,In_488);
nand U1686 (N_1686,In_1830,In_495);
or U1687 (N_1687,In_48,In_1856);
or U1688 (N_1688,In_1582,In_1941);
or U1689 (N_1689,In_42,In_1246);
xnor U1690 (N_1690,In_1438,In_299);
and U1691 (N_1691,In_680,In_723);
nor U1692 (N_1692,In_67,In_234);
nand U1693 (N_1693,In_209,In_1424);
and U1694 (N_1694,In_31,In_1854);
or U1695 (N_1695,In_961,In_1070);
and U1696 (N_1696,In_404,In_149);
nor U1697 (N_1697,In_439,In_1993);
or U1698 (N_1698,In_240,In_1572);
nand U1699 (N_1699,In_1168,In_968);
nor U1700 (N_1700,In_79,In_9);
and U1701 (N_1701,In_11,In_733);
or U1702 (N_1702,In_386,In_1986);
nor U1703 (N_1703,In_1012,In_62);
nor U1704 (N_1704,In_1038,In_388);
xor U1705 (N_1705,In_229,In_678);
nand U1706 (N_1706,In_1223,In_580);
or U1707 (N_1707,In_383,In_940);
or U1708 (N_1708,In_1927,In_74);
nor U1709 (N_1709,In_1932,In_1091);
and U1710 (N_1710,In_1196,In_1139);
and U1711 (N_1711,In_1872,In_44);
nor U1712 (N_1712,In_1630,In_1852);
nand U1713 (N_1713,In_500,In_1296);
xnor U1714 (N_1714,In_1384,In_1609);
nand U1715 (N_1715,In_220,In_1756);
nand U1716 (N_1716,In_856,In_1768);
and U1717 (N_1717,In_363,In_574);
nand U1718 (N_1718,In_1132,In_1097);
nor U1719 (N_1719,In_1297,In_899);
nand U1720 (N_1720,In_1879,In_1007);
nand U1721 (N_1721,In_1426,In_510);
nor U1722 (N_1722,In_526,In_40);
nand U1723 (N_1723,In_1147,In_1262);
xnor U1724 (N_1724,In_629,In_1013);
xor U1725 (N_1725,In_1124,In_205);
nand U1726 (N_1726,In_479,In_1544);
xnor U1727 (N_1727,In_1123,In_1687);
or U1728 (N_1728,In_269,In_56);
nand U1729 (N_1729,In_266,In_622);
nand U1730 (N_1730,In_167,In_1457);
or U1731 (N_1731,In_1117,In_901);
and U1732 (N_1732,In_58,In_1382);
nor U1733 (N_1733,In_1441,In_769);
nand U1734 (N_1734,In_250,In_1690);
and U1735 (N_1735,In_377,In_1408);
or U1736 (N_1736,In_1410,In_1480);
xor U1737 (N_1737,In_49,In_462);
nor U1738 (N_1738,In_808,In_7);
and U1739 (N_1739,In_1827,In_299);
nor U1740 (N_1740,In_1492,In_1759);
or U1741 (N_1741,In_1667,In_868);
or U1742 (N_1742,In_213,In_1350);
or U1743 (N_1743,In_617,In_1758);
and U1744 (N_1744,In_436,In_1116);
xnor U1745 (N_1745,In_397,In_1704);
nor U1746 (N_1746,In_57,In_973);
nor U1747 (N_1747,In_1751,In_327);
nand U1748 (N_1748,In_969,In_1716);
nor U1749 (N_1749,In_916,In_1422);
nor U1750 (N_1750,In_307,In_613);
and U1751 (N_1751,In_1637,In_173);
and U1752 (N_1752,In_1358,In_1701);
nor U1753 (N_1753,In_158,In_1288);
nor U1754 (N_1754,In_688,In_1060);
nand U1755 (N_1755,In_1805,In_1320);
and U1756 (N_1756,In_968,In_1619);
nand U1757 (N_1757,In_1209,In_634);
nor U1758 (N_1758,In_1823,In_689);
and U1759 (N_1759,In_1857,In_768);
nand U1760 (N_1760,In_902,In_1827);
nand U1761 (N_1761,In_543,In_461);
nor U1762 (N_1762,In_1544,In_517);
nor U1763 (N_1763,In_1426,In_305);
nand U1764 (N_1764,In_1547,In_1015);
or U1765 (N_1765,In_799,In_1827);
nand U1766 (N_1766,In_390,In_1711);
or U1767 (N_1767,In_1661,In_1829);
and U1768 (N_1768,In_849,In_1236);
nand U1769 (N_1769,In_1059,In_647);
nand U1770 (N_1770,In_711,In_1324);
nand U1771 (N_1771,In_532,In_1267);
nand U1772 (N_1772,In_1032,In_1163);
nor U1773 (N_1773,In_1503,In_1691);
and U1774 (N_1774,In_1986,In_593);
and U1775 (N_1775,In_721,In_792);
and U1776 (N_1776,In_1910,In_221);
xnor U1777 (N_1777,In_352,In_225);
or U1778 (N_1778,In_991,In_1118);
xor U1779 (N_1779,In_114,In_1335);
nand U1780 (N_1780,In_1384,In_1529);
and U1781 (N_1781,In_1556,In_244);
nand U1782 (N_1782,In_1282,In_309);
or U1783 (N_1783,In_1220,In_591);
nand U1784 (N_1784,In_809,In_683);
nand U1785 (N_1785,In_1889,In_497);
and U1786 (N_1786,In_1700,In_154);
nor U1787 (N_1787,In_1041,In_554);
and U1788 (N_1788,In_1057,In_107);
nor U1789 (N_1789,In_952,In_668);
and U1790 (N_1790,In_1707,In_18);
and U1791 (N_1791,In_1815,In_778);
xnor U1792 (N_1792,In_605,In_907);
and U1793 (N_1793,In_349,In_1445);
and U1794 (N_1794,In_1346,In_1684);
nand U1795 (N_1795,In_618,In_339);
nand U1796 (N_1796,In_938,In_92);
and U1797 (N_1797,In_74,In_109);
or U1798 (N_1798,In_163,In_993);
nor U1799 (N_1799,In_1090,In_1459);
or U1800 (N_1800,In_1269,In_292);
nor U1801 (N_1801,In_1162,In_696);
or U1802 (N_1802,In_836,In_846);
nand U1803 (N_1803,In_144,In_338);
or U1804 (N_1804,In_419,In_1060);
nor U1805 (N_1805,In_783,In_203);
or U1806 (N_1806,In_1277,In_518);
nand U1807 (N_1807,In_643,In_1722);
and U1808 (N_1808,In_1862,In_643);
nor U1809 (N_1809,In_1248,In_1956);
nor U1810 (N_1810,In_1789,In_1494);
nor U1811 (N_1811,In_1055,In_570);
nand U1812 (N_1812,In_1111,In_270);
xnor U1813 (N_1813,In_1783,In_672);
or U1814 (N_1814,In_317,In_249);
nand U1815 (N_1815,In_1733,In_4);
nand U1816 (N_1816,In_1428,In_1444);
nand U1817 (N_1817,In_552,In_575);
nor U1818 (N_1818,In_1285,In_600);
nor U1819 (N_1819,In_1671,In_1372);
nand U1820 (N_1820,In_535,In_1155);
and U1821 (N_1821,In_1461,In_252);
xnor U1822 (N_1822,In_120,In_1696);
or U1823 (N_1823,In_1719,In_238);
or U1824 (N_1824,In_895,In_1002);
and U1825 (N_1825,In_1835,In_1374);
or U1826 (N_1826,In_1794,In_1399);
or U1827 (N_1827,In_1577,In_1272);
nand U1828 (N_1828,In_261,In_650);
or U1829 (N_1829,In_242,In_295);
or U1830 (N_1830,In_242,In_1667);
and U1831 (N_1831,In_1501,In_1405);
nand U1832 (N_1832,In_1434,In_670);
nor U1833 (N_1833,In_681,In_313);
nor U1834 (N_1834,In_972,In_1251);
or U1835 (N_1835,In_1165,In_1674);
or U1836 (N_1836,In_1238,In_575);
or U1837 (N_1837,In_1149,In_766);
nand U1838 (N_1838,In_227,In_1398);
xnor U1839 (N_1839,In_291,In_568);
nor U1840 (N_1840,In_1572,In_425);
nor U1841 (N_1841,In_1764,In_237);
or U1842 (N_1842,In_1350,In_937);
nand U1843 (N_1843,In_1988,In_1199);
nand U1844 (N_1844,In_1697,In_2);
and U1845 (N_1845,In_1164,In_1305);
nor U1846 (N_1846,In_234,In_116);
nor U1847 (N_1847,In_1944,In_1488);
xnor U1848 (N_1848,In_843,In_1166);
nor U1849 (N_1849,In_679,In_1030);
nand U1850 (N_1850,In_1683,In_1327);
or U1851 (N_1851,In_835,In_1170);
nand U1852 (N_1852,In_1849,In_363);
nor U1853 (N_1853,In_1843,In_1667);
nor U1854 (N_1854,In_1977,In_54);
xnor U1855 (N_1855,In_857,In_877);
nor U1856 (N_1856,In_1512,In_181);
xor U1857 (N_1857,In_228,In_895);
and U1858 (N_1858,In_1819,In_1049);
xnor U1859 (N_1859,In_733,In_1242);
nand U1860 (N_1860,In_1975,In_892);
xor U1861 (N_1861,In_1846,In_1549);
and U1862 (N_1862,In_1204,In_1909);
nand U1863 (N_1863,In_472,In_1676);
nor U1864 (N_1864,In_904,In_80);
nand U1865 (N_1865,In_462,In_444);
nand U1866 (N_1866,In_117,In_294);
xnor U1867 (N_1867,In_1298,In_522);
or U1868 (N_1868,In_1655,In_445);
or U1869 (N_1869,In_1110,In_955);
nand U1870 (N_1870,In_1684,In_566);
or U1871 (N_1871,In_518,In_869);
xor U1872 (N_1872,In_1515,In_1944);
and U1873 (N_1873,In_1282,In_937);
xnor U1874 (N_1874,In_1164,In_258);
nand U1875 (N_1875,In_111,In_659);
or U1876 (N_1876,In_705,In_416);
nor U1877 (N_1877,In_229,In_1376);
xor U1878 (N_1878,In_252,In_340);
and U1879 (N_1879,In_1892,In_1485);
xor U1880 (N_1880,In_708,In_707);
or U1881 (N_1881,In_606,In_737);
and U1882 (N_1882,In_538,In_287);
nor U1883 (N_1883,In_1344,In_344);
nor U1884 (N_1884,In_879,In_1500);
nor U1885 (N_1885,In_1445,In_796);
or U1886 (N_1886,In_1893,In_915);
nand U1887 (N_1887,In_168,In_310);
xor U1888 (N_1888,In_1883,In_103);
nor U1889 (N_1889,In_517,In_1211);
and U1890 (N_1890,In_535,In_584);
or U1891 (N_1891,In_1348,In_464);
nor U1892 (N_1892,In_972,In_1159);
nor U1893 (N_1893,In_1833,In_1581);
and U1894 (N_1894,In_998,In_1973);
nor U1895 (N_1895,In_222,In_1388);
or U1896 (N_1896,In_1941,In_962);
and U1897 (N_1897,In_167,In_1517);
and U1898 (N_1898,In_1159,In_2);
or U1899 (N_1899,In_1056,In_163);
and U1900 (N_1900,In_1726,In_1311);
nand U1901 (N_1901,In_757,In_554);
nor U1902 (N_1902,In_1154,In_1597);
and U1903 (N_1903,In_140,In_321);
or U1904 (N_1904,In_574,In_293);
nor U1905 (N_1905,In_1270,In_840);
nor U1906 (N_1906,In_1581,In_325);
and U1907 (N_1907,In_617,In_960);
nor U1908 (N_1908,In_270,In_683);
and U1909 (N_1909,In_257,In_804);
nor U1910 (N_1910,In_1214,In_1941);
and U1911 (N_1911,In_146,In_1879);
nand U1912 (N_1912,In_1821,In_566);
and U1913 (N_1913,In_278,In_973);
or U1914 (N_1914,In_1096,In_1557);
nand U1915 (N_1915,In_76,In_1973);
nor U1916 (N_1916,In_17,In_1548);
and U1917 (N_1917,In_1173,In_87);
nand U1918 (N_1918,In_1230,In_1147);
or U1919 (N_1919,In_580,In_1317);
and U1920 (N_1920,In_1589,In_466);
and U1921 (N_1921,In_1547,In_277);
nand U1922 (N_1922,In_1407,In_1644);
or U1923 (N_1923,In_196,In_606);
or U1924 (N_1924,In_622,In_772);
nand U1925 (N_1925,In_754,In_1555);
xnor U1926 (N_1926,In_1677,In_1761);
nor U1927 (N_1927,In_733,In_1661);
nand U1928 (N_1928,In_355,In_244);
nand U1929 (N_1929,In_1614,In_669);
nand U1930 (N_1930,In_1722,In_76);
nor U1931 (N_1931,In_1045,In_1178);
nand U1932 (N_1932,In_70,In_655);
or U1933 (N_1933,In_1795,In_1387);
and U1934 (N_1934,In_654,In_1337);
xor U1935 (N_1935,In_743,In_246);
or U1936 (N_1936,In_1510,In_987);
and U1937 (N_1937,In_1657,In_1170);
nor U1938 (N_1938,In_591,In_976);
or U1939 (N_1939,In_1788,In_1220);
nand U1940 (N_1940,In_626,In_1700);
or U1941 (N_1941,In_1040,In_1599);
nand U1942 (N_1942,In_1681,In_1309);
nor U1943 (N_1943,In_497,In_1496);
nor U1944 (N_1944,In_1001,In_119);
or U1945 (N_1945,In_92,In_1471);
and U1946 (N_1946,In_129,In_642);
xor U1947 (N_1947,In_1032,In_1803);
nand U1948 (N_1948,In_1931,In_181);
and U1949 (N_1949,In_1311,In_550);
or U1950 (N_1950,In_1005,In_1972);
nand U1951 (N_1951,In_715,In_293);
or U1952 (N_1952,In_762,In_554);
nand U1953 (N_1953,In_783,In_347);
and U1954 (N_1954,In_1728,In_1831);
nor U1955 (N_1955,In_101,In_1475);
and U1956 (N_1956,In_1933,In_1683);
and U1957 (N_1957,In_218,In_1268);
or U1958 (N_1958,In_406,In_877);
nor U1959 (N_1959,In_1161,In_906);
xnor U1960 (N_1960,In_731,In_1490);
nand U1961 (N_1961,In_1653,In_852);
or U1962 (N_1962,In_1078,In_1607);
nor U1963 (N_1963,In_826,In_991);
nand U1964 (N_1964,In_531,In_161);
or U1965 (N_1965,In_659,In_1203);
nand U1966 (N_1966,In_667,In_1073);
nand U1967 (N_1967,In_717,In_980);
nand U1968 (N_1968,In_1715,In_1668);
nand U1969 (N_1969,In_535,In_1714);
or U1970 (N_1970,In_578,In_1206);
or U1971 (N_1971,In_1669,In_1126);
or U1972 (N_1972,In_1025,In_353);
nor U1973 (N_1973,In_1317,In_1536);
xor U1974 (N_1974,In_143,In_741);
nand U1975 (N_1975,In_1981,In_201);
and U1976 (N_1976,In_301,In_457);
nor U1977 (N_1977,In_462,In_1149);
xnor U1978 (N_1978,In_1011,In_864);
nand U1979 (N_1979,In_1071,In_351);
nand U1980 (N_1980,In_1484,In_1418);
or U1981 (N_1981,In_1663,In_1097);
nor U1982 (N_1982,In_1997,In_1231);
xnor U1983 (N_1983,In_1847,In_526);
or U1984 (N_1984,In_502,In_361);
nand U1985 (N_1985,In_1648,In_1112);
xnor U1986 (N_1986,In_1920,In_920);
nand U1987 (N_1987,In_414,In_1973);
or U1988 (N_1988,In_319,In_741);
or U1989 (N_1989,In_1058,In_1968);
and U1990 (N_1990,In_1310,In_295);
nor U1991 (N_1991,In_161,In_1130);
and U1992 (N_1992,In_1957,In_513);
and U1993 (N_1993,In_1406,In_1059);
nor U1994 (N_1994,In_330,In_1961);
nor U1995 (N_1995,In_169,In_1984);
nand U1996 (N_1996,In_545,In_1290);
nor U1997 (N_1997,In_1458,In_1356);
nor U1998 (N_1998,In_332,In_1005);
nor U1999 (N_1999,In_339,In_632);
or U2000 (N_2000,In_501,In_1352);
and U2001 (N_2001,In_1671,In_1584);
or U2002 (N_2002,In_871,In_1333);
and U2003 (N_2003,In_1359,In_1425);
and U2004 (N_2004,In_407,In_401);
and U2005 (N_2005,In_1001,In_861);
nor U2006 (N_2006,In_547,In_1009);
or U2007 (N_2007,In_289,In_1164);
xor U2008 (N_2008,In_855,In_1237);
nand U2009 (N_2009,In_211,In_737);
and U2010 (N_2010,In_1222,In_727);
or U2011 (N_2011,In_471,In_1045);
nand U2012 (N_2012,In_1955,In_410);
nand U2013 (N_2013,In_685,In_1271);
and U2014 (N_2014,In_1583,In_529);
xnor U2015 (N_2015,In_1602,In_1600);
nor U2016 (N_2016,In_392,In_4);
nand U2017 (N_2017,In_62,In_412);
nor U2018 (N_2018,In_1149,In_59);
xor U2019 (N_2019,In_804,In_201);
xnor U2020 (N_2020,In_30,In_1596);
or U2021 (N_2021,In_1387,In_1542);
and U2022 (N_2022,In_43,In_932);
nand U2023 (N_2023,In_1674,In_44);
and U2024 (N_2024,In_1736,In_654);
nor U2025 (N_2025,In_1570,In_316);
nor U2026 (N_2026,In_244,In_1005);
nor U2027 (N_2027,In_1543,In_1331);
nand U2028 (N_2028,In_1897,In_121);
and U2029 (N_2029,In_862,In_186);
nand U2030 (N_2030,In_566,In_1824);
nand U2031 (N_2031,In_476,In_407);
and U2032 (N_2032,In_1355,In_1882);
nand U2033 (N_2033,In_1217,In_118);
or U2034 (N_2034,In_1404,In_881);
nor U2035 (N_2035,In_436,In_549);
and U2036 (N_2036,In_1569,In_1305);
or U2037 (N_2037,In_830,In_1943);
nor U2038 (N_2038,In_872,In_1496);
or U2039 (N_2039,In_339,In_1932);
and U2040 (N_2040,In_851,In_1220);
nand U2041 (N_2041,In_823,In_1389);
and U2042 (N_2042,In_1217,In_544);
and U2043 (N_2043,In_1089,In_869);
nand U2044 (N_2044,In_823,In_1558);
or U2045 (N_2045,In_1667,In_1983);
or U2046 (N_2046,In_1095,In_130);
nor U2047 (N_2047,In_1752,In_1242);
nand U2048 (N_2048,In_1466,In_106);
nand U2049 (N_2049,In_713,In_1118);
and U2050 (N_2050,In_413,In_1966);
nor U2051 (N_2051,In_145,In_1937);
nor U2052 (N_2052,In_1982,In_1524);
and U2053 (N_2053,In_97,In_1812);
xnor U2054 (N_2054,In_877,In_1028);
or U2055 (N_2055,In_1853,In_803);
nand U2056 (N_2056,In_1405,In_1072);
and U2057 (N_2057,In_354,In_1271);
and U2058 (N_2058,In_1118,In_977);
nor U2059 (N_2059,In_1548,In_1174);
or U2060 (N_2060,In_1260,In_306);
and U2061 (N_2061,In_877,In_752);
or U2062 (N_2062,In_1294,In_390);
nor U2063 (N_2063,In_785,In_1119);
or U2064 (N_2064,In_1831,In_899);
or U2065 (N_2065,In_309,In_1983);
and U2066 (N_2066,In_1409,In_615);
and U2067 (N_2067,In_1074,In_1393);
nand U2068 (N_2068,In_1934,In_1824);
or U2069 (N_2069,In_1844,In_31);
nand U2070 (N_2070,In_820,In_1969);
nand U2071 (N_2071,In_684,In_105);
xnor U2072 (N_2072,In_1611,In_414);
nor U2073 (N_2073,In_656,In_1646);
nor U2074 (N_2074,In_628,In_181);
nor U2075 (N_2075,In_893,In_1220);
and U2076 (N_2076,In_112,In_337);
nand U2077 (N_2077,In_1026,In_421);
nand U2078 (N_2078,In_1715,In_817);
nor U2079 (N_2079,In_604,In_1376);
nor U2080 (N_2080,In_95,In_1247);
nand U2081 (N_2081,In_996,In_262);
nor U2082 (N_2082,In_797,In_1067);
and U2083 (N_2083,In_26,In_807);
nand U2084 (N_2084,In_1056,In_311);
and U2085 (N_2085,In_1361,In_1273);
nor U2086 (N_2086,In_1532,In_682);
nor U2087 (N_2087,In_213,In_1450);
or U2088 (N_2088,In_1773,In_1358);
nand U2089 (N_2089,In_705,In_377);
nand U2090 (N_2090,In_1422,In_558);
xor U2091 (N_2091,In_195,In_41);
nor U2092 (N_2092,In_1921,In_1402);
nor U2093 (N_2093,In_722,In_1526);
or U2094 (N_2094,In_1260,In_1795);
or U2095 (N_2095,In_710,In_1659);
nor U2096 (N_2096,In_6,In_633);
nor U2097 (N_2097,In_1828,In_1016);
nand U2098 (N_2098,In_1057,In_40);
xor U2099 (N_2099,In_690,In_1204);
or U2100 (N_2100,In_1320,In_558);
nor U2101 (N_2101,In_1148,In_1193);
xnor U2102 (N_2102,In_499,In_83);
nand U2103 (N_2103,In_848,In_895);
or U2104 (N_2104,In_123,In_34);
and U2105 (N_2105,In_648,In_1141);
nand U2106 (N_2106,In_1136,In_1041);
or U2107 (N_2107,In_1756,In_369);
and U2108 (N_2108,In_1781,In_1768);
xor U2109 (N_2109,In_1566,In_1556);
or U2110 (N_2110,In_43,In_520);
or U2111 (N_2111,In_991,In_1635);
nor U2112 (N_2112,In_926,In_1877);
nor U2113 (N_2113,In_1242,In_872);
nand U2114 (N_2114,In_858,In_1135);
or U2115 (N_2115,In_1650,In_1170);
nand U2116 (N_2116,In_296,In_1485);
nand U2117 (N_2117,In_510,In_148);
and U2118 (N_2118,In_369,In_1708);
nand U2119 (N_2119,In_283,In_849);
or U2120 (N_2120,In_1282,In_1188);
and U2121 (N_2121,In_1819,In_612);
or U2122 (N_2122,In_243,In_307);
nor U2123 (N_2123,In_1955,In_1041);
or U2124 (N_2124,In_207,In_552);
or U2125 (N_2125,In_237,In_449);
nand U2126 (N_2126,In_222,In_131);
nor U2127 (N_2127,In_782,In_1341);
nor U2128 (N_2128,In_1068,In_1227);
nor U2129 (N_2129,In_1894,In_446);
or U2130 (N_2130,In_1129,In_1310);
and U2131 (N_2131,In_740,In_165);
or U2132 (N_2132,In_50,In_1986);
and U2133 (N_2133,In_821,In_1089);
and U2134 (N_2134,In_968,In_289);
and U2135 (N_2135,In_830,In_681);
nand U2136 (N_2136,In_1185,In_1259);
xor U2137 (N_2137,In_1865,In_112);
or U2138 (N_2138,In_590,In_529);
and U2139 (N_2139,In_1384,In_640);
or U2140 (N_2140,In_831,In_1853);
nor U2141 (N_2141,In_1932,In_651);
xnor U2142 (N_2142,In_424,In_246);
nor U2143 (N_2143,In_1331,In_528);
and U2144 (N_2144,In_779,In_955);
and U2145 (N_2145,In_136,In_1003);
and U2146 (N_2146,In_53,In_185);
or U2147 (N_2147,In_1899,In_951);
and U2148 (N_2148,In_1428,In_1364);
nand U2149 (N_2149,In_160,In_1199);
and U2150 (N_2150,In_1107,In_1646);
xnor U2151 (N_2151,In_1712,In_685);
or U2152 (N_2152,In_1849,In_1048);
or U2153 (N_2153,In_858,In_1142);
nand U2154 (N_2154,In_1036,In_503);
nand U2155 (N_2155,In_1138,In_1966);
and U2156 (N_2156,In_1137,In_191);
and U2157 (N_2157,In_37,In_1222);
and U2158 (N_2158,In_1102,In_678);
xor U2159 (N_2159,In_1681,In_1930);
or U2160 (N_2160,In_1433,In_1998);
nor U2161 (N_2161,In_195,In_1463);
and U2162 (N_2162,In_1541,In_436);
and U2163 (N_2163,In_1789,In_1077);
or U2164 (N_2164,In_1341,In_1228);
nand U2165 (N_2165,In_105,In_1670);
xor U2166 (N_2166,In_863,In_1839);
or U2167 (N_2167,In_1952,In_1160);
nor U2168 (N_2168,In_968,In_297);
nand U2169 (N_2169,In_1194,In_1950);
xnor U2170 (N_2170,In_968,In_960);
nand U2171 (N_2171,In_687,In_1260);
xor U2172 (N_2172,In_1116,In_1081);
xor U2173 (N_2173,In_127,In_87);
and U2174 (N_2174,In_1732,In_1336);
and U2175 (N_2175,In_1772,In_1133);
and U2176 (N_2176,In_1014,In_454);
and U2177 (N_2177,In_549,In_1437);
and U2178 (N_2178,In_474,In_36);
nand U2179 (N_2179,In_1756,In_813);
nand U2180 (N_2180,In_81,In_1073);
or U2181 (N_2181,In_1995,In_1515);
or U2182 (N_2182,In_701,In_1172);
xnor U2183 (N_2183,In_624,In_126);
xnor U2184 (N_2184,In_1937,In_713);
nor U2185 (N_2185,In_1983,In_327);
xnor U2186 (N_2186,In_487,In_834);
or U2187 (N_2187,In_341,In_1095);
or U2188 (N_2188,In_489,In_576);
nand U2189 (N_2189,In_1927,In_1598);
nor U2190 (N_2190,In_1282,In_605);
and U2191 (N_2191,In_191,In_1620);
and U2192 (N_2192,In_1896,In_1034);
nand U2193 (N_2193,In_946,In_624);
and U2194 (N_2194,In_1885,In_399);
nand U2195 (N_2195,In_1442,In_1815);
or U2196 (N_2196,In_1225,In_1722);
and U2197 (N_2197,In_1948,In_257);
nor U2198 (N_2198,In_1018,In_427);
and U2199 (N_2199,In_263,In_292);
nor U2200 (N_2200,In_272,In_612);
or U2201 (N_2201,In_1593,In_716);
and U2202 (N_2202,In_994,In_1733);
and U2203 (N_2203,In_1322,In_1768);
nor U2204 (N_2204,In_229,In_1719);
xnor U2205 (N_2205,In_1515,In_731);
or U2206 (N_2206,In_325,In_1350);
xor U2207 (N_2207,In_315,In_1794);
and U2208 (N_2208,In_1036,In_1271);
or U2209 (N_2209,In_647,In_1792);
nand U2210 (N_2210,In_1676,In_1779);
and U2211 (N_2211,In_467,In_983);
xnor U2212 (N_2212,In_1791,In_1130);
nand U2213 (N_2213,In_188,In_1517);
and U2214 (N_2214,In_388,In_1778);
and U2215 (N_2215,In_192,In_1210);
xor U2216 (N_2216,In_1586,In_133);
and U2217 (N_2217,In_73,In_1158);
and U2218 (N_2218,In_1457,In_1159);
nor U2219 (N_2219,In_309,In_743);
xor U2220 (N_2220,In_1930,In_1885);
nand U2221 (N_2221,In_1712,In_1120);
xor U2222 (N_2222,In_1306,In_1895);
and U2223 (N_2223,In_1045,In_1248);
nand U2224 (N_2224,In_1483,In_90);
nand U2225 (N_2225,In_1012,In_1812);
xnor U2226 (N_2226,In_56,In_1873);
and U2227 (N_2227,In_670,In_806);
nand U2228 (N_2228,In_90,In_1760);
nor U2229 (N_2229,In_1252,In_680);
nand U2230 (N_2230,In_573,In_1559);
or U2231 (N_2231,In_1359,In_1490);
nand U2232 (N_2232,In_25,In_1988);
nor U2233 (N_2233,In_1122,In_375);
and U2234 (N_2234,In_883,In_1415);
nand U2235 (N_2235,In_1533,In_1402);
nand U2236 (N_2236,In_10,In_1036);
or U2237 (N_2237,In_941,In_1635);
nor U2238 (N_2238,In_1856,In_1138);
nand U2239 (N_2239,In_1833,In_1843);
nor U2240 (N_2240,In_535,In_733);
nor U2241 (N_2241,In_1197,In_795);
nand U2242 (N_2242,In_1093,In_1486);
nand U2243 (N_2243,In_1866,In_496);
nor U2244 (N_2244,In_868,In_437);
nand U2245 (N_2245,In_181,In_1868);
nand U2246 (N_2246,In_606,In_1793);
or U2247 (N_2247,In_683,In_13);
nor U2248 (N_2248,In_1315,In_714);
nor U2249 (N_2249,In_707,In_1713);
nand U2250 (N_2250,In_1847,In_1708);
nand U2251 (N_2251,In_371,In_1211);
xor U2252 (N_2252,In_562,In_1756);
nand U2253 (N_2253,In_686,In_1340);
nand U2254 (N_2254,In_1062,In_1691);
nor U2255 (N_2255,In_1711,In_1663);
and U2256 (N_2256,In_1291,In_792);
nand U2257 (N_2257,In_1231,In_879);
nand U2258 (N_2258,In_1446,In_1436);
or U2259 (N_2259,In_289,In_152);
nor U2260 (N_2260,In_1949,In_779);
and U2261 (N_2261,In_639,In_389);
or U2262 (N_2262,In_330,In_1924);
nor U2263 (N_2263,In_980,In_1139);
and U2264 (N_2264,In_1342,In_1014);
nand U2265 (N_2265,In_1784,In_610);
nand U2266 (N_2266,In_219,In_178);
nor U2267 (N_2267,In_1984,In_542);
and U2268 (N_2268,In_266,In_460);
and U2269 (N_2269,In_540,In_115);
nand U2270 (N_2270,In_289,In_627);
nand U2271 (N_2271,In_1468,In_1801);
nand U2272 (N_2272,In_1220,In_426);
nor U2273 (N_2273,In_1093,In_683);
and U2274 (N_2274,In_1609,In_1197);
nand U2275 (N_2275,In_606,In_565);
nor U2276 (N_2276,In_994,In_1128);
nand U2277 (N_2277,In_146,In_420);
nor U2278 (N_2278,In_926,In_1661);
xnor U2279 (N_2279,In_1077,In_905);
nor U2280 (N_2280,In_858,In_637);
nand U2281 (N_2281,In_931,In_414);
or U2282 (N_2282,In_789,In_1145);
or U2283 (N_2283,In_164,In_422);
nor U2284 (N_2284,In_558,In_1266);
nor U2285 (N_2285,In_966,In_1246);
and U2286 (N_2286,In_1277,In_1362);
or U2287 (N_2287,In_644,In_957);
xnor U2288 (N_2288,In_214,In_1709);
nor U2289 (N_2289,In_1627,In_466);
and U2290 (N_2290,In_1079,In_1773);
and U2291 (N_2291,In_323,In_1178);
nor U2292 (N_2292,In_1534,In_1171);
nor U2293 (N_2293,In_1547,In_1251);
or U2294 (N_2294,In_466,In_1006);
nand U2295 (N_2295,In_663,In_1232);
nand U2296 (N_2296,In_1459,In_360);
or U2297 (N_2297,In_50,In_1233);
and U2298 (N_2298,In_1339,In_59);
nor U2299 (N_2299,In_172,In_491);
and U2300 (N_2300,In_674,In_1101);
nand U2301 (N_2301,In_1732,In_450);
and U2302 (N_2302,In_826,In_15);
and U2303 (N_2303,In_643,In_590);
and U2304 (N_2304,In_1296,In_699);
and U2305 (N_2305,In_363,In_1725);
or U2306 (N_2306,In_1870,In_1510);
or U2307 (N_2307,In_94,In_714);
xnor U2308 (N_2308,In_1568,In_1033);
xnor U2309 (N_2309,In_1013,In_349);
and U2310 (N_2310,In_335,In_136);
nor U2311 (N_2311,In_1514,In_1574);
nor U2312 (N_2312,In_1293,In_1160);
or U2313 (N_2313,In_34,In_324);
and U2314 (N_2314,In_502,In_1553);
nand U2315 (N_2315,In_1182,In_1150);
nand U2316 (N_2316,In_735,In_1419);
nor U2317 (N_2317,In_538,In_1716);
nor U2318 (N_2318,In_935,In_1069);
or U2319 (N_2319,In_1899,In_1686);
nor U2320 (N_2320,In_225,In_1076);
xor U2321 (N_2321,In_417,In_640);
xnor U2322 (N_2322,In_1922,In_579);
nand U2323 (N_2323,In_1972,In_864);
nor U2324 (N_2324,In_1432,In_1990);
or U2325 (N_2325,In_1553,In_265);
and U2326 (N_2326,In_463,In_309);
nand U2327 (N_2327,In_234,In_834);
nand U2328 (N_2328,In_539,In_1515);
nor U2329 (N_2329,In_1245,In_1277);
and U2330 (N_2330,In_1103,In_94);
nor U2331 (N_2331,In_1636,In_1325);
and U2332 (N_2332,In_1277,In_1168);
nor U2333 (N_2333,In_1216,In_1826);
nand U2334 (N_2334,In_50,In_284);
or U2335 (N_2335,In_425,In_847);
nor U2336 (N_2336,In_915,In_188);
nor U2337 (N_2337,In_1024,In_225);
or U2338 (N_2338,In_1215,In_986);
nand U2339 (N_2339,In_182,In_1901);
nor U2340 (N_2340,In_1262,In_238);
xor U2341 (N_2341,In_39,In_891);
and U2342 (N_2342,In_59,In_339);
or U2343 (N_2343,In_1445,In_1123);
xor U2344 (N_2344,In_269,In_815);
nor U2345 (N_2345,In_1927,In_1593);
and U2346 (N_2346,In_1123,In_1141);
or U2347 (N_2347,In_1169,In_15);
nor U2348 (N_2348,In_345,In_6);
xor U2349 (N_2349,In_664,In_92);
or U2350 (N_2350,In_1801,In_1444);
xnor U2351 (N_2351,In_85,In_848);
or U2352 (N_2352,In_1886,In_327);
nor U2353 (N_2353,In_1753,In_188);
and U2354 (N_2354,In_1176,In_1793);
or U2355 (N_2355,In_228,In_1494);
nor U2356 (N_2356,In_1662,In_251);
nor U2357 (N_2357,In_15,In_1361);
and U2358 (N_2358,In_205,In_18);
or U2359 (N_2359,In_1477,In_688);
nand U2360 (N_2360,In_1951,In_1309);
nor U2361 (N_2361,In_1737,In_1485);
xor U2362 (N_2362,In_483,In_1632);
and U2363 (N_2363,In_1282,In_427);
nand U2364 (N_2364,In_1424,In_84);
or U2365 (N_2365,In_116,In_719);
nor U2366 (N_2366,In_251,In_1420);
xor U2367 (N_2367,In_827,In_1115);
nor U2368 (N_2368,In_1601,In_993);
and U2369 (N_2369,In_833,In_1914);
or U2370 (N_2370,In_1142,In_595);
and U2371 (N_2371,In_1870,In_188);
nor U2372 (N_2372,In_447,In_1171);
and U2373 (N_2373,In_1041,In_1232);
nor U2374 (N_2374,In_1362,In_1428);
or U2375 (N_2375,In_1406,In_1313);
and U2376 (N_2376,In_1423,In_1174);
nor U2377 (N_2377,In_916,In_630);
or U2378 (N_2378,In_680,In_628);
and U2379 (N_2379,In_91,In_522);
nand U2380 (N_2380,In_534,In_497);
xnor U2381 (N_2381,In_1015,In_1320);
and U2382 (N_2382,In_731,In_908);
and U2383 (N_2383,In_1149,In_1874);
and U2384 (N_2384,In_1847,In_1945);
or U2385 (N_2385,In_1432,In_790);
xor U2386 (N_2386,In_597,In_1159);
nand U2387 (N_2387,In_1706,In_1103);
nand U2388 (N_2388,In_1943,In_139);
or U2389 (N_2389,In_1636,In_1104);
or U2390 (N_2390,In_670,In_1822);
nand U2391 (N_2391,In_1310,In_421);
nor U2392 (N_2392,In_1880,In_445);
and U2393 (N_2393,In_937,In_1060);
or U2394 (N_2394,In_1864,In_13);
xnor U2395 (N_2395,In_1067,In_235);
nand U2396 (N_2396,In_1871,In_240);
nand U2397 (N_2397,In_999,In_1251);
and U2398 (N_2398,In_1602,In_300);
xnor U2399 (N_2399,In_901,In_1831);
nand U2400 (N_2400,In_1708,In_602);
nand U2401 (N_2401,In_530,In_1760);
and U2402 (N_2402,In_1605,In_344);
xnor U2403 (N_2403,In_1671,In_51);
and U2404 (N_2404,In_591,In_1222);
and U2405 (N_2405,In_310,In_329);
and U2406 (N_2406,In_1108,In_275);
or U2407 (N_2407,In_1670,In_911);
nor U2408 (N_2408,In_1441,In_1772);
nor U2409 (N_2409,In_1597,In_1347);
xnor U2410 (N_2410,In_625,In_226);
and U2411 (N_2411,In_48,In_1127);
or U2412 (N_2412,In_118,In_416);
nand U2413 (N_2413,In_1522,In_439);
or U2414 (N_2414,In_1096,In_1549);
and U2415 (N_2415,In_1016,In_1313);
xnor U2416 (N_2416,In_1129,In_1400);
and U2417 (N_2417,In_1330,In_1446);
and U2418 (N_2418,In_333,In_1583);
and U2419 (N_2419,In_1891,In_885);
nor U2420 (N_2420,In_307,In_1551);
xnor U2421 (N_2421,In_286,In_514);
nand U2422 (N_2422,In_214,In_1030);
nor U2423 (N_2423,In_348,In_90);
nand U2424 (N_2424,In_1445,In_1742);
and U2425 (N_2425,In_1015,In_31);
or U2426 (N_2426,In_840,In_48);
and U2427 (N_2427,In_1561,In_1253);
and U2428 (N_2428,In_111,In_275);
and U2429 (N_2429,In_1709,In_523);
nand U2430 (N_2430,In_261,In_182);
or U2431 (N_2431,In_1947,In_1745);
nand U2432 (N_2432,In_643,In_855);
nor U2433 (N_2433,In_1997,In_654);
or U2434 (N_2434,In_590,In_162);
and U2435 (N_2435,In_1133,In_17);
xor U2436 (N_2436,In_611,In_1510);
and U2437 (N_2437,In_1908,In_1148);
nor U2438 (N_2438,In_1308,In_1187);
nand U2439 (N_2439,In_1816,In_1397);
nand U2440 (N_2440,In_176,In_14);
and U2441 (N_2441,In_431,In_179);
xor U2442 (N_2442,In_650,In_730);
and U2443 (N_2443,In_90,In_1472);
and U2444 (N_2444,In_1126,In_634);
or U2445 (N_2445,In_680,In_1301);
nand U2446 (N_2446,In_424,In_1768);
and U2447 (N_2447,In_1654,In_1140);
and U2448 (N_2448,In_1075,In_352);
nand U2449 (N_2449,In_1056,In_20);
or U2450 (N_2450,In_307,In_856);
nand U2451 (N_2451,In_1095,In_1293);
or U2452 (N_2452,In_363,In_1169);
nor U2453 (N_2453,In_1550,In_1708);
nand U2454 (N_2454,In_665,In_150);
and U2455 (N_2455,In_865,In_1096);
xnor U2456 (N_2456,In_1336,In_176);
nand U2457 (N_2457,In_884,In_1574);
or U2458 (N_2458,In_338,In_1455);
or U2459 (N_2459,In_1845,In_1398);
nand U2460 (N_2460,In_344,In_1294);
or U2461 (N_2461,In_945,In_988);
or U2462 (N_2462,In_1107,In_1506);
nor U2463 (N_2463,In_1918,In_777);
nand U2464 (N_2464,In_141,In_46);
nand U2465 (N_2465,In_1309,In_1407);
or U2466 (N_2466,In_1758,In_237);
nand U2467 (N_2467,In_1682,In_38);
or U2468 (N_2468,In_1063,In_1816);
or U2469 (N_2469,In_606,In_1493);
nor U2470 (N_2470,In_1259,In_586);
nor U2471 (N_2471,In_1081,In_471);
xor U2472 (N_2472,In_135,In_658);
nand U2473 (N_2473,In_60,In_1666);
and U2474 (N_2474,In_1769,In_1657);
or U2475 (N_2475,In_1502,In_1819);
xor U2476 (N_2476,In_1698,In_805);
nor U2477 (N_2477,In_228,In_1269);
and U2478 (N_2478,In_439,In_250);
xnor U2479 (N_2479,In_910,In_253);
nor U2480 (N_2480,In_167,In_731);
and U2481 (N_2481,In_1836,In_233);
and U2482 (N_2482,In_170,In_371);
nor U2483 (N_2483,In_365,In_1522);
and U2484 (N_2484,In_1857,In_444);
or U2485 (N_2485,In_146,In_1334);
and U2486 (N_2486,In_1968,In_361);
nand U2487 (N_2487,In_1336,In_260);
nor U2488 (N_2488,In_1861,In_1541);
nand U2489 (N_2489,In_183,In_984);
nand U2490 (N_2490,In_1290,In_713);
nand U2491 (N_2491,In_1861,In_647);
xnor U2492 (N_2492,In_1735,In_1225);
nor U2493 (N_2493,In_1607,In_1061);
nor U2494 (N_2494,In_1988,In_896);
and U2495 (N_2495,In_1052,In_84);
nor U2496 (N_2496,In_514,In_1802);
and U2497 (N_2497,In_276,In_1903);
and U2498 (N_2498,In_956,In_1416);
nand U2499 (N_2499,In_1947,In_866);
nand U2500 (N_2500,In_56,In_1487);
xor U2501 (N_2501,In_338,In_141);
and U2502 (N_2502,In_1814,In_568);
and U2503 (N_2503,In_1375,In_620);
nor U2504 (N_2504,In_1744,In_1060);
and U2505 (N_2505,In_742,In_1546);
and U2506 (N_2506,In_795,In_1986);
nor U2507 (N_2507,In_1804,In_1765);
or U2508 (N_2508,In_1426,In_1784);
nor U2509 (N_2509,In_1048,In_1333);
nand U2510 (N_2510,In_1308,In_1401);
nand U2511 (N_2511,In_1309,In_1719);
xnor U2512 (N_2512,In_1768,In_1063);
or U2513 (N_2513,In_1829,In_1120);
xor U2514 (N_2514,In_756,In_1651);
and U2515 (N_2515,In_235,In_310);
nand U2516 (N_2516,In_419,In_244);
nor U2517 (N_2517,In_567,In_293);
and U2518 (N_2518,In_816,In_479);
nand U2519 (N_2519,In_267,In_690);
or U2520 (N_2520,In_1843,In_1304);
and U2521 (N_2521,In_1810,In_389);
or U2522 (N_2522,In_963,In_484);
nor U2523 (N_2523,In_1472,In_417);
nand U2524 (N_2524,In_628,In_1661);
nor U2525 (N_2525,In_1481,In_1840);
nor U2526 (N_2526,In_262,In_886);
and U2527 (N_2527,In_656,In_1230);
nor U2528 (N_2528,In_560,In_1763);
or U2529 (N_2529,In_1302,In_1536);
xnor U2530 (N_2530,In_1431,In_461);
nor U2531 (N_2531,In_1167,In_1847);
nand U2532 (N_2532,In_1355,In_919);
and U2533 (N_2533,In_155,In_344);
nor U2534 (N_2534,In_1953,In_754);
or U2535 (N_2535,In_503,In_744);
nand U2536 (N_2536,In_806,In_1025);
or U2537 (N_2537,In_1901,In_451);
or U2538 (N_2538,In_20,In_1376);
nor U2539 (N_2539,In_1678,In_999);
and U2540 (N_2540,In_274,In_1783);
and U2541 (N_2541,In_193,In_1957);
nor U2542 (N_2542,In_1808,In_689);
and U2543 (N_2543,In_175,In_291);
or U2544 (N_2544,In_1877,In_544);
and U2545 (N_2545,In_1675,In_1858);
xor U2546 (N_2546,In_939,In_731);
or U2547 (N_2547,In_1752,In_272);
nand U2548 (N_2548,In_445,In_955);
nor U2549 (N_2549,In_739,In_307);
and U2550 (N_2550,In_861,In_980);
or U2551 (N_2551,In_217,In_445);
nor U2552 (N_2552,In_1428,In_1439);
and U2553 (N_2553,In_1963,In_1476);
nand U2554 (N_2554,In_1803,In_225);
nand U2555 (N_2555,In_92,In_814);
and U2556 (N_2556,In_922,In_1795);
and U2557 (N_2557,In_4,In_1656);
nor U2558 (N_2558,In_277,In_157);
or U2559 (N_2559,In_993,In_1679);
or U2560 (N_2560,In_1919,In_1753);
xnor U2561 (N_2561,In_877,In_910);
nand U2562 (N_2562,In_1913,In_704);
nor U2563 (N_2563,In_1459,In_1679);
or U2564 (N_2564,In_1777,In_1830);
nor U2565 (N_2565,In_749,In_1660);
or U2566 (N_2566,In_853,In_235);
nand U2567 (N_2567,In_1354,In_207);
or U2568 (N_2568,In_67,In_1627);
or U2569 (N_2569,In_1535,In_1547);
or U2570 (N_2570,In_279,In_1934);
and U2571 (N_2571,In_1016,In_950);
or U2572 (N_2572,In_722,In_1954);
or U2573 (N_2573,In_1477,In_1969);
xnor U2574 (N_2574,In_1912,In_562);
nor U2575 (N_2575,In_1286,In_1252);
nor U2576 (N_2576,In_1561,In_283);
or U2577 (N_2577,In_940,In_1149);
nand U2578 (N_2578,In_1873,In_847);
nor U2579 (N_2579,In_1769,In_1976);
or U2580 (N_2580,In_1348,In_1598);
or U2581 (N_2581,In_114,In_538);
nor U2582 (N_2582,In_1933,In_291);
nor U2583 (N_2583,In_1829,In_1591);
nor U2584 (N_2584,In_1882,In_499);
or U2585 (N_2585,In_1238,In_483);
or U2586 (N_2586,In_1550,In_1062);
or U2587 (N_2587,In_1475,In_79);
nand U2588 (N_2588,In_381,In_1927);
nor U2589 (N_2589,In_591,In_1042);
nor U2590 (N_2590,In_1905,In_1410);
xor U2591 (N_2591,In_1596,In_1435);
and U2592 (N_2592,In_480,In_397);
or U2593 (N_2593,In_1620,In_718);
nor U2594 (N_2594,In_1614,In_1386);
nand U2595 (N_2595,In_149,In_836);
nand U2596 (N_2596,In_929,In_34);
xnor U2597 (N_2597,In_723,In_1905);
and U2598 (N_2598,In_251,In_372);
xnor U2599 (N_2599,In_1541,In_579);
xor U2600 (N_2600,In_907,In_1824);
or U2601 (N_2601,In_177,In_209);
or U2602 (N_2602,In_1350,In_728);
xor U2603 (N_2603,In_152,In_890);
xor U2604 (N_2604,In_343,In_67);
nor U2605 (N_2605,In_1583,In_369);
nor U2606 (N_2606,In_489,In_328);
and U2607 (N_2607,In_547,In_549);
and U2608 (N_2608,In_728,In_1284);
nand U2609 (N_2609,In_1594,In_848);
nor U2610 (N_2610,In_520,In_1039);
nand U2611 (N_2611,In_408,In_1285);
nand U2612 (N_2612,In_1634,In_1262);
nor U2613 (N_2613,In_1896,In_1436);
nor U2614 (N_2614,In_674,In_342);
nand U2615 (N_2615,In_237,In_240);
and U2616 (N_2616,In_826,In_1451);
and U2617 (N_2617,In_1582,In_1460);
and U2618 (N_2618,In_780,In_898);
nand U2619 (N_2619,In_735,In_836);
nor U2620 (N_2620,In_1088,In_702);
and U2621 (N_2621,In_1645,In_1758);
or U2622 (N_2622,In_533,In_343);
nand U2623 (N_2623,In_1419,In_1279);
xnor U2624 (N_2624,In_1741,In_28);
nor U2625 (N_2625,In_592,In_1303);
nor U2626 (N_2626,In_1123,In_245);
nor U2627 (N_2627,In_1029,In_1924);
or U2628 (N_2628,In_1710,In_81);
nand U2629 (N_2629,In_956,In_1233);
and U2630 (N_2630,In_1234,In_665);
and U2631 (N_2631,In_135,In_1322);
or U2632 (N_2632,In_1788,In_1132);
or U2633 (N_2633,In_1317,In_63);
nor U2634 (N_2634,In_688,In_787);
nor U2635 (N_2635,In_24,In_1844);
nand U2636 (N_2636,In_798,In_1379);
or U2637 (N_2637,In_1617,In_1925);
nor U2638 (N_2638,In_340,In_1200);
or U2639 (N_2639,In_1312,In_909);
or U2640 (N_2640,In_1680,In_1913);
or U2641 (N_2641,In_1368,In_911);
or U2642 (N_2642,In_1468,In_301);
or U2643 (N_2643,In_136,In_423);
nand U2644 (N_2644,In_1312,In_1305);
nand U2645 (N_2645,In_725,In_435);
or U2646 (N_2646,In_778,In_883);
and U2647 (N_2647,In_366,In_1558);
nand U2648 (N_2648,In_1160,In_612);
or U2649 (N_2649,In_957,In_1881);
nor U2650 (N_2650,In_1304,In_345);
nand U2651 (N_2651,In_571,In_1718);
or U2652 (N_2652,In_1849,In_847);
nor U2653 (N_2653,In_1780,In_1776);
nand U2654 (N_2654,In_1657,In_1876);
nor U2655 (N_2655,In_829,In_1922);
nand U2656 (N_2656,In_1088,In_1975);
nand U2657 (N_2657,In_688,In_1499);
nand U2658 (N_2658,In_990,In_648);
or U2659 (N_2659,In_1610,In_149);
xnor U2660 (N_2660,In_262,In_1179);
nand U2661 (N_2661,In_297,In_1442);
xor U2662 (N_2662,In_1141,In_854);
nand U2663 (N_2663,In_1642,In_517);
nor U2664 (N_2664,In_152,In_892);
xor U2665 (N_2665,In_229,In_704);
nand U2666 (N_2666,In_1626,In_1112);
and U2667 (N_2667,In_1442,In_1354);
nand U2668 (N_2668,In_1212,In_1768);
and U2669 (N_2669,In_445,In_210);
nand U2670 (N_2670,In_730,In_1404);
or U2671 (N_2671,In_1933,In_1598);
nor U2672 (N_2672,In_1193,In_914);
nand U2673 (N_2673,In_679,In_1051);
nor U2674 (N_2674,In_1950,In_1784);
or U2675 (N_2675,In_43,In_1494);
xnor U2676 (N_2676,In_137,In_279);
nand U2677 (N_2677,In_379,In_393);
and U2678 (N_2678,In_221,In_922);
nor U2679 (N_2679,In_1323,In_1447);
xor U2680 (N_2680,In_1942,In_377);
and U2681 (N_2681,In_1139,In_416);
nor U2682 (N_2682,In_1290,In_1628);
xor U2683 (N_2683,In_1503,In_1586);
or U2684 (N_2684,In_747,In_1245);
nand U2685 (N_2685,In_458,In_1604);
nor U2686 (N_2686,In_708,In_1462);
or U2687 (N_2687,In_722,In_734);
and U2688 (N_2688,In_1412,In_706);
xor U2689 (N_2689,In_814,In_789);
or U2690 (N_2690,In_693,In_209);
nand U2691 (N_2691,In_311,In_1300);
nor U2692 (N_2692,In_848,In_939);
or U2693 (N_2693,In_1632,In_905);
nor U2694 (N_2694,In_861,In_302);
nor U2695 (N_2695,In_299,In_348);
or U2696 (N_2696,In_1054,In_61);
or U2697 (N_2697,In_1176,In_1186);
nand U2698 (N_2698,In_721,In_1672);
and U2699 (N_2699,In_1169,In_1192);
and U2700 (N_2700,In_1503,In_321);
and U2701 (N_2701,In_181,In_1044);
or U2702 (N_2702,In_1218,In_23);
or U2703 (N_2703,In_1733,In_50);
nor U2704 (N_2704,In_716,In_539);
nor U2705 (N_2705,In_314,In_957);
or U2706 (N_2706,In_1436,In_471);
xnor U2707 (N_2707,In_767,In_1099);
nand U2708 (N_2708,In_775,In_1244);
and U2709 (N_2709,In_601,In_961);
nor U2710 (N_2710,In_756,In_1471);
and U2711 (N_2711,In_1573,In_273);
or U2712 (N_2712,In_31,In_894);
nor U2713 (N_2713,In_1407,In_129);
nand U2714 (N_2714,In_1768,In_1783);
nand U2715 (N_2715,In_1184,In_561);
or U2716 (N_2716,In_599,In_1103);
xor U2717 (N_2717,In_1533,In_848);
or U2718 (N_2718,In_781,In_966);
nand U2719 (N_2719,In_790,In_1020);
or U2720 (N_2720,In_1082,In_576);
nand U2721 (N_2721,In_512,In_1854);
or U2722 (N_2722,In_34,In_483);
and U2723 (N_2723,In_830,In_421);
or U2724 (N_2724,In_1822,In_870);
nor U2725 (N_2725,In_1018,In_485);
nand U2726 (N_2726,In_553,In_278);
or U2727 (N_2727,In_654,In_1262);
xnor U2728 (N_2728,In_172,In_398);
or U2729 (N_2729,In_1544,In_630);
and U2730 (N_2730,In_461,In_1416);
xor U2731 (N_2731,In_1605,In_1917);
nor U2732 (N_2732,In_552,In_1799);
or U2733 (N_2733,In_1277,In_891);
or U2734 (N_2734,In_1685,In_1912);
and U2735 (N_2735,In_589,In_802);
or U2736 (N_2736,In_289,In_418);
nand U2737 (N_2737,In_657,In_1474);
nand U2738 (N_2738,In_354,In_504);
nor U2739 (N_2739,In_1124,In_65);
nand U2740 (N_2740,In_307,In_816);
and U2741 (N_2741,In_5,In_51);
or U2742 (N_2742,In_1963,In_1236);
and U2743 (N_2743,In_387,In_404);
or U2744 (N_2744,In_1065,In_1644);
or U2745 (N_2745,In_1306,In_1845);
or U2746 (N_2746,In_1667,In_664);
or U2747 (N_2747,In_1180,In_1908);
or U2748 (N_2748,In_476,In_140);
nor U2749 (N_2749,In_677,In_1056);
nor U2750 (N_2750,In_1261,In_1361);
nand U2751 (N_2751,In_1854,In_150);
or U2752 (N_2752,In_1701,In_1869);
nand U2753 (N_2753,In_1041,In_1873);
nand U2754 (N_2754,In_774,In_1637);
nand U2755 (N_2755,In_994,In_1039);
nor U2756 (N_2756,In_1333,In_368);
nand U2757 (N_2757,In_1191,In_270);
or U2758 (N_2758,In_396,In_1348);
nor U2759 (N_2759,In_1160,In_246);
nor U2760 (N_2760,In_1917,In_275);
or U2761 (N_2761,In_465,In_345);
nor U2762 (N_2762,In_1339,In_497);
nand U2763 (N_2763,In_226,In_1845);
nor U2764 (N_2764,In_1769,In_128);
and U2765 (N_2765,In_1786,In_1398);
nor U2766 (N_2766,In_1222,In_1869);
xnor U2767 (N_2767,In_234,In_712);
xnor U2768 (N_2768,In_977,In_1148);
or U2769 (N_2769,In_1682,In_54);
nand U2770 (N_2770,In_1160,In_1228);
nor U2771 (N_2771,In_1620,In_1907);
nor U2772 (N_2772,In_139,In_892);
nor U2773 (N_2773,In_922,In_316);
xnor U2774 (N_2774,In_298,In_987);
nand U2775 (N_2775,In_1450,In_549);
and U2776 (N_2776,In_1562,In_1211);
xor U2777 (N_2777,In_69,In_1946);
nand U2778 (N_2778,In_1,In_712);
or U2779 (N_2779,In_1188,In_1458);
nand U2780 (N_2780,In_874,In_409);
nor U2781 (N_2781,In_486,In_1567);
and U2782 (N_2782,In_92,In_1745);
and U2783 (N_2783,In_25,In_214);
nor U2784 (N_2784,In_1888,In_1466);
nand U2785 (N_2785,In_140,In_901);
nand U2786 (N_2786,In_1941,In_556);
nand U2787 (N_2787,In_604,In_1911);
nor U2788 (N_2788,In_194,In_315);
nand U2789 (N_2789,In_868,In_1825);
xnor U2790 (N_2790,In_178,In_1408);
xor U2791 (N_2791,In_1676,In_506);
xnor U2792 (N_2792,In_225,In_422);
xor U2793 (N_2793,In_874,In_1544);
and U2794 (N_2794,In_718,In_1730);
nor U2795 (N_2795,In_1645,In_1851);
xor U2796 (N_2796,In_156,In_776);
or U2797 (N_2797,In_710,In_1333);
or U2798 (N_2798,In_1898,In_1900);
or U2799 (N_2799,In_1456,In_567);
and U2800 (N_2800,In_1870,In_252);
and U2801 (N_2801,In_1659,In_143);
nand U2802 (N_2802,In_667,In_761);
nor U2803 (N_2803,In_865,In_1355);
nand U2804 (N_2804,In_1192,In_1929);
nor U2805 (N_2805,In_1967,In_1921);
and U2806 (N_2806,In_1179,In_202);
or U2807 (N_2807,In_125,In_341);
or U2808 (N_2808,In_967,In_1173);
nand U2809 (N_2809,In_1513,In_1148);
nand U2810 (N_2810,In_1621,In_446);
nand U2811 (N_2811,In_1244,In_1421);
or U2812 (N_2812,In_908,In_207);
or U2813 (N_2813,In_792,In_46);
nand U2814 (N_2814,In_572,In_1185);
nor U2815 (N_2815,In_600,In_566);
nor U2816 (N_2816,In_815,In_1518);
and U2817 (N_2817,In_1905,In_670);
nor U2818 (N_2818,In_1782,In_1176);
xnor U2819 (N_2819,In_1393,In_1216);
and U2820 (N_2820,In_67,In_1111);
xor U2821 (N_2821,In_1371,In_362);
xor U2822 (N_2822,In_183,In_1502);
or U2823 (N_2823,In_1577,In_1928);
nand U2824 (N_2824,In_297,In_1425);
and U2825 (N_2825,In_1393,In_1347);
nand U2826 (N_2826,In_676,In_1846);
nor U2827 (N_2827,In_1655,In_596);
nand U2828 (N_2828,In_863,In_230);
nand U2829 (N_2829,In_1228,In_1601);
nand U2830 (N_2830,In_501,In_222);
nor U2831 (N_2831,In_308,In_932);
and U2832 (N_2832,In_241,In_984);
nor U2833 (N_2833,In_1542,In_1700);
nand U2834 (N_2834,In_1901,In_1575);
nand U2835 (N_2835,In_10,In_245);
xor U2836 (N_2836,In_1365,In_722);
and U2837 (N_2837,In_71,In_499);
nor U2838 (N_2838,In_930,In_234);
nand U2839 (N_2839,In_1440,In_952);
nor U2840 (N_2840,In_613,In_1363);
or U2841 (N_2841,In_1434,In_1370);
and U2842 (N_2842,In_1998,In_1505);
nor U2843 (N_2843,In_706,In_828);
and U2844 (N_2844,In_1715,In_455);
nand U2845 (N_2845,In_1268,In_1117);
nor U2846 (N_2846,In_1862,In_446);
nor U2847 (N_2847,In_1493,In_518);
nand U2848 (N_2848,In_68,In_62);
and U2849 (N_2849,In_1580,In_1388);
nand U2850 (N_2850,In_1329,In_1984);
xnor U2851 (N_2851,In_633,In_1384);
or U2852 (N_2852,In_1532,In_581);
and U2853 (N_2853,In_1864,In_1753);
nor U2854 (N_2854,In_1005,In_1537);
and U2855 (N_2855,In_1302,In_191);
nand U2856 (N_2856,In_1913,In_1606);
or U2857 (N_2857,In_721,In_318);
nand U2858 (N_2858,In_623,In_751);
xor U2859 (N_2859,In_616,In_1070);
nor U2860 (N_2860,In_384,In_1045);
or U2861 (N_2861,In_1885,In_9);
xnor U2862 (N_2862,In_1920,In_1044);
nor U2863 (N_2863,In_892,In_1833);
or U2864 (N_2864,In_249,In_1167);
nor U2865 (N_2865,In_280,In_503);
nor U2866 (N_2866,In_1285,In_420);
nand U2867 (N_2867,In_398,In_1016);
and U2868 (N_2868,In_20,In_128);
or U2869 (N_2869,In_608,In_1213);
nand U2870 (N_2870,In_279,In_1357);
nand U2871 (N_2871,In_671,In_1769);
and U2872 (N_2872,In_1988,In_1457);
nor U2873 (N_2873,In_1579,In_1021);
and U2874 (N_2874,In_801,In_1543);
nor U2875 (N_2875,In_505,In_36);
nand U2876 (N_2876,In_1501,In_720);
and U2877 (N_2877,In_1423,In_26);
nand U2878 (N_2878,In_1459,In_491);
and U2879 (N_2879,In_1197,In_295);
xor U2880 (N_2880,In_139,In_1415);
and U2881 (N_2881,In_543,In_1152);
and U2882 (N_2882,In_467,In_1581);
and U2883 (N_2883,In_1688,In_1117);
or U2884 (N_2884,In_1668,In_377);
nand U2885 (N_2885,In_481,In_632);
nor U2886 (N_2886,In_291,In_1517);
nor U2887 (N_2887,In_1180,In_64);
or U2888 (N_2888,In_283,In_1118);
or U2889 (N_2889,In_1203,In_585);
or U2890 (N_2890,In_246,In_1262);
and U2891 (N_2891,In_227,In_1975);
nand U2892 (N_2892,In_1421,In_526);
nand U2893 (N_2893,In_109,In_1964);
and U2894 (N_2894,In_374,In_1173);
nand U2895 (N_2895,In_264,In_688);
or U2896 (N_2896,In_647,In_1199);
and U2897 (N_2897,In_87,In_644);
nand U2898 (N_2898,In_1083,In_908);
nand U2899 (N_2899,In_749,In_288);
nand U2900 (N_2900,In_1322,In_864);
and U2901 (N_2901,In_1654,In_1153);
nor U2902 (N_2902,In_1606,In_1507);
or U2903 (N_2903,In_1284,In_944);
nand U2904 (N_2904,In_134,In_1056);
nand U2905 (N_2905,In_830,In_1416);
nand U2906 (N_2906,In_1558,In_481);
nor U2907 (N_2907,In_717,In_710);
nor U2908 (N_2908,In_1290,In_556);
nand U2909 (N_2909,In_1794,In_1466);
or U2910 (N_2910,In_1422,In_579);
nor U2911 (N_2911,In_976,In_484);
or U2912 (N_2912,In_317,In_1360);
nor U2913 (N_2913,In_1552,In_952);
and U2914 (N_2914,In_817,In_894);
xor U2915 (N_2915,In_1001,In_1708);
or U2916 (N_2916,In_1748,In_886);
nand U2917 (N_2917,In_275,In_1933);
nor U2918 (N_2918,In_1572,In_1396);
or U2919 (N_2919,In_590,In_1527);
or U2920 (N_2920,In_322,In_1663);
and U2921 (N_2921,In_1925,In_89);
xor U2922 (N_2922,In_188,In_1802);
or U2923 (N_2923,In_450,In_1693);
nor U2924 (N_2924,In_1016,In_486);
and U2925 (N_2925,In_475,In_131);
nand U2926 (N_2926,In_1312,In_1888);
nor U2927 (N_2927,In_715,In_1482);
nand U2928 (N_2928,In_1026,In_1594);
and U2929 (N_2929,In_1269,In_607);
nand U2930 (N_2930,In_1552,In_1599);
or U2931 (N_2931,In_1661,In_1972);
or U2932 (N_2932,In_1227,In_1904);
and U2933 (N_2933,In_837,In_1326);
nor U2934 (N_2934,In_901,In_532);
or U2935 (N_2935,In_1084,In_1596);
or U2936 (N_2936,In_345,In_968);
nand U2937 (N_2937,In_1458,In_609);
or U2938 (N_2938,In_513,In_188);
nor U2939 (N_2939,In_1419,In_1120);
nor U2940 (N_2940,In_1288,In_1064);
or U2941 (N_2941,In_114,In_959);
nand U2942 (N_2942,In_936,In_384);
and U2943 (N_2943,In_1394,In_1730);
nand U2944 (N_2944,In_1331,In_1675);
or U2945 (N_2945,In_1690,In_945);
nor U2946 (N_2946,In_118,In_567);
or U2947 (N_2947,In_1533,In_1786);
nor U2948 (N_2948,In_72,In_1678);
or U2949 (N_2949,In_1013,In_1711);
nor U2950 (N_2950,In_1472,In_1920);
xor U2951 (N_2951,In_1020,In_1704);
or U2952 (N_2952,In_1185,In_915);
nand U2953 (N_2953,In_1850,In_1244);
nand U2954 (N_2954,In_782,In_1312);
and U2955 (N_2955,In_1077,In_644);
nor U2956 (N_2956,In_1852,In_198);
xor U2957 (N_2957,In_307,In_519);
or U2958 (N_2958,In_750,In_447);
and U2959 (N_2959,In_795,In_600);
and U2960 (N_2960,In_758,In_1731);
nor U2961 (N_2961,In_1367,In_1912);
and U2962 (N_2962,In_1251,In_924);
nand U2963 (N_2963,In_436,In_437);
or U2964 (N_2964,In_1211,In_520);
or U2965 (N_2965,In_153,In_291);
nor U2966 (N_2966,In_1844,In_1316);
nand U2967 (N_2967,In_1975,In_1582);
xor U2968 (N_2968,In_103,In_165);
xor U2969 (N_2969,In_1927,In_1054);
xnor U2970 (N_2970,In_711,In_1108);
nor U2971 (N_2971,In_1355,In_506);
nor U2972 (N_2972,In_589,In_1365);
nor U2973 (N_2973,In_284,In_339);
and U2974 (N_2974,In_167,In_1918);
or U2975 (N_2975,In_1250,In_1047);
nor U2976 (N_2976,In_1380,In_127);
or U2977 (N_2977,In_1278,In_1326);
nand U2978 (N_2978,In_900,In_1932);
nor U2979 (N_2979,In_525,In_1855);
and U2980 (N_2980,In_518,In_1917);
nor U2981 (N_2981,In_1461,In_1153);
and U2982 (N_2982,In_1069,In_493);
nand U2983 (N_2983,In_1112,In_1064);
and U2984 (N_2984,In_1991,In_688);
nand U2985 (N_2985,In_1339,In_1080);
and U2986 (N_2986,In_10,In_1218);
and U2987 (N_2987,In_1729,In_1244);
and U2988 (N_2988,In_1009,In_650);
nand U2989 (N_2989,In_730,In_603);
and U2990 (N_2990,In_1376,In_1442);
nand U2991 (N_2991,In_1416,In_1705);
or U2992 (N_2992,In_1346,In_395);
nor U2993 (N_2993,In_895,In_105);
nor U2994 (N_2994,In_1523,In_323);
nand U2995 (N_2995,In_1302,In_1303);
nor U2996 (N_2996,In_1749,In_673);
and U2997 (N_2997,In_1320,In_828);
nor U2998 (N_2998,In_1176,In_1756);
nor U2999 (N_2999,In_421,In_1746);
and U3000 (N_3000,In_1158,In_1381);
nor U3001 (N_3001,In_932,In_1043);
nor U3002 (N_3002,In_1836,In_1516);
nor U3003 (N_3003,In_334,In_206);
nor U3004 (N_3004,In_972,In_1275);
xnor U3005 (N_3005,In_991,In_1493);
xor U3006 (N_3006,In_1326,In_82);
nor U3007 (N_3007,In_880,In_449);
and U3008 (N_3008,In_842,In_1550);
nand U3009 (N_3009,In_1776,In_411);
nor U3010 (N_3010,In_1810,In_653);
or U3011 (N_3011,In_1016,In_95);
nor U3012 (N_3012,In_2,In_1352);
and U3013 (N_3013,In_321,In_1559);
xor U3014 (N_3014,In_1193,In_1365);
and U3015 (N_3015,In_1088,In_310);
nand U3016 (N_3016,In_1085,In_36);
nor U3017 (N_3017,In_430,In_1654);
or U3018 (N_3018,In_1965,In_531);
nor U3019 (N_3019,In_1306,In_1804);
and U3020 (N_3020,In_1587,In_786);
nand U3021 (N_3021,In_293,In_744);
nand U3022 (N_3022,In_876,In_1890);
nand U3023 (N_3023,In_1521,In_1434);
or U3024 (N_3024,In_191,In_355);
or U3025 (N_3025,In_659,In_401);
nand U3026 (N_3026,In_1917,In_744);
nand U3027 (N_3027,In_532,In_231);
and U3028 (N_3028,In_20,In_1641);
or U3029 (N_3029,In_841,In_95);
and U3030 (N_3030,In_933,In_253);
and U3031 (N_3031,In_1238,In_634);
xnor U3032 (N_3032,In_321,In_102);
nand U3033 (N_3033,In_1493,In_633);
nor U3034 (N_3034,In_1871,In_394);
or U3035 (N_3035,In_374,In_1417);
or U3036 (N_3036,In_451,In_1329);
and U3037 (N_3037,In_741,In_1184);
and U3038 (N_3038,In_1160,In_1985);
xnor U3039 (N_3039,In_935,In_1245);
or U3040 (N_3040,In_757,In_1512);
or U3041 (N_3041,In_1066,In_48);
nor U3042 (N_3042,In_1825,In_1671);
nand U3043 (N_3043,In_1267,In_902);
nand U3044 (N_3044,In_1361,In_1624);
and U3045 (N_3045,In_707,In_1301);
nand U3046 (N_3046,In_1698,In_1990);
and U3047 (N_3047,In_829,In_671);
and U3048 (N_3048,In_18,In_696);
or U3049 (N_3049,In_1020,In_1630);
or U3050 (N_3050,In_690,In_209);
and U3051 (N_3051,In_571,In_1951);
nor U3052 (N_3052,In_356,In_314);
nor U3053 (N_3053,In_1366,In_403);
and U3054 (N_3054,In_1921,In_1327);
or U3055 (N_3055,In_36,In_1581);
nand U3056 (N_3056,In_206,In_1339);
nor U3057 (N_3057,In_888,In_1853);
and U3058 (N_3058,In_1173,In_1414);
nand U3059 (N_3059,In_746,In_79);
nor U3060 (N_3060,In_103,In_1304);
and U3061 (N_3061,In_1157,In_1620);
or U3062 (N_3062,In_92,In_323);
nor U3063 (N_3063,In_1963,In_359);
nand U3064 (N_3064,In_1454,In_1201);
or U3065 (N_3065,In_425,In_1193);
nand U3066 (N_3066,In_1908,In_413);
nor U3067 (N_3067,In_1293,In_57);
and U3068 (N_3068,In_326,In_1306);
or U3069 (N_3069,In_296,In_1316);
xor U3070 (N_3070,In_1815,In_268);
or U3071 (N_3071,In_398,In_30);
nand U3072 (N_3072,In_488,In_631);
nand U3073 (N_3073,In_1154,In_827);
nand U3074 (N_3074,In_1328,In_18);
and U3075 (N_3075,In_832,In_1552);
nand U3076 (N_3076,In_1412,In_1593);
xor U3077 (N_3077,In_845,In_1362);
nor U3078 (N_3078,In_1671,In_1970);
and U3079 (N_3079,In_280,In_921);
and U3080 (N_3080,In_994,In_871);
nand U3081 (N_3081,In_1766,In_215);
nor U3082 (N_3082,In_1687,In_1853);
or U3083 (N_3083,In_1814,In_1743);
nor U3084 (N_3084,In_1079,In_511);
nand U3085 (N_3085,In_1673,In_285);
xor U3086 (N_3086,In_716,In_1516);
nor U3087 (N_3087,In_912,In_984);
and U3088 (N_3088,In_1715,In_1866);
and U3089 (N_3089,In_1783,In_1513);
nand U3090 (N_3090,In_291,In_1502);
xor U3091 (N_3091,In_852,In_1474);
or U3092 (N_3092,In_1017,In_741);
nand U3093 (N_3093,In_1464,In_1836);
nand U3094 (N_3094,In_1688,In_690);
and U3095 (N_3095,In_975,In_1721);
nand U3096 (N_3096,In_1479,In_1594);
nor U3097 (N_3097,In_1770,In_1741);
nand U3098 (N_3098,In_1629,In_521);
nand U3099 (N_3099,In_1884,In_970);
or U3100 (N_3100,In_1124,In_235);
nor U3101 (N_3101,In_988,In_1106);
nor U3102 (N_3102,In_1456,In_824);
nand U3103 (N_3103,In_769,In_177);
and U3104 (N_3104,In_298,In_661);
nor U3105 (N_3105,In_1956,In_1716);
nand U3106 (N_3106,In_516,In_1265);
nor U3107 (N_3107,In_885,In_1414);
nor U3108 (N_3108,In_1401,In_239);
or U3109 (N_3109,In_1758,In_1220);
nor U3110 (N_3110,In_905,In_1303);
or U3111 (N_3111,In_1763,In_132);
and U3112 (N_3112,In_1674,In_1453);
nor U3113 (N_3113,In_596,In_12);
or U3114 (N_3114,In_1815,In_1253);
nor U3115 (N_3115,In_1999,In_1506);
xor U3116 (N_3116,In_915,In_1443);
or U3117 (N_3117,In_780,In_954);
or U3118 (N_3118,In_46,In_295);
or U3119 (N_3119,In_1052,In_1562);
or U3120 (N_3120,In_614,In_1299);
nor U3121 (N_3121,In_482,In_837);
and U3122 (N_3122,In_1799,In_361);
or U3123 (N_3123,In_450,In_1613);
xnor U3124 (N_3124,In_406,In_649);
or U3125 (N_3125,In_879,In_1316);
and U3126 (N_3126,In_1258,In_1455);
or U3127 (N_3127,In_988,In_1278);
and U3128 (N_3128,In_1424,In_1512);
xor U3129 (N_3129,In_124,In_575);
or U3130 (N_3130,In_53,In_998);
xor U3131 (N_3131,In_1417,In_34);
nor U3132 (N_3132,In_231,In_488);
nor U3133 (N_3133,In_1795,In_972);
nand U3134 (N_3134,In_238,In_525);
nand U3135 (N_3135,In_1862,In_348);
and U3136 (N_3136,In_1308,In_801);
nand U3137 (N_3137,In_1685,In_891);
nand U3138 (N_3138,In_1045,In_285);
and U3139 (N_3139,In_1457,In_1447);
xnor U3140 (N_3140,In_562,In_451);
nand U3141 (N_3141,In_764,In_1754);
or U3142 (N_3142,In_1656,In_398);
xor U3143 (N_3143,In_1018,In_1514);
or U3144 (N_3144,In_420,In_793);
or U3145 (N_3145,In_578,In_641);
or U3146 (N_3146,In_399,In_1569);
or U3147 (N_3147,In_498,In_1399);
or U3148 (N_3148,In_1764,In_849);
and U3149 (N_3149,In_1079,In_1701);
or U3150 (N_3150,In_1873,In_1726);
nand U3151 (N_3151,In_138,In_141);
nor U3152 (N_3152,In_1811,In_43);
or U3153 (N_3153,In_1699,In_861);
xor U3154 (N_3154,In_1999,In_267);
nor U3155 (N_3155,In_1941,In_911);
nand U3156 (N_3156,In_1029,In_1361);
or U3157 (N_3157,In_1727,In_449);
nor U3158 (N_3158,In_747,In_375);
nand U3159 (N_3159,In_1468,In_1211);
and U3160 (N_3160,In_160,In_1555);
or U3161 (N_3161,In_565,In_1354);
and U3162 (N_3162,In_1032,In_431);
or U3163 (N_3163,In_1847,In_665);
nand U3164 (N_3164,In_248,In_158);
nand U3165 (N_3165,In_624,In_324);
nand U3166 (N_3166,In_233,In_584);
nor U3167 (N_3167,In_253,In_757);
nor U3168 (N_3168,In_807,In_1628);
nand U3169 (N_3169,In_1549,In_1309);
nor U3170 (N_3170,In_1130,In_432);
and U3171 (N_3171,In_1460,In_1610);
nand U3172 (N_3172,In_133,In_1544);
or U3173 (N_3173,In_344,In_1097);
or U3174 (N_3174,In_110,In_645);
xor U3175 (N_3175,In_1234,In_887);
and U3176 (N_3176,In_1597,In_1435);
nor U3177 (N_3177,In_1804,In_698);
and U3178 (N_3178,In_443,In_485);
and U3179 (N_3179,In_1019,In_1731);
and U3180 (N_3180,In_517,In_171);
or U3181 (N_3181,In_1713,In_1300);
or U3182 (N_3182,In_459,In_1463);
nand U3183 (N_3183,In_1859,In_510);
nand U3184 (N_3184,In_1137,In_445);
or U3185 (N_3185,In_756,In_40);
nand U3186 (N_3186,In_675,In_1675);
nor U3187 (N_3187,In_1679,In_1783);
nand U3188 (N_3188,In_1502,In_731);
nand U3189 (N_3189,In_1164,In_123);
or U3190 (N_3190,In_850,In_246);
and U3191 (N_3191,In_98,In_1048);
and U3192 (N_3192,In_1730,In_989);
nor U3193 (N_3193,In_1658,In_1613);
nor U3194 (N_3194,In_975,In_735);
and U3195 (N_3195,In_1515,In_388);
nor U3196 (N_3196,In_106,In_851);
or U3197 (N_3197,In_1129,In_57);
nor U3198 (N_3198,In_854,In_1723);
or U3199 (N_3199,In_1470,In_684);
nand U3200 (N_3200,In_406,In_1257);
xor U3201 (N_3201,In_1665,In_1989);
and U3202 (N_3202,In_929,In_459);
xor U3203 (N_3203,In_1332,In_1068);
nand U3204 (N_3204,In_470,In_1522);
or U3205 (N_3205,In_1183,In_1199);
or U3206 (N_3206,In_438,In_1168);
nand U3207 (N_3207,In_1704,In_1573);
nor U3208 (N_3208,In_942,In_1974);
nand U3209 (N_3209,In_586,In_820);
nor U3210 (N_3210,In_1806,In_1899);
nand U3211 (N_3211,In_589,In_1316);
nand U3212 (N_3212,In_124,In_122);
nand U3213 (N_3213,In_1749,In_1113);
and U3214 (N_3214,In_1727,In_1925);
xnor U3215 (N_3215,In_689,In_1243);
nand U3216 (N_3216,In_1627,In_598);
and U3217 (N_3217,In_188,In_1187);
nor U3218 (N_3218,In_1735,In_622);
and U3219 (N_3219,In_135,In_1482);
or U3220 (N_3220,In_1544,In_914);
xnor U3221 (N_3221,In_754,In_1212);
and U3222 (N_3222,In_958,In_1597);
nor U3223 (N_3223,In_1947,In_1213);
nand U3224 (N_3224,In_944,In_1496);
nor U3225 (N_3225,In_581,In_109);
xor U3226 (N_3226,In_1770,In_826);
or U3227 (N_3227,In_1496,In_1068);
and U3228 (N_3228,In_79,In_1601);
and U3229 (N_3229,In_441,In_256);
and U3230 (N_3230,In_834,In_792);
or U3231 (N_3231,In_1140,In_1358);
or U3232 (N_3232,In_294,In_1567);
and U3233 (N_3233,In_115,In_468);
nor U3234 (N_3234,In_657,In_315);
or U3235 (N_3235,In_1682,In_1520);
nand U3236 (N_3236,In_1985,In_1707);
nand U3237 (N_3237,In_644,In_1068);
nor U3238 (N_3238,In_1120,In_733);
nor U3239 (N_3239,In_1617,In_1764);
xor U3240 (N_3240,In_1867,In_1236);
and U3241 (N_3241,In_667,In_360);
nor U3242 (N_3242,In_35,In_1706);
nand U3243 (N_3243,In_297,In_1011);
or U3244 (N_3244,In_825,In_830);
nor U3245 (N_3245,In_1323,In_357);
xor U3246 (N_3246,In_1494,In_1447);
nand U3247 (N_3247,In_1466,In_1048);
or U3248 (N_3248,In_913,In_1766);
nand U3249 (N_3249,In_1802,In_881);
or U3250 (N_3250,In_679,In_748);
and U3251 (N_3251,In_1407,In_324);
nand U3252 (N_3252,In_1132,In_1045);
or U3253 (N_3253,In_1117,In_710);
nor U3254 (N_3254,In_1220,In_852);
xnor U3255 (N_3255,In_1511,In_1182);
nand U3256 (N_3256,In_128,In_1113);
nand U3257 (N_3257,In_297,In_1335);
nor U3258 (N_3258,In_1751,In_1673);
xor U3259 (N_3259,In_276,In_1922);
and U3260 (N_3260,In_1994,In_1080);
nor U3261 (N_3261,In_1230,In_1288);
and U3262 (N_3262,In_44,In_824);
or U3263 (N_3263,In_464,In_742);
xnor U3264 (N_3264,In_1732,In_1817);
and U3265 (N_3265,In_504,In_1889);
or U3266 (N_3266,In_1530,In_68);
nand U3267 (N_3267,In_48,In_1910);
or U3268 (N_3268,In_1047,In_1256);
nand U3269 (N_3269,In_413,In_1082);
nand U3270 (N_3270,In_572,In_1557);
nor U3271 (N_3271,In_332,In_1324);
nand U3272 (N_3272,In_1711,In_1430);
xor U3273 (N_3273,In_401,In_1451);
xnor U3274 (N_3274,In_1936,In_1078);
xor U3275 (N_3275,In_475,In_15);
or U3276 (N_3276,In_1724,In_408);
or U3277 (N_3277,In_1894,In_1948);
and U3278 (N_3278,In_1404,In_1648);
or U3279 (N_3279,In_1470,In_1391);
and U3280 (N_3280,In_1186,In_1839);
and U3281 (N_3281,In_785,In_410);
nand U3282 (N_3282,In_804,In_1464);
nor U3283 (N_3283,In_1411,In_1444);
or U3284 (N_3284,In_232,In_1890);
nor U3285 (N_3285,In_30,In_894);
and U3286 (N_3286,In_743,In_371);
nand U3287 (N_3287,In_1695,In_1087);
nand U3288 (N_3288,In_1748,In_1097);
or U3289 (N_3289,In_1221,In_1222);
or U3290 (N_3290,In_719,In_1412);
and U3291 (N_3291,In_395,In_1528);
and U3292 (N_3292,In_147,In_1492);
or U3293 (N_3293,In_1425,In_954);
nor U3294 (N_3294,In_1152,In_1125);
nor U3295 (N_3295,In_1096,In_279);
nand U3296 (N_3296,In_690,In_530);
and U3297 (N_3297,In_1599,In_461);
xnor U3298 (N_3298,In_1815,In_1512);
nand U3299 (N_3299,In_910,In_114);
or U3300 (N_3300,In_831,In_1177);
or U3301 (N_3301,In_394,In_1179);
and U3302 (N_3302,In_1541,In_365);
nor U3303 (N_3303,In_253,In_626);
nor U3304 (N_3304,In_1729,In_1303);
nand U3305 (N_3305,In_1087,In_123);
and U3306 (N_3306,In_135,In_1016);
or U3307 (N_3307,In_435,In_1775);
or U3308 (N_3308,In_1359,In_1869);
nand U3309 (N_3309,In_1604,In_1484);
nand U3310 (N_3310,In_607,In_1152);
nor U3311 (N_3311,In_767,In_795);
nand U3312 (N_3312,In_204,In_1241);
nand U3313 (N_3313,In_1794,In_281);
or U3314 (N_3314,In_1661,In_848);
nand U3315 (N_3315,In_1944,In_614);
nand U3316 (N_3316,In_669,In_1672);
or U3317 (N_3317,In_1042,In_890);
and U3318 (N_3318,In_225,In_152);
and U3319 (N_3319,In_374,In_1552);
nand U3320 (N_3320,In_1476,In_888);
nand U3321 (N_3321,In_287,In_1599);
and U3322 (N_3322,In_900,In_1833);
or U3323 (N_3323,In_1556,In_1658);
nand U3324 (N_3324,In_703,In_923);
or U3325 (N_3325,In_1336,In_1365);
and U3326 (N_3326,In_1474,In_779);
nand U3327 (N_3327,In_1262,In_1625);
xor U3328 (N_3328,In_1809,In_628);
nor U3329 (N_3329,In_346,In_551);
nor U3330 (N_3330,In_1013,In_541);
nand U3331 (N_3331,In_1136,In_166);
and U3332 (N_3332,In_460,In_1407);
or U3333 (N_3333,In_769,In_1088);
and U3334 (N_3334,In_783,In_1808);
nor U3335 (N_3335,In_335,In_1135);
and U3336 (N_3336,In_1284,In_1030);
and U3337 (N_3337,In_945,In_1070);
or U3338 (N_3338,In_1693,In_1739);
and U3339 (N_3339,In_151,In_747);
nor U3340 (N_3340,In_910,In_448);
and U3341 (N_3341,In_333,In_1477);
and U3342 (N_3342,In_1811,In_1175);
nor U3343 (N_3343,In_462,In_1905);
nor U3344 (N_3344,In_928,In_1096);
nand U3345 (N_3345,In_1667,In_125);
and U3346 (N_3346,In_288,In_905);
or U3347 (N_3347,In_1194,In_717);
nand U3348 (N_3348,In_258,In_328);
and U3349 (N_3349,In_316,In_2);
nand U3350 (N_3350,In_901,In_298);
nand U3351 (N_3351,In_1337,In_619);
nor U3352 (N_3352,In_1812,In_1231);
nor U3353 (N_3353,In_464,In_687);
nor U3354 (N_3354,In_499,In_704);
and U3355 (N_3355,In_350,In_152);
nand U3356 (N_3356,In_455,In_1403);
or U3357 (N_3357,In_1204,In_725);
and U3358 (N_3358,In_1281,In_1824);
nand U3359 (N_3359,In_1907,In_1712);
and U3360 (N_3360,In_1999,In_913);
nand U3361 (N_3361,In_460,In_1524);
and U3362 (N_3362,In_678,In_341);
nand U3363 (N_3363,In_400,In_687);
nand U3364 (N_3364,In_1598,In_1338);
nand U3365 (N_3365,In_290,In_1190);
or U3366 (N_3366,In_466,In_1304);
and U3367 (N_3367,In_554,In_684);
and U3368 (N_3368,In_84,In_325);
nor U3369 (N_3369,In_317,In_335);
xor U3370 (N_3370,In_1132,In_177);
nand U3371 (N_3371,In_1852,In_88);
nand U3372 (N_3372,In_98,In_1158);
nand U3373 (N_3373,In_1074,In_263);
nand U3374 (N_3374,In_1489,In_328);
and U3375 (N_3375,In_666,In_1382);
nor U3376 (N_3376,In_1535,In_246);
nand U3377 (N_3377,In_520,In_1414);
nor U3378 (N_3378,In_417,In_49);
and U3379 (N_3379,In_485,In_736);
nor U3380 (N_3380,In_301,In_1387);
or U3381 (N_3381,In_1072,In_234);
or U3382 (N_3382,In_1894,In_1210);
and U3383 (N_3383,In_793,In_423);
nand U3384 (N_3384,In_1693,In_181);
or U3385 (N_3385,In_219,In_1889);
nor U3386 (N_3386,In_1680,In_1055);
and U3387 (N_3387,In_225,In_845);
or U3388 (N_3388,In_1160,In_944);
nor U3389 (N_3389,In_1474,In_707);
or U3390 (N_3390,In_1964,In_1476);
or U3391 (N_3391,In_15,In_1576);
nand U3392 (N_3392,In_755,In_1289);
nor U3393 (N_3393,In_974,In_322);
or U3394 (N_3394,In_890,In_502);
or U3395 (N_3395,In_561,In_752);
nor U3396 (N_3396,In_44,In_870);
or U3397 (N_3397,In_228,In_482);
nor U3398 (N_3398,In_1504,In_67);
nor U3399 (N_3399,In_1856,In_385);
nor U3400 (N_3400,In_477,In_933);
nand U3401 (N_3401,In_288,In_654);
nand U3402 (N_3402,In_342,In_1060);
nand U3403 (N_3403,In_1862,In_1180);
nor U3404 (N_3404,In_1392,In_1814);
nand U3405 (N_3405,In_1608,In_1961);
nand U3406 (N_3406,In_1522,In_1526);
and U3407 (N_3407,In_1560,In_787);
or U3408 (N_3408,In_63,In_765);
nand U3409 (N_3409,In_1917,In_406);
nand U3410 (N_3410,In_531,In_819);
nor U3411 (N_3411,In_1655,In_557);
nand U3412 (N_3412,In_298,In_206);
nand U3413 (N_3413,In_924,In_1712);
or U3414 (N_3414,In_1144,In_1169);
and U3415 (N_3415,In_1136,In_668);
nor U3416 (N_3416,In_1424,In_1745);
nand U3417 (N_3417,In_359,In_1249);
or U3418 (N_3418,In_1148,In_1504);
and U3419 (N_3419,In_1578,In_394);
nor U3420 (N_3420,In_865,In_734);
and U3421 (N_3421,In_1856,In_826);
nor U3422 (N_3422,In_1310,In_781);
xnor U3423 (N_3423,In_1939,In_809);
and U3424 (N_3424,In_347,In_261);
nor U3425 (N_3425,In_651,In_1877);
nor U3426 (N_3426,In_1172,In_1927);
or U3427 (N_3427,In_805,In_1746);
xor U3428 (N_3428,In_1285,In_433);
nand U3429 (N_3429,In_1727,In_1884);
or U3430 (N_3430,In_929,In_345);
and U3431 (N_3431,In_633,In_394);
xnor U3432 (N_3432,In_1407,In_933);
nand U3433 (N_3433,In_512,In_1059);
xor U3434 (N_3434,In_1859,In_1863);
and U3435 (N_3435,In_69,In_68);
nand U3436 (N_3436,In_42,In_706);
nand U3437 (N_3437,In_1788,In_1524);
and U3438 (N_3438,In_1360,In_1422);
and U3439 (N_3439,In_875,In_327);
nand U3440 (N_3440,In_28,In_1425);
or U3441 (N_3441,In_727,In_675);
or U3442 (N_3442,In_1334,In_1926);
nor U3443 (N_3443,In_758,In_350);
nand U3444 (N_3444,In_1298,In_1782);
xnor U3445 (N_3445,In_1409,In_109);
or U3446 (N_3446,In_634,In_1588);
nor U3447 (N_3447,In_1883,In_285);
nand U3448 (N_3448,In_1571,In_1755);
xnor U3449 (N_3449,In_1352,In_1767);
nor U3450 (N_3450,In_708,In_1269);
and U3451 (N_3451,In_953,In_219);
nand U3452 (N_3452,In_1967,In_1525);
or U3453 (N_3453,In_1104,In_1527);
nand U3454 (N_3454,In_1715,In_603);
or U3455 (N_3455,In_1320,In_883);
nor U3456 (N_3456,In_32,In_719);
or U3457 (N_3457,In_275,In_1986);
nand U3458 (N_3458,In_799,In_1006);
nor U3459 (N_3459,In_1672,In_508);
nor U3460 (N_3460,In_1399,In_525);
or U3461 (N_3461,In_852,In_1016);
nand U3462 (N_3462,In_465,In_127);
xnor U3463 (N_3463,In_117,In_1466);
nor U3464 (N_3464,In_1363,In_1718);
and U3465 (N_3465,In_799,In_856);
and U3466 (N_3466,In_358,In_1947);
or U3467 (N_3467,In_662,In_787);
or U3468 (N_3468,In_1088,In_1587);
and U3469 (N_3469,In_1308,In_850);
or U3470 (N_3470,In_1503,In_1142);
or U3471 (N_3471,In_1161,In_1229);
or U3472 (N_3472,In_1940,In_1259);
nor U3473 (N_3473,In_1617,In_912);
nor U3474 (N_3474,In_562,In_1208);
or U3475 (N_3475,In_1894,In_1416);
nor U3476 (N_3476,In_1522,In_1353);
nor U3477 (N_3477,In_1606,In_573);
nor U3478 (N_3478,In_122,In_1728);
and U3479 (N_3479,In_1023,In_412);
nand U3480 (N_3480,In_1662,In_943);
and U3481 (N_3481,In_169,In_1371);
nand U3482 (N_3482,In_823,In_1323);
and U3483 (N_3483,In_386,In_1966);
and U3484 (N_3484,In_1131,In_1947);
or U3485 (N_3485,In_794,In_1886);
or U3486 (N_3486,In_1212,In_257);
xor U3487 (N_3487,In_1554,In_1697);
nand U3488 (N_3488,In_1080,In_319);
or U3489 (N_3489,In_1844,In_1651);
or U3490 (N_3490,In_1623,In_53);
or U3491 (N_3491,In_1423,In_886);
nand U3492 (N_3492,In_1958,In_135);
nor U3493 (N_3493,In_781,In_1957);
nand U3494 (N_3494,In_1996,In_1075);
nor U3495 (N_3495,In_1284,In_537);
nand U3496 (N_3496,In_72,In_1630);
or U3497 (N_3497,In_1042,In_51);
nand U3498 (N_3498,In_1600,In_455);
nor U3499 (N_3499,In_250,In_1434);
nor U3500 (N_3500,In_31,In_927);
nand U3501 (N_3501,In_1024,In_559);
xnor U3502 (N_3502,In_182,In_767);
and U3503 (N_3503,In_1055,In_672);
and U3504 (N_3504,In_444,In_1381);
nand U3505 (N_3505,In_1788,In_1935);
nor U3506 (N_3506,In_1941,In_897);
xnor U3507 (N_3507,In_945,In_1875);
nand U3508 (N_3508,In_1211,In_1929);
and U3509 (N_3509,In_1353,In_438);
nor U3510 (N_3510,In_1887,In_1110);
nand U3511 (N_3511,In_1516,In_973);
nor U3512 (N_3512,In_1034,In_804);
and U3513 (N_3513,In_305,In_1110);
nand U3514 (N_3514,In_896,In_747);
nand U3515 (N_3515,In_88,In_1694);
or U3516 (N_3516,In_749,In_989);
and U3517 (N_3517,In_141,In_114);
and U3518 (N_3518,In_1650,In_1276);
xnor U3519 (N_3519,In_1693,In_1567);
nand U3520 (N_3520,In_235,In_1220);
or U3521 (N_3521,In_63,In_107);
or U3522 (N_3522,In_964,In_733);
nor U3523 (N_3523,In_1674,In_346);
nor U3524 (N_3524,In_1219,In_378);
nor U3525 (N_3525,In_104,In_906);
nand U3526 (N_3526,In_1746,In_1251);
nor U3527 (N_3527,In_601,In_795);
and U3528 (N_3528,In_1902,In_187);
and U3529 (N_3529,In_1579,In_730);
xnor U3530 (N_3530,In_20,In_337);
and U3531 (N_3531,In_1929,In_1308);
nor U3532 (N_3532,In_26,In_1034);
or U3533 (N_3533,In_951,In_1662);
and U3534 (N_3534,In_1790,In_1145);
or U3535 (N_3535,In_724,In_1342);
or U3536 (N_3536,In_1760,In_1343);
nand U3537 (N_3537,In_107,In_1564);
or U3538 (N_3538,In_1106,In_1284);
and U3539 (N_3539,In_1083,In_1485);
or U3540 (N_3540,In_62,In_961);
or U3541 (N_3541,In_561,In_290);
and U3542 (N_3542,In_1970,In_1526);
nor U3543 (N_3543,In_1133,In_1410);
and U3544 (N_3544,In_746,In_1223);
nand U3545 (N_3545,In_123,In_1921);
and U3546 (N_3546,In_1497,In_872);
and U3547 (N_3547,In_1495,In_1870);
nand U3548 (N_3548,In_983,In_1499);
or U3549 (N_3549,In_491,In_183);
and U3550 (N_3550,In_1033,In_1833);
nand U3551 (N_3551,In_857,In_328);
nor U3552 (N_3552,In_1791,In_744);
nand U3553 (N_3553,In_719,In_130);
xor U3554 (N_3554,In_497,In_974);
and U3555 (N_3555,In_1293,In_654);
and U3556 (N_3556,In_1517,In_1425);
xnor U3557 (N_3557,In_1164,In_1330);
nor U3558 (N_3558,In_1689,In_892);
nand U3559 (N_3559,In_1153,In_943);
and U3560 (N_3560,In_1487,In_1145);
or U3561 (N_3561,In_1738,In_836);
xnor U3562 (N_3562,In_1747,In_542);
and U3563 (N_3563,In_1885,In_357);
nand U3564 (N_3564,In_45,In_759);
or U3565 (N_3565,In_660,In_230);
nor U3566 (N_3566,In_649,In_736);
and U3567 (N_3567,In_1575,In_213);
or U3568 (N_3568,In_1529,In_1549);
and U3569 (N_3569,In_315,In_91);
or U3570 (N_3570,In_415,In_1041);
and U3571 (N_3571,In_204,In_212);
and U3572 (N_3572,In_625,In_963);
nor U3573 (N_3573,In_14,In_1630);
nor U3574 (N_3574,In_1905,In_1899);
nor U3575 (N_3575,In_1879,In_654);
or U3576 (N_3576,In_1371,In_234);
nor U3577 (N_3577,In_119,In_248);
or U3578 (N_3578,In_1490,In_504);
or U3579 (N_3579,In_1517,In_1568);
and U3580 (N_3580,In_524,In_1374);
and U3581 (N_3581,In_1527,In_1080);
nor U3582 (N_3582,In_1569,In_306);
nand U3583 (N_3583,In_1740,In_437);
or U3584 (N_3584,In_1438,In_1109);
and U3585 (N_3585,In_266,In_593);
xnor U3586 (N_3586,In_312,In_1987);
nor U3587 (N_3587,In_1892,In_38);
and U3588 (N_3588,In_1731,In_1561);
or U3589 (N_3589,In_1034,In_965);
xnor U3590 (N_3590,In_1396,In_664);
and U3591 (N_3591,In_82,In_1028);
or U3592 (N_3592,In_1395,In_162);
or U3593 (N_3593,In_500,In_1957);
or U3594 (N_3594,In_839,In_1969);
or U3595 (N_3595,In_741,In_958);
and U3596 (N_3596,In_381,In_1760);
nand U3597 (N_3597,In_53,In_1792);
or U3598 (N_3598,In_1337,In_1518);
and U3599 (N_3599,In_1811,In_1690);
nor U3600 (N_3600,In_397,In_1003);
xor U3601 (N_3601,In_886,In_666);
nand U3602 (N_3602,In_1299,In_1671);
nand U3603 (N_3603,In_1474,In_1267);
and U3604 (N_3604,In_588,In_1296);
or U3605 (N_3605,In_907,In_1607);
nor U3606 (N_3606,In_153,In_253);
and U3607 (N_3607,In_874,In_1409);
and U3608 (N_3608,In_1367,In_1087);
and U3609 (N_3609,In_526,In_8);
or U3610 (N_3610,In_1326,In_853);
nor U3611 (N_3611,In_1667,In_629);
nor U3612 (N_3612,In_323,In_1023);
and U3613 (N_3613,In_1384,In_275);
nand U3614 (N_3614,In_946,In_1504);
nor U3615 (N_3615,In_56,In_1060);
and U3616 (N_3616,In_1552,In_476);
nand U3617 (N_3617,In_339,In_1209);
nor U3618 (N_3618,In_1790,In_1151);
and U3619 (N_3619,In_584,In_879);
or U3620 (N_3620,In_498,In_1139);
and U3621 (N_3621,In_1281,In_1603);
or U3622 (N_3622,In_855,In_1576);
nor U3623 (N_3623,In_1329,In_864);
nand U3624 (N_3624,In_375,In_1253);
nor U3625 (N_3625,In_883,In_351);
and U3626 (N_3626,In_1594,In_395);
and U3627 (N_3627,In_831,In_516);
and U3628 (N_3628,In_1795,In_1460);
and U3629 (N_3629,In_440,In_590);
and U3630 (N_3630,In_1671,In_1297);
nor U3631 (N_3631,In_447,In_320);
and U3632 (N_3632,In_49,In_53);
or U3633 (N_3633,In_700,In_1331);
nand U3634 (N_3634,In_1164,In_416);
and U3635 (N_3635,In_1795,In_1718);
nor U3636 (N_3636,In_948,In_151);
xor U3637 (N_3637,In_1033,In_414);
nand U3638 (N_3638,In_592,In_1238);
nor U3639 (N_3639,In_1423,In_722);
nor U3640 (N_3640,In_271,In_1507);
and U3641 (N_3641,In_204,In_1739);
nand U3642 (N_3642,In_1516,In_1752);
and U3643 (N_3643,In_486,In_953);
and U3644 (N_3644,In_496,In_650);
or U3645 (N_3645,In_11,In_442);
xnor U3646 (N_3646,In_1608,In_603);
xnor U3647 (N_3647,In_1163,In_1382);
xor U3648 (N_3648,In_1248,In_1638);
or U3649 (N_3649,In_652,In_1632);
nand U3650 (N_3650,In_1696,In_1603);
nand U3651 (N_3651,In_105,In_704);
and U3652 (N_3652,In_1204,In_986);
or U3653 (N_3653,In_1749,In_527);
and U3654 (N_3654,In_463,In_304);
nand U3655 (N_3655,In_848,In_1921);
or U3656 (N_3656,In_1171,In_1264);
nor U3657 (N_3657,In_1138,In_146);
nor U3658 (N_3658,In_1706,In_1776);
or U3659 (N_3659,In_834,In_1887);
or U3660 (N_3660,In_1874,In_550);
or U3661 (N_3661,In_1809,In_1212);
and U3662 (N_3662,In_236,In_682);
nand U3663 (N_3663,In_339,In_112);
nand U3664 (N_3664,In_670,In_1075);
nor U3665 (N_3665,In_167,In_699);
or U3666 (N_3666,In_1688,In_1481);
or U3667 (N_3667,In_493,In_1626);
xnor U3668 (N_3668,In_659,In_1737);
or U3669 (N_3669,In_453,In_1991);
xor U3670 (N_3670,In_145,In_1325);
nor U3671 (N_3671,In_770,In_1596);
nor U3672 (N_3672,In_1442,In_555);
and U3673 (N_3673,In_822,In_485);
nor U3674 (N_3674,In_1734,In_235);
or U3675 (N_3675,In_413,In_1542);
nand U3676 (N_3676,In_674,In_376);
nand U3677 (N_3677,In_8,In_1031);
nor U3678 (N_3678,In_1271,In_570);
nand U3679 (N_3679,In_1022,In_753);
nor U3680 (N_3680,In_389,In_1613);
and U3681 (N_3681,In_1223,In_538);
nor U3682 (N_3682,In_1106,In_480);
and U3683 (N_3683,In_39,In_1400);
nand U3684 (N_3684,In_1004,In_219);
nand U3685 (N_3685,In_979,In_453);
or U3686 (N_3686,In_1240,In_1194);
nand U3687 (N_3687,In_715,In_878);
nand U3688 (N_3688,In_1337,In_1722);
or U3689 (N_3689,In_1558,In_946);
or U3690 (N_3690,In_206,In_1724);
xnor U3691 (N_3691,In_455,In_492);
nand U3692 (N_3692,In_1214,In_704);
nand U3693 (N_3693,In_616,In_948);
nand U3694 (N_3694,In_281,In_1712);
or U3695 (N_3695,In_1537,In_1857);
and U3696 (N_3696,In_855,In_1993);
xnor U3697 (N_3697,In_552,In_599);
and U3698 (N_3698,In_1361,In_1539);
nor U3699 (N_3699,In_49,In_334);
nor U3700 (N_3700,In_1388,In_1158);
and U3701 (N_3701,In_930,In_1685);
nand U3702 (N_3702,In_1817,In_1658);
and U3703 (N_3703,In_572,In_54);
nand U3704 (N_3704,In_545,In_1808);
nor U3705 (N_3705,In_1673,In_169);
nand U3706 (N_3706,In_549,In_229);
and U3707 (N_3707,In_1373,In_1860);
and U3708 (N_3708,In_1085,In_1202);
or U3709 (N_3709,In_1675,In_36);
and U3710 (N_3710,In_1621,In_813);
xnor U3711 (N_3711,In_976,In_1791);
or U3712 (N_3712,In_270,In_1536);
xnor U3713 (N_3713,In_59,In_319);
nand U3714 (N_3714,In_739,In_1523);
and U3715 (N_3715,In_784,In_254);
or U3716 (N_3716,In_1984,In_741);
nand U3717 (N_3717,In_1258,In_792);
or U3718 (N_3718,In_819,In_1709);
xnor U3719 (N_3719,In_266,In_448);
nand U3720 (N_3720,In_1423,In_279);
or U3721 (N_3721,In_729,In_228);
nand U3722 (N_3722,In_1076,In_1086);
or U3723 (N_3723,In_21,In_1579);
or U3724 (N_3724,In_1238,In_166);
and U3725 (N_3725,In_804,In_706);
nor U3726 (N_3726,In_799,In_1009);
nand U3727 (N_3727,In_1756,In_1482);
and U3728 (N_3728,In_1465,In_1219);
and U3729 (N_3729,In_1305,In_1958);
and U3730 (N_3730,In_614,In_249);
nor U3731 (N_3731,In_1367,In_895);
and U3732 (N_3732,In_1247,In_1161);
or U3733 (N_3733,In_642,In_1997);
and U3734 (N_3734,In_171,In_1596);
nand U3735 (N_3735,In_1119,In_814);
and U3736 (N_3736,In_227,In_1942);
nand U3737 (N_3737,In_1779,In_1059);
nor U3738 (N_3738,In_709,In_1803);
xor U3739 (N_3739,In_418,In_1807);
nand U3740 (N_3740,In_571,In_208);
and U3741 (N_3741,In_1453,In_1720);
and U3742 (N_3742,In_992,In_1637);
and U3743 (N_3743,In_1163,In_62);
and U3744 (N_3744,In_270,In_1109);
or U3745 (N_3745,In_1510,In_882);
nor U3746 (N_3746,In_178,In_897);
nor U3747 (N_3747,In_1091,In_841);
and U3748 (N_3748,In_257,In_160);
and U3749 (N_3749,In_1440,In_592);
and U3750 (N_3750,In_1438,In_1637);
and U3751 (N_3751,In_785,In_803);
nor U3752 (N_3752,In_1111,In_1140);
nand U3753 (N_3753,In_1777,In_939);
nor U3754 (N_3754,In_1727,In_814);
nor U3755 (N_3755,In_1353,In_236);
and U3756 (N_3756,In_389,In_670);
nand U3757 (N_3757,In_1802,In_1399);
nand U3758 (N_3758,In_128,In_974);
and U3759 (N_3759,In_519,In_408);
and U3760 (N_3760,In_1400,In_1335);
or U3761 (N_3761,In_323,In_894);
or U3762 (N_3762,In_986,In_267);
nor U3763 (N_3763,In_1503,In_1898);
xnor U3764 (N_3764,In_1786,In_1430);
and U3765 (N_3765,In_1614,In_895);
or U3766 (N_3766,In_146,In_1625);
nor U3767 (N_3767,In_323,In_186);
nor U3768 (N_3768,In_1444,In_1578);
and U3769 (N_3769,In_1014,In_81);
nor U3770 (N_3770,In_872,In_121);
and U3771 (N_3771,In_1516,In_528);
or U3772 (N_3772,In_868,In_997);
or U3773 (N_3773,In_748,In_1602);
nor U3774 (N_3774,In_443,In_1400);
and U3775 (N_3775,In_859,In_1792);
or U3776 (N_3776,In_17,In_391);
or U3777 (N_3777,In_1276,In_1772);
and U3778 (N_3778,In_1293,In_1180);
or U3779 (N_3779,In_468,In_1869);
nand U3780 (N_3780,In_648,In_628);
or U3781 (N_3781,In_125,In_984);
nand U3782 (N_3782,In_326,In_1302);
or U3783 (N_3783,In_1485,In_1544);
and U3784 (N_3784,In_1499,In_11);
and U3785 (N_3785,In_116,In_1671);
xor U3786 (N_3786,In_738,In_159);
nand U3787 (N_3787,In_1058,In_1281);
nor U3788 (N_3788,In_79,In_1192);
nor U3789 (N_3789,In_231,In_1266);
or U3790 (N_3790,In_1268,In_287);
and U3791 (N_3791,In_333,In_233);
nand U3792 (N_3792,In_1187,In_678);
nand U3793 (N_3793,In_1540,In_1111);
nor U3794 (N_3794,In_907,In_1351);
nand U3795 (N_3795,In_730,In_741);
and U3796 (N_3796,In_1500,In_1618);
or U3797 (N_3797,In_1198,In_628);
or U3798 (N_3798,In_837,In_1737);
and U3799 (N_3799,In_1930,In_899);
nor U3800 (N_3800,In_1515,In_504);
and U3801 (N_3801,In_450,In_1257);
nand U3802 (N_3802,In_965,In_1755);
nor U3803 (N_3803,In_1267,In_588);
and U3804 (N_3804,In_412,In_1493);
nor U3805 (N_3805,In_1379,In_908);
nor U3806 (N_3806,In_717,In_1906);
and U3807 (N_3807,In_1863,In_1402);
nand U3808 (N_3808,In_1898,In_1822);
xor U3809 (N_3809,In_1113,In_779);
or U3810 (N_3810,In_1976,In_1467);
nor U3811 (N_3811,In_1944,In_477);
nor U3812 (N_3812,In_1362,In_205);
xor U3813 (N_3813,In_1577,In_1480);
nand U3814 (N_3814,In_865,In_1432);
nand U3815 (N_3815,In_570,In_1478);
xor U3816 (N_3816,In_933,In_99);
and U3817 (N_3817,In_220,In_1150);
or U3818 (N_3818,In_533,In_1086);
xor U3819 (N_3819,In_1907,In_1292);
nand U3820 (N_3820,In_1346,In_213);
and U3821 (N_3821,In_1637,In_1631);
or U3822 (N_3822,In_356,In_594);
and U3823 (N_3823,In_1624,In_214);
and U3824 (N_3824,In_51,In_147);
nand U3825 (N_3825,In_1121,In_159);
nor U3826 (N_3826,In_491,In_1722);
and U3827 (N_3827,In_1898,In_1153);
nor U3828 (N_3828,In_268,In_56);
and U3829 (N_3829,In_1747,In_1324);
or U3830 (N_3830,In_1847,In_1940);
and U3831 (N_3831,In_174,In_1513);
or U3832 (N_3832,In_643,In_1704);
or U3833 (N_3833,In_869,In_1638);
nand U3834 (N_3834,In_1876,In_1879);
nand U3835 (N_3835,In_1497,In_124);
and U3836 (N_3836,In_1340,In_744);
nand U3837 (N_3837,In_1104,In_413);
xnor U3838 (N_3838,In_1620,In_1418);
xnor U3839 (N_3839,In_1547,In_1811);
and U3840 (N_3840,In_202,In_1287);
or U3841 (N_3841,In_619,In_419);
or U3842 (N_3842,In_1147,In_1604);
nor U3843 (N_3843,In_1175,In_1357);
nand U3844 (N_3844,In_1327,In_1340);
nand U3845 (N_3845,In_1797,In_1609);
xor U3846 (N_3846,In_617,In_1821);
xor U3847 (N_3847,In_1242,In_1942);
or U3848 (N_3848,In_680,In_138);
nor U3849 (N_3849,In_0,In_1539);
nand U3850 (N_3850,In_1393,In_1848);
and U3851 (N_3851,In_1139,In_847);
or U3852 (N_3852,In_1332,In_747);
and U3853 (N_3853,In_1773,In_467);
nor U3854 (N_3854,In_1864,In_1481);
or U3855 (N_3855,In_253,In_1004);
and U3856 (N_3856,In_43,In_700);
nor U3857 (N_3857,In_381,In_167);
nand U3858 (N_3858,In_1681,In_1789);
and U3859 (N_3859,In_941,In_962);
or U3860 (N_3860,In_1378,In_1919);
or U3861 (N_3861,In_1629,In_723);
nor U3862 (N_3862,In_832,In_1927);
and U3863 (N_3863,In_667,In_1004);
nand U3864 (N_3864,In_172,In_78);
nand U3865 (N_3865,In_398,In_1378);
nor U3866 (N_3866,In_1746,In_1196);
and U3867 (N_3867,In_1525,In_1503);
nor U3868 (N_3868,In_1154,In_1352);
nand U3869 (N_3869,In_383,In_546);
xor U3870 (N_3870,In_443,In_843);
nand U3871 (N_3871,In_1493,In_923);
nor U3872 (N_3872,In_894,In_272);
or U3873 (N_3873,In_819,In_1917);
and U3874 (N_3874,In_1110,In_1296);
nor U3875 (N_3875,In_1628,In_690);
xnor U3876 (N_3876,In_1638,In_429);
or U3877 (N_3877,In_388,In_1716);
or U3878 (N_3878,In_653,In_545);
or U3879 (N_3879,In_733,In_1964);
nor U3880 (N_3880,In_2,In_856);
or U3881 (N_3881,In_834,In_526);
nand U3882 (N_3882,In_1991,In_1760);
and U3883 (N_3883,In_1074,In_1949);
and U3884 (N_3884,In_86,In_1625);
and U3885 (N_3885,In_623,In_471);
and U3886 (N_3886,In_164,In_1763);
or U3887 (N_3887,In_752,In_1378);
nor U3888 (N_3888,In_1321,In_1747);
or U3889 (N_3889,In_1407,In_1865);
nor U3890 (N_3890,In_1107,In_32);
nand U3891 (N_3891,In_829,In_616);
or U3892 (N_3892,In_863,In_1593);
and U3893 (N_3893,In_482,In_291);
nand U3894 (N_3894,In_1154,In_114);
and U3895 (N_3895,In_693,In_1316);
or U3896 (N_3896,In_1572,In_542);
xnor U3897 (N_3897,In_1480,In_340);
and U3898 (N_3898,In_1104,In_1398);
or U3899 (N_3899,In_965,In_1655);
or U3900 (N_3900,In_1713,In_242);
nor U3901 (N_3901,In_38,In_1314);
and U3902 (N_3902,In_1604,In_1589);
or U3903 (N_3903,In_241,In_705);
and U3904 (N_3904,In_622,In_1818);
nor U3905 (N_3905,In_827,In_186);
and U3906 (N_3906,In_417,In_218);
and U3907 (N_3907,In_1856,In_1196);
or U3908 (N_3908,In_856,In_1953);
and U3909 (N_3909,In_172,In_702);
or U3910 (N_3910,In_852,In_1469);
or U3911 (N_3911,In_1507,In_1247);
xnor U3912 (N_3912,In_1880,In_1094);
nand U3913 (N_3913,In_1378,In_1620);
or U3914 (N_3914,In_1736,In_1541);
nor U3915 (N_3915,In_1915,In_322);
nand U3916 (N_3916,In_1239,In_1649);
nor U3917 (N_3917,In_1879,In_1968);
and U3918 (N_3918,In_738,In_1503);
nand U3919 (N_3919,In_1318,In_795);
and U3920 (N_3920,In_1201,In_951);
nand U3921 (N_3921,In_522,In_1033);
xnor U3922 (N_3922,In_1966,In_1851);
nor U3923 (N_3923,In_1393,In_1869);
nor U3924 (N_3924,In_67,In_248);
xnor U3925 (N_3925,In_969,In_897);
nand U3926 (N_3926,In_604,In_1555);
nand U3927 (N_3927,In_1862,In_1409);
nor U3928 (N_3928,In_988,In_687);
and U3929 (N_3929,In_1221,In_1307);
and U3930 (N_3930,In_206,In_1822);
nand U3931 (N_3931,In_773,In_1669);
and U3932 (N_3932,In_1344,In_1391);
and U3933 (N_3933,In_345,In_969);
nand U3934 (N_3934,In_1450,In_1808);
nor U3935 (N_3935,In_1552,In_737);
and U3936 (N_3936,In_1419,In_911);
or U3937 (N_3937,In_1746,In_1780);
xnor U3938 (N_3938,In_791,In_1488);
or U3939 (N_3939,In_1200,In_859);
nor U3940 (N_3940,In_1190,In_1874);
xnor U3941 (N_3941,In_1617,In_812);
nand U3942 (N_3942,In_921,In_427);
nand U3943 (N_3943,In_499,In_653);
xnor U3944 (N_3944,In_920,In_1112);
or U3945 (N_3945,In_12,In_1899);
nor U3946 (N_3946,In_530,In_1233);
nor U3947 (N_3947,In_1303,In_1594);
xor U3948 (N_3948,In_519,In_1127);
xnor U3949 (N_3949,In_478,In_1704);
or U3950 (N_3950,In_634,In_1135);
nor U3951 (N_3951,In_1549,In_524);
nand U3952 (N_3952,In_1789,In_1980);
xnor U3953 (N_3953,In_613,In_1474);
nand U3954 (N_3954,In_1617,In_492);
nor U3955 (N_3955,In_1341,In_232);
and U3956 (N_3956,In_659,In_1956);
and U3957 (N_3957,In_272,In_1555);
and U3958 (N_3958,In_1234,In_1513);
or U3959 (N_3959,In_1633,In_1762);
nor U3960 (N_3960,In_1749,In_864);
nand U3961 (N_3961,In_1473,In_258);
and U3962 (N_3962,In_784,In_557);
or U3963 (N_3963,In_236,In_1888);
and U3964 (N_3964,In_1595,In_1710);
and U3965 (N_3965,In_1423,In_217);
xnor U3966 (N_3966,In_785,In_632);
and U3967 (N_3967,In_146,In_467);
nand U3968 (N_3968,In_222,In_1410);
or U3969 (N_3969,In_1208,In_482);
or U3970 (N_3970,In_1128,In_89);
and U3971 (N_3971,In_1895,In_866);
nor U3972 (N_3972,In_26,In_1876);
nor U3973 (N_3973,In_1443,In_1931);
and U3974 (N_3974,In_970,In_1820);
or U3975 (N_3975,In_1673,In_412);
nor U3976 (N_3976,In_1336,In_1509);
nor U3977 (N_3977,In_935,In_1283);
xnor U3978 (N_3978,In_1747,In_117);
xnor U3979 (N_3979,In_1293,In_282);
and U3980 (N_3980,In_1005,In_693);
and U3981 (N_3981,In_385,In_97);
and U3982 (N_3982,In_142,In_1781);
nand U3983 (N_3983,In_1498,In_1671);
nor U3984 (N_3984,In_923,In_691);
nor U3985 (N_3985,In_494,In_1042);
nor U3986 (N_3986,In_170,In_490);
and U3987 (N_3987,In_87,In_868);
xor U3988 (N_3988,In_864,In_1245);
nor U3989 (N_3989,In_287,In_1787);
nand U3990 (N_3990,In_555,In_1701);
or U3991 (N_3991,In_45,In_1254);
and U3992 (N_3992,In_1548,In_1300);
or U3993 (N_3993,In_453,In_1641);
xor U3994 (N_3994,In_1905,In_1431);
and U3995 (N_3995,In_721,In_1533);
and U3996 (N_3996,In_1355,In_897);
nand U3997 (N_3997,In_303,In_1963);
nand U3998 (N_3998,In_1637,In_464);
or U3999 (N_3999,In_1722,In_124);
or U4000 (N_4000,N_188,N_3305);
and U4001 (N_4001,N_3092,N_3590);
xor U4002 (N_4002,N_2736,N_1896);
nand U4003 (N_4003,N_682,N_850);
and U4004 (N_4004,N_2397,N_3224);
nand U4005 (N_4005,N_24,N_2528);
nor U4006 (N_4006,N_2877,N_3094);
nand U4007 (N_4007,N_201,N_2704);
nand U4008 (N_4008,N_3902,N_732);
nor U4009 (N_4009,N_1966,N_2266);
or U4010 (N_4010,N_1234,N_2104);
and U4011 (N_4011,N_1099,N_274);
or U4012 (N_4012,N_3886,N_1963);
nor U4013 (N_4013,N_2468,N_913);
nor U4014 (N_4014,N_2093,N_1331);
or U4015 (N_4015,N_1066,N_2676);
and U4016 (N_4016,N_3301,N_2047);
nor U4017 (N_4017,N_510,N_2150);
and U4018 (N_4018,N_1822,N_3551);
nor U4019 (N_4019,N_1904,N_1807);
xnor U4020 (N_4020,N_2957,N_1696);
nor U4021 (N_4021,N_2671,N_1200);
nor U4022 (N_4022,N_2503,N_731);
nor U4023 (N_4023,N_1558,N_1);
or U4024 (N_4024,N_1713,N_3166);
nor U4025 (N_4025,N_2342,N_55);
or U4026 (N_4026,N_2247,N_1054);
xnor U4027 (N_4027,N_1702,N_2937);
nor U4028 (N_4028,N_3350,N_3736);
nand U4029 (N_4029,N_1447,N_1420);
and U4030 (N_4030,N_215,N_1813);
nor U4031 (N_4031,N_887,N_1092);
and U4032 (N_4032,N_1164,N_2315);
nor U4033 (N_4033,N_1529,N_3307);
and U4034 (N_4034,N_2183,N_507);
nor U4035 (N_4035,N_3270,N_3329);
nand U4036 (N_4036,N_189,N_515);
nor U4037 (N_4037,N_2445,N_1943);
and U4038 (N_4038,N_1658,N_1568);
nor U4039 (N_4039,N_2823,N_284);
nand U4040 (N_4040,N_1586,N_404);
and U4041 (N_4041,N_3624,N_3968);
and U4042 (N_4042,N_569,N_1498);
nand U4043 (N_4043,N_3415,N_2885);
nand U4044 (N_4044,N_1839,N_1353);
or U4045 (N_4045,N_3703,N_3868);
and U4046 (N_4046,N_2152,N_1992);
or U4047 (N_4047,N_2238,N_2112);
or U4048 (N_4048,N_499,N_3744);
nand U4049 (N_4049,N_1470,N_1442);
or U4050 (N_4050,N_1081,N_1358);
xnor U4051 (N_4051,N_2624,N_167);
and U4052 (N_4052,N_3107,N_1743);
nand U4053 (N_4053,N_344,N_2506);
xnor U4054 (N_4054,N_2589,N_1874);
and U4055 (N_4055,N_30,N_103);
nor U4056 (N_4056,N_3017,N_3198);
nand U4057 (N_4057,N_3487,N_2322);
and U4058 (N_4058,N_1112,N_2904);
and U4059 (N_4059,N_3405,N_1968);
and U4060 (N_4060,N_1138,N_2526);
and U4061 (N_4061,N_2870,N_2893);
nor U4062 (N_4062,N_593,N_3413);
and U4063 (N_4063,N_2961,N_3796);
or U4064 (N_4064,N_1335,N_3163);
nand U4065 (N_4065,N_3167,N_3569);
xnor U4066 (N_4066,N_2006,N_793);
nand U4067 (N_4067,N_2082,N_2107);
and U4068 (N_4068,N_1569,N_3374);
or U4069 (N_4069,N_2387,N_3943);
nand U4070 (N_4070,N_2162,N_3820);
and U4071 (N_4071,N_2921,N_3354);
xor U4072 (N_4072,N_3843,N_203);
or U4073 (N_4073,N_31,N_1545);
or U4074 (N_4074,N_478,N_843);
or U4075 (N_4075,N_1387,N_1903);
nor U4076 (N_4076,N_3225,N_3472);
or U4077 (N_4077,N_1394,N_1119);
or U4078 (N_4078,N_2631,N_2802);
nand U4079 (N_4079,N_3102,N_3561);
nand U4080 (N_4080,N_763,N_3360);
or U4081 (N_4081,N_2625,N_3383);
or U4082 (N_4082,N_2177,N_3040);
xor U4083 (N_4083,N_1067,N_3719);
nand U4084 (N_4084,N_559,N_2700);
nand U4085 (N_4085,N_1158,N_2778);
nor U4086 (N_4086,N_3372,N_3461);
and U4087 (N_4087,N_749,N_1727);
nor U4088 (N_4088,N_3620,N_1267);
or U4089 (N_4089,N_2829,N_3190);
and U4090 (N_4090,N_3099,N_2358);
nand U4091 (N_4091,N_3189,N_3644);
nor U4092 (N_4092,N_1539,N_3481);
or U4093 (N_4093,N_3257,N_1315);
nand U4094 (N_4094,N_2556,N_2500);
nand U4095 (N_4095,N_3809,N_1153);
nand U4096 (N_4096,N_3647,N_3860);
or U4097 (N_4097,N_759,N_3815);
nand U4098 (N_4098,N_906,N_597);
xnor U4099 (N_4099,N_3835,N_2081);
and U4100 (N_4100,N_3291,N_1742);
xnor U4101 (N_4101,N_2760,N_464);
or U4102 (N_4102,N_3712,N_1374);
or U4103 (N_4103,N_1795,N_1564);
nand U4104 (N_4104,N_3451,N_821);
and U4105 (N_4105,N_3641,N_3739);
nor U4106 (N_4106,N_3687,N_1176);
nand U4107 (N_4107,N_350,N_3955);
and U4108 (N_4108,N_17,N_2030);
and U4109 (N_4109,N_3020,N_1731);
nor U4110 (N_4110,N_1383,N_3759);
nand U4111 (N_4111,N_1068,N_85);
xor U4112 (N_4112,N_1243,N_2057);
nor U4113 (N_4113,N_3885,N_514);
or U4114 (N_4114,N_1484,N_931);
nor U4115 (N_4115,N_1403,N_1320);
and U4116 (N_4116,N_3090,N_1427);
and U4117 (N_4117,N_1690,N_156);
nor U4118 (N_4118,N_3573,N_3169);
nand U4119 (N_4119,N_1371,N_2175);
nand U4120 (N_4120,N_1299,N_2723);
or U4121 (N_4121,N_526,N_2211);
nor U4122 (N_4122,N_865,N_3227);
nand U4123 (N_4123,N_2910,N_3807);
or U4124 (N_4124,N_208,N_1030);
or U4125 (N_4125,N_390,N_500);
or U4126 (N_4126,N_3001,N_3850);
or U4127 (N_4127,N_2043,N_2301);
and U4128 (N_4128,N_3531,N_2703);
and U4129 (N_4129,N_2362,N_2552);
and U4130 (N_4130,N_1302,N_3164);
nand U4131 (N_4131,N_2989,N_3332);
nor U4132 (N_4132,N_2965,N_3865);
and U4133 (N_4133,N_2694,N_2742);
nor U4134 (N_4134,N_1217,N_198);
and U4135 (N_4135,N_445,N_3116);
nor U4136 (N_4136,N_577,N_1973);
and U4137 (N_4137,N_3370,N_3022);
nand U4138 (N_4138,N_2109,N_448);
nand U4139 (N_4139,N_3373,N_3580);
nor U4140 (N_4140,N_1009,N_567);
or U4141 (N_4141,N_1046,N_2633);
or U4142 (N_4142,N_549,N_1750);
or U4143 (N_4143,N_439,N_565);
or U4144 (N_4144,N_989,N_3987);
or U4145 (N_4145,N_2472,N_3948);
nor U4146 (N_4146,N_1824,N_742);
nor U4147 (N_4147,N_1974,N_592);
or U4148 (N_4148,N_886,N_2602);
xnor U4149 (N_4149,N_1666,N_1191);
and U4150 (N_4150,N_3312,N_1855);
and U4151 (N_4151,N_1058,N_585);
xor U4152 (N_4152,N_1579,N_3658);
nand U4153 (N_4153,N_1525,N_3394);
and U4154 (N_4154,N_1537,N_3000);
nor U4155 (N_4155,N_2309,N_2771);
or U4156 (N_4156,N_3606,N_2600);
xor U4157 (N_4157,N_2966,N_3345);
nand U4158 (N_4158,N_3651,N_2350);
xnor U4159 (N_4159,N_3664,N_1803);
nand U4160 (N_4160,N_1983,N_2592);
nor U4161 (N_4161,N_3371,N_456);
and U4162 (N_4162,N_3236,N_287);
and U4163 (N_4163,N_3926,N_626);
or U4164 (N_4164,N_3366,N_303);
nand U4165 (N_4165,N_2680,N_229);
and U4166 (N_4166,N_3592,N_286);
or U4167 (N_4167,N_880,N_2594);
nand U4168 (N_4168,N_957,N_2292);
or U4169 (N_4169,N_3696,N_87);
nand U4170 (N_4170,N_300,N_1951);
xnor U4171 (N_4171,N_368,N_3051);
nor U4172 (N_4172,N_107,N_1155);
and U4173 (N_4173,N_1179,N_1082);
or U4174 (N_4174,N_2856,N_3155);
or U4175 (N_4175,N_81,N_2151);
nor U4176 (N_4176,N_1532,N_3384);
and U4177 (N_4177,N_3336,N_283);
or U4178 (N_4178,N_1031,N_102);
and U4179 (N_4179,N_1755,N_681);
and U4180 (N_4180,N_2487,N_863);
or U4181 (N_4181,N_3258,N_1481);
or U4182 (N_4182,N_2812,N_135);
nor U4183 (N_4183,N_1825,N_3381);
and U4184 (N_4184,N_1362,N_105);
and U4185 (N_4185,N_3134,N_3513);
nor U4186 (N_4186,N_1310,N_1608);
and U4187 (N_4187,N_2347,N_3724);
nand U4188 (N_4188,N_3053,N_940);
nor U4189 (N_4189,N_1661,N_1655);
nand U4190 (N_4190,N_1872,N_1754);
xnor U4191 (N_4191,N_777,N_830);
and U4192 (N_4192,N_19,N_1469);
xnor U4193 (N_4193,N_463,N_3057);
nand U4194 (N_4194,N_2629,N_438);
or U4195 (N_4195,N_2719,N_2400);
nand U4196 (N_4196,N_823,N_1053);
nand U4197 (N_4197,N_2750,N_1132);
or U4198 (N_4198,N_3672,N_1706);
or U4199 (N_4199,N_612,N_1207);
and U4200 (N_4200,N_2765,N_934);
and U4201 (N_4201,N_651,N_3816);
or U4202 (N_4202,N_1664,N_222);
and U4203 (N_4203,N_2832,N_190);
and U4204 (N_4204,N_3254,N_1865);
and U4205 (N_4205,N_1926,N_2690);
or U4206 (N_4206,N_2618,N_3996);
nand U4207 (N_4207,N_1039,N_477);
and U4208 (N_4208,N_1329,N_178);
nand U4209 (N_4209,N_1256,N_3694);
or U4210 (N_4210,N_3993,N_1739);
nand U4211 (N_4211,N_2681,N_3362);
or U4212 (N_4212,N_3125,N_2311);
and U4213 (N_4213,N_2155,N_2191);
nand U4214 (N_4214,N_774,N_538);
and U4215 (N_4215,N_124,N_2094);
nor U4216 (N_4216,N_3699,N_3516);
nor U4217 (N_4217,N_3443,N_1952);
or U4218 (N_4218,N_2406,N_688);
or U4219 (N_4219,N_1154,N_2022);
nor U4220 (N_4220,N_154,N_45);
xnor U4221 (N_4221,N_3289,N_2337);
xnor U4222 (N_4222,N_2981,N_485);
nor U4223 (N_4223,N_2115,N_2188);
or U4224 (N_4224,N_2903,N_3033);
or U4225 (N_4225,N_1915,N_722);
and U4226 (N_4226,N_2139,N_648);
nand U4227 (N_4227,N_3014,N_3842);
or U4228 (N_4228,N_795,N_2161);
nand U4229 (N_4229,N_2687,N_3386);
nand U4230 (N_4230,N_753,N_840);
nor U4231 (N_4231,N_1546,N_762);
and U4232 (N_4232,N_3088,N_2834);
or U4233 (N_4233,N_995,N_2665);
xor U4234 (N_4234,N_3859,N_3610);
nor U4235 (N_4235,N_486,N_3091);
and U4236 (N_4236,N_816,N_436);
and U4237 (N_4237,N_2697,N_3806);
nor U4238 (N_4238,N_1863,N_1991);
or U4239 (N_4239,N_3547,N_1404);
and U4240 (N_4240,N_1467,N_3075);
nand U4241 (N_4241,N_2086,N_3940);
and U4242 (N_4242,N_1388,N_3441);
nand U4243 (N_4243,N_1004,N_1185);
or U4244 (N_4244,N_1471,N_2270);
nand U4245 (N_4245,N_726,N_1715);
or U4246 (N_4246,N_721,N_406);
and U4247 (N_4247,N_1245,N_1604);
and U4248 (N_4248,N_3751,N_3660);
or U4249 (N_4249,N_433,N_956);
xor U4250 (N_4250,N_2553,N_2546);
or U4251 (N_4251,N_2414,N_3553);
nand U4252 (N_4252,N_217,N_3630);
or U4253 (N_4253,N_1137,N_3789);
nor U4254 (N_4254,N_1761,N_2100);
or U4255 (N_4255,N_2875,N_750);
or U4256 (N_4256,N_733,N_2853);
or U4257 (N_4257,N_3283,N_3844);
or U4258 (N_4258,N_2088,N_2340);
and U4259 (N_4259,N_3450,N_2717);
xor U4260 (N_4260,N_2864,N_2193);
nand U4261 (N_4261,N_2336,N_2729);
nand U4262 (N_4262,N_1492,N_3783);
nor U4263 (N_4263,N_1878,N_3463);
xor U4264 (N_4264,N_973,N_2579);
nand U4265 (N_4265,N_134,N_320);
nor U4266 (N_4266,N_389,N_1305);
nand U4267 (N_4267,N_645,N_3454);
nor U4268 (N_4268,N_233,N_37);
nor U4269 (N_4269,N_3087,N_1435);
nor U4270 (N_4270,N_1291,N_1444);
and U4271 (N_4271,N_64,N_2627);
nor U4272 (N_4272,N_2999,N_2324);
or U4273 (N_4273,N_3201,N_3890);
xnor U4274 (N_4274,N_114,N_836);
nor U4275 (N_4275,N_4,N_2686);
nor U4276 (N_4276,N_79,N_1107);
xor U4277 (N_4277,N_3064,N_3595);
and U4278 (N_4278,N_2805,N_677);
or U4279 (N_4279,N_2172,N_26);
xor U4280 (N_4280,N_2,N_555);
nor U4281 (N_4281,N_981,N_318);
and U4282 (N_4282,N_1889,N_1100);
or U4283 (N_4283,N_2262,N_3012);
or U4284 (N_4284,N_2170,N_1180);
or U4285 (N_4285,N_3863,N_3168);
nand U4286 (N_4286,N_2210,N_1847);
and U4287 (N_4287,N_1640,N_1900);
xnor U4288 (N_4288,N_3275,N_2016);
nor U4289 (N_4289,N_987,N_2245);
nand U4290 (N_4290,N_3156,N_2648);
nand U4291 (N_4291,N_480,N_3929);
nor U4292 (N_4292,N_1965,N_3839);
nor U4293 (N_4293,N_652,N_1653);
xnor U4294 (N_4294,N_2833,N_2300);
or U4295 (N_4295,N_59,N_2126);
and U4296 (N_4296,N_3294,N_2939);
nor U4297 (N_4297,N_548,N_1593);
nor U4298 (N_4298,N_686,N_2450);
or U4299 (N_4299,N_768,N_2221);
nor U4300 (N_4300,N_3388,N_1919);
nand U4301 (N_4301,N_504,N_988);
nand U4302 (N_4302,N_925,N_3627);
and U4303 (N_4303,N_3858,N_3027);
nor U4304 (N_4304,N_892,N_3532);
or U4305 (N_4305,N_3741,N_1766);
or U4306 (N_4306,N_1065,N_3032);
and U4307 (N_4307,N_1748,N_2695);
nor U4308 (N_4308,N_1596,N_3105);
or U4309 (N_4309,N_2424,N_3436);
nor U4310 (N_4310,N_251,N_1946);
and U4311 (N_4311,N_2174,N_3278);
and U4312 (N_4312,N_3976,N_1478);
and U4313 (N_4313,N_2233,N_2169);
nor U4314 (N_4314,N_2576,N_473);
and U4315 (N_4315,N_3262,N_3591);
and U4316 (N_4316,N_1248,N_226);
or U4317 (N_4317,N_3625,N_3315);
xnor U4318 (N_4318,N_3206,N_3133);
nor U4319 (N_4319,N_361,N_2940);
nor U4320 (N_4320,N_3805,N_3674);
nand U4321 (N_4321,N_815,N_88);
nor U4322 (N_4322,N_2960,N_3678);
nand U4323 (N_4323,N_2838,N_2458);
and U4324 (N_4324,N_334,N_3306);
or U4325 (N_4325,N_3086,N_496);
nor U4326 (N_4326,N_2845,N_2715);
and U4327 (N_4327,N_2105,N_2048);
and U4328 (N_4328,N_1543,N_1511);
nand U4329 (N_4329,N_3251,N_1028);
and U4330 (N_4330,N_1106,N_370);
or U4331 (N_4331,N_3477,N_3212);
xnor U4332 (N_4332,N_2754,N_838);
and U4333 (N_4333,N_3565,N_2316);
nor U4334 (N_4334,N_2840,N_1105);
or U4335 (N_4335,N_2947,N_275);
nor U4336 (N_4336,N_2140,N_308);
nor U4337 (N_4337,N_2120,N_2741);
nor U4338 (N_4338,N_3135,N_50);
and U4339 (N_4339,N_3395,N_595);
nand U4340 (N_4340,N_2611,N_183);
and U4341 (N_4341,N_961,N_3072);
and U4342 (N_4342,N_2605,N_1140);
or U4343 (N_4343,N_1981,N_3946);
or U4344 (N_4344,N_978,N_125);
and U4345 (N_4345,N_2413,N_980);
nor U4346 (N_4346,N_3442,N_185);
or U4347 (N_4347,N_2938,N_1408);
nor U4348 (N_4348,N_3083,N_2251);
nand U4349 (N_4349,N_3872,N_2705);
and U4350 (N_4350,N_348,N_2523);
nand U4351 (N_4351,N_2720,N_3958);
nor U4352 (N_4352,N_2612,N_802);
nand U4353 (N_4353,N_2144,N_1202);
nand U4354 (N_4354,N_3473,N_3879);
or U4355 (N_4355,N_455,N_2917);
xor U4356 (N_4356,N_740,N_1641);
nand U4357 (N_4357,N_950,N_2492);
or U4358 (N_4358,N_1225,N_3884);
and U4359 (N_4359,N_3002,N_527);
or U4360 (N_4360,N_1113,N_798);
and U4361 (N_4361,N_946,N_1259);
nand U4362 (N_4362,N_3145,N_1769);
xnor U4363 (N_4363,N_1483,N_3279);
nor U4364 (N_4364,N_3732,N_3512);
nor U4365 (N_4365,N_3813,N_3605);
nand U4366 (N_4366,N_674,N_3338);
or U4367 (N_4367,N_1345,N_3855);
nand U4368 (N_4368,N_1798,N_3132);
or U4369 (N_4369,N_498,N_1728);
and U4370 (N_4370,N_2606,N_2601);
nand U4371 (N_4371,N_1506,N_191);
or U4372 (N_4372,N_3136,N_3418);
nor U4373 (N_4373,N_1232,N_2257);
or U4374 (N_4374,N_1346,N_3552);
xor U4375 (N_4375,N_773,N_3024);
or U4376 (N_4376,N_1687,N_714);
and U4377 (N_4377,N_3250,N_930);
nand U4378 (N_4378,N_2025,N_2465);
nand U4379 (N_4379,N_2452,N_3670);
nor U4380 (N_4380,N_1920,N_2329);
nor U4381 (N_4381,N_1209,N_3753);
nor U4382 (N_4382,N_1573,N_708);
xor U4383 (N_4383,N_262,N_2933);
nand U4384 (N_4384,N_3713,N_709);
and U4385 (N_4385,N_2099,N_1917);
or U4386 (N_4386,N_2352,N_3247);
and U4387 (N_4387,N_1227,N_3389);
and U4388 (N_4388,N_1826,N_2818);
or U4389 (N_4389,N_1147,N_2872);
nand U4390 (N_4390,N_2032,N_809);
and U4391 (N_4391,N_482,N_3424);
nor U4392 (N_4392,N_2843,N_1022);
nor U4393 (N_4393,N_3339,N_3676);
nand U4394 (N_4394,N_3937,N_1665);
nand U4395 (N_4395,N_3367,N_285);
nand U4396 (N_4396,N_517,N_864);
or U4397 (N_4397,N_3080,N_2454);
nor U4398 (N_4398,N_2216,N_2573);
or U4399 (N_4399,N_3823,N_3705);
nand U4400 (N_4400,N_3439,N_571);
or U4401 (N_4401,N_1636,N_1675);
xnor U4402 (N_4402,N_2357,N_1434);
and U4403 (N_4403,N_2411,N_3607);
xnor U4404 (N_4404,N_1454,N_718);
or U4405 (N_4405,N_1458,N_2461);
or U4406 (N_4406,N_2020,N_547);
and U4407 (N_4407,N_2936,N_1941);
nand U4408 (N_4408,N_1990,N_2319);
nand U4409 (N_4409,N_3071,N_1521);
and U4410 (N_4410,N_535,N_2683);
and U4411 (N_4411,N_1544,N_1133);
nand U4412 (N_4412,N_2998,N_2429);
or U4413 (N_4413,N_634,N_2739);
nor U4414 (N_4414,N_1489,N_831);
nand U4415 (N_4415,N_3750,N_76);
or U4416 (N_4416,N_2133,N_2136);
nor U4417 (N_4417,N_74,N_1491);
xor U4418 (N_4418,N_926,N_2249);
and U4419 (N_4419,N_33,N_1777);
and U4420 (N_4420,N_399,N_945);
and U4421 (N_4421,N_2967,N_2428);
and U4422 (N_4422,N_3414,N_3347);
xnor U4423 (N_4423,N_1479,N_2031);
and U4424 (N_4424,N_1954,N_1349);
nor U4425 (N_4425,N_3947,N_174);
xnor U4426 (N_4426,N_2444,N_1765);
or U4427 (N_4427,N_2163,N_1311);
and U4428 (N_4428,N_3335,N_66);
nand U4429 (N_4429,N_600,N_1504);
nor U4430 (N_4430,N_2184,N_3488);
or U4431 (N_4431,N_860,N_3470);
or U4432 (N_4432,N_1007,N_1985);
and U4433 (N_4433,N_935,N_2083);
xor U4434 (N_4434,N_1413,N_411);
nand U4435 (N_4435,N_146,N_413);
or U4436 (N_4436,N_3710,N_2649);
and U4437 (N_4437,N_2531,N_1286);
nand U4438 (N_4438,N_1307,N_1197);
or U4439 (N_4439,N_3469,N_1018);
and U4440 (N_4440,N_893,N_2287);
nor U4441 (N_4441,N_84,N_173);
and U4442 (N_4442,N_3096,N_3941);
xor U4443 (N_4443,N_542,N_3542);
nand U4444 (N_4444,N_888,N_2095);
nor U4445 (N_4445,N_2436,N_3861);
xnor U4446 (N_4446,N_457,N_966);
nand U4447 (N_4447,N_1339,N_2603);
nor U4448 (N_4448,N_3044,N_1588);
nand U4449 (N_4449,N_3587,N_1669);
nor U4450 (N_4450,N_3284,N_3921);
nor U4451 (N_4451,N_964,N_1476);
nand U4452 (N_4452,N_611,N_2534);
or U4453 (N_4453,N_2376,N_3453);
nand U4454 (N_4454,N_965,N_126);
nor U4455 (N_4455,N_2326,N_1123);
xor U4456 (N_4456,N_3277,N_3160);
and U4457 (N_4457,N_3503,N_1297);
or U4458 (N_4458,N_2747,N_2632);
and U4459 (N_4459,N_2228,N_1707);
nand U4460 (N_4460,N_193,N_1783);
nand U4461 (N_4461,N_1396,N_1401);
or U4462 (N_4462,N_1314,N_1948);
or U4463 (N_4463,N_3927,N_354);
nand U4464 (N_4464,N_884,N_3799);
xnor U4465 (N_4465,N_3998,N_2770);
xnor U4466 (N_4466,N_3034,N_3965);
nand U4467 (N_4467,N_1689,N_3458);
nand U4468 (N_4468,N_2550,N_1277);
xnor U4469 (N_4469,N_557,N_280);
nand U4470 (N_4470,N_3103,N_1437);
nand U4471 (N_4471,N_3304,N_2525);
xor U4472 (N_4472,N_2306,N_3060);
nor U4473 (N_4473,N_1522,N_2499);
nand U4474 (N_4474,N_2970,N_2551);
nor U4475 (N_4475,N_866,N_3500);
xor U4476 (N_4476,N_18,N_469);
nand U4477 (N_4477,N_2246,N_1460);
or U4478 (N_4478,N_78,N_2056);
nor U4479 (N_4479,N_3120,N_3777);
nand U4480 (N_4480,N_1841,N_1221);
and U4481 (N_4481,N_631,N_2619);
or U4482 (N_4482,N_3497,N_138);
or U4483 (N_4483,N_494,N_282);
nor U4484 (N_4484,N_3269,N_1862);
nor U4485 (N_4485,N_147,N_954);
and U4486 (N_4486,N_1814,N_2673);
xnor U4487 (N_4487,N_3158,N_2331);
nand U4488 (N_4488,N_637,N_2263);
nor U4489 (N_4489,N_3889,N_1016);
or U4490 (N_4490,N_2637,N_3485);
and U4491 (N_4491,N_1587,N_3646);
or U4492 (N_4492,N_3334,N_3085);
and U4493 (N_4493,N_1617,N_3717);
nand U4494 (N_4494,N_2344,N_1024);
nand U4495 (N_4495,N_2621,N_2023);
xnor U4496 (N_4496,N_2467,N_1231);
nand U4497 (N_4497,N_1885,N_417);
nand U4498 (N_4498,N_249,N_705);
nor U4499 (N_4499,N_220,N_771);
nand U4500 (N_4500,N_2691,N_2761);
nand U4501 (N_4501,N_1226,N_3042);
nor U4502 (N_4502,N_3008,N_3808);
nor U4503 (N_4503,N_3084,N_969);
xor U4504 (N_4504,N_3242,N_2808);
nand U4505 (N_4505,N_2494,N_661);
or U4506 (N_4506,N_1561,N_1117);
nor U4507 (N_4507,N_3364,N_2814);
and U4508 (N_4508,N_1073,N_3772);
nand U4509 (N_4509,N_1169,N_1052);
and U4510 (N_4510,N_2973,N_1908);
and U4511 (N_4511,N_1412,N_2563);
or U4512 (N_4512,N_1927,N_1737);
nor U4513 (N_4513,N_2635,N_3931);
and U4514 (N_4514,N_1167,N_3194);
nand U4515 (N_4515,N_405,N_2491);
nor U4516 (N_4516,N_2407,N_1050);
nor U4517 (N_4517,N_898,N_1255);
nand U4518 (N_4518,N_1338,N_3975);
nor U4519 (N_4519,N_2071,N_2979);
nand U4520 (N_4520,N_349,N_927);
and U4521 (N_4521,N_3738,N_1429);
or U4522 (N_4522,N_2574,N_3535);
nand U4523 (N_4523,N_505,N_1375);
nor U4524 (N_4524,N_3711,N_3208);
or U4525 (N_4525,N_1061,N_2386);
or U4526 (N_4526,N_1982,N_2154);
nor U4527 (N_4527,N_1772,N_2220);
nor U4528 (N_4528,N_649,N_1567);
or U4529 (N_4529,N_1271,N_403);
or U4530 (N_4530,N_1260,N_3895);
and U4531 (N_4531,N_3368,N_804);
or U4532 (N_4532,N_1125,N_3121);
and U4533 (N_4533,N_1163,N_671);
or U4534 (N_4534,N_2328,N_181);
nor U4535 (N_4535,N_1290,N_3474);
xnor U4536 (N_4536,N_1222,N_1647);
nand U4537 (N_4537,N_32,N_171);
nand U4538 (N_4538,N_1809,N_824);
nand U4539 (N_4539,N_3175,N_1205);
nor U4540 (N_4540,N_3237,N_2102);
nor U4541 (N_4541,N_1723,N_2433);
and U4542 (N_4542,N_2272,N_1497);
nand U4543 (N_4543,N_1352,N_44);
nand U4544 (N_4544,N_3721,N_2945);
and U4545 (N_4545,N_594,N_822);
nand U4546 (N_4546,N_3583,N_3186);
xnor U4547 (N_4547,N_2268,N_536);
nor U4548 (N_4548,N_2069,N_3907);
nor U4549 (N_4549,N_449,N_2724);
nand U4550 (N_4550,N_1688,N_393);
and U4551 (N_4551,N_148,N_342);
nor U4552 (N_4552,N_164,N_3011);
or U4553 (N_4553,N_916,N_2207);
or U4554 (N_4554,N_1400,N_72);
or U4555 (N_4555,N_3814,N_1663);
or U4556 (N_4556,N_3144,N_1350);
nor U4557 (N_4557,N_1601,N_3046);
or U4558 (N_4558,N_108,N_1936);
nand U4559 (N_4559,N_1235,N_3392);
and U4560 (N_4560,N_3904,N_415);
nor U4561 (N_4561,N_3459,N_1410);
or U4562 (N_4562,N_3616,N_1281);
or U4563 (N_4563,N_835,N_2439);
or U4564 (N_4564,N_698,N_3421);
nor U4565 (N_4565,N_2914,N_1402);
or U4566 (N_4566,N_3852,N_1378);
nor U4567 (N_4567,N_2423,N_3101);
or U4568 (N_4568,N_3666,N_2469);
xor U4569 (N_4569,N_650,N_2405);
nand U4570 (N_4570,N_1372,N_3762);
and U4571 (N_4571,N_3431,N_2905);
nand U4572 (N_4572,N_744,N_3893);
nand U4573 (N_4573,N_587,N_3337);
nor U4574 (N_4574,N_2524,N_2751);
xnor U4575 (N_4575,N_3296,N_2888);
nand U4576 (N_4576,N_2176,N_1421);
nand U4577 (N_4577,N_2532,N_3429);
nor U4578 (N_4578,N_2447,N_116);
nor U4579 (N_4579,N_3986,N_3936);
nand U4580 (N_4580,N_590,N_1868);
and U4581 (N_4581,N_1716,N_2291);
nor U4582 (N_4582,N_2559,N_269);
nor U4583 (N_4583,N_1048,N_1553);
and U4584 (N_4584,N_1284,N_2488);
or U4585 (N_4585,N_2348,N_1070);
nor U4586 (N_4586,N_3643,N_3077);
nor U4587 (N_4587,N_2854,N_132);
or U4588 (N_4588,N_1683,N_1363);
nand U4589 (N_4589,N_781,N_3141);
nand U4590 (N_4590,N_46,N_2587);
or U4591 (N_4591,N_2733,N_1997);
nand U4592 (N_4592,N_1942,N_3661);
and U4593 (N_4593,N_1064,N_2243);
nand U4594 (N_4594,N_2641,N_3114);
or U4595 (N_4595,N_2430,N_2213);
xor U4596 (N_4596,N_920,N_56);
nand U4597 (N_4597,N_3745,N_3508);
nand U4598 (N_4598,N_471,N_3264);
or U4599 (N_4599,N_1294,N_1357);
or U4600 (N_4600,N_1932,N_172);
and U4601 (N_4601,N_416,N_3427);
and U4602 (N_4602,N_1779,N_1898);
and U4603 (N_4603,N_2415,N_3478);
nand U4604 (N_4604,N_1725,N_2726);
or U4605 (N_4605,N_2642,N_3361);
or U4606 (N_4606,N_2137,N_2209);
nor U4607 (N_4607,N_3891,N_2816);
and U4608 (N_4608,N_2302,N_1619);
nor U4609 (N_4609,N_101,N_2652);
and U4610 (N_4610,N_985,N_2855);
nand U4611 (N_4611,N_3455,N_992);
nand U4612 (N_4612,N_503,N_3667);
nor U4613 (N_4613,N_1577,N_3793);
nand U4614 (N_4614,N_2643,N_2768);
nor U4615 (N_4615,N_3862,N_423);
and U4616 (N_4616,N_1626,N_3098);
and U4617 (N_4617,N_2886,N_2568);
nand U4618 (N_4618,N_3391,N_2501);
and U4619 (N_4619,N_2237,N_3545);
nand U4620 (N_4620,N_1502,N_1930);
nand U4621 (N_4621,N_1673,N_1369);
nand U4622 (N_4622,N_2135,N_2283);
nand U4623 (N_4623,N_1589,N_414);
nor U4624 (N_4624,N_3310,N_829);
or U4625 (N_4625,N_3558,N_430);
xnor U4626 (N_4626,N_1215,N_218);
and U4627 (N_4627,N_3233,N_2992);
and U4628 (N_4628,N_3273,N_2475);
xor U4629 (N_4629,N_2712,N_1890);
xor U4630 (N_4630,N_3523,N_861);
or U4631 (N_4631,N_2395,N_2173);
or U4632 (N_4632,N_3548,N_3185);
nor U4633 (N_4633,N_2274,N_3460);
nor U4634 (N_4634,N_1088,N_2264);
nor U4635 (N_4635,N_578,N_936);
or U4636 (N_4636,N_2837,N_2485);
nand U4637 (N_4637,N_2219,N_3137);
or U4638 (N_4638,N_410,N_839);
or U4639 (N_4639,N_1323,N_3636);
or U4640 (N_4640,N_144,N_2464);
nor U4641 (N_4641,N_2985,N_3492);
nor U4642 (N_4642,N_1474,N_80);
nor U4643 (N_4643,N_3089,N_1439);
and U4644 (N_4644,N_2062,N_680);
or U4645 (N_4645,N_3702,N_3566);
nor U4646 (N_4646,N_790,N_1480);
or U4647 (N_4647,N_679,N_3196);
nor U4648 (N_4648,N_528,N_212);
or U4649 (N_4649,N_3322,N_1832);
nand U4650 (N_4650,N_3271,N_2497);
and U4651 (N_4651,N_2258,N_2752);
nand U4652 (N_4652,N_1275,N_3397);
and U4653 (N_4653,N_2013,N_2544);
and U4654 (N_4654,N_2335,N_1786);
nor U4655 (N_4655,N_375,N_1089);
xor U4656 (N_4656,N_3490,N_810);
and U4657 (N_4657,N_152,N_2659);
and U4658 (N_4658,N_638,N_2054);
nor U4659 (N_4659,N_785,N_3790);
xor U4660 (N_4660,N_976,N_1833);
nand U4661 (N_4661,N_3292,N_1762);
and U4662 (N_4662,N_211,N_2644);
nand U4663 (N_4663,N_1940,N_2675);
nor U4664 (N_4664,N_1220,N_1817);
nand U4665 (N_4665,N_3864,N_519);
nor U4666 (N_4666,N_3841,N_1916);
nor U4667 (N_4667,N_1679,N_2884);
nor U4668 (N_4668,N_1893,N_1041);
or U4669 (N_4669,N_1806,N_2284);
nand U4670 (N_4670,N_2014,N_3798);
or U4671 (N_4671,N_764,N_738);
nor U4672 (N_4672,N_1414,N_908);
nor U4673 (N_4673,N_673,N_290);
nor U4674 (N_4674,N_1918,N_1194);
and U4675 (N_4675,N_1615,N_794);
nand U4676 (N_4676,N_2008,N_2732);
and U4677 (N_4677,N_803,N_533);
and U4678 (N_4678,N_511,N_3061);
nand U4679 (N_4679,N_1599,N_3274);
or U4680 (N_4680,N_1272,N_2529);
and U4681 (N_4681,N_3426,N_3821);
or U4682 (N_4682,N_2798,N_2953);
and U4683 (N_4683,N_2096,N_1103);
nand U4684 (N_4684,N_41,N_938);
or U4685 (N_4685,N_1241,N_112);
nor U4686 (N_4686,N_1780,N_2748);
nor U4687 (N_4687,N_28,N_2129);
and U4688 (N_4688,N_2634,N_2230);
xnor U4689 (N_4689,N_3677,N_2995);
nor U4690 (N_4690,N_3131,N_1901);
xnor U4691 (N_4691,N_1978,N_221);
or U4692 (N_4692,N_1459,N_2543);
or U4693 (N_4693,N_1751,N_3681);
nor U4694 (N_4694,N_1616,N_2359);
and U4695 (N_4695,N_481,N_3228);
nor U4696 (N_4696,N_3496,N_663);
nor U4697 (N_4697,N_2607,N_1559);
and U4698 (N_4698,N_851,N_224);
xnor U4699 (N_4699,N_1306,N_3901);
nor U4700 (N_4700,N_206,N_264);
and U4701 (N_4701,N_3363,N_3288);
nor U4702 (N_4702,N_1888,N_3159);
xor U4703 (N_4703,N_730,N_2507);
nor U4704 (N_4704,N_2709,N_2004);
nand U4705 (N_4705,N_307,N_3897);
or U4706 (N_4706,N_163,N_1287);
nand U4707 (N_4707,N_1160,N_60);
xor U4708 (N_4708,N_2891,N_1876);
nand U4709 (N_4709,N_2178,N_2225);
or U4710 (N_4710,N_3430,N_2731);
and U4711 (N_4711,N_2323,N_3097);
or U4712 (N_4712,N_3143,N_3540);
and U4713 (N_4713,N_3445,N_306);
nor U4714 (N_4714,N_1671,N_3760);
nand U4715 (N_4715,N_1846,N_3867);
and U4716 (N_4716,N_2570,N_1449);
nand U4717 (N_4717,N_2639,N_2145);
and U4718 (N_4718,N_1468,N_51);
xnor U4719 (N_4719,N_1152,N_3050);
xor U4720 (N_4720,N_1457,N_1367);
nand U4721 (N_4721,N_1810,N_472);
nand U4722 (N_4722,N_832,N_3448);
nor U4723 (N_4723,N_2518,N_2663);
and U4724 (N_4724,N_2034,N_1212);
and U4725 (N_4725,N_3903,N_170);
nand U4726 (N_4726,N_1446,N_2810);
or U4727 (N_4727,N_3776,N_1043);
and U4728 (N_4728,N_3659,N_1431);
and U4729 (N_4729,N_490,N_3079);
nor U4730 (N_4730,N_1720,N_2075);
and U4731 (N_4731,N_2002,N_659);
nand U4732 (N_4732,N_3874,N_3124);
and U4733 (N_4733,N_1711,N_1584);
and U4734 (N_4734,N_635,N_86);
and U4735 (N_4735,N_3650,N_1101);
nand U4736 (N_4736,N_2339,N_3489);
and U4737 (N_4737,N_534,N_739);
nand U4738 (N_4738,N_169,N_345);
nand U4739 (N_4739,N_2913,N_3675);
and U4740 (N_4740,N_3549,N_706);
or U4741 (N_4741,N_3857,N_2153);
nand U4742 (N_4742,N_2988,N_2822);
nand U4743 (N_4743,N_3309,N_2111);
nand U4744 (N_4744,N_3204,N_1590);
or U4745 (N_4745,N_3142,N_1203);
or U4746 (N_4746,N_1691,N_2061);
or U4747 (N_4747,N_3544,N_3231);
nand U4748 (N_4748,N_2636,N_639);
and U4749 (N_4749,N_3645,N_1211);
and U4750 (N_4750,N_3556,N_3295);
and U4751 (N_4751,N_1334,N_2522);
nor U4752 (N_4752,N_3416,N_2481);
nand U4753 (N_4753,N_943,N_2078);
nor U4754 (N_4754,N_3218,N_3311);
nand U4755 (N_4755,N_2236,N_2206);
or U4756 (N_4756,N_1538,N_3265);
nand U4757 (N_4757,N_39,N_475);
or U4758 (N_4758,N_1818,N_2035);
nand U4759 (N_4759,N_1891,N_3953);
xor U4760 (N_4760,N_2349,N_3526);
and U4761 (N_4761,N_3297,N_2560);
nor U4762 (N_4762,N_3021,N_3393);
or U4763 (N_4763,N_2926,N_3520);
xnor U4764 (N_4764,N_1907,N_1288);
or U4765 (N_4765,N_242,N_1768);
nor U4766 (N_4766,N_2882,N_3457);
or U4767 (N_4767,N_2585,N_939);
nor U4768 (N_4768,N_2897,N_3404);
xor U4769 (N_4769,N_2108,N_2354);
and U4770 (N_4770,N_2363,N_1834);
and U4771 (N_4771,N_2502,N_2867);
nand U4772 (N_4772,N_1764,N_58);
nor U4773 (N_4773,N_629,N_2053);
nor U4774 (N_4774,N_3849,N_70);
and U4775 (N_4775,N_2125,N_3058);
nor U4776 (N_4776,N_952,N_784);
and U4777 (N_4777,N_2647,N_951);
or U4778 (N_4778,N_371,N_2171);
and U4779 (N_4779,N_613,N_543);
nand U4780 (N_4780,N_570,N_1516);
and U4781 (N_4781,N_3570,N_3505);
and U4782 (N_4782,N_2156,N_2842);
or U4783 (N_4783,N_701,N_3748);
or U4784 (N_4784,N_3165,N_1109);
or U4785 (N_4785,N_3932,N_1042);
and U4786 (N_4786,N_1273,N_622);
or U4787 (N_4787,N_3533,N_1598);
or U4788 (N_4788,N_3599,N_2929);
nand U4789 (N_4789,N_3263,N_336);
nand U4790 (N_4790,N_2044,N_2595);
nand U4791 (N_4791,N_1292,N_3045);
or U4792 (N_4792,N_1634,N_3752);
or U4793 (N_4793,N_1301,N_628);
or U4794 (N_4794,N_735,N_1303);
or U4795 (N_4795,N_168,N_3234);
nor U4796 (N_4796,N_219,N_3486);
xnor U4797 (N_4797,N_3148,N_319);
and U4798 (N_4798,N_1703,N_2655);
or U4799 (N_4799,N_2725,N_3716);
or U4800 (N_4800,N_1632,N_2416);
nor U4801 (N_4801,N_1121,N_1455);
xnor U4802 (N_4802,N_1120,N_3232);
and U4803 (N_4803,N_501,N_1738);
or U4804 (N_4804,N_1097,N_1034);
xor U4805 (N_4805,N_872,N_580);
nand U4806 (N_4806,N_1600,N_3435);
nand U4807 (N_4807,N_1988,N_1370);
nand U4808 (N_4808,N_2441,N_2583);
and U4809 (N_4809,N_1721,N_1488);
or U4810 (N_4810,N_2041,N_3272);
and U4811 (N_4811,N_71,N_665);
or U4812 (N_4812,N_2201,N_1409);
nand U4813 (N_4813,N_3216,N_1850);
nand U4814 (N_4814,N_3112,N_576);
nor U4815 (N_4815,N_3377,N_922);
and U4816 (N_4816,N_2982,N_1613);
nand U4817 (N_4817,N_1017,N_3108);
or U4818 (N_4818,N_115,N_955);
nand U4819 (N_4819,N_3640,N_2745);
nand U4820 (N_4820,N_1079,N_2539);
and U4821 (N_4821,N_1283,N_2575);
nand U4822 (N_4822,N_1989,N_1642);
and U4823 (N_4823,N_263,N_476);
or U4824 (N_4824,N_2866,N_1971);
nor U4825 (N_4825,N_2915,N_2367);
or U4826 (N_4826,N_351,N_3846);
or U4827 (N_4827,N_1757,N_1708);
or U4828 (N_4828,N_3151,N_2473);
nand U4829 (N_4829,N_2353,N_3192);
nand U4830 (N_4830,N_2828,N_2685);
and U4831 (N_4831,N_1631,N_751);
or U4832 (N_4832,N_3161,N_3018);
nor U4833 (N_4833,N_2773,N_2758);
nor U4834 (N_4834,N_1312,N_2110);
and U4835 (N_4835,N_1678,N_591);
or U4836 (N_4836,N_3950,N_75);
nand U4837 (N_4837,N_377,N_244);
and U4838 (N_4838,N_2696,N_2097);
or U4839 (N_4839,N_1265,N_255);
nor U4840 (N_4840,N_1745,N_797);
xnor U4841 (N_4841,N_3313,N_2811);
and U4842 (N_4842,N_465,N_2256);
nand U4843 (N_4843,N_3199,N_1380);
xnor U4844 (N_4844,N_531,N_1247);
nand U4845 (N_4845,N_1712,N_702);
or U4846 (N_4846,N_3239,N_603);
nand U4847 (N_4847,N_3631,N_2131);
and U4848 (N_4848,N_3803,N_572);
xnor U4849 (N_4849,N_2118,N_231);
and U4850 (N_4850,N_2516,N_1851);
nand U4851 (N_4851,N_509,N_2508);
nor U4852 (N_4852,N_1263,N_2401);
and U4853 (N_4853,N_1956,N_1417);
nand U4854 (N_4854,N_3130,N_2426);
nor U4855 (N_4855,N_783,N_895);
nand U4856 (N_4856,N_137,N_49);
or U4857 (N_4857,N_253,N_2588);
or U4858 (N_4858,N_658,N_487);
nand U4859 (N_4859,N_346,N_1969);
or U4860 (N_4860,N_2657,N_380);
xnor U4861 (N_4861,N_2645,N_1293);
nor U4862 (N_4862,N_3506,N_376);
and U4863 (N_4863,N_2200,N_1976);
nor U4864 (N_4864,N_1475,N_563);
and U4865 (N_4865,N_3619,N_3564);
nor U4866 (N_4866,N_3200,N_2271);
nand U4867 (N_4867,N_1060,N_34);
and U4868 (N_4868,N_2558,N_3476);
nand U4869 (N_4869,N_3966,N_1680);
nor U4870 (N_4870,N_161,N_717);
and U4871 (N_4871,N_3210,N_2463);
xnor U4872 (N_4872,N_1622,N_2670);
and U4873 (N_4873,N_3568,N_699);
or U4874 (N_4874,N_3346,N_2141);
or U4875 (N_4875,N_3626,N_2333);
nand U4876 (N_4876,N_1800,N_3764);
or U4877 (N_4877,N_1912,N_3656);
nand U4878 (N_4878,N_3562,N_2050);
and U4879 (N_4879,N_3538,N_1925);
and U4880 (N_4880,N_941,N_521);
or U4881 (N_4881,N_1808,N_160);
nand U4882 (N_4882,N_2789,N_1332);
or U4883 (N_4883,N_347,N_2478);
nor U4884 (N_4884,N_3883,N_2067);
and U4885 (N_4885,N_68,N_2231);
nor U4886 (N_4886,N_901,N_1580);
or U4887 (N_4887,N_1318,N_2295);
xor U4888 (N_4888,N_313,N_2011);
or U4889 (N_4889,N_2943,N_352);
nor U4890 (N_4890,N_1262,N_1785);
nor U4891 (N_4891,N_826,N_619);
or U4892 (N_4892,N_820,N_796);
or U4893 (N_4893,N_800,N_315);
and U4894 (N_4894,N_725,N_204);
and U4895 (N_4895,N_2782,N_2134);
and U4896 (N_4896,N_849,N_1026);
nor U4897 (N_4897,N_1151,N_2265);
nor U4898 (N_4898,N_3356,N_97);
xor U4899 (N_4899,N_450,N_944);
nor U4900 (N_4900,N_1790,N_1198);
xor U4901 (N_4901,N_3028,N_1436);
or U4902 (N_4902,N_3780,N_158);
and U4903 (N_4903,N_3994,N_2380);
xnor U4904 (N_4904,N_1835,N_2743);
nand U4905 (N_4905,N_1719,N_2571);
nor U4906 (N_4906,N_873,N_2749);
nand U4907 (N_4907,N_687,N_1298);
xor U4908 (N_4908,N_2418,N_606);
or U4909 (N_4909,N_182,N_3817);
or U4910 (N_4910,N_337,N_150);
or U4911 (N_4911,N_2296,N_1487);
nor U4912 (N_4912,N_2527,N_2549);
and U4913 (N_4913,N_2003,N_903);
nor U4914 (N_4914,N_402,N_1508);
xnor U4915 (N_4915,N_2058,N_523);
or U4916 (N_4916,N_3387,N_1882);
nand U4917 (N_4917,N_1049,N_400);
xnor U4918 (N_4918,N_2285,N_3006);
xnor U4919 (N_4919,N_2991,N_25);
nor U4920 (N_4920,N_3259,N_2898);
nor U4921 (N_4921,N_605,N_799);
xnor U4922 (N_4922,N_568,N_583);
and U4923 (N_4923,N_2846,N_3684);
xnor U4924 (N_4924,N_2956,N_968);
or U4925 (N_4925,N_2005,N_2616);
nand U4926 (N_4926,N_1914,N_2474);
nor U4927 (N_4927,N_3819,N_420);
xor U4928 (N_4928,N_2325,N_2127);
or U4929 (N_4929,N_243,N_630);
nand U4930 (N_4930,N_2975,N_2159);
nor U4931 (N_4931,N_3298,N_2693);
or U4932 (N_4932,N_1530,N_3357);
and U4933 (N_4933,N_200,N_3880);
or U4934 (N_4934,N_2369,N_3119);
nor U4935 (N_4935,N_716,N_1858);
and U4936 (N_4936,N_746,N_713);
nor U4937 (N_4937,N_1285,N_3109);
xnor U4938 (N_4938,N_3173,N_3340);
nand U4939 (N_4939,N_1110,N_1962);
and U4940 (N_4940,N_3695,N_133);
nor U4941 (N_4941,N_194,N_1141);
xor U4942 (N_4942,N_2651,N_1006);
nor U4943 (N_4943,N_353,N_846);
nand U4944 (N_4944,N_801,N_129);
nor U4945 (N_4945,N_668,N_3220);
or U4946 (N_4946,N_3869,N_1253);
xnor U4947 (N_4947,N_43,N_12);
nand U4948 (N_4948,N_3589,N_2431);
nor U4949 (N_4949,N_366,N_3241);
xnor U4950 (N_4950,N_1570,N_252);
nand U4951 (N_4951,N_2654,N_1122);
or U4952 (N_4952,N_1257,N_2626);
nand U4953 (N_4953,N_1044,N_3826);
or U4954 (N_4954,N_2646,N_977);
nand U4955 (N_4955,N_2668,N_870);
nor U4956 (N_4956,N_3688,N_647);
nor U4957 (N_4957,N_151,N_660);
nor U4958 (N_4958,N_640,N_1223);
nor U4959 (N_4959,N_2451,N_3727);
nor U4960 (N_4960,N_878,N_3693);
or U4961 (N_4961,N_2373,N_2519);
or U4962 (N_4962,N_765,N_1085);
or U4963 (N_4963,N_1077,N_1274);
nor U4964 (N_4964,N_1463,N_3930);
or U4965 (N_4965,N_525,N_3106);
nor U4966 (N_4966,N_2781,N_3074);
nor U4967 (N_4967,N_2241,N_3691);
nor U4968 (N_4968,N_1933,N_894);
nor U4969 (N_4969,N_3981,N_3709);
or U4970 (N_4970,N_3697,N_2364);
nor U4971 (N_4971,N_1433,N_1415);
nand U4972 (N_4972,N_2132,N_2968);
and U4973 (N_4973,N_2734,N_819);
or U4974 (N_4974,N_2239,N_230);
nand U4975 (N_4975,N_432,N_1002);
nor U4976 (N_4976,N_3554,N_959);
nor U4977 (N_4977,N_3327,N_1607);
or U4978 (N_4978,N_1650,N_919);
nand U4979 (N_4979,N_3179,N_3482);
nand U4980 (N_4980,N_3153,N_2799);
nand U4981 (N_4981,N_2567,N_656);
nor U4982 (N_4982,N_761,N_729);
nand U4983 (N_4983,N_3905,N_3603);
or U4984 (N_4984,N_561,N_2821);
and U4985 (N_4985,N_2776,N_2242);
nand U4986 (N_4986,N_3343,N_327);
nand U4987 (N_4987,N_484,N_3248);
and U4988 (N_4988,N_2505,N_1849);
nand U4989 (N_4989,N_22,N_2453);
nand U4990 (N_4990,N_3054,N_1407);
nand U4991 (N_4991,N_3682,N_696);
nor U4992 (N_4992,N_1652,N_2613);
and U4993 (N_4993,N_3766,N_1922);
or U4994 (N_4994,N_1210,N_2288);
nor U4995 (N_4995,N_2334,N_3437);
nand U4996 (N_4996,N_461,N_1950);
nand U4997 (N_4997,N_3041,N_329);
nand U4998 (N_4998,N_3828,N_268);
xor U4999 (N_4999,N_844,N_3983);
nand U5000 (N_5000,N_2623,N_128);
and U5001 (N_5001,N_1887,N_780);
nor U5002 (N_5002,N_1639,N_1270);
or U5003 (N_5003,N_246,N_3519);
and U5004 (N_5004,N_3768,N_1554);
nand U5005 (N_5005,N_991,N_1500);
nor U5006 (N_5006,N_1326,N_2969);
nor U5007 (N_5007,N_602,N_2425);
or U5008 (N_5008,N_566,N_122);
nand U5009 (N_5009,N_6,N_970);
or U5010 (N_5010,N_385,N_378);
xor U5011 (N_5011,N_2935,N_2919);
nand U5012 (N_5012,N_3635,N_1732);
nor U5013 (N_5013,N_3972,N_2138);
xnor U5014 (N_5014,N_271,N_2950);
nand U5015 (N_5015,N_601,N_3344);
or U5016 (N_5016,N_3588,N_2598);
nor U5017 (N_5017,N_2158,N_3172);
xnor U5018 (N_5018,N_1199,N_1391);
xor U5019 (N_5019,N_3333,N_3911);
and U5020 (N_5020,N_427,N_2545);
nor U5021 (N_5021,N_2847,N_2861);
nor U5022 (N_5022,N_2198,N_2772);
nand U5023 (N_5023,N_2775,N_3898);
or U5024 (N_5024,N_1381,N_2806);
or U5025 (N_5025,N_3801,N_2388);
nand U5026 (N_5026,N_1237,N_842);
and U5027 (N_5027,N_1752,N_2863);
xnor U5028 (N_5028,N_1124,N_3685);
nand U5029 (N_5029,N_518,N_237);
or U5030 (N_5030,N_2774,N_1033);
or U5031 (N_5031,N_792,N_1242);
nand U5032 (N_5032,N_3596,N_564);
and U5033 (N_5033,N_1791,N_3854);
and U5034 (N_5034,N_2202,N_2820);
xor U5035 (N_5035,N_140,N_2455);
and U5036 (N_5036,N_2640,N_3615);
nand U5037 (N_5037,N_2282,N_3649);
and U5038 (N_5038,N_723,N_2409);
nor U5039 (N_5039,N_3731,N_3026);
and U5040 (N_5040,N_3055,N_2448);
nand U5041 (N_5041,N_1514,N_1093);
and U5042 (N_5042,N_3479,N_1937);
and U5043 (N_5043,N_1224,N_1555);
nor U5044 (N_5044,N_460,N_2276);
nand U5045 (N_5045,N_3530,N_1695);
nor U5046 (N_5046,N_3341,N_1359);
or U5047 (N_5047,N_3456,N_470);
and U5048 (N_5048,N_374,N_3253);
and U5049 (N_5049,N_2437,N_2996);
and U5050 (N_5050,N_1333,N_2858);
nor U5051 (N_5051,N_1045,N_3837);
or U5052 (N_5052,N_971,N_664);
xor U5053 (N_5053,N_841,N_2801);
nor U5054 (N_5054,N_3214,N_267);
or U5055 (N_5055,N_339,N_83);
nor U5056 (N_5056,N_1337,N_2941);
nor U5057 (N_5057,N_23,N_3870);
nor U5058 (N_5058,N_710,N_972);
nor U5059 (N_5059,N_1377,N_1204);
or U5060 (N_5060,N_2064,N_3662);
nor U5061 (N_5061,N_1637,N_1884);
nand U5062 (N_5062,N_3938,N_1356);
xor U5063 (N_5063,N_1386,N_1819);
and U5064 (N_5064,N_2240,N_669);
nor U5065 (N_5065,N_1156,N_2763);
xnor U5066 (N_5066,N_3952,N_690);
nand U5067 (N_5067,N_3601,N_2604);
or U5068 (N_5068,N_2449,N_1838);
nand U5069 (N_5069,N_216,N_2142);
nor U5070 (N_5070,N_2018,N_2227);
or U5071 (N_5071,N_94,N_3420);
nor U5072 (N_5072,N_2059,N_1694);
nand U5073 (N_5073,N_1341,N_3742);
nand U5074 (N_5074,N_2490,N_1801);
and U5075 (N_5075,N_3733,N_259);
and U5076 (N_5076,N_2457,N_2327);
nor U5077 (N_5077,N_3840,N_633);
nand U5078 (N_5078,N_3238,N_1953);
or U5079 (N_5079,N_110,N_1899);
nand U5080 (N_5080,N_1911,N_805);
xor U5081 (N_5081,N_2710,N_586);
and U5082 (N_5082,N_489,N_2383);
nand U5083 (N_5083,N_2599,N_1361);
nand U5084 (N_5084,N_3671,N_845);
nor U5085 (N_5085,N_2381,N_3330);
or U5086 (N_5086,N_236,N_3081);
and U5087 (N_5087,N_1960,N_3961);
or U5088 (N_5088,N_724,N_3990);
and U5089 (N_5089,N_3916,N_142);
nor U5090 (N_5090,N_2908,N_2958);
nor U5091 (N_5091,N_1660,N_2214);
or U5092 (N_5092,N_2756,N_245);
nor U5093 (N_5093,N_15,N_2630);
xnor U5094 (N_5094,N_3673,N_1347);
or U5095 (N_5095,N_1551,N_513);
xor U5096 (N_5096,N_1794,N_1354);
and U5097 (N_5097,N_1360,N_812);
or U5098 (N_5098,N_431,N_998);
or U5099 (N_5099,N_1998,N_614);
and U5100 (N_5100,N_3539,N_1685);
xnor U5101 (N_5101,N_196,N_2250);
nor U5102 (N_5102,N_1928,N_3755);
or U5103 (N_5103,N_3359,N_391);
nand U5104 (N_5104,N_394,N_3375);
nor U5105 (N_5105,N_2557,N_382);
or U5106 (N_5106,N_2707,N_2804);
and U5107 (N_5107,N_550,N_2548);
or U5108 (N_5108,N_2389,N_3811);
xnor U5109 (N_5109,N_1827,N_1422);
nor U5110 (N_5110,N_3637,N_3577);
or U5111 (N_5111,N_707,N_2826);
or U5112 (N_5112,N_3207,N_2385);
or U5113 (N_5113,N_1684,N_1756);
nor U5114 (N_5114,N_1343,N_2180);
xor U5115 (N_5115,N_2714,N_3528);
nand U5116 (N_5116,N_3623,N_1251);
or U5117 (N_5117,N_91,N_2959);
xnor U5118 (N_5118,N_363,N_479);
xnor U5119 (N_5119,N_1623,N_532);
xnor U5120 (N_5120,N_1510,N_3786);
and U5121 (N_5121,N_2012,N_694);
and U5122 (N_5122,N_2894,N_2711);
xor U5123 (N_5123,N_1879,N_1011);
nor U5124 (N_5124,N_2515,N_715);
nor U5125 (N_5125,N_2620,N_2590);
nand U5126 (N_5126,N_2420,N_3586);
or U5127 (N_5127,N_2356,N_881);
and U5128 (N_5128,N_1036,N_644);
nor U5129 (N_5129,N_3049,N_1520);
xnor U5130 (N_5130,N_1842,N_1236);
nor U5131 (N_5131,N_869,N_2290);
or U5132 (N_5132,N_1556,N_2931);
or U5133 (N_5133,N_3524,N_1787);
xnor U5134 (N_5134,N_3914,N_2713);
nor U5135 (N_5135,N_3316,N_2317);
nor U5136 (N_5136,N_3193,N_1485);
nor U5137 (N_5137,N_2314,N_1098);
and U5138 (N_5138,N_109,N_2857);
or U5139 (N_5139,N_3319,N_3434);
and U5140 (N_5140,N_3300,N_2074);
and U5141 (N_5141,N_2851,N_2435);
or U5142 (N_5142,N_3504,N_859);
nand U5143 (N_5143,N_1698,N_1609);
nand U5144 (N_5144,N_468,N_3222);
nor U5145 (N_5145,N_3639,N_1804);
xnor U5146 (N_5146,N_1184,N_3609);
nand U5147 (N_5147,N_856,N_2702);
or U5148 (N_5148,N_2661,N_2850);
or U5149 (N_5149,N_205,N_372);
and U5150 (N_5150,N_2477,N_910);
or U5151 (N_5151,N_2664,N_2375);
nor U5152 (N_5152,N_2410,N_1005);
and U5153 (N_5153,N_3400,N_3498);
nor U5154 (N_5154,N_1659,N_2672);
and U5155 (N_5155,N_295,N_1240);
nand U5156 (N_5156,N_2901,N_3791);
xor U5157 (N_5157,N_333,N_149);
xor U5158 (N_5158,N_444,N_2308);
or U5159 (N_5159,N_2224,N_2143);
or U5160 (N_5160,N_1844,N_2614);
nor U5161 (N_5161,N_3899,N_529);
and U5162 (N_5162,N_1518,N_1466);
nor U5163 (N_5163,N_3266,N_2993);
nand U5164 (N_5164,N_3412,N_1126);
xnor U5165 (N_5165,N_2980,N_579);
nor U5166 (N_5166,N_3446,N_697);
nand U5167 (N_5167,N_1705,N_1441);
nor U5168 (N_5168,N_3183,N_3223);
nor U5169 (N_5169,N_875,N_98);
or U5170 (N_5170,N_516,N_2521);
nand U5171 (N_5171,N_745,N_3632);
or U5172 (N_5172,N_3634,N_1550);
nand U5173 (N_5173,N_57,N_667);
or U5174 (N_5174,N_3122,N_3910);
xnor U5175 (N_5175,N_2909,N_446);
and U5176 (N_5176,N_3977,N_755);
and U5177 (N_5177,N_1395,N_2650);
nand U5178 (N_5178,N_3382,N_891);
nand U5179 (N_5179,N_1692,N_2366);
and U5180 (N_5180,N_2722,N_3365);
nor U5181 (N_5181,N_2304,N_2116);
nor U5182 (N_5182,N_1195,N_3725);
nor U5183 (N_5183,N_3118,N_3714);
or U5184 (N_5184,N_2504,N_2015);
or U5185 (N_5185,N_537,N_1578);
or U5186 (N_5186,N_2399,N_827);
nand U5187 (N_5187,N_1701,N_2819);
or U5188 (N_5188,N_2080,N_3019);
nor U5189 (N_5189,N_1078,N_3720);
or U5190 (N_5190,N_99,N_3836);
nand U5191 (N_5191,N_3698,N_3795);
nor U5192 (N_5192,N_2060,N_3452);
nand U5193 (N_5193,N_727,N_1432);
xnor U5194 (N_5194,N_422,N_558);
or U5195 (N_5195,N_2160,N_1710);
nand U5196 (N_5196,N_2997,N_1515);
or U5197 (N_5197,N_1540,N_2382);
or U5198 (N_5198,N_3317,N_3171);
or U5199 (N_5199,N_2924,N_889);
and U5200 (N_5200,N_1086,N_426);
and U5201 (N_5201,N_2197,N_5);
nor U5202 (N_5202,N_3059,N_187);
nand U5203 (N_5203,N_250,N_1135);
nand U5204 (N_5204,N_1854,N_111);
nor U5205 (N_5205,N_3286,N_855);
nand U5206 (N_5206,N_1758,N_3942);
nor U5207 (N_5207,N_2596,N_2343);
xor U5208 (N_5208,N_3440,N_2113);
or U5209 (N_5209,N_3226,N_2796);
or U5210 (N_5210,N_3152,N_451);
and U5211 (N_5211,N_2951,N_42);
nand U5212 (N_5212,N_120,N_541);
nand U5213 (N_5213,N_837,N_458);
or U5214 (N_5214,N_1526,N_1490);
or U5215 (N_5215,N_3068,N_3707);
nor U5216 (N_5216,N_1709,N_1729);
and U5217 (N_5217,N_2277,N_3501);
nand U5218 (N_5218,N_1228,N_1594);
nand U5219 (N_5219,N_1159,N_1428);
nor U5220 (N_5220,N_2783,N_2976);
or U5221 (N_5221,N_1486,N_3995);
and U5222 (N_5222,N_2628,N_1456);
nand U5223 (N_5223,N_1945,N_1574);
nand U5224 (N_5224,N_3480,N_2815);
or U5225 (N_5225,N_2942,N_314);
nand U5226 (N_5226,N_607,N_1192);
and U5227 (N_5227,N_2677,N_3070);
nand U5228 (N_5228,N_2755,N_2880);
nand U5229 (N_5229,N_2701,N_3906);
xor U5230 (N_5230,N_1507,N_2148);
nand U5231 (N_5231,N_2024,N_2949);
nand U5232 (N_5232,N_1646,N_442);
and U5233 (N_5233,N_1069,N_2391);
nand U5234 (N_5234,N_1165,N_3403);
and U5235 (N_5235,N_261,N_1127);
and U5236 (N_5236,N_3973,N_3612);
nand U5237 (N_5237,N_2807,N_2338);
and U5238 (N_5238,N_3878,N_1144);
nor U5239 (N_5239,N_704,N_3281);
and U5240 (N_5240,N_3013,N_767);
and U5241 (N_5241,N_984,N_2223);
nor U5242 (N_5242,N_1857,N_2540);
and U5243 (N_5243,N_932,N_2147);
nor U5244 (N_5244,N_1206,N_573);
nor U5245 (N_5245,N_1268,N_1672);
nor U5246 (N_5246,N_388,N_990);
nor U5247 (N_5247,N_2536,N_904);
or U5248 (N_5248,N_1802,N_3522);
xor U5249 (N_5249,N_1651,N_1495);
nor U5250 (N_5250,N_2565,N_2797);
nand U5251 (N_5251,N_335,N_2609);
nor U5252 (N_5252,N_248,N_3462);
and U5253 (N_5253,N_1866,N_296);
nand U5254 (N_5254,N_2076,N_176);
or U5255 (N_5255,N_3686,N_902);
nand U5256 (N_5256,N_2103,N_3997);
and U5257 (N_5257,N_409,N_2365);
xor U5258 (N_5258,N_3900,N_3529);
nand U5259 (N_5259,N_3881,N_3598);
nor U5260 (N_5260,N_2179,N_911);
or U5261 (N_5261,N_2123,N_2622);
and U5262 (N_5262,N_3877,N_3988);
nand U5263 (N_5263,N_719,N_522);
or U5264 (N_5264,N_847,N_3617);
nand U5265 (N_5265,N_3765,N_1010);
xnor U5266 (N_5266,N_921,N_2852);
or U5267 (N_5267,N_2617,N_3982);
or U5268 (N_5268,N_1714,N_2278);
or U5269 (N_5269,N_2037,N_1139);
or U5270 (N_5270,N_1216,N_1430);
nor U5271 (N_5271,N_1254,N_2215);
nand U5272 (N_5272,N_3618,N_3909);
nor U5273 (N_5273,N_1905,N_1581);
nand U5274 (N_5274,N_3888,N_1771);
nor U5275 (N_5275,N_3761,N_2900);
nor U5276 (N_5276,N_2124,N_1503);
or U5277 (N_5277,N_736,N_2860);
xnor U5278 (N_5278,N_2669,N_1788);
nand U5279 (N_5279,N_3773,N_232);
nand U5280 (N_5280,N_1448,N_3056);
xnor U5281 (N_5281,N_811,N_2396);
and U5282 (N_5282,N_2718,N_1423);
nand U5283 (N_5283,N_1451,N_3692);
or U5284 (N_5284,N_1399,N_2706);
xnor U5285 (N_5285,N_3030,N_758);
or U5286 (N_5286,N_2289,N_1071);
and U5287 (N_5287,N_1012,N_1261);
nand U5288 (N_5288,N_703,N_929);
nand U5289 (N_5289,N_2608,N_2117);
nor U5290 (N_5290,N_3423,N_928);
nor U5291 (N_5291,N_2922,N_1186);
nand U5292 (N_5292,N_3302,N_3038);
nor U5293 (N_5293,N_179,N_3991);
and U5294 (N_5294,N_2417,N_239);
or U5295 (N_5295,N_539,N_2408);
and U5296 (N_5296,N_3464,N_1881);
xor U5297 (N_5297,N_257,N_867);
nand U5298 (N_5298,N_1464,N_1183);
and U5299 (N_5299,N_14,N_3170);
nor U5300 (N_5300,N_1793,N_3575);
nor U5301 (N_5301,N_3919,N_0);
nor U5302 (N_5302,N_1674,N_3680);
or U5303 (N_5303,N_2873,N_1967);
and U5304 (N_5304,N_2371,N_676);
or U5305 (N_5305,N_38,N_852);
xnor U5306 (N_5306,N_1096,N_1025);
or U5307 (N_5307,N_1513,N_279);
or U5308 (N_5308,N_1450,N_3177);
or U5309 (N_5309,N_1336,N_3110);
or U5310 (N_5310,N_2784,N_421);
and U5311 (N_5311,N_3396,N_3256);
or U5312 (N_5312,N_1670,N_256);
and U5313 (N_5313,N_2438,N_2566);
or U5314 (N_5314,N_3406,N_2537);
and U5315 (N_5315,N_82,N_3229);
or U5316 (N_5316,N_3432,N_2165);
xnor U5317 (N_5317,N_2046,N_2346);
nand U5318 (N_5318,N_1477,N_1445);
or U5319 (N_5319,N_2222,N_1175);
or U5320 (N_5320,N_1880,N_2708);
nand U5321 (N_5321,N_1667,N_2780);
nand U5322 (N_5322,N_2281,N_1744);
and U5323 (N_5323,N_2026,N_1797);
and U5324 (N_5324,N_641,N_355);
nor U5325 (N_5325,N_3737,N_2930);
nor U5326 (N_5326,N_143,N_3611);
nand U5327 (N_5327,N_3466,N_1625);
nor U5328 (N_5328,N_734,N_1276);
nand U5329 (N_5329,N_1784,N_2902);
nand U5330 (N_5330,N_325,N_1662);
nor U5331 (N_5331,N_3920,N_912);
nor U5332 (N_5332,N_3908,N_3576);
nand U5333 (N_5333,N_604,N_874);
xor U5334 (N_5334,N_2164,N_2928);
or U5335 (N_5335,N_1934,N_1136);
nand U5336 (N_5336,N_13,N_2261);
nor U5337 (N_5337,N_786,N_3648);
nand U5338 (N_5338,N_1606,N_1173);
nor U5339 (N_5339,N_67,N_407);
or U5340 (N_5340,N_3629,N_130);
nor U5341 (N_5341,N_1390,N_2859);
xnor U5342 (N_5342,N_2584,N_1384);
nand U5343 (N_5343,N_2009,N_197);
and U5344 (N_5344,N_1062,N_1187);
nand U5345 (N_5345,N_2896,N_2101);
nand U5346 (N_5346,N_3348,N_502);
or U5347 (N_5347,N_2195,N_2398);
nor U5348 (N_5348,N_2513,N_3211);
nand U5349 (N_5349,N_387,N_118);
and U5350 (N_5350,N_3037,N_1493);
or U5351 (N_5351,N_3174,N_2986);
or U5352 (N_5352,N_186,N_2638);
or U5353 (N_5353,N_317,N_588);
and U5354 (N_5354,N_2994,N_452);
nand U5355 (N_5355,N_1704,N_3299);
or U5356 (N_5356,N_1724,N_1047);
nor U5357 (N_5357,N_2581,N_2248);
nand U5358 (N_5358,N_1523,N_949);
or U5359 (N_5359,N_2535,N_2964);
nand U5360 (N_5360,N_2055,N_1278);
and U5361 (N_5361,N_3683,N_3005);
or U5362 (N_5362,N_2542,N_153);
nor U5363 (N_5363,N_373,N_1929);
or U5364 (N_5364,N_3743,N_2456);
or U5365 (N_5365,N_293,N_1351);
and U5366 (N_5366,N_1171,N_2345);
nor U5367 (N_5367,N_575,N_1519);
nor U5368 (N_5368,N_3833,N_2051);
and U5369 (N_5369,N_2298,N_2332);
nand U5370 (N_5370,N_1792,N_1781);
nand U5371 (N_5371,N_1244,N_1572);
or U5372 (N_5372,N_395,N_1763);
and U5373 (N_5373,N_1717,N_1773);
and U5374 (N_5374,N_1309,N_885);
and U5375 (N_5375,N_1322,N_1560);
nand U5376 (N_5376,N_2114,N_1583);
xnor U5377 (N_5377,N_1829,N_1090);
and U5378 (N_5378,N_276,N_1032);
nor U5379 (N_5379,N_328,N_209);
or U5380 (N_5380,N_3853,N_2512);
or U5381 (N_5381,N_1533,N_551);
nand U5382 (N_5382,N_3822,N_1114);
and U5383 (N_5383,N_3104,N_788);
xnor U5384 (N_5384,N_918,N_1148);
or U5385 (N_5385,N_1193,N_3933);
and U5386 (N_5386,N_3303,N_675);
or U5387 (N_5387,N_1527,N_915);
and U5388 (N_5388,N_3770,N_3138);
nand U5389 (N_5389,N_1214,N_3276);
and U5390 (N_5390,N_2001,N_1638);
nor U5391 (N_5391,N_3875,N_1935);
nor U5392 (N_5392,N_1548,N_1534);
nor U5393 (N_5393,N_1020,N_1972);
nor U5394 (N_5394,N_2466,N_3475);
nand U5395 (N_5395,N_562,N_2779);
nor U5396 (N_5396,N_2735,N_1870);
and U5397 (N_5397,N_3127,N_1999);
and U5398 (N_5398,N_3408,N_2442);
or U5399 (N_5399,N_3514,N_1735);
and U5400 (N_5400,N_963,N_1393);
nand U5401 (N_5401,N_3959,N_1964);
and U5402 (N_5402,N_1102,N_1775);
and U5403 (N_5403,N_210,N_817);
and U5404 (N_5404,N_2790,N_425);
or U5405 (N_5405,N_3729,N_1321);
and U5406 (N_5406,N_3924,N_324);
and U5407 (N_5407,N_2422,N_1161);
xnor U5408 (N_5408,N_2927,N_119);
or U5409 (N_5409,N_3555,N_2189);
nor U5410 (N_5410,N_3078,N_3180);
and U5411 (N_5411,N_876,N_1837);
nor U5412 (N_5412,N_1104,N_3410);
nand U5413 (N_5413,N_2483,N_3989);
and U5414 (N_5414,N_1059,N_2087);
nor U5415 (N_5415,N_3036,N_1902);
nor U5416 (N_5416,N_2186,N_2460);
xor U5417 (N_5417,N_1365,N_3353);
nor U5418 (N_5418,N_175,N_2767);
nor U5419 (N_5419,N_299,N_3062);
nand U5420 (N_5420,N_2591,N_40);
nor U5421 (N_5421,N_2698,N_3043);
nor U5422 (N_5422,N_1628,N_3654);
nor U5423 (N_5423,N_3502,N_3411);
xnor U5424 (N_5424,N_1258,N_1886);
or U5425 (N_5425,N_2684,N_1056);
and U5426 (N_5426,N_776,N_397);
or U5427 (N_5427,N_260,N_589);
and U5428 (N_5428,N_2421,N_3812);
or U5429 (N_5429,N_907,N_3581);
nor U5430 (N_5430,N_8,N_1382);
or U5431 (N_5431,N_1629,N_2962);
nor U5432 (N_5432,N_1871,N_1799);
xnor U5433 (N_5433,N_711,N_1462);
nand U5434 (N_5434,N_3851,N_506);
and U5435 (N_5435,N_3409,N_2393);
and U5436 (N_5436,N_270,N_258);
or U5437 (N_5437,N_3621,N_747);
or U5438 (N_5438,N_1700,N_1535);
and U5439 (N_5439,N_608,N_2785);
nand U5440 (N_5440,N_1740,N_3093);
nand U5441 (N_5441,N_2273,N_1482);
nand U5442 (N_5442,N_2689,N_3963);
or U5443 (N_5443,N_3594,N_2404);
nor U5444 (N_5444,N_540,N_1859);
nor U5445 (N_5445,N_3,N_454);
and U5446 (N_5446,N_2070,N_3754);
and U5447 (N_5447,N_2572,N_1465);
nor U5448 (N_5448,N_3527,N_1340);
or U5449 (N_5449,N_748,N_235);
nor U5450 (N_5450,N_2212,N_289);
nor U5451 (N_5451,N_2753,N_365);
nor U5452 (N_5452,N_806,N_3493);
and U5453 (N_5453,N_1196,N_974);
nand U5454 (N_5454,N_2392,N_466);
nor U5455 (N_5455,N_2166,N_462);
and U5456 (N_5456,N_1189,N_3191);
nor U5457 (N_5457,N_766,N_778);
or U5458 (N_5458,N_369,N_3471);
nor U5459 (N_5459,N_316,N_27);
or U5460 (N_5460,N_2484,N_2038);
nor U5461 (N_5461,N_2871,N_392);
and U5462 (N_5462,N_298,N_2403);
xnor U5463 (N_5463,N_3779,N_2321);
xor U5464 (N_5464,N_2275,N_2977);
xor U5465 (N_5465,N_1753,N_2027);
and U5466 (N_5466,N_3992,N_3376);
xnor U5467 (N_5467,N_2052,N_1000);
xnor U5468 (N_5468,N_1828,N_3240);
or U5469 (N_5469,N_791,N_1979);
nor U5470 (N_5470,N_1602,N_3985);
nor U5471 (N_5471,N_3358,N_814);
or U5472 (N_5472,N_3342,N_3572);
and U5473 (N_5473,N_2377,N_383);
and U5474 (N_5474,N_3140,N_3856);
or U5475 (N_5475,N_3700,N_999);
nand U5476 (N_5476,N_1517,N_360);
xnor U5477 (N_5477,N_530,N_2090);
xor U5478 (N_5478,N_2881,N_3622);
nand U5479 (N_5479,N_1923,N_2547);
xor U5480 (N_5480,N_858,N_1324);
nor U5481 (N_5481,N_3379,N_3267);
nand U5482 (N_5482,N_2666,N_2865);
or U5483 (N_5483,N_2226,N_2259);
nand U5484 (N_5484,N_3100,N_2744);
nor U5485 (N_5485,N_1128,N_359);
or U5486 (N_5486,N_1592,N_1591);
nor U5487 (N_5487,N_997,N_3126);
nand U5488 (N_5488,N_1376,N_3962);
xnor U5489 (N_5489,N_1986,N_1250);
nor U5490 (N_5490,N_1722,N_1355);
and U5491 (N_5491,N_3390,N_241);
nand U5492 (N_5492,N_2330,N_3268);
nor U5493 (N_5493,N_2509,N_598);
and U5494 (N_5494,N_2678,N_2844);
or U5495 (N_5495,N_3261,N_1931);
nor U5496 (N_5496,N_2963,N_623);
xor U5497 (N_5497,N_254,N_1512);
and U5498 (N_5498,N_3655,N_435);
and U5499 (N_5499,N_2462,N_2520);
nor U5500 (N_5500,N_93,N_712);
and U5501 (N_5501,N_2181,N_3559);
nor U5502 (N_5502,N_3608,N_3425);
nand U5503 (N_5503,N_909,N_434);
and U5504 (N_5504,N_2495,N_1473);
xnor U5505 (N_5505,N_20,N_1643);
nand U5506 (N_5506,N_1562,N_3585);
nand U5507 (N_5507,N_96,N_1509);
or U5508 (N_5508,N_2827,N_1815);
nor U5509 (N_5509,N_2434,N_3876);
or U5510 (N_5510,N_618,N_195);
nand U5511 (N_5511,N_2255,N_265);
nor U5512 (N_5512,N_1230,N_2800);
and U5513 (N_5513,N_1252,N_900);
or U5514 (N_5514,N_73,N_104);
or U5515 (N_5515,N_2092,N_3964);
and U5516 (N_5516,N_1373,N_1975);
or U5517 (N_5517,N_443,N_2971);
nor U5518 (N_5518,N_3510,N_3578);
nand U5519 (N_5519,N_3115,N_1633);
nor U5520 (N_5520,N_3290,N_2586);
or U5521 (N_5521,N_2786,N_2787);
nand U5522 (N_5522,N_47,N_2091);
xnor U5523 (N_5523,N_1621,N_3557);
and U5524 (N_5524,N_440,N_3730);
nand U5525 (N_5525,N_2313,N_2932);
and U5526 (N_5526,N_3633,N_1496);
or U5527 (N_5527,N_127,N_1368);
nor U5528 (N_5528,N_1416,N_1875);
and U5529 (N_5529,N_1438,N_2232);
and U5530 (N_5530,N_678,N_1693);
nand U5531 (N_5531,N_1681,N_3320);
nor U5532 (N_5532,N_3657,N_3593);
xnor U5533 (N_5533,N_1289,N_621);
or U5534 (N_5534,N_1994,N_1668);
or U5535 (N_5535,N_1038,N_1906);
and U5536 (N_5536,N_1921,N_2699);
and U5537 (N_5537,N_2868,N_3401);
nor U5538 (N_5538,N_1816,N_947);
nor U5539 (N_5539,N_3255,N_3679);
and U5540 (N_5540,N_2167,N_1304);
or U5541 (N_5541,N_3536,N_3378);
or U5542 (N_5542,N_1142,N_1037);
xor U5543 (N_5543,N_3939,N_1611);
nand U5544 (N_5544,N_166,N_2656);
nand U5545 (N_5545,N_3467,N_2593);
nor U5546 (N_5546,N_1389,N_180);
nand U5547 (N_5547,N_3029,N_3818);
nor U5548 (N_5548,N_3447,N_273);
and U5549 (N_5549,N_3951,N_853);
nor U5550 (N_5550,N_1892,N_447);
xor U5551 (N_5551,N_2564,N_2899);
or U5552 (N_5552,N_16,N_2889);
nor U5553 (N_5553,N_3521,N_2762);
nor U5554 (N_5554,N_1563,N_3847);
and U5555 (N_5555,N_2068,N_1282);
nand U5556 (N_5556,N_1630,N_3369);
or U5557 (N_5557,N_1697,N_3150);
nand U5558 (N_5558,N_1055,N_1760);
or U5559 (N_5559,N_2916,N_1531);
xnor U5560 (N_5560,N_3331,N_2229);
nand U5561 (N_5561,N_2305,N_3747);
and U5562 (N_5562,N_1618,N_1397);
and U5563 (N_5563,N_2063,N_807);
nand U5564 (N_5564,N_3484,N_1734);
and U5565 (N_5565,N_862,N_3735);
or U5566 (N_5566,N_1014,N_958);
nand U5567 (N_5567,N_610,N_3563);
nand U5568 (N_5568,N_560,N_617);
nand U5569 (N_5569,N_3794,N_1040);
nand U5570 (N_5570,N_1342,N_627);
or U5571 (N_5571,N_1452,N_453);
nor U5572 (N_5572,N_1730,N_2066);
or U5573 (N_5573,N_288,N_1970);
or U5574 (N_5574,N_1741,N_294);
nand U5575 (N_5575,N_1172,N_2489);
or U5576 (N_5576,N_2045,N_1649);
xnor U5577 (N_5577,N_1736,N_145);
or U5578 (N_5578,N_2817,N_983);
nor U5579 (N_5579,N_3571,N_3638);
nand U5580 (N_5580,N_2084,N_202);
nand U5581 (N_5581,N_3244,N_1181);
nor U5582 (N_5582,N_157,N_3787);
nor U5583 (N_5583,N_655,N_1094);
or U5584 (N_5584,N_92,N_1811);
nor U5585 (N_5585,N_3491,N_3746);
or U5586 (N_5586,N_1645,N_2878);
nand U5587 (N_5587,N_3202,N_396);
xor U5588 (N_5588,N_323,N_692);
nor U5589 (N_5589,N_933,N_1295);
nor U5590 (N_5590,N_2911,N_21);
xnor U5591 (N_5591,N_3449,N_2253);
nand U5592 (N_5592,N_654,N_2267);
and U5593 (N_5593,N_3957,N_3934);
nor U5594 (N_5594,N_1861,N_3515);
nor U5595 (N_5595,N_877,N_1718);
or U5596 (N_5596,N_90,N_3063);
xor U5597 (N_5597,N_2692,N_1993);
or U5598 (N_5598,N_743,N_2208);
and U5599 (N_5599,N_1190,N_1676);
and U5600 (N_5600,N_1726,N_3715);
and U5601 (N_5601,N_1131,N_2848);
and U5602 (N_5602,N_3873,N_2809);
nand U5603 (N_5603,N_1542,N_332);
nor U5604 (N_5604,N_2974,N_1080);
or U5605 (N_5605,N_1614,N_1843);
xor U5606 (N_5606,N_1411,N_1648);
or U5607 (N_5607,N_228,N_994);
or U5608 (N_5608,N_100,N_497);
nor U5609 (N_5609,N_1883,N_3325);
or U5610 (N_5610,N_769,N_3249);
nor U5611 (N_5611,N_1576,N_3047);
or U5612 (N_5612,N_3243,N_2217);
or U5613 (N_5613,N_2476,N_424);
and U5614 (N_5614,N_1501,N_1461);
nand U5615 (N_5615,N_3128,N_1472);
nand U5616 (N_5616,N_1406,N_1239);
nand U5617 (N_5617,N_1328,N_9);
or U5618 (N_5618,N_1836,N_3543);
nor U5619 (N_5619,N_3775,N_139);
nand U5620 (N_5620,N_1188,N_3197);
and U5621 (N_5621,N_3848,N_1201);
xor U5622 (N_5622,N_2269,N_2835);
or U5623 (N_5623,N_3922,N_379);
xnor U5624 (N_5624,N_1170,N_3960);
nor U5625 (N_5625,N_2597,N_2533);
or U5626 (N_5626,N_240,N_685);
nor U5627 (N_5627,N_1823,N_3728);
or U5628 (N_5628,N_2355,N_636);
or U5629 (N_5629,N_2017,N_340);
and U5630 (N_5630,N_3956,N_1366);
nand U5631 (N_5631,N_291,N_2839);
nand U5632 (N_5632,N_3781,N_3004);
xnor U5633 (N_5633,N_1108,N_1313);
nor U5634 (N_5634,N_2769,N_3537);
and U5635 (N_5635,N_1853,N_330);
nor U5636 (N_5636,N_3918,N_2580);
nand U5637 (N_5637,N_1939,N_3784);
and U5638 (N_5638,N_3065,N_666);
and U5639 (N_5639,N_1279,N_1300);
nand U5640 (N_5640,N_53,N_311);
nand U5641 (N_5641,N_833,N_177);
and U5642 (N_5642,N_1443,N_2402);
or U5643 (N_5643,N_199,N_574);
or U5644 (N_5644,N_1269,N_3541);
nand U5645 (N_5645,N_3215,N_3550);
nand U5646 (N_5646,N_2496,N_3800);
nor U5647 (N_5647,N_3015,N_1095);
nand U5648 (N_5648,N_207,N_3066);
or U5649 (N_5649,N_3221,N_3653);
nor U5650 (N_5650,N_818,N_1524);
nor U5651 (N_5651,N_141,N_3984);
and U5652 (N_5652,N_272,N_1063);
or U5653 (N_5653,N_278,N_2372);
or U5654 (N_5654,N_670,N_2286);
and U5655 (N_5655,N_1536,N_223);
and U5656 (N_5656,N_1419,N_2658);
and U5657 (N_5657,N_429,N_2299);
or U5658 (N_5658,N_871,N_1770);
nand U5659 (N_5659,N_2813,N_3546);
nor U5660 (N_5660,N_1091,N_3518);
xor U5661 (N_5661,N_1860,N_11);
or U5662 (N_5662,N_899,N_1796);
nand U5663 (N_5663,N_3954,N_1182);
xor U5664 (N_5664,N_3829,N_2254);
or U5665 (N_5665,N_412,N_2541);
nor U5666 (N_5666,N_1296,N_225);
or U5667 (N_5667,N_789,N_2049);
nand U5668 (N_5668,N_2157,N_657);
or U5669 (N_5669,N_2759,N_1129);
or U5670 (N_5670,N_3417,N_1867);
nor U5671 (N_5671,N_584,N_1958);
nand U5672 (N_5672,N_3892,N_3213);
or U5673 (N_5673,N_2987,N_441);
nand U5674 (N_5674,N_1035,N_672);
nor U5675 (N_5675,N_1877,N_937);
nor U5676 (N_5676,N_2555,N_1848);
nor U5677 (N_5677,N_1325,N_3614);
and U5678 (N_5678,N_2374,N_3280);
nand U5679 (N_5679,N_419,N_2777);
or U5680 (N_5680,N_512,N_3162);
nand U5681 (N_5681,N_1130,N_1980);
nor U5682 (N_5682,N_3668,N_2479);
xor U5683 (N_5683,N_3602,N_123);
and U5684 (N_5684,N_1995,N_3025);
nand U5685 (N_5685,N_3825,N_1610);
nor U5686 (N_5686,N_2737,N_3511);
nand U5687 (N_5687,N_1656,N_2493);
or U5688 (N_5688,N_1733,N_3246);
nand U5689 (N_5689,N_54,N_2042);
nor U5690 (N_5690,N_1015,N_2119);
nor U5691 (N_5691,N_3763,N_643);
nor U5692 (N_5692,N_1840,N_3704);
and U5693 (N_5693,N_3495,N_227);
nand U5694 (N_5694,N_3399,N_2895);
nor U5695 (N_5695,N_459,N_1327);
and U5696 (N_5696,N_277,N_2470);
or U5697 (N_5697,N_3349,N_2918);
and U5698 (N_5698,N_1541,N_2746);
and U5699 (N_5699,N_362,N_2766);
nor U5700 (N_5700,N_3582,N_2688);
nor U5701 (N_5701,N_1620,N_3402);
and U5702 (N_5702,N_408,N_3613);
nand U5703 (N_5703,N_896,N_1654);
xnor U5704 (N_5704,N_3534,N_3525);
nand U5705 (N_5705,N_2019,N_1603);
and U5706 (N_5706,N_1547,N_3007);
nand U5707 (N_5707,N_552,N_1774);
nand U5708 (N_5708,N_1864,N_3321);
nor U5709 (N_5709,N_3701,N_2946);
nor U5710 (N_5710,N_1494,N_3663);
and U5711 (N_5711,N_1213,N_310);
and U5712 (N_5712,N_1996,N_162);
nor U5713 (N_5713,N_3285,N_3468);
nand U5714 (N_5714,N_1897,N_1624);
or U5715 (N_5715,N_770,N_2361);
and U5716 (N_5716,N_2793,N_3749);
nor U5717 (N_5717,N_3871,N_1146);
nand U5718 (N_5718,N_2795,N_615);
or U5719 (N_5719,N_2089,N_77);
nor U5720 (N_5720,N_1505,N_3722);
and U5721 (N_5721,N_2033,N_36);
and U5722 (N_5722,N_923,N_1075);
and U5723 (N_5723,N_2310,N_493);
nand U5724 (N_5724,N_782,N_2660);
nand U5725 (N_5725,N_2028,N_1008);
or U5726 (N_5726,N_3147,N_2791);
and U5727 (N_5727,N_3802,N_3896);
or U5728 (N_5728,N_3188,N_1385);
nand U5729 (N_5729,N_3230,N_326);
and U5730 (N_5730,N_848,N_756);
and U5731 (N_5731,N_3970,N_700);
nor U5732 (N_5732,N_3154,N_625);
or U5733 (N_5733,N_3095,N_3023);
or U5734 (N_5734,N_1959,N_3579);
and U5735 (N_5735,N_2955,N_1961);
nand U5736 (N_5736,N_2912,N_3035);
nor U5737 (N_5737,N_1145,N_1682);
and U5738 (N_5738,N_1566,N_398);
nor U5739 (N_5739,N_1057,N_1575);
nor U5740 (N_5740,N_2972,N_3282);
and U5741 (N_5741,N_2482,N_2368);
nand U5742 (N_5742,N_1453,N_2244);
nor U5743 (N_5743,N_2836,N_238);
or U5744 (N_5744,N_2196,N_358);
or U5745 (N_5745,N_2869,N_492);
or U5746 (N_5746,N_1072,N_2007);
nand U5747 (N_5747,N_3967,N_3734);
nor U5748 (N_5748,N_63,N_3178);
and U5749 (N_5749,N_3009,N_3690);
or U5750 (N_5750,N_1424,N_1873);
nand U5751 (N_5751,N_1894,N_1657);
nand U5752 (N_5752,N_3969,N_3203);
and U5753 (N_5753,N_1266,N_3076);
nand U5754 (N_5754,N_1499,N_3385);
or U5755 (N_5755,N_3971,N_2653);
xor U5756 (N_5756,N_2318,N_302);
nor U5757 (N_5757,N_993,N_2128);
and U5758 (N_5758,N_2582,N_2379);
or U5759 (N_5759,N_1869,N_3804);
nor U5760 (N_5760,N_467,N_2190);
and U5761 (N_5761,N_967,N_1582);
nor U5762 (N_5762,N_808,N_3999);
nand U5763 (N_5763,N_1585,N_1027);
nor U5764 (N_5764,N_2831,N_3831);
nand U5765 (N_5765,N_775,N_1418);
nor U5766 (N_5766,N_3767,N_155);
or U5767 (N_5767,N_281,N_1947);
or U5768 (N_5768,N_3669,N_616);
or U5769 (N_5769,N_2890,N_3149);
nand U5770 (N_5770,N_2907,N_720);
nor U5771 (N_5771,N_1747,N_1426);
and U5772 (N_5772,N_1831,N_3146);
and U5773 (N_5773,N_52,N_3494);
nand U5774 (N_5774,N_2021,N_2730);
or U5775 (N_5775,N_953,N_3380);
nand U5776 (N_5776,N_653,N_2194);
or U5777 (N_5777,N_2887,N_2146);
nand U5778 (N_5778,N_3782,N_1812);
xnor U5779 (N_5779,N_642,N_3323);
nor U5780 (N_5780,N_2615,N_61);
or U5781 (N_5781,N_1789,N_2514);
and U5782 (N_5782,N_2235,N_3517);
and U5783 (N_5783,N_3407,N_689);
nor U5784 (N_5784,N_1549,N_914);
xor U5785 (N_5785,N_322,N_2260);
xor U5786 (N_5786,N_2394,N_3917);
nor U5787 (N_5787,N_3326,N_924);
and U5788 (N_5788,N_2279,N_2036);
or U5789 (N_5789,N_3740,N_1820);
nor U5790 (N_5790,N_1856,N_1845);
nor U5791 (N_5791,N_760,N_1910);
xor U5792 (N_5792,N_897,N_2440);
xnor U5793 (N_5793,N_3845,N_2517);
nor U5794 (N_5794,N_3774,N_691);
nand U5795 (N_5795,N_553,N_3176);
xor U5796 (N_5796,N_3935,N_3726);
and U5797 (N_5797,N_825,N_752);
and U5798 (N_5798,N_384,N_1440);
nor U5799 (N_5799,N_1895,N_1984);
or U5800 (N_5800,N_1379,N_2562);
and U5801 (N_5801,N_3706,N_3433);
and U5802 (N_5802,N_3048,N_2610);
and U5803 (N_5803,N_3642,N_1776);
xor U5804 (N_5804,N_1178,N_2073);
nand U5805 (N_5805,N_2794,N_2471);
or U5806 (N_5806,N_1699,N_386);
nand U5807 (N_5807,N_2360,N_3419);
nand U5808 (N_5808,N_2234,N_545);
nor U5809 (N_5809,N_69,N_7);
nor U5810 (N_5810,N_184,N_596);
and U5811 (N_5811,N_2192,N_3756);
or U5812 (N_5812,N_2674,N_3499);
or U5813 (N_5813,N_2944,N_2106);
nor U5814 (N_5814,N_2486,N_772);
xnor U5815 (N_5815,N_828,N_3925);
nand U5816 (N_5816,N_305,N_917);
nand U5817 (N_5817,N_2662,N_95);
or U5818 (N_5818,N_1074,N_1957);
xnor U5819 (N_5819,N_1364,N_3507);
xor U5820 (N_5820,N_1029,N_1021);
nor U5821 (N_5821,N_2727,N_1557);
or U5822 (N_5822,N_779,N_868);
xor U5823 (N_5823,N_3483,N_2149);
nand U5824 (N_5824,N_883,N_2307);
nand U5825 (N_5825,N_2538,N_1595);
and U5826 (N_5826,N_2297,N_948);
and U5827 (N_5827,N_1398,N_1913);
nand U5828 (N_5828,N_3560,N_2923);
nand U5829 (N_5829,N_309,N_3182);
and U5830 (N_5830,N_2419,N_3708);
nand U5831 (N_5831,N_3428,N_737);
or U5832 (N_5832,N_741,N_2569);
nor U5833 (N_5833,N_2716,N_1677);
nor U5834 (N_5834,N_960,N_491);
or U5835 (N_5835,N_544,N_2187);
and U5836 (N_5836,N_2667,N_3252);
or U5837 (N_5837,N_2432,N_1218);
or U5838 (N_5838,N_2952,N_3652);
nand U5839 (N_5839,N_418,N_2498);
and U5840 (N_5840,N_1319,N_582);
nand U5841 (N_5841,N_2303,N_2098);
and U5842 (N_5842,N_3184,N_1805);
and U5843 (N_5843,N_2000,N_3785);
or U5844 (N_5844,N_3797,N_3830);
or U5845 (N_5845,N_3723,N_3509);
or U5846 (N_5846,N_3628,N_3129);
xor U5847 (N_5847,N_1749,N_3195);
and U5848 (N_5848,N_2874,N_1280);
and U5849 (N_5849,N_1134,N_662);
nor U5850 (N_5850,N_2121,N_3915);
nor U5851 (N_5851,N_3039,N_524);
or U5852 (N_5852,N_556,N_2876);
or U5853 (N_5853,N_165,N_2446);
or U5854 (N_5854,N_2841,N_3827);
or U5855 (N_5855,N_343,N_3778);
xnor U5856 (N_5856,N_1759,N_2954);
or U5857 (N_5857,N_3139,N_3117);
or U5858 (N_5858,N_1116,N_834);
or U5859 (N_5859,N_3031,N_1308);
and U5860 (N_5860,N_757,N_1013);
and U5861 (N_5861,N_554,N_2920);
nand U5862 (N_5862,N_1782,N_1944);
xnor U5863 (N_5863,N_3758,N_3073);
or U5864 (N_5864,N_292,N_1168);
nand U5865 (N_5865,N_3217,N_2577);
nor U5866 (N_5866,N_2480,N_3718);
and U5867 (N_5867,N_2280,N_1317);
nor U5868 (N_5868,N_1246,N_304);
and U5869 (N_5869,N_367,N_2378);
nand U5870 (N_5870,N_684,N_2370);
or U5871 (N_5871,N_266,N_3352);
or U5872 (N_5872,N_1571,N_3574);
nor U5873 (N_5873,N_624,N_2764);
nand U5874 (N_5874,N_3003,N_483);
nand U5875 (N_5875,N_106,N_975);
nor U5876 (N_5876,N_2990,N_1238);
nand U5877 (N_5877,N_3324,N_1644);
and U5878 (N_5878,N_35,N_1157);
nor U5879 (N_5879,N_62,N_1166);
nand U5880 (N_5880,N_3838,N_2721);
nor U5881 (N_5881,N_3069,N_3444);
or U5882 (N_5882,N_2934,N_1552);
and U5883 (N_5883,N_1977,N_646);
nand U5884 (N_5884,N_2185,N_1686);
or U5885 (N_5885,N_247,N_10);
nor U5886 (N_5886,N_3438,N_882);
nand U5887 (N_5887,N_2320,N_2459);
or U5888 (N_5888,N_3157,N_136);
nand U5889 (N_5889,N_979,N_1143);
xnor U5890 (N_5890,N_1528,N_3351);
or U5891 (N_5891,N_2824,N_65);
nor U5892 (N_5892,N_3810,N_2412);
xnor U5893 (N_5893,N_3792,N_3422);
or U5894 (N_5894,N_117,N_2029);
or U5895 (N_5895,N_1565,N_48);
nand U5896 (N_5896,N_214,N_728);
nor U5897 (N_5897,N_2948,N_508);
or U5898 (N_5898,N_1118,N_1955);
nand U5899 (N_5899,N_3769,N_2792);
and U5900 (N_5900,N_2122,N_1605);
or U5901 (N_5901,N_986,N_3824);
xor U5902 (N_5902,N_3866,N_2130);
and U5903 (N_5903,N_234,N_488);
nor U5904 (N_5904,N_3600,N_3010);
nand U5905 (N_5905,N_2906,N_297);
or U5906 (N_5906,N_2072,N_1150);
and U5907 (N_5907,N_3832,N_1344);
xor U5908 (N_5908,N_2182,N_2010);
nor U5909 (N_5909,N_609,N_1083);
nand U5910 (N_5910,N_3882,N_437);
nand U5911 (N_5911,N_3974,N_1174);
nor U5912 (N_5912,N_1778,N_581);
nor U5913 (N_5913,N_813,N_2788);
xnor U5914 (N_5914,N_3113,N_1924);
xnor U5915 (N_5915,N_857,N_3209);
nand U5916 (N_5916,N_3355,N_2341);
or U5917 (N_5917,N_982,N_401);
nand U5918 (N_5918,N_356,N_1162);
nand U5919 (N_5919,N_2925,N_2199);
nor U5920 (N_5920,N_3771,N_312);
and U5921 (N_5921,N_1051,N_3757);
and U5922 (N_5922,N_2218,N_1084);
or U5923 (N_5923,N_3923,N_131);
or U5924 (N_5924,N_213,N_3894);
xnor U5925 (N_5925,N_3067,N_2168);
xor U5926 (N_5926,N_159,N_2803);
or U5927 (N_5927,N_2682,N_2204);
nor U5928 (N_5928,N_3205,N_632);
or U5929 (N_5929,N_1316,N_1612);
or U5930 (N_5930,N_905,N_1177);
and U5931 (N_5931,N_962,N_3665);
nor U5932 (N_5932,N_3945,N_3287);
or U5933 (N_5933,N_1149,N_754);
nand U5934 (N_5934,N_1019,N_1627);
nor U5935 (N_5935,N_1229,N_996);
xor U5936 (N_5936,N_3111,N_599);
nand U5937 (N_5937,N_3949,N_2293);
xor U5938 (N_5938,N_879,N_2530);
or U5939 (N_5939,N_1767,N_2862);
and U5940 (N_5940,N_2065,N_2830);
nand U5941 (N_5941,N_2510,N_3465);
nor U5942 (N_5942,N_3052,N_2294);
xnor U5943 (N_5943,N_3260,N_1405);
nand U5944 (N_5944,N_2203,N_787);
xor U5945 (N_5945,N_2757,N_3567);
nor U5946 (N_5946,N_2578,N_89);
nor U5947 (N_5947,N_3398,N_2883);
nand U5948 (N_5948,N_3928,N_693);
and U5949 (N_5949,N_2983,N_1392);
xor U5950 (N_5950,N_1219,N_3318);
or U5951 (N_5951,N_3181,N_1264);
nand U5952 (N_5952,N_1330,N_113);
nor U5953 (N_5953,N_3980,N_2039);
nand U5954 (N_5954,N_301,N_3016);
nand U5955 (N_5955,N_683,N_192);
or U5956 (N_5956,N_1938,N_3944);
nor U5957 (N_5957,N_121,N_3689);
and U5958 (N_5958,N_2079,N_495);
or U5959 (N_5959,N_1087,N_3219);
nand U5960 (N_5960,N_2384,N_2443);
or U5961 (N_5961,N_3979,N_2984);
or U5962 (N_5962,N_2427,N_3604);
nand U5963 (N_5963,N_695,N_3293);
nand U5964 (N_5964,N_29,N_2892);
nor U5965 (N_5965,N_546,N_1003);
or U5966 (N_5966,N_2351,N_2077);
nand U5967 (N_5967,N_1233,N_2205);
nand U5968 (N_5968,N_1023,N_341);
nand U5969 (N_5969,N_2390,N_3978);
nand U5970 (N_5970,N_3834,N_2728);
or U5971 (N_5971,N_338,N_2825);
or U5972 (N_5972,N_428,N_1076);
or U5973 (N_5973,N_2252,N_357);
nand U5974 (N_5974,N_3187,N_1111);
and U5975 (N_5975,N_3912,N_2978);
nand U5976 (N_5976,N_2738,N_331);
or U5977 (N_5977,N_2561,N_1425);
nand U5978 (N_5978,N_3597,N_2554);
xor U5979 (N_5979,N_854,N_3308);
or U5980 (N_5980,N_2740,N_1348);
or U5981 (N_5981,N_3245,N_3328);
xor U5982 (N_5982,N_620,N_1830);
xor U5983 (N_5983,N_520,N_3887);
nand U5984 (N_5984,N_1249,N_1949);
or U5985 (N_5985,N_1746,N_2040);
nor U5986 (N_5986,N_1597,N_942);
nor U5987 (N_5987,N_890,N_3082);
nand U5988 (N_5988,N_3584,N_1001);
and U5989 (N_5989,N_2879,N_1987);
and U5990 (N_5990,N_1852,N_3235);
nor U5991 (N_5991,N_2085,N_1635);
nor U5992 (N_5992,N_3788,N_2849);
and U5993 (N_5993,N_381,N_2312);
nand U5994 (N_5994,N_2679,N_1821);
and U5995 (N_5995,N_321,N_3913);
or U5996 (N_5996,N_1208,N_364);
nand U5997 (N_5997,N_474,N_1909);
nand U5998 (N_5998,N_2511,N_3123);
xor U5999 (N_5999,N_3314,N_1115);
and U6000 (N_6000,N_2193,N_617);
nor U6001 (N_6001,N_117,N_3173);
or U6002 (N_6002,N_2157,N_2370);
nor U6003 (N_6003,N_2622,N_916);
nand U6004 (N_6004,N_1886,N_1401);
nand U6005 (N_6005,N_2871,N_2865);
or U6006 (N_6006,N_1534,N_2510);
or U6007 (N_6007,N_1503,N_2226);
xnor U6008 (N_6008,N_305,N_1183);
and U6009 (N_6009,N_3311,N_3700);
and U6010 (N_6010,N_1151,N_2089);
nor U6011 (N_6011,N_431,N_2329);
or U6012 (N_6012,N_777,N_3942);
nand U6013 (N_6013,N_1528,N_3772);
and U6014 (N_6014,N_1273,N_2882);
nand U6015 (N_6015,N_1043,N_2959);
or U6016 (N_6016,N_1952,N_2843);
nand U6017 (N_6017,N_2360,N_2816);
nor U6018 (N_6018,N_3338,N_1027);
or U6019 (N_6019,N_1917,N_2116);
or U6020 (N_6020,N_432,N_3996);
or U6021 (N_6021,N_2913,N_2764);
and U6022 (N_6022,N_3838,N_2804);
or U6023 (N_6023,N_1876,N_3932);
nor U6024 (N_6024,N_138,N_2991);
and U6025 (N_6025,N_721,N_2478);
nand U6026 (N_6026,N_3335,N_292);
or U6027 (N_6027,N_1385,N_2052);
nand U6028 (N_6028,N_239,N_1992);
nor U6029 (N_6029,N_3649,N_3630);
or U6030 (N_6030,N_1638,N_216);
nor U6031 (N_6031,N_2962,N_2456);
or U6032 (N_6032,N_774,N_1291);
nor U6033 (N_6033,N_3993,N_2689);
nand U6034 (N_6034,N_1389,N_2487);
nand U6035 (N_6035,N_3483,N_148);
or U6036 (N_6036,N_3201,N_132);
nand U6037 (N_6037,N_2221,N_3273);
and U6038 (N_6038,N_1589,N_678);
nor U6039 (N_6039,N_128,N_3834);
and U6040 (N_6040,N_3580,N_3075);
or U6041 (N_6041,N_1144,N_3967);
and U6042 (N_6042,N_1528,N_2296);
and U6043 (N_6043,N_2175,N_3804);
and U6044 (N_6044,N_3456,N_3828);
and U6045 (N_6045,N_1085,N_345);
and U6046 (N_6046,N_344,N_386);
xnor U6047 (N_6047,N_2280,N_549);
and U6048 (N_6048,N_3504,N_1284);
or U6049 (N_6049,N_1073,N_571);
nor U6050 (N_6050,N_1570,N_3889);
nand U6051 (N_6051,N_681,N_2903);
and U6052 (N_6052,N_6,N_104);
nor U6053 (N_6053,N_3135,N_1911);
and U6054 (N_6054,N_1880,N_1628);
or U6055 (N_6055,N_433,N_1905);
nand U6056 (N_6056,N_1432,N_295);
xor U6057 (N_6057,N_3869,N_2434);
nand U6058 (N_6058,N_1651,N_2740);
nor U6059 (N_6059,N_1626,N_764);
nor U6060 (N_6060,N_3067,N_2681);
nor U6061 (N_6061,N_3414,N_2030);
nor U6062 (N_6062,N_1623,N_1301);
and U6063 (N_6063,N_2106,N_747);
and U6064 (N_6064,N_1784,N_923);
nor U6065 (N_6065,N_1216,N_3980);
nor U6066 (N_6066,N_3046,N_3529);
xnor U6067 (N_6067,N_989,N_3437);
nand U6068 (N_6068,N_1184,N_3308);
xnor U6069 (N_6069,N_3042,N_2883);
nor U6070 (N_6070,N_3042,N_2643);
nand U6071 (N_6071,N_3748,N_1595);
or U6072 (N_6072,N_1515,N_1530);
or U6073 (N_6073,N_208,N_2978);
and U6074 (N_6074,N_51,N_2565);
nand U6075 (N_6075,N_3565,N_3922);
nand U6076 (N_6076,N_2637,N_3120);
nand U6077 (N_6077,N_2892,N_591);
xor U6078 (N_6078,N_1715,N_3718);
nor U6079 (N_6079,N_2005,N_664);
or U6080 (N_6080,N_3683,N_183);
or U6081 (N_6081,N_2774,N_3240);
nor U6082 (N_6082,N_585,N_1824);
and U6083 (N_6083,N_3353,N_1724);
nor U6084 (N_6084,N_779,N_2039);
nor U6085 (N_6085,N_2462,N_2630);
and U6086 (N_6086,N_2782,N_3692);
and U6087 (N_6087,N_3058,N_3012);
nand U6088 (N_6088,N_326,N_3856);
or U6089 (N_6089,N_3168,N_3949);
or U6090 (N_6090,N_2158,N_1945);
xnor U6091 (N_6091,N_2973,N_1433);
xor U6092 (N_6092,N_1886,N_3254);
nor U6093 (N_6093,N_3403,N_533);
and U6094 (N_6094,N_928,N_904);
and U6095 (N_6095,N_738,N_2889);
or U6096 (N_6096,N_2652,N_1416);
nor U6097 (N_6097,N_3056,N_3614);
or U6098 (N_6098,N_1666,N_3861);
nand U6099 (N_6099,N_994,N_3734);
or U6100 (N_6100,N_2813,N_2371);
nor U6101 (N_6101,N_1437,N_580);
nor U6102 (N_6102,N_754,N_3623);
and U6103 (N_6103,N_2418,N_3316);
or U6104 (N_6104,N_2595,N_2680);
and U6105 (N_6105,N_425,N_69);
and U6106 (N_6106,N_3757,N_1763);
nor U6107 (N_6107,N_940,N_3386);
nand U6108 (N_6108,N_3549,N_1590);
xnor U6109 (N_6109,N_2089,N_3930);
nor U6110 (N_6110,N_2123,N_3534);
nand U6111 (N_6111,N_1499,N_3442);
xor U6112 (N_6112,N_2122,N_2177);
and U6113 (N_6113,N_2558,N_641);
nand U6114 (N_6114,N_3655,N_3806);
and U6115 (N_6115,N_2186,N_627);
or U6116 (N_6116,N_2029,N_3303);
nand U6117 (N_6117,N_1720,N_1475);
nor U6118 (N_6118,N_1710,N_444);
or U6119 (N_6119,N_3538,N_3793);
nand U6120 (N_6120,N_3840,N_1545);
nand U6121 (N_6121,N_3350,N_1284);
and U6122 (N_6122,N_578,N_2891);
and U6123 (N_6123,N_2408,N_62);
and U6124 (N_6124,N_2937,N_3767);
and U6125 (N_6125,N_1236,N_2093);
and U6126 (N_6126,N_624,N_3271);
xnor U6127 (N_6127,N_1618,N_2877);
and U6128 (N_6128,N_335,N_3997);
xnor U6129 (N_6129,N_2050,N_1499);
and U6130 (N_6130,N_1383,N_3574);
or U6131 (N_6131,N_3658,N_3544);
nor U6132 (N_6132,N_151,N_71);
nand U6133 (N_6133,N_81,N_2075);
or U6134 (N_6134,N_2311,N_1389);
and U6135 (N_6135,N_3093,N_370);
and U6136 (N_6136,N_2877,N_821);
and U6137 (N_6137,N_715,N_2586);
nor U6138 (N_6138,N_90,N_2395);
or U6139 (N_6139,N_3766,N_91);
nand U6140 (N_6140,N_1666,N_3265);
nand U6141 (N_6141,N_1120,N_3880);
nor U6142 (N_6142,N_3051,N_1018);
or U6143 (N_6143,N_2842,N_3360);
xnor U6144 (N_6144,N_3753,N_1746);
nor U6145 (N_6145,N_1186,N_1348);
and U6146 (N_6146,N_2482,N_433);
and U6147 (N_6147,N_2824,N_2004);
nand U6148 (N_6148,N_1924,N_3190);
or U6149 (N_6149,N_286,N_1393);
nor U6150 (N_6150,N_2264,N_687);
and U6151 (N_6151,N_3363,N_2886);
nand U6152 (N_6152,N_178,N_3728);
nor U6153 (N_6153,N_956,N_691);
nor U6154 (N_6154,N_2020,N_1421);
or U6155 (N_6155,N_662,N_2328);
nand U6156 (N_6156,N_3950,N_115);
and U6157 (N_6157,N_3957,N_2863);
and U6158 (N_6158,N_2809,N_3696);
xor U6159 (N_6159,N_1486,N_3889);
or U6160 (N_6160,N_1938,N_1490);
and U6161 (N_6161,N_1458,N_2588);
nand U6162 (N_6162,N_2163,N_3505);
nor U6163 (N_6163,N_1023,N_1879);
xor U6164 (N_6164,N_3277,N_1353);
or U6165 (N_6165,N_317,N_471);
and U6166 (N_6166,N_202,N_2908);
or U6167 (N_6167,N_2326,N_914);
or U6168 (N_6168,N_2214,N_1154);
and U6169 (N_6169,N_670,N_1592);
and U6170 (N_6170,N_2836,N_3929);
and U6171 (N_6171,N_3486,N_2453);
nor U6172 (N_6172,N_2019,N_2432);
nor U6173 (N_6173,N_1779,N_2574);
nor U6174 (N_6174,N_1984,N_3599);
xor U6175 (N_6175,N_1744,N_621);
or U6176 (N_6176,N_3460,N_2220);
or U6177 (N_6177,N_2105,N_393);
and U6178 (N_6178,N_1834,N_2457);
xnor U6179 (N_6179,N_2992,N_516);
nor U6180 (N_6180,N_3070,N_2327);
and U6181 (N_6181,N_2594,N_379);
nand U6182 (N_6182,N_1628,N_2714);
xor U6183 (N_6183,N_2257,N_2576);
nand U6184 (N_6184,N_2854,N_1150);
nand U6185 (N_6185,N_373,N_1438);
nor U6186 (N_6186,N_1236,N_3527);
nor U6187 (N_6187,N_319,N_1581);
nor U6188 (N_6188,N_3268,N_780);
or U6189 (N_6189,N_3018,N_860);
nor U6190 (N_6190,N_2869,N_3134);
nor U6191 (N_6191,N_2328,N_605);
and U6192 (N_6192,N_2379,N_694);
nand U6193 (N_6193,N_434,N_53);
nor U6194 (N_6194,N_2726,N_1916);
nand U6195 (N_6195,N_2428,N_2990);
nor U6196 (N_6196,N_2994,N_3453);
or U6197 (N_6197,N_1677,N_222);
nand U6198 (N_6198,N_1000,N_2141);
xor U6199 (N_6199,N_751,N_3168);
or U6200 (N_6200,N_3478,N_961);
or U6201 (N_6201,N_1263,N_1816);
and U6202 (N_6202,N_3297,N_3575);
nand U6203 (N_6203,N_2936,N_3232);
or U6204 (N_6204,N_1777,N_3341);
nand U6205 (N_6205,N_408,N_2687);
nor U6206 (N_6206,N_1406,N_487);
nand U6207 (N_6207,N_1243,N_285);
and U6208 (N_6208,N_3285,N_2744);
xnor U6209 (N_6209,N_2993,N_639);
nand U6210 (N_6210,N_1483,N_199);
and U6211 (N_6211,N_2177,N_3307);
and U6212 (N_6212,N_3969,N_1403);
and U6213 (N_6213,N_3816,N_3077);
nand U6214 (N_6214,N_3605,N_2144);
xor U6215 (N_6215,N_2719,N_2111);
nand U6216 (N_6216,N_673,N_2089);
xor U6217 (N_6217,N_1691,N_2307);
or U6218 (N_6218,N_3726,N_800);
nor U6219 (N_6219,N_327,N_455);
nor U6220 (N_6220,N_3679,N_1745);
or U6221 (N_6221,N_3298,N_2771);
and U6222 (N_6222,N_2857,N_2802);
nand U6223 (N_6223,N_430,N_1192);
or U6224 (N_6224,N_1597,N_3248);
and U6225 (N_6225,N_2053,N_1868);
nand U6226 (N_6226,N_2659,N_2967);
nor U6227 (N_6227,N_786,N_3193);
nor U6228 (N_6228,N_840,N_634);
xnor U6229 (N_6229,N_1335,N_1148);
or U6230 (N_6230,N_3347,N_2676);
and U6231 (N_6231,N_2160,N_3932);
nor U6232 (N_6232,N_3165,N_2717);
nor U6233 (N_6233,N_3027,N_3393);
and U6234 (N_6234,N_3635,N_1958);
nand U6235 (N_6235,N_3968,N_2984);
nand U6236 (N_6236,N_621,N_978);
nor U6237 (N_6237,N_2752,N_3307);
nor U6238 (N_6238,N_538,N_1169);
xnor U6239 (N_6239,N_713,N_2153);
nor U6240 (N_6240,N_3584,N_1759);
xor U6241 (N_6241,N_3067,N_2585);
or U6242 (N_6242,N_3060,N_3201);
xor U6243 (N_6243,N_3893,N_825);
xor U6244 (N_6244,N_1823,N_593);
and U6245 (N_6245,N_441,N_971);
or U6246 (N_6246,N_2912,N_858);
xnor U6247 (N_6247,N_2516,N_1217);
nand U6248 (N_6248,N_2658,N_3730);
xnor U6249 (N_6249,N_3299,N_590);
xnor U6250 (N_6250,N_3691,N_911);
nor U6251 (N_6251,N_1831,N_2344);
and U6252 (N_6252,N_1141,N_469);
nor U6253 (N_6253,N_3556,N_2097);
or U6254 (N_6254,N_1898,N_3980);
nand U6255 (N_6255,N_589,N_1288);
nor U6256 (N_6256,N_2114,N_3677);
or U6257 (N_6257,N_3004,N_274);
nor U6258 (N_6258,N_2509,N_1816);
nor U6259 (N_6259,N_3475,N_1325);
and U6260 (N_6260,N_1613,N_1686);
or U6261 (N_6261,N_2108,N_97);
nor U6262 (N_6262,N_1618,N_583);
or U6263 (N_6263,N_1114,N_3791);
xnor U6264 (N_6264,N_2553,N_2118);
xnor U6265 (N_6265,N_2333,N_870);
nor U6266 (N_6266,N_3918,N_3834);
nand U6267 (N_6267,N_1419,N_3793);
xnor U6268 (N_6268,N_1470,N_556);
and U6269 (N_6269,N_266,N_3146);
nand U6270 (N_6270,N_268,N_577);
or U6271 (N_6271,N_2205,N_2618);
and U6272 (N_6272,N_2839,N_2442);
or U6273 (N_6273,N_2762,N_2559);
nor U6274 (N_6274,N_370,N_396);
or U6275 (N_6275,N_3498,N_570);
or U6276 (N_6276,N_3062,N_1345);
and U6277 (N_6277,N_1781,N_1570);
and U6278 (N_6278,N_508,N_1533);
nor U6279 (N_6279,N_1717,N_3935);
nand U6280 (N_6280,N_2943,N_3995);
and U6281 (N_6281,N_532,N_2956);
or U6282 (N_6282,N_3550,N_13);
or U6283 (N_6283,N_3544,N_379);
nand U6284 (N_6284,N_3214,N_414);
or U6285 (N_6285,N_1588,N_2617);
or U6286 (N_6286,N_702,N_2389);
xor U6287 (N_6287,N_1028,N_2662);
xnor U6288 (N_6288,N_3474,N_3182);
nor U6289 (N_6289,N_2695,N_1182);
nand U6290 (N_6290,N_2582,N_290);
nand U6291 (N_6291,N_2482,N_1843);
nand U6292 (N_6292,N_371,N_2123);
or U6293 (N_6293,N_1486,N_249);
or U6294 (N_6294,N_984,N_1979);
and U6295 (N_6295,N_2048,N_1443);
or U6296 (N_6296,N_1919,N_3982);
and U6297 (N_6297,N_1764,N_2403);
or U6298 (N_6298,N_92,N_689);
and U6299 (N_6299,N_2352,N_3198);
and U6300 (N_6300,N_842,N_1172);
nor U6301 (N_6301,N_3587,N_3645);
xor U6302 (N_6302,N_2846,N_87);
nor U6303 (N_6303,N_2530,N_2002);
or U6304 (N_6304,N_677,N_3687);
or U6305 (N_6305,N_3619,N_3554);
xor U6306 (N_6306,N_2835,N_983);
nand U6307 (N_6307,N_1616,N_3150);
nand U6308 (N_6308,N_701,N_6);
nand U6309 (N_6309,N_2786,N_3271);
nand U6310 (N_6310,N_1424,N_3371);
and U6311 (N_6311,N_573,N_3568);
xnor U6312 (N_6312,N_3215,N_2624);
or U6313 (N_6313,N_11,N_3638);
nor U6314 (N_6314,N_2723,N_966);
or U6315 (N_6315,N_3482,N_1178);
nor U6316 (N_6316,N_1269,N_2794);
nor U6317 (N_6317,N_2853,N_608);
and U6318 (N_6318,N_1365,N_797);
xor U6319 (N_6319,N_1384,N_1874);
and U6320 (N_6320,N_2192,N_3502);
and U6321 (N_6321,N_3812,N_3832);
nor U6322 (N_6322,N_2154,N_2799);
and U6323 (N_6323,N_2664,N_394);
and U6324 (N_6324,N_144,N_2141);
nand U6325 (N_6325,N_3,N_3077);
nor U6326 (N_6326,N_573,N_2954);
nor U6327 (N_6327,N_1451,N_3992);
or U6328 (N_6328,N_1152,N_943);
xor U6329 (N_6329,N_483,N_507);
and U6330 (N_6330,N_2235,N_307);
and U6331 (N_6331,N_3060,N_1460);
nor U6332 (N_6332,N_1027,N_3410);
or U6333 (N_6333,N_491,N_1243);
and U6334 (N_6334,N_1944,N_3761);
nand U6335 (N_6335,N_3062,N_733);
and U6336 (N_6336,N_2114,N_3911);
nand U6337 (N_6337,N_1586,N_2377);
and U6338 (N_6338,N_3308,N_3504);
or U6339 (N_6339,N_1841,N_2938);
or U6340 (N_6340,N_2885,N_3749);
or U6341 (N_6341,N_1758,N_902);
and U6342 (N_6342,N_3321,N_3690);
xor U6343 (N_6343,N_3329,N_1234);
nor U6344 (N_6344,N_89,N_1979);
nor U6345 (N_6345,N_3107,N_3438);
or U6346 (N_6346,N_1879,N_357);
or U6347 (N_6347,N_3012,N_1026);
and U6348 (N_6348,N_96,N_601);
nor U6349 (N_6349,N_640,N_742);
nand U6350 (N_6350,N_246,N_545);
nand U6351 (N_6351,N_562,N_3598);
or U6352 (N_6352,N_3802,N_229);
nand U6353 (N_6353,N_2715,N_3098);
nand U6354 (N_6354,N_721,N_1077);
nand U6355 (N_6355,N_2697,N_866);
nand U6356 (N_6356,N_2119,N_3339);
and U6357 (N_6357,N_2345,N_862);
and U6358 (N_6358,N_1827,N_3622);
or U6359 (N_6359,N_832,N_2102);
and U6360 (N_6360,N_3225,N_3812);
nor U6361 (N_6361,N_461,N_1340);
nor U6362 (N_6362,N_1992,N_1024);
nand U6363 (N_6363,N_3182,N_1600);
nand U6364 (N_6364,N_3532,N_2601);
and U6365 (N_6365,N_3611,N_1702);
and U6366 (N_6366,N_2054,N_2917);
nand U6367 (N_6367,N_1691,N_3191);
and U6368 (N_6368,N_1075,N_3325);
or U6369 (N_6369,N_184,N_3782);
and U6370 (N_6370,N_255,N_3848);
and U6371 (N_6371,N_2951,N_1259);
nor U6372 (N_6372,N_1723,N_2604);
nor U6373 (N_6373,N_1175,N_1531);
or U6374 (N_6374,N_2532,N_1698);
nand U6375 (N_6375,N_2560,N_938);
or U6376 (N_6376,N_2354,N_2516);
nand U6377 (N_6377,N_2610,N_1916);
and U6378 (N_6378,N_1594,N_2840);
xor U6379 (N_6379,N_3589,N_1610);
xor U6380 (N_6380,N_1426,N_1395);
xor U6381 (N_6381,N_1931,N_65);
nand U6382 (N_6382,N_2335,N_2444);
nand U6383 (N_6383,N_3409,N_3722);
xor U6384 (N_6384,N_492,N_3806);
or U6385 (N_6385,N_953,N_3270);
nand U6386 (N_6386,N_2023,N_3546);
and U6387 (N_6387,N_2154,N_3433);
and U6388 (N_6388,N_1841,N_3886);
or U6389 (N_6389,N_2494,N_166);
nand U6390 (N_6390,N_1958,N_2117);
nor U6391 (N_6391,N_36,N_319);
nor U6392 (N_6392,N_3735,N_3750);
nand U6393 (N_6393,N_1910,N_3157);
nor U6394 (N_6394,N_3629,N_1355);
or U6395 (N_6395,N_570,N_3458);
or U6396 (N_6396,N_2364,N_302);
or U6397 (N_6397,N_2678,N_3317);
nand U6398 (N_6398,N_1347,N_351);
or U6399 (N_6399,N_525,N_3369);
nor U6400 (N_6400,N_3338,N_2940);
or U6401 (N_6401,N_553,N_2806);
or U6402 (N_6402,N_3426,N_478);
nor U6403 (N_6403,N_361,N_681);
and U6404 (N_6404,N_3945,N_2215);
nor U6405 (N_6405,N_2121,N_1660);
and U6406 (N_6406,N_1994,N_3963);
nor U6407 (N_6407,N_798,N_679);
xnor U6408 (N_6408,N_3857,N_1082);
nand U6409 (N_6409,N_686,N_374);
nand U6410 (N_6410,N_2016,N_2482);
and U6411 (N_6411,N_2980,N_2753);
or U6412 (N_6412,N_2111,N_2067);
nor U6413 (N_6413,N_2274,N_1238);
nand U6414 (N_6414,N_3854,N_2725);
nand U6415 (N_6415,N_3984,N_22);
nand U6416 (N_6416,N_568,N_1345);
and U6417 (N_6417,N_3784,N_2751);
or U6418 (N_6418,N_1765,N_3572);
or U6419 (N_6419,N_1027,N_1535);
nor U6420 (N_6420,N_1471,N_2268);
nand U6421 (N_6421,N_1720,N_1326);
nand U6422 (N_6422,N_2193,N_2559);
nor U6423 (N_6423,N_3032,N_696);
nor U6424 (N_6424,N_1014,N_1671);
and U6425 (N_6425,N_2408,N_848);
nand U6426 (N_6426,N_1734,N_810);
nor U6427 (N_6427,N_674,N_857);
nor U6428 (N_6428,N_1216,N_2452);
nor U6429 (N_6429,N_3733,N_3011);
xor U6430 (N_6430,N_2800,N_232);
or U6431 (N_6431,N_2722,N_3701);
or U6432 (N_6432,N_1303,N_2020);
and U6433 (N_6433,N_3315,N_928);
and U6434 (N_6434,N_3845,N_1699);
and U6435 (N_6435,N_1714,N_3762);
and U6436 (N_6436,N_3756,N_3158);
or U6437 (N_6437,N_836,N_415);
nor U6438 (N_6438,N_166,N_3869);
or U6439 (N_6439,N_3890,N_660);
nor U6440 (N_6440,N_2860,N_327);
and U6441 (N_6441,N_977,N_481);
or U6442 (N_6442,N_3380,N_2021);
nor U6443 (N_6443,N_2594,N_383);
nor U6444 (N_6444,N_842,N_1351);
nor U6445 (N_6445,N_3708,N_1545);
and U6446 (N_6446,N_3240,N_3706);
nor U6447 (N_6447,N_1273,N_2909);
nand U6448 (N_6448,N_1284,N_1063);
nor U6449 (N_6449,N_2075,N_387);
nor U6450 (N_6450,N_2517,N_3668);
xnor U6451 (N_6451,N_3830,N_37);
nor U6452 (N_6452,N_2228,N_3980);
or U6453 (N_6453,N_1426,N_1095);
nand U6454 (N_6454,N_2979,N_3167);
or U6455 (N_6455,N_3699,N_1921);
nor U6456 (N_6456,N_2110,N_1341);
nand U6457 (N_6457,N_919,N_1706);
or U6458 (N_6458,N_2355,N_2910);
nand U6459 (N_6459,N_2537,N_1943);
and U6460 (N_6460,N_3438,N_1486);
nor U6461 (N_6461,N_2759,N_30);
and U6462 (N_6462,N_38,N_3524);
and U6463 (N_6463,N_1807,N_3501);
or U6464 (N_6464,N_3688,N_3829);
and U6465 (N_6465,N_1847,N_2997);
nor U6466 (N_6466,N_492,N_2229);
or U6467 (N_6467,N_3717,N_2495);
nand U6468 (N_6468,N_521,N_1892);
and U6469 (N_6469,N_3470,N_1238);
nand U6470 (N_6470,N_1062,N_3177);
and U6471 (N_6471,N_3070,N_3243);
or U6472 (N_6472,N_1934,N_3272);
xor U6473 (N_6473,N_361,N_2584);
nor U6474 (N_6474,N_3175,N_1949);
and U6475 (N_6475,N_1124,N_2809);
and U6476 (N_6476,N_2081,N_3067);
and U6477 (N_6477,N_3397,N_3829);
or U6478 (N_6478,N_873,N_2016);
nand U6479 (N_6479,N_3006,N_3562);
xor U6480 (N_6480,N_2809,N_151);
and U6481 (N_6481,N_1578,N_3714);
or U6482 (N_6482,N_1593,N_1573);
and U6483 (N_6483,N_3815,N_3822);
nand U6484 (N_6484,N_3356,N_801);
and U6485 (N_6485,N_607,N_304);
and U6486 (N_6486,N_3403,N_1642);
and U6487 (N_6487,N_2020,N_3173);
and U6488 (N_6488,N_2935,N_1763);
nand U6489 (N_6489,N_3252,N_3981);
nor U6490 (N_6490,N_3431,N_2917);
nand U6491 (N_6491,N_3097,N_1084);
and U6492 (N_6492,N_1380,N_2596);
or U6493 (N_6493,N_2443,N_3860);
and U6494 (N_6494,N_1059,N_505);
and U6495 (N_6495,N_2689,N_3698);
xnor U6496 (N_6496,N_3405,N_623);
or U6497 (N_6497,N_2704,N_2293);
or U6498 (N_6498,N_312,N_3064);
and U6499 (N_6499,N_1789,N_3646);
and U6500 (N_6500,N_3555,N_3242);
nand U6501 (N_6501,N_2765,N_1956);
nand U6502 (N_6502,N_1565,N_1986);
and U6503 (N_6503,N_2524,N_169);
nand U6504 (N_6504,N_1955,N_2162);
or U6505 (N_6505,N_2577,N_3496);
and U6506 (N_6506,N_172,N_497);
and U6507 (N_6507,N_2780,N_3859);
and U6508 (N_6508,N_1879,N_1656);
nand U6509 (N_6509,N_2584,N_2518);
nand U6510 (N_6510,N_3118,N_645);
and U6511 (N_6511,N_999,N_3279);
nor U6512 (N_6512,N_3030,N_2084);
and U6513 (N_6513,N_1087,N_361);
nand U6514 (N_6514,N_523,N_228);
or U6515 (N_6515,N_2931,N_2791);
and U6516 (N_6516,N_216,N_1568);
nor U6517 (N_6517,N_2010,N_2788);
nor U6518 (N_6518,N_2548,N_2597);
nand U6519 (N_6519,N_1219,N_1597);
or U6520 (N_6520,N_2873,N_1202);
nand U6521 (N_6521,N_2857,N_896);
nand U6522 (N_6522,N_3342,N_3022);
and U6523 (N_6523,N_3218,N_612);
or U6524 (N_6524,N_2205,N_1700);
nand U6525 (N_6525,N_2863,N_2178);
or U6526 (N_6526,N_627,N_594);
xnor U6527 (N_6527,N_1904,N_2719);
and U6528 (N_6528,N_2176,N_2816);
or U6529 (N_6529,N_3601,N_3047);
and U6530 (N_6530,N_3894,N_538);
nor U6531 (N_6531,N_3695,N_931);
or U6532 (N_6532,N_1501,N_1369);
or U6533 (N_6533,N_3730,N_2550);
nor U6534 (N_6534,N_1024,N_1447);
nor U6535 (N_6535,N_2179,N_3827);
and U6536 (N_6536,N_1543,N_1599);
or U6537 (N_6537,N_1507,N_2626);
nor U6538 (N_6538,N_1096,N_342);
nand U6539 (N_6539,N_1940,N_3379);
nand U6540 (N_6540,N_3972,N_2014);
or U6541 (N_6541,N_1918,N_3044);
and U6542 (N_6542,N_3605,N_2681);
or U6543 (N_6543,N_3118,N_3800);
nand U6544 (N_6544,N_1974,N_1553);
nand U6545 (N_6545,N_3636,N_3132);
or U6546 (N_6546,N_1594,N_3103);
and U6547 (N_6547,N_2862,N_2329);
or U6548 (N_6548,N_814,N_2583);
or U6549 (N_6549,N_558,N_2686);
nand U6550 (N_6550,N_2365,N_1731);
or U6551 (N_6551,N_420,N_10);
nand U6552 (N_6552,N_2795,N_2638);
xnor U6553 (N_6553,N_556,N_548);
or U6554 (N_6554,N_393,N_3577);
or U6555 (N_6555,N_1759,N_3435);
and U6556 (N_6556,N_893,N_3410);
and U6557 (N_6557,N_1204,N_1946);
nor U6558 (N_6558,N_1386,N_2856);
xor U6559 (N_6559,N_2622,N_2929);
or U6560 (N_6560,N_479,N_1568);
xor U6561 (N_6561,N_2923,N_1758);
xor U6562 (N_6562,N_497,N_2117);
nand U6563 (N_6563,N_348,N_2080);
xnor U6564 (N_6564,N_634,N_668);
nand U6565 (N_6565,N_2314,N_559);
nand U6566 (N_6566,N_2902,N_1258);
nor U6567 (N_6567,N_475,N_2071);
nand U6568 (N_6568,N_2421,N_714);
nor U6569 (N_6569,N_101,N_1088);
or U6570 (N_6570,N_535,N_2862);
nand U6571 (N_6571,N_2495,N_1628);
or U6572 (N_6572,N_1307,N_1955);
and U6573 (N_6573,N_1221,N_2377);
or U6574 (N_6574,N_800,N_1419);
nand U6575 (N_6575,N_2554,N_14);
and U6576 (N_6576,N_2519,N_1681);
or U6577 (N_6577,N_858,N_2434);
or U6578 (N_6578,N_87,N_1881);
and U6579 (N_6579,N_981,N_3188);
nand U6580 (N_6580,N_1291,N_2602);
nand U6581 (N_6581,N_3388,N_3343);
or U6582 (N_6582,N_3088,N_2692);
nand U6583 (N_6583,N_2833,N_3366);
or U6584 (N_6584,N_3198,N_2062);
nand U6585 (N_6585,N_2404,N_1227);
nand U6586 (N_6586,N_1160,N_237);
nand U6587 (N_6587,N_290,N_2728);
nand U6588 (N_6588,N_1348,N_970);
or U6589 (N_6589,N_1351,N_532);
nor U6590 (N_6590,N_582,N_1412);
nand U6591 (N_6591,N_470,N_2308);
and U6592 (N_6592,N_3951,N_974);
nor U6593 (N_6593,N_1489,N_1302);
or U6594 (N_6594,N_3373,N_3724);
xor U6595 (N_6595,N_1877,N_134);
nor U6596 (N_6596,N_556,N_654);
nor U6597 (N_6597,N_864,N_1689);
xnor U6598 (N_6598,N_3723,N_2780);
or U6599 (N_6599,N_3917,N_522);
xor U6600 (N_6600,N_586,N_3235);
and U6601 (N_6601,N_959,N_3270);
xnor U6602 (N_6602,N_3433,N_2635);
nand U6603 (N_6603,N_545,N_528);
nor U6604 (N_6604,N_3568,N_2068);
nand U6605 (N_6605,N_2097,N_3546);
and U6606 (N_6606,N_1135,N_3118);
or U6607 (N_6607,N_2534,N_1691);
nor U6608 (N_6608,N_1896,N_149);
and U6609 (N_6609,N_2003,N_592);
or U6610 (N_6610,N_2830,N_1817);
or U6611 (N_6611,N_2743,N_1282);
xor U6612 (N_6612,N_916,N_1136);
nand U6613 (N_6613,N_2074,N_2717);
or U6614 (N_6614,N_3680,N_1459);
nand U6615 (N_6615,N_2146,N_805);
or U6616 (N_6616,N_2428,N_2756);
or U6617 (N_6617,N_3571,N_1964);
nor U6618 (N_6618,N_1504,N_886);
nor U6619 (N_6619,N_1253,N_1193);
nor U6620 (N_6620,N_1724,N_341);
and U6621 (N_6621,N_3435,N_3310);
nor U6622 (N_6622,N_2468,N_3455);
nand U6623 (N_6623,N_3243,N_442);
or U6624 (N_6624,N_1114,N_3452);
xnor U6625 (N_6625,N_505,N_1481);
nor U6626 (N_6626,N_1516,N_1995);
nand U6627 (N_6627,N_3628,N_85);
nand U6628 (N_6628,N_1226,N_3180);
xnor U6629 (N_6629,N_2550,N_413);
or U6630 (N_6630,N_2758,N_1662);
or U6631 (N_6631,N_2505,N_2846);
xor U6632 (N_6632,N_133,N_3844);
nor U6633 (N_6633,N_282,N_9);
nor U6634 (N_6634,N_3303,N_3269);
and U6635 (N_6635,N_313,N_1784);
nand U6636 (N_6636,N_122,N_47);
nand U6637 (N_6637,N_2034,N_2121);
nor U6638 (N_6638,N_3818,N_1692);
nand U6639 (N_6639,N_802,N_3112);
nand U6640 (N_6640,N_2801,N_1715);
nand U6641 (N_6641,N_3140,N_3308);
or U6642 (N_6642,N_1668,N_3978);
nor U6643 (N_6643,N_3281,N_1785);
nand U6644 (N_6644,N_1726,N_3237);
xor U6645 (N_6645,N_3874,N_1168);
or U6646 (N_6646,N_3743,N_2264);
nand U6647 (N_6647,N_2612,N_3771);
nand U6648 (N_6648,N_1985,N_492);
nor U6649 (N_6649,N_804,N_1900);
nand U6650 (N_6650,N_3893,N_2222);
nor U6651 (N_6651,N_1311,N_2760);
nand U6652 (N_6652,N_3485,N_1743);
or U6653 (N_6653,N_3536,N_2195);
nand U6654 (N_6654,N_3554,N_3577);
nor U6655 (N_6655,N_2931,N_16);
or U6656 (N_6656,N_1932,N_959);
or U6657 (N_6657,N_3182,N_1697);
and U6658 (N_6658,N_840,N_1393);
nor U6659 (N_6659,N_562,N_3254);
or U6660 (N_6660,N_2729,N_3966);
and U6661 (N_6661,N_1811,N_2311);
or U6662 (N_6662,N_3157,N_466);
nor U6663 (N_6663,N_784,N_207);
nand U6664 (N_6664,N_188,N_1816);
or U6665 (N_6665,N_3236,N_3333);
nand U6666 (N_6666,N_481,N_1046);
and U6667 (N_6667,N_1322,N_1801);
and U6668 (N_6668,N_2483,N_2898);
nor U6669 (N_6669,N_2727,N_1806);
or U6670 (N_6670,N_1023,N_674);
nand U6671 (N_6671,N_2106,N_317);
and U6672 (N_6672,N_1421,N_897);
nor U6673 (N_6673,N_1989,N_3395);
and U6674 (N_6674,N_3991,N_486);
nor U6675 (N_6675,N_2939,N_3043);
nand U6676 (N_6676,N_2965,N_1023);
and U6677 (N_6677,N_3298,N_2529);
nor U6678 (N_6678,N_1494,N_3670);
xnor U6679 (N_6679,N_1373,N_2085);
nor U6680 (N_6680,N_3501,N_1438);
nand U6681 (N_6681,N_664,N_1016);
nor U6682 (N_6682,N_90,N_2874);
and U6683 (N_6683,N_3011,N_604);
nand U6684 (N_6684,N_657,N_1374);
or U6685 (N_6685,N_1271,N_3915);
and U6686 (N_6686,N_3528,N_1787);
and U6687 (N_6687,N_2648,N_301);
and U6688 (N_6688,N_3885,N_1954);
or U6689 (N_6689,N_2402,N_3635);
xnor U6690 (N_6690,N_2587,N_1320);
or U6691 (N_6691,N_3818,N_2438);
and U6692 (N_6692,N_1205,N_2668);
nor U6693 (N_6693,N_949,N_1781);
nor U6694 (N_6694,N_880,N_1665);
nand U6695 (N_6695,N_3388,N_3005);
and U6696 (N_6696,N_1943,N_1194);
and U6697 (N_6697,N_1876,N_50);
nor U6698 (N_6698,N_3174,N_559);
xnor U6699 (N_6699,N_3153,N_1471);
and U6700 (N_6700,N_3844,N_3456);
nand U6701 (N_6701,N_345,N_1974);
or U6702 (N_6702,N_2876,N_1815);
xnor U6703 (N_6703,N_2717,N_3010);
or U6704 (N_6704,N_557,N_342);
nand U6705 (N_6705,N_2792,N_1617);
nor U6706 (N_6706,N_40,N_1743);
nor U6707 (N_6707,N_3246,N_2765);
or U6708 (N_6708,N_2517,N_1050);
and U6709 (N_6709,N_429,N_1678);
nand U6710 (N_6710,N_3245,N_841);
xnor U6711 (N_6711,N_3434,N_1648);
nand U6712 (N_6712,N_2841,N_661);
nand U6713 (N_6713,N_3608,N_285);
xnor U6714 (N_6714,N_1653,N_3500);
or U6715 (N_6715,N_3890,N_2260);
or U6716 (N_6716,N_3604,N_3777);
or U6717 (N_6717,N_3298,N_164);
nand U6718 (N_6718,N_948,N_1793);
nand U6719 (N_6719,N_1877,N_3084);
xor U6720 (N_6720,N_3943,N_31);
nor U6721 (N_6721,N_2093,N_3627);
xor U6722 (N_6722,N_2073,N_3248);
nor U6723 (N_6723,N_1078,N_2150);
nand U6724 (N_6724,N_2678,N_185);
and U6725 (N_6725,N_1188,N_3590);
or U6726 (N_6726,N_99,N_3489);
nand U6727 (N_6727,N_2545,N_1778);
and U6728 (N_6728,N_146,N_713);
nand U6729 (N_6729,N_1411,N_601);
and U6730 (N_6730,N_658,N_1956);
nor U6731 (N_6731,N_1594,N_231);
and U6732 (N_6732,N_718,N_808);
or U6733 (N_6733,N_2426,N_146);
nand U6734 (N_6734,N_2429,N_2311);
nor U6735 (N_6735,N_2449,N_3347);
and U6736 (N_6736,N_3119,N_2669);
xor U6737 (N_6737,N_3547,N_3388);
or U6738 (N_6738,N_3433,N_1794);
xnor U6739 (N_6739,N_3937,N_2097);
and U6740 (N_6740,N_2958,N_1268);
nor U6741 (N_6741,N_3136,N_286);
nor U6742 (N_6742,N_219,N_565);
nor U6743 (N_6743,N_2500,N_1533);
xor U6744 (N_6744,N_392,N_1822);
nand U6745 (N_6745,N_3298,N_1857);
nor U6746 (N_6746,N_1242,N_1442);
nand U6747 (N_6747,N_1976,N_364);
or U6748 (N_6748,N_3430,N_208);
xnor U6749 (N_6749,N_1260,N_1952);
nor U6750 (N_6750,N_2215,N_579);
or U6751 (N_6751,N_1246,N_3180);
or U6752 (N_6752,N_3414,N_2335);
nand U6753 (N_6753,N_1083,N_3265);
and U6754 (N_6754,N_3126,N_2727);
and U6755 (N_6755,N_2988,N_2617);
and U6756 (N_6756,N_1073,N_1239);
or U6757 (N_6757,N_545,N_2593);
or U6758 (N_6758,N_227,N_2483);
nand U6759 (N_6759,N_200,N_1233);
xnor U6760 (N_6760,N_1493,N_172);
nor U6761 (N_6761,N_2176,N_266);
or U6762 (N_6762,N_3905,N_3844);
and U6763 (N_6763,N_1997,N_3770);
nand U6764 (N_6764,N_3661,N_218);
nor U6765 (N_6765,N_2097,N_2474);
nor U6766 (N_6766,N_3087,N_1361);
nand U6767 (N_6767,N_1215,N_1156);
and U6768 (N_6768,N_2547,N_1991);
xnor U6769 (N_6769,N_712,N_1289);
nor U6770 (N_6770,N_628,N_1815);
nor U6771 (N_6771,N_368,N_951);
nand U6772 (N_6772,N_777,N_3578);
nor U6773 (N_6773,N_2915,N_2356);
and U6774 (N_6774,N_2494,N_1598);
and U6775 (N_6775,N_365,N_3826);
nand U6776 (N_6776,N_1102,N_1347);
and U6777 (N_6777,N_3292,N_928);
nand U6778 (N_6778,N_3444,N_364);
or U6779 (N_6779,N_1554,N_1584);
or U6780 (N_6780,N_2906,N_1216);
and U6781 (N_6781,N_3603,N_179);
or U6782 (N_6782,N_582,N_1941);
and U6783 (N_6783,N_1672,N_713);
nor U6784 (N_6784,N_3007,N_1973);
and U6785 (N_6785,N_827,N_31);
nor U6786 (N_6786,N_660,N_1702);
or U6787 (N_6787,N_2439,N_2294);
nand U6788 (N_6788,N_2828,N_3169);
or U6789 (N_6789,N_3179,N_1276);
nor U6790 (N_6790,N_3768,N_3000);
nor U6791 (N_6791,N_1759,N_2415);
xor U6792 (N_6792,N_3707,N_2409);
and U6793 (N_6793,N_731,N_1925);
nand U6794 (N_6794,N_3617,N_2695);
xnor U6795 (N_6795,N_1698,N_3306);
or U6796 (N_6796,N_2540,N_457);
nand U6797 (N_6797,N_2152,N_830);
or U6798 (N_6798,N_449,N_553);
nand U6799 (N_6799,N_2810,N_3897);
nand U6800 (N_6800,N_1751,N_3588);
and U6801 (N_6801,N_2952,N_668);
or U6802 (N_6802,N_3084,N_2327);
xnor U6803 (N_6803,N_3415,N_1732);
nand U6804 (N_6804,N_1414,N_2485);
nand U6805 (N_6805,N_174,N_2606);
xor U6806 (N_6806,N_2247,N_1973);
nor U6807 (N_6807,N_270,N_67);
and U6808 (N_6808,N_1112,N_2485);
or U6809 (N_6809,N_568,N_3791);
and U6810 (N_6810,N_2973,N_1806);
nor U6811 (N_6811,N_1323,N_3110);
and U6812 (N_6812,N_1894,N_1021);
and U6813 (N_6813,N_239,N_1707);
nor U6814 (N_6814,N_2057,N_2073);
and U6815 (N_6815,N_1357,N_2897);
nand U6816 (N_6816,N_2101,N_3757);
nor U6817 (N_6817,N_866,N_531);
nor U6818 (N_6818,N_1864,N_3258);
and U6819 (N_6819,N_3703,N_1731);
or U6820 (N_6820,N_2046,N_3118);
or U6821 (N_6821,N_100,N_729);
nor U6822 (N_6822,N_1680,N_367);
nor U6823 (N_6823,N_777,N_2648);
nor U6824 (N_6824,N_2626,N_336);
and U6825 (N_6825,N_2954,N_775);
nor U6826 (N_6826,N_449,N_1557);
and U6827 (N_6827,N_1166,N_3200);
and U6828 (N_6828,N_2226,N_3776);
xor U6829 (N_6829,N_1284,N_887);
xnor U6830 (N_6830,N_3704,N_2917);
or U6831 (N_6831,N_2682,N_3447);
nand U6832 (N_6832,N_406,N_2952);
nand U6833 (N_6833,N_865,N_1947);
xnor U6834 (N_6834,N_271,N_1091);
and U6835 (N_6835,N_3057,N_985);
nand U6836 (N_6836,N_1908,N_3544);
and U6837 (N_6837,N_399,N_1934);
xnor U6838 (N_6838,N_972,N_3440);
nand U6839 (N_6839,N_253,N_3803);
and U6840 (N_6840,N_1789,N_131);
nand U6841 (N_6841,N_1672,N_1244);
and U6842 (N_6842,N_3049,N_2715);
nand U6843 (N_6843,N_3384,N_3914);
and U6844 (N_6844,N_971,N_1565);
or U6845 (N_6845,N_232,N_3942);
or U6846 (N_6846,N_2377,N_3660);
nand U6847 (N_6847,N_2372,N_3217);
nor U6848 (N_6848,N_3486,N_225);
nor U6849 (N_6849,N_1593,N_476);
or U6850 (N_6850,N_2187,N_2822);
or U6851 (N_6851,N_2571,N_827);
xnor U6852 (N_6852,N_1803,N_3712);
and U6853 (N_6853,N_1251,N_1645);
nor U6854 (N_6854,N_15,N_2711);
nand U6855 (N_6855,N_3893,N_3268);
nor U6856 (N_6856,N_2683,N_38);
nor U6857 (N_6857,N_226,N_187);
nor U6858 (N_6858,N_3330,N_1604);
nand U6859 (N_6859,N_2067,N_2317);
and U6860 (N_6860,N_3368,N_1329);
and U6861 (N_6861,N_3403,N_233);
nand U6862 (N_6862,N_1221,N_2820);
and U6863 (N_6863,N_897,N_1733);
and U6864 (N_6864,N_3260,N_2196);
or U6865 (N_6865,N_263,N_1003);
or U6866 (N_6866,N_1564,N_2989);
and U6867 (N_6867,N_3847,N_3462);
and U6868 (N_6868,N_3065,N_3818);
nor U6869 (N_6869,N_658,N_2125);
or U6870 (N_6870,N_247,N_3286);
nor U6871 (N_6871,N_3337,N_1594);
or U6872 (N_6872,N_2478,N_3010);
and U6873 (N_6873,N_174,N_3638);
and U6874 (N_6874,N_607,N_2664);
or U6875 (N_6875,N_1859,N_900);
nor U6876 (N_6876,N_2985,N_2147);
nor U6877 (N_6877,N_1131,N_1030);
or U6878 (N_6878,N_3173,N_3412);
and U6879 (N_6879,N_3856,N_2637);
or U6880 (N_6880,N_2816,N_3768);
and U6881 (N_6881,N_3170,N_3737);
nor U6882 (N_6882,N_3575,N_3371);
xor U6883 (N_6883,N_1605,N_184);
or U6884 (N_6884,N_3461,N_703);
and U6885 (N_6885,N_1387,N_2437);
and U6886 (N_6886,N_2156,N_2615);
nand U6887 (N_6887,N_389,N_1103);
nand U6888 (N_6888,N_3004,N_2627);
or U6889 (N_6889,N_3389,N_855);
nand U6890 (N_6890,N_1160,N_3555);
xnor U6891 (N_6891,N_3215,N_2165);
nor U6892 (N_6892,N_3853,N_1076);
nor U6893 (N_6893,N_1432,N_122);
and U6894 (N_6894,N_1746,N_2398);
nor U6895 (N_6895,N_2313,N_3500);
nand U6896 (N_6896,N_1146,N_1461);
and U6897 (N_6897,N_513,N_3377);
or U6898 (N_6898,N_351,N_2570);
and U6899 (N_6899,N_143,N_3963);
and U6900 (N_6900,N_947,N_1110);
nor U6901 (N_6901,N_809,N_2587);
and U6902 (N_6902,N_855,N_3791);
and U6903 (N_6903,N_943,N_478);
nor U6904 (N_6904,N_309,N_1585);
or U6905 (N_6905,N_3919,N_1058);
xor U6906 (N_6906,N_2500,N_1280);
and U6907 (N_6907,N_2884,N_877);
nand U6908 (N_6908,N_2317,N_125);
nor U6909 (N_6909,N_3530,N_2462);
or U6910 (N_6910,N_2021,N_1348);
nor U6911 (N_6911,N_3854,N_2947);
nor U6912 (N_6912,N_1361,N_209);
nand U6913 (N_6913,N_2563,N_1436);
and U6914 (N_6914,N_742,N_677);
or U6915 (N_6915,N_2066,N_1406);
or U6916 (N_6916,N_939,N_1673);
and U6917 (N_6917,N_2801,N_1099);
or U6918 (N_6918,N_853,N_1061);
xnor U6919 (N_6919,N_796,N_3269);
or U6920 (N_6920,N_1319,N_3095);
or U6921 (N_6921,N_1462,N_1263);
nand U6922 (N_6922,N_1332,N_2803);
and U6923 (N_6923,N_3584,N_670);
nor U6924 (N_6924,N_1242,N_207);
nor U6925 (N_6925,N_1494,N_2556);
nor U6926 (N_6926,N_1728,N_400);
or U6927 (N_6927,N_1948,N_3092);
xor U6928 (N_6928,N_805,N_3116);
nand U6929 (N_6929,N_3008,N_2257);
and U6930 (N_6930,N_727,N_1008);
xnor U6931 (N_6931,N_562,N_2876);
and U6932 (N_6932,N_1548,N_3891);
or U6933 (N_6933,N_493,N_3060);
and U6934 (N_6934,N_954,N_1417);
nor U6935 (N_6935,N_1230,N_3032);
and U6936 (N_6936,N_608,N_2262);
or U6937 (N_6937,N_687,N_3993);
nand U6938 (N_6938,N_3444,N_1097);
nand U6939 (N_6939,N_3254,N_1864);
or U6940 (N_6940,N_1081,N_2094);
and U6941 (N_6941,N_2828,N_1688);
and U6942 (N_6942,N_1899,N_1702);
nand U6943 (N_6943,N_2899,N_2171);
nor U6944 (N_6944,N_2331,N_683);
nand U6945 (N_6945,N_282,N_3451);
nor U6946 (N_6946,N_3180,N_399);
and U6947 (N_6947,N_3165,N_1525);
xor U6948 (N_6948,N_3511,N_1903);
or U6949 (N_6949,N_3836,N_2493);
or U6950 (N_6950,N_1781,N_1954);
xnor U6951 (N_6951,N_493,N_3329);
or U6952 (N_6952,N_3495,N_1416);
and U6953 (N_6953,N_34,N_1930);
nor U6954 (N_6954,N_3010,N_1602);
xnor U6955 (N_6955,N_3088,N_655);
or U6956 (N_6956,N_3664,N_1474);
nor U6957 (N_6957,N_968,N_3993);
and U6958 (N_6958,N_3656,N_3523);
nand U6959 (N_6959,N_2052,N_1035);
or U6960 (N_6960,N_1441,N_2167);
nor U6961 (N_6961,N_3921,N_3510);
and U6962 (N_6962,N_776,N_1693);
xnor U6963 (N_6963,N_2118,N_1359);
or U6964 (N_6964,N_2224,N_1723);
nand U6965 (N_6965,N_1733,N_2688);
nand U6966 (N_6966,N_721,N_655);
and U6967 (N_6967,N_562,N_3279);
nor U6968 (N_6968,N_218,N_2563);
and U6969 (N_6969,N_3443,N_1403);
nor U6970 (N_6970,N_1701,N_443);
and U6971 (N_6971,N_1829,N_2190);
nor U6972 (N_6972,N_2227,N_1479);
xnor U6973 (N_6973,N_2786,N_2147);
and U6974 (N_6974,N_1837,N_516);
nand U6975 (N_6975,N_3167,N_3420);
nand U6976 (N_6976,N_1492,N_762);
or U6977 (N_6977,N_3052,N_1453);
or U6978 (N_6978,N_1047,N_572);
or U6979 (N_6979,N_3277,N_299);
or U6980 (N_6980,N_1895,N_3051);
and U6981 (N_6981,N_3010,N_1029);
or U6982 (N_6982,N_1633,N_3193);
nand U6983 (N_6983,N_323,N_543);
nand U6984 (N_6984,N_3156,N_1066);
and U6985 (N_6985,N_1305,N_143);
or U6986 (N_6986,N_3071,N_3365);
nor U6987 (N_6987,N_3265,N_306);
nand U6988 (N_6988,N_2253,N_2725);
xnor U6989 (N_6989,N_632,N_992);
nor U6990 (N_6990,N_2424,N_3017);
nor U6991 (N_6991,N_640,N_377);
xor U6992 (N_6992,N_1449,N_3155);
nand U6993 (N_6993,N_1731,N_3984);
nor U6994 (N_6994,N_722,N_2660);
xor U6995 (N_6995,N_3268,N_809);
xor U6996 (N_6996,N_2362,N_2257);
or U6997 (N_6997,N_1113,N_2132);
nand U6998 (N_6998,N_2990,N_2446);
nand U6999 (N_6999,N_1397,N_1574);
xor U7000 (N_7000,N_224,N_3908);
or U7001 (N_7001,N_540,N_3526);
xnor U7002 (N_7002,N_1461,N_2775);
or U7003 (N_7003,N_3904,N_933);
nor U7004 (N_7004,N_1738,N_1888);
and U7005 (N_7005,N_3817,N_2135);
nand U7006 (N_7006,N_1816,N_3844);
nand U7007 (N_7007,N_906,N_3993);
and U7008 (N_7008,N_793,N_839);
or U7009 (N_7009,N_346,N_198);
xnor U7010 (N_7010,N_904,N_3711);
nor U7011 (N_7011,N_637,N_1614);
nor U7012 (N_7012,N_150,N_420);
or U7013 (N_7013,N_3572,N_3606);
or U7014 (N_7014,N_2504,N_1199);
nand U7015 (N_7015,N_2721,N_503);
nand U7016 (N_7016,N_3655,N_3795);
or U7017 (N_7017,N_2458,N_1046);
nand U7018 (N_7018,N_885,N_190);
and U7019 (N_7019,N_378,N_156);
and U7020 (N_7020,N_3103,N_54);
and U7021 (N_7021,N_1216,N_587);
xor U7022 (N_7022,N_974,N_2979);
xnor U7023 (N_7023,N_3465,N_2034);
nor U7024 (N_7024,N_341,N_2280);
nand U7025 (N_7025,N_1084,N_2904);
or U7026 (N_7026,N_3521,N_227);
nor U7027 (N_7027,N_393,N_1935);
and U7028 (N_7028,N_3854,N_1287);
nor U7029 (N_7029,N_3912,N_3871);
or U7030 (N_7030,N_3935,N_1516);
or U7031 (N_7031,N_3886,N_2847);
nor U7032 (N_7032,N_413,N_345);
nand U7033 (N_7033,N_236,N_3343);
and U7034 (N_7034,N_3690,N_16);
or U7035 (N_7035,N_2674,N_3975);
nor U7036 (N_7036,N_1960,N_1002);
nand U7037 (N_7037,N_2002,N_3346);
nand U7038 (N_7038,N_2664,N_2706);
and U7039 (N_7039,N_828,N_3918);
nor U7040 (N_7040,N_1875,N_3283);
and U7041 (N_7041,N_3825,N_2138);
nand U7042 (N_7042,N_1175,N_406);
and U7043 (N_7043,N_1901,N_1755);
or U7044 (N_7044,N_3291,N_3035);
nor U7045 (N_7045,N_3061,N_1119);
nor U7046 (N_7046,N_2723,N_3019);
nor U7047 (N_7047,N_1282,N_2067);
and U7048 (N_7048,N_3356,N_2296);
nand U7049 (N_7049,N_2867,N_2054);
xnor U7050 (N_7050,N_3286,N_620);
or U7051 (N_7051,N_3121,N_2663);
and U7052 (N_7052,N_1040,N_1702);
and U7053 (N_7053,N_1233,N_3025);
nand U7054 (N_7054,N_951,N_2465);
or U7055 (N_7055,N_3490,N_2800);
nor U7056 (N_7056,N_185,N_991);
and U7057 (N_7057,N_1059,N_365);
and U7058 (N_7058,N_1839,N_781);
and U7059 (N_7059,N_2581,N_457);
and U7060 (N_7060,N_1522,N_1506);
nor U7061 (N_7061,N_295,N_752);
or U7062 (N_7062,N_1906,N_1539);
nand U7063 (N_7063,N_606,N_2474);
and U7064 (N_7064,N_1594,N_1318);
or U7065 (N_7065,N_3778,N_3640);
nand U7066 (N_7066,N_3222,N_3755);
nand U7067 (N_7067,N_1123,N_803);
nand U7068 (N_7068,N_3025,N_3241);
and U7069 (N_7069,N_3139,N_1178);
nand U7070 (N_7070,N_2452,N_1437);
xor U7071 (N_7071,N_497,N_577);
xnor U7072 (N_7072,N_2933,N_528);
and U7073 (N_7073,N_2189,N_996);
nand U7074 (N_7074,N_223,N_1444);
and U7075 (N_7075,N_761,N_1989);
and U7076 (N_7076,N_3676,N_2422);
xor U7077 (N_7077,N_2328,N_1984);
and U7078 (N_7078,N_2890,N_1151);
or U7079 (N_7079,N_330,N_3952);
and U7080 (N_7080,N_3347,N_489);
and U7081 (N_7081,N_3843,N_1563);
nand U7082 (N_7082,N_798,N_3926);
xor U7083 (N_7083,N_1098,N_3177);
or U7084 (N_7084,N_2320,N_2484);
or U7085 (N_7085,N_2474,N_3561);
or U7086 (N_7086,N_679,N_2873);
or U7087 (N_7087,N_1307,N_1487);
nor U7088 (N_7088,N_343,N_2758);
xor U7089 (N_7089,N_1822,N_906);
or U7090 (N_7090,N_1888,N_131);
nand U7091 (N_7091,N_49,N_491);
nor U7092 (N_7092,N_1826,N_3733);
or U7093 (N_7093,N_944,N_1851);
nor U7094 (N_7094,N_3972,N_3562);
nand U7095 (N_7095,N_3396,N_1146);
nor U7096 (N_7096,N_1679,N_1179);
nor U7097 (N_7097,N_2004,N_3842);
nand U7098 (N_7098,N_721,N_2790);
nor U7099 (N_7099,N_3507,N_2914);
xnor U7100 (N_7100,N_1404,N_3784);
nor U7101 (N_7101,N_3347,N_1245);
nor U7102 (N_7102,N_1574,N_3689);
and U7103 (N_7103,N_1215,N_1002);
or U7104 (N_7104,N_914,N_3563);
xor U7105 (N_7105,N_303,N_3188);
xnor U7106 (N_7106,N_3403,N_3923);
and U7107 (N_7107,N_2590,N_1185);
nand U7108 (N_7108,N_3223,N_1309);
or U7109 (N_7109,N_1347,N_2937);
xor U7110 (N_7110,N_3693,N_1807);
and U7111 (N_7111,N_845,N_321);
nand U7112 (N_7112,N_414,N_1651);
and U7113 (N_7113,N_757,N_2739);
or U7114 (N_7114,N_2856,N_2300);
nand U7115 (N_7115,N_3786,N_586);
and U7116 (N_7116,N_1010,N_1645);
xnor U7117 (N_7117,N_1178,N_482);
nor U7118 (N_7118,N_3282,N_3983);
nor U7119 (N_7119,N_1819,N_3522);
and U7120 (N_7120,N_3756,N_2394);
or U7121 (N_7121,N_1540,N_3401);
nor U7122 (N_7122,N_1470,N_2782);
xnor U7123 (N_7123,N_861,N_1296);
or U7124 (N_7124,N_3067,N_180);
xnor U7125 (N_7125,N_1012,N_556);
xnor U7126 (N_7126,N_8,N_3766);
nor U7127 (N_7127,N_1488,N_3777);
and U7128 (N_7128,N_3769,N_3756);
and U7129 (N_7129,N_2425,N_1554);
and U7130 (N_7130,N_2128,N_3125);
nor U7131 (N_7131,N_2291,N_417);
nor U7132 (N_7132,N_2807,N_675);
and U7133 (N_7133,N_3456,N_776);
and U7134 (N_7134,N_1683,N_3687);
nand U7135 (N_7135,N_2046,N_2122);
and U7136 (N_7136,N_2838,N_2466);
nor U7137 (N_7137,N_1228,N_3445);
or U7138 (N_7138,N_2481,N_2768);
or U7139 (N_7139,N_3232,N_115);
and U7140 (N_7140,N_3824,N_3689);
xor U7141 (N_7141,N_3424,N_1995);
and U7142 (N_7142,N_645,N_2020);
nand U7143 (N_7143,N_1535,N_563);
nor U7144 (N_7144,N_240,N_423);
nand U7145 (N_7145,N_2135,N_3482);
or U7146 (N_7146,N_2833,N_2621);
and U7147 (N_7147,N_545,N_1556);
nand U7148 (N_7148,N_2821,N_576);
nor U7149 (N_7149,N_2373,N_3005);
and U7150 (N_7150,N_1944,N_465);
nor U7151 (N_7151,N_681,N_2088);
nor U7152 (N_7152,N_743,N_935);
nand U7153 (N_7153,N_353,N_3532);
and U7154 (N_7154,N_3257,N_2036);
or U7155 (N_7155,N_635,N_2067);
xnor U7156 (N_7156,N_1389,N_1217);
and U7157 (N_7157,N_2241,N_181);
xnor U7158 (N_7158,N_2381,N_2473);
and U7159 (N_7159,N_37,N_2050);
and U7160 (N_7160,N_3462,N_388);
xnor U7161 (N_7161,N_176,N_617);
and U7162 (N_7162,N_2696,N_2689);
nor U7163 (N_7163,N_1725,N_1271);
xor U7164 (N_7164,N_3007,N_2334);
nand U7165 (N_7165,N_1912,N_3899);
and U7166 (N_7166,N_1689,N_3985);
nand U7167 (N_7167,N_3323,N_520);
and U7168 (N_7168,N_2162,N_2302);
and U7169 (N_7169,N_1686,N_1846);
xor U7170 (N_7170,N_2732,N_3201);
nand U7171 (N_7171,N_2027,N_3019);
or U7172 (N_7172,N_2804,N_2290);
and U7173 (N_7173,N_3124,N_421);
and U7174 (N_7174,N_2434,N_872);
nor U7175 (N_7175,N_619,N_2304);
nor U7176 (N_7176,N_1198,N_1161);
and U7177 (N_7177,N_136,N_3776);
or U7178 (N_7178,N_1821,N_1602);
nor U7179 (N_7179,N_2794,N_113);
nor U7180 (N_7180,N_1523,N_650);
and U7181 (N_7181,N_2063,N_1879);
and U7182 (N_7182,N_1709,N_411);
xnor U7183 (N_7183,N_2309,N_1822);
nor U7184 (N_7184,N_1514,N_2489);
or U7185 (N_7185,N_2247,N_443);
or U7186 (N_7186,N_3310,N_2074);
and U7187 (N_7187,N_1412,N_3226);
nor U7188 (N_7188,N_498,N_1882);
and U7189 (N_7189,N_2477,N_1392);
and U7190 (N_7190,N_3496,N_511);
nand U7191 (N_7191,N_466,N_686);
nor U7192 (N_7192,N_2524,N_1462);
and U7193 (N_7193,N_124,N_3793);
or U7194 (N_7194,N_476,N_1933);
nand U7195 (N_7195,N_1654,N_3613);
nor U7196 (N_7196,N_2838,N_1144);
and U7197 (N_7197,N_2662,N_3754);
or U7198 (N_7198,N_2528,N_2407);
nor U7199 (N_7199,N_2746,N_1837);
nor U7200 (N_7200,N_2141,N_1252);
and U7201 (N_7201,N_685,N_1961);
or U7202 (N_7202,N_668,N_2349);
and U7203 (N_7203,N_32,N_2575);
nand U7204 (N_7204,N_1546,N_3854);
nor U7205 (N_7205,N_3988,N_2099);
or U7206 (N_7206,N_890,N_1086);
and U7207 (N_7207,N_1505,N_1829);
or U7208 (N_7208,N_3200,N_1759);
or U7209 (N_7209,N_1399,N_2000);
nor U7210 (N_7210,N_711,N_646);
and U7211 (N_7211,N_1009,N_3050);
nand U7212 (N_7212,N_3880,N_3891);
nand U7213 (N_7213,N_3225,N_3095);
nand U7214 (N_7214,N_3375,N_1072);
nor U7215 (N_7215,N_497,N_2670);
and U7216 (N_7216,N_115,N_1499);
and U7217 (N_7217,N_3082,N_3779);
nand U7218 (N_7218,N_818,N_1427);
xnor U7219 (N_7219,N_3192,N_2105);
nor U7220 (N_7220,N_1371,N_329);
xor U7221 (N_7221,N_1310,N_1406);
nand U7222 (N_7222,N_167,N_2675);
nand U7223 (N_7223,N_2501,N_3262);
and U7224 (N_7224,N_2198,N_45);
or U7225 (N_7225,N_1363,N_117);
nor U7226 (N_7226,N_3885,N_2937);
nor U7227 (N_7227,N_681,N_1626);
xor U7228 (N_7228,N_3865,N_2247);
nor U7229 (N_7229,N_2325,N_2106);
and U7230 (N_7230,N_465,N_1895);
nand U7231 (N_7231,N_1686,N_932);
or U7232 (N_7232,N_1776,N_2328);
nand U7233 (N_7233,N_1831,N_268);
or U7234 (N_7234,N_461,N_25);
xnor U7235 (N_7235,N_2683,N_750);
and U7236 (N_7236,N_3741,N_3541);
nand U7237 (N_7237,N_3466,N_1265);
nand U7238 (N_7238,N_2133,N_1457);
and U7239 (N_7239,N_116,N_3681);
and U7240 (N_7240,N_1006,N_118);
nand U7241 (N_7241,N_1138,N_3959);
and U7242 (N_7242,N_871,N_910);
nor U7243 (N_7243,N_1066,N_3786);
nor U7244 (N_7244,N_3724,N_2964);
nand U7245 (N_7245,N_1321,N_1625);
nor U7246 (N_7246,N_1200,N_2745);
nand U7247 (N_7247,N_1318,N_2225);
and U7248 (N_7248,N_1370,N_3597);
or U7249 (N_7249,N_898,N_1838);
nand U7250 (N_7250,N_1466,N_2010);
or U7251 (N_7251,N_1117,N_552);
nor U7252 (N_7252,N_2297,N_3219);
or U7253 (N_7253,N_2672,N_2962);
nor U7254 (N_7254,N_2270,N_1677);
or U7255 (N_7255,N_3950,N_2003);
nor U7256 (N_7256,N_2281,N_762);
nor U7257 (N_7257,N_1354,N_749);
nor U7258 (N_7258,N_2889,N_437);
nand U7259 (N_7259,N_1473,N_427);
nor U7260 (N_7260,N_3127,N_3302);
nor U7261 (N_7261,N_3847,N_3911);
nand U7262 (N_7262,N_330,N_2649);
nand U7263 (N_7263,N_2038,N_1380);
nor U7264 (N_7264,N_2039,N_1555);
and U7265 (N_7265,N_321,N_2816);
and U7266 (N_7266,N_1729,N_3817);
and U7267 (N_7267,N_1736,N_2907);
and U7268 (N_7268,N_3375,N_1261);
nor U7269 (N_7269,N_2517,N_2994);
nand U7270 (N_7270,N_1740,N_70);
nor U7271 (N_7271,N_1743,N_1117);
or U7272 (N_7272,N_2454,N_977);
and U7273 (N_7273,N_3710,N_2589);
and U7274 (N_7274,N_1639,N_2932);
nor U7275 (N_7275,N_2232,N_3990);
and U7276 (N_7276,N_3726,N_1249);
or U7277 (N_7277,N_3272,N_3038);
or U7278 (N_7278,N_801,N_524);
nand U7279 (N_7279,N_472,N_646);
nand U7280 (N_7280,N_3552,N_505);
and U7281 (N_7281,N_820,N_3537);
or U7282 (N_7282,N_2032,N_930);
or U7283 (N_7283,N_1682,N_27);
xnor U7284 (N_7284,N_2156,N_1041);
nor U7285 (N_7285,N_1121,N_501);
and U7286 (N_7286,N_3407,N_2544);
or U7287 (N_7287,N_3272,N_2639);
and U7288 (N_7288,N_2115,N_632);
or U7289 (N_7289,N_2784,N_3347);
nand U7290 (N_7290,N_3650,N_911);
or U7291 (N_7291,N_416,N_3249);
xnor U7292 (N_7292,N_3316,N_1596);
nand U7293 (N_7293,N_2014,N_3139);
or U7294 (N_7294,N_1416,N_3952);
and U7295 (N_7295,N_735,N_2723);
and U7296 (N_7296,N_773,N_3440);
or U7297 (N_7297,N_2382,N_3039);
nor U7298 (N_7298,N_132,N_0);
or U7299 (N_7299,N_1125,N_281);
nand U7300 (N_7300,N_2679,N_819);
and U7301 (N_7301,N_1177,N_1152);
and U7302 (N_7302,N_3230,N_3488);
and U7303 (N_7303,N_1498,N_3226);
nand U7304 (N_7304,N_225,N_237);
nand U7305 (N_7305,N_2476,N_3141);
or U7306 (N_7306,N_3327,N_3360);
xor U7307 (N_7307,N_3633,N_1907);
and U7308 (N_7308,N_3342,N_3914);
nor U7309 (N_7309,N_1761,N_1246);
nand U7310 (N_7310,N_349,N_663);
or U7311 (N_7311,N_3937,N_2761);
or U7312 (N_7312,N_799,N_878);
and U7313 (N_7313,N_1637,N_3339);
nand U7314 (N_7314,N_910,N_1124);
nor U7315 (N_7315,N_511,N_2121);
and U7316 (N_7316,N_1323,N_134);
and U7317 (N_7317,N_65,N_1543);
nor U7318 (N_7318,N_107,N_3718);
and U7319 (N_7319,N_2064,N_2519);
and U7320 (N_7320,N_1265,N_1048);
and U7321 (N_7321,N_2532,N_3554);
and U7322 (N_7322,N_2476,N_331);
and U7323 (N_7323,N_1994,N_1046);
or U7324 (N_7324,N_2564,N_1767);
xnor U7325 (N_7325,N_429,N_944);
xnor U7326 (N_7326,N_1382,N_3056);
or U7327 (N_7327,N_2892,N_2332);
nand U7328 (N_7328,N_24,N_2262);
nor U7329 (N_7329,N_992,N_798);
and U7330 (N_7330,N_3719,N_382);
and U7331 (N_7331,N_1837,N_2654);
nand U7332 (N_7332,N_1484,N_1810);
or U7333 (N_7333,N_1450,N_2900);
and U7334 (N_7334,N_1382,N_1069);
nand U7335 (N_7335,N_1695,N_1152);
or U7336 (N_7336,N_1684,N_2346);
nand U7337 (N_7337,N_3451,N_2605);
nor U7338 (N_7338,N_1453,N_1544);
xnor U7339 (N_7339,N_1641,N_1753);
and U7340 (N_7340,N_3757,N_464);
xor U7341 (N_7341,N_2816,N_1364);
or U7342 (N_7342,N_2117,N_270);
nand U7343 (N_7343,N_1119,N_288);
or U7344 (N_7344,N_1171,N_2816);
nor U7345 (N_7345,N_3319,N_1270);
or U7346 (N_7346,N_949,N_2002);
or U7347 (N_7347,N_2449,N_3368);
and U7348 (N_7348,N_2415,N_3955);
nor U7349 (N_7349,N_3667,N_97);
or U7350 (N_7350,N_3701,N_236);
nor U7351 (N_7351,N_711,N_1491);
or U7352 (N_7352,N_170,N_1149);
xnor U7353 (N_7353,N_1185,N_2477);
xnor U7354 (N_7354,N_2879,N_1330);
and U7355 (N_7355,N_1004,N_1080);
or U7356 (N_7356,N_2520,N_2842);
nand U7357 (N_7357,N_1221,N_3335);
or U7358 (N_7358,N_634,N_1817);
or U7359 (N_7359,N_191,N_2562);
nand U7360 (N_7360,N_433,N_3484);
nand U7361 (N_7361,N_1852,N_1094);
nor U7362 (N_7362,N_3848,N_1714);
nor U7363 (N_7363,N_3302,N_3344);
nor U7364 (N_7364,N_2563,N_1320);
xnor U7365 (N_7365,N_1406,N_3001);
and U7366 (N_7366,N_2643,N_2209);
and U7367 (N_7367,N_6,N_316);
nor U7368 (N_7368,N_3282,N_952);
nand U7369 (N_7369,N_3105,N_809);
and U7370 (N_7370,N_2538,N_2665);
or U7371 (N_7371,N_1086,N_2857);
nor U7372 (N_7372,N_1310,N_1593);
nand U7373 (N_7373,N_536,N_300);
and U7374 (N_7374,N_2275,N_1794);
and U7375 (N_7375,N_535,N_3038);
nand U7376 (N_7376,N_2109,N_1772);
and U7377 (N_7377,N_2899,N_3783);
xor U7378 (N_7378,N_1184,N_1054);
or U7379 (N_7379,N_1430,N_2051);
xor U7380 (N_7380,N_1036,N_2762);
nor U7381 (N_7381,N_2398,N_319);
and U7382 (N_7382,N_3964,N_1330);
nand U7383 (N_7383,N_1970,N_3820);
or U7384 (N_7384,N_2860,N_1306);
and U7385 (N_7385,N_1582,N_2745);
xnor U7386 (N_7386,N_1875,N_521);
and U7387 (N_7387,N_2648,N_2078);
or U7388 (N_7388,N_1691,N_490);
nor U7389 (N_7389,N_311,N_3072);
and U7390 (N_7390,N_3326,N_526);
and U7391 (N_7391,N_1363,N_1679);
xor U7392 (N_7392,N_58,N_1347);
nor U7393 (N_7393,N_2574,N_1821);
and U7394 (N_7394,N_436,N_2759);
or U7395 (N_7395,N_805,N_2992);
and U7396 (N_7396,N_3589,N_2387);
and U7397 (N_7397,N_307,N_2382);
and U7398 (N_7398,N_1160,N_767);
or U7399 (N_7399,N_589,N_3043);
nand U7400 (N_7400,N_435,N_1587);
and U7401 (N_7401,N_2745,N_1416);
nand U7402 (N_7402,N_3906,N_3232);
and U7403 (N_7403,N_456,N_2305);
nand U7404 (N_7404,N_3,N_1903);
nand U7405 (N_7405,N_2921,N_524);
or U7406 (N_7406,N_3365,N_274);
nor U7407 (N_7407,N_194,N_500);
or U7408 (N_7408,N_1415,N_1522);
and U7409 (N_7409,N_784,N_3862);
or U7410 (N_7410,N_2740,N_335);
nand U7411 (N_7411,N_561,N_3002);
nand U7412 (N_7412,N_2701,N_554);
or U7413 (N_7413,N_3393,N_2931);
or U7414 (N_7414,N_3011,N_3914);
and U7415 (N_7415,N_1697,N_2855);
nand U7416 (N_7416,N_2976,N_2080);
nor U7417 (N_7417,N_182,N_2649);
nor U7418 (N_7418,N_3557,N_3380);
or U7419 (N_7419,N_470,N_1937);
nand U7420 (N_7420,N_652,N_164);
nor U7421 (N_7421,N_2476,N_2670);
nor U7422 (N_7422,N_2960,N_3022);
or U7423 (N_7423,N_3385,N_2430);
nand U7424 (N_7424,N_2823,N_3940);
or U7425 (N_7425,N_411,N_3985);
nand U7426 (N_7426,N_1607,N_348);
xnor U7427 (N_7427,N_1744,N_647);
nor U7428 (N_7428,N_2347,N_259);
or U7429 (N_7429,N_2390,N_1757);
nand U7430 (N_7430,N_1670,N_649);
or U7431 (N_7431,N_2127,N_655);
or U7432 (N_7432,N_1356,N_1593);
or U7433 (N_7433,N_3648,N_2341);
nor U7434 (N_7434,N_220,N_3805);
or U7435 (N_7435,N_2839,N_3152);
nor U7436 (N_7436,N_1424,N_1505);
nor U7437 (N_7437,N_3056,N_345);
nor U7438 (N_7438,N_2864,N_753);
nand U7439 (N_7439,N_1724,N_1583);
nor U7440 (N_7440,N_3037,N_2529);
and U7441 (N_7441,N_269,N_81);
xnor U7442 (N_7442,N_3986,N_1848);
nand U7443 (N_7443,N_2779,N_327);
and U7444 (N_7444,N_3042,N_2484);
nand U7445 (N_7445,N_516,N_1729);
or U7446 (N_7446,N_3643,N_2384);
or U7447 (N_7447,N_439,N_154);
or U7448 (N_7448,N_3490,N_1957);
nor U7449 (N_7449,N_2606,N_1947);
nand U7450 (N_7450,N_3520,N_692);
nand U7451 (N_7451,N_2505,N_1998);
nor U7452 (N_7452,N_508,N_906);
or U7453 (N_7453,N_1788,N_960);
nor U7454 (N_7454,N_1448,N_3612);
nor U7455 (N_7455,N_6,N_2386);
nand U7456 (N_7456,N_1138,N_797);
nand U7457 (N_7457,N_947,N_404);
xor U7458 (N_7458,N_2919,N_2157);
and U7459 (N_7459,N_3183,N_3384);
or U7460 (N_7460,N_2484,N_1178);
nand U7461 (N_7461,N_64,N_1534);
nand U7462 (N_7462,N_3352,N_1220);
and U7463 (N_7463,N_3384,N_3171);
nand U7464 (N_7464,N_2917,N_2728);
nor U7465 (N_7465,N_1575,N_2475);
and U7466 (N_7466,N_3274,N_455);
nor U7467 (N_7467,N_3220,N_1251);
or U7468 (N_7468,N_843,N_1454);
and U7469 (N_7469,N_2332,N_723);
and U7470 (N_7470,N_3458,N_1089);
xnor U7471 (N_7471,N_2540,N_2832);
and U7472 (N_7472,N_1312,N_2062);
xnor U7473 (N_7473,N_3095,N_1102);
or U7474 (N_7474,N_791,N_3098);
or U7475 (N_7475,N_2145,N_1392);
nor U7476 (N_7476,N_2405,N_2430);
and U7477 (N_7477,N_3416,N_981);
xor U7478 (N_7478,N_345,N_1152);
and U7479 (N_7479,N_1888,N_1394);
or U7480 (N_7480,N_3258,N_1839);
and U7481 (N_7481,N_2839,N_3305);
nand U7482 (N_7482,N_3088,N_2032);
xnor U7483 (N_7483,N_1842,N_2073);
nand U7484 (N_7484,N_3495,N_3382);
xnor U7485 (N_7485,N_276,N_3938);
or U7486 (N_7486,N_2680,N_2002);
nand U7487 (N_7487,N_3201,N_1007);
and U7488 (N_7488,N_3224,N_1068);
nand U7489 (N_7489,N_178,N_3242);
nand U7490 (N_7490,N_2733,N_3215);
and U7491 (N_7491,N_1000,N_2350);
nor U7492 (N_7492,N_332,N_2877);
xnor U7493 (N_7493,N_631,N_1382);
and U7494 (N_7494,N_444,N_865);
xnor U7495 (N_7495,N_1799,N_76);
and U7496 (N_7496,N_2064,N_2165);
and U7497 (N_7497,N_3096,N_2970);
and U7498 (N_7498,N_2725,N_758);
and U7499 (N_7499,N_3925,N_2176);
and U7500 (N_7500,N_1320,N_3912);
and U7501 (N_7501,N_2113,N_977);
nand U7502 (N_7502,N_3317,N_1168);
and U7503 (N_7503,N_597,N_2428);
or U7504 (N_7504,N_459,N_2813);
and U7505 (N_7505,N_946,N_2492);
and U7506 (N_7506,N_1061,N_1410);
nand U7507 (N_7507,N_662,N_374);
nand U7508 (N_7508,N_989,N_3823);
and U7509 (N_7509,N_2106,N_683);
nand U7510 (N_7510,N_1052,N_820);
and U7511 (N_7511,N_520,N_2786);
or U7512 (N_7512,N_38,N_3045);
and U7513 (N_7513,N_3633,N_50);
nand U7514 (N_7514,N_528,N_3931);
nor U7515 (N_7515,N_731,N_3622);
nand U7516 (N_7516,N_2785,N_1916);
nand U7517 (N_7517,N_836,N_3053);
nor U7518 (N_7518,N_3646,N_3598);
xor U7519 (N_7519,N_404,N_1004);
or U7520 (N_7520,N_2523,N_3732);
and U7521 (N_7521,N_2382,N_3229);
nand U7522 (N_7522,N_427,N_2076);
and U7523 (N_7523,N_3806,N_1266);
and U7524 (N_7524,N_3190,N_1875);
or U7525 (N_7525,N_2617,N_618);
nand U7526 (N_7526,N_2647,N_2683);
or U7527 (N_7527,N_2043,N_1638);
nor U7528 (N_7528,N_3908,N_1094);
nor U7529 (N_7529,N_1819,N_3992);
nand U7530 (N_7530,N_1509,N_3294);
nor U7531 (N_7531,N_2723,N_167);
or U7532 (N_7532,N_3066,N_2643);
nor U7533 (N_7533,N_2015,N_1396);
or U7534 (N_7534,N_3074,N_3949);
or U7535 (N_7535,N_40,N_2396);
nand U7536 (N_7536,N_2668,N_343);
nand U7537 (N_7537,N_3061,N_293);
or U7538 (N_7538,N_3133,N_3343);
xor U7539 (N_7539,N_2101,N_10);
nand U7540 (N_7540,N_2781,N_764);
nor U7541 (N_7541,N_2054,N_1274);
and U7542 (N_7542,N_3486,N_1819);
nor U7543 (N_7543,N_512,N_2884);
nor U7544 (N_7544,N_683,N_82);
nand U7545 (N_7545,N_3992,N_2265);
and U7546 (N_7546,N_3362,N_2009);
nand U7547 (N_7547,N_3640,N_3461);
or U7548 (N_7548,N_1492,N_1227);
xnor U7549 (N_7549,N_2938,N_606);
and U7550 (N_7550,N_3211,N_2582);
nand U7551 (N_7551,N_3205,N_2827);
or U7552 (N_7552,N_554,N_2416);
nor U7553 (N_7553,N_2510,N_2698);
nand U7554 (N_7554,N_2311,N_2399);
xor U7555 (N_7555,N_1245,N_2817);
and U7556 (N_7556,N_3169,N_2864);
and U7557 (N_7557,N_316,N_3851);
and U7558 (N_7558,N_652,N_1660);
or U7559 (N_7559,N_2099,N_2954);
and U7560 (N_7560,N_71,N_3407);
nand U7561 (N_7561,N_3943,N_3542);
xnor U7562 (N_7562,N_3818,N_3903);
nand U7563 (N_7563,N_2169,N_1506);
nor U7564 (N_7564,N_75,N_1619);
nand U7565 (N_7565,N_2297,N_2838);
nand U7566 (N_7566,N_318,N_1863);
xor U7567 (N_7567,N_2809,N_2046);
or U7568 (N_7568,N_269,N_3871);
nor U7569 (N_7569,N_2182,N_3481);
xnor U7570 (N_7570,N_128,N_3753);
or U7571 (N_7571,N_430,N_3199);
and U7572 (N_7572,N_1821,N_3138);
nor U7573 (N_7573,N_2513,N_133);
nand U7574 (N_7574,N_1371,N_2899);
or U7575 (N_7575,N_2007,N_150);
and U7576 (N_7576,N_1535,N_3238);
nand U7577 (N_7577,N_3701,N_2693);
and U7578 (N_7578,N_2094,N_840);
or U7579 (N_7579,N_1759,N_89);
nor U7580 (N_7580,N_1951,N_3079);
nand U7581 (N_7581,N_3766,N_704);
and U7582 (N_7582,N_3980,N_794);
xor U7583 (N_7583,N_1441,N_3667);
and U7584 (N_7584,N_2949,N_562);
nor U7585 (N_7585,N_1648,N_501);
nand U7586 (N_7586,N_2126,N_772);
nand U7587 (N_7587,N_3267,N_3596);
or U7588 (N_7588,N_2586,N_1480);
and U7589 (N_7589,N_978,N_110);
nor U7590 (N_7590,N_2782,N_3779);
xor U7591 (N_7591,N_595,N_2654);
and U7592 (N_7592,N_388,N_2776);
and U7593 (N_7593,N_2160,N_1228);
and U7594 (N_7594,N_3915,N_3367);
nor U7595 (N_7595,N_1256,N_369);
nand U7596 (N_7596,N_3635,N_2394);
or U7597 (N_7597,N_2395,N_1072);
xor U7598 (N_7598,N_3583,N_1077);
nand U7599 (N_7599,N_1618,N_1644);
and U7600 (N_7600,N_2280,N_3922);
xnor U7601 (N_7601,N_1795,N_3073);
nor U7602 (N_7602,N_3794,N_3311);
nor U7603 (N_7603,N_2187,N_2534);
nand U7604 (N_7604,N_2818,N_3247);
nor U7605 (N_7605,N_2584,N_3508);
and U7606 (N_7606,N_1551,N_910);
and U7607 (N_7607,N_658,N_3606);
and U7608 (N_7608,N_954,N_1715);
nand U7609 (N_7609,N_2216,N_1533);
or U7610 (N_7610,N_2731,N_966);
and U7611 (N_7611,N_3139,N_768);
or U7612 (N_7612,N_3505,N_2825);
nand U7613 (N_7613,N_2312,N_3458);
nand U7614 (N_7614,N_1128,N_2901);
nor U7615 (N_7615,N_1121,N_1564);
nand U7616 (N_7616,N_707,N_2548);
nor U7617 (N_7617,N_1945,N_451);
and U7618 (N_7618,N_1285,N_2618);
and U7619 (N_7619,N_1422,N_3341);
nand U7620 (N_7620,N_665,N_2371);
and U7621 (N_7621,N_2553,N_2726);
nor U7622 (N_7622,N_427,N_548);
nand U7623 (N_7623,N_1593,N_2536);
or U7624 (N_7624,N_2939,N_3527);
xnor U7625 (N_7625,N_1468,N_2098);
nor U7626 (N_7626,N_878,N_3271);
nand U7627 (N_7627,N_3812,N_2233);
nor U7628 (N_7628,N_3629,N_396);
nand U7629 (N_7629,N_3175,N_1669);
nor U7630 (N_7630,N_2739,N_2736);
nand U7631 (N_7631,N_1180,N_1448);
nor U7632 (N_7632,N_3726,N_3031);
nor U7633 (N_7633,N_1019,N_339);
and U7634 (N_7634,N_3302,N_1044);
nor U7635 (N_7635,N_1614,N_3636);
nor U7636 (N_7636,N_3821,N_2976);
and U7637 (N_7637,N_2216,N_1055);
or U7638 (N_7638,N_2146,N_645);
nor U7639 (N_7639,N_3276,N_21);
nor U7640 (N_7640,N_1911,N_2660);
and U7641 (N_7641,N_2287,N_3643);
nand U7642 (N_7642,N_1150,N_2891);
and U7643 (N_7643,N_2500,N_3424);
and U7644 (N_7644,N_2382,N_3114);
and U7645 (N_7645,N_1559,N_150);
nand U7646 (N_7646,N_2814,N_3586);
nand U7647 (N_7647,N_588,N_3356);
or U7648 (N_7648,N_1303,N_1588);
or U7649 (N_7649,N_2156,N_2276);
nand U7650 (N_7650,N_2285,N_2193);
nor U7651 (N_7651,N_1270,N_3403);
or U7652 (N_7652,N_2072,N_2728);
nand U7653 (N_7653,N_2850,N_3992);
nand U7654 (N_7654,N_1206,N_3571);
or U7655 (N_7655,N_2915,N_2538);
or U7656 (N_7656,N_1536,N_1969);
nor U7657 (N_7657,N_807,N_1345);
or U7658 (N_7658,N_3687,N_2929);
and U7659 (N_7659,N_1991,N_2973);
nor U7660 (N_7660,N_3367,N_3428);
nor U7661 (N_7661,N_3695,N_3828);
or U7662 (N_7662,N_3020,N_503);
or U7663 (N_7663,N_339,N_713);
or U7664 (N_7664,N_1061,N_1205);
nand U7665 (N_7665,N_2716,N_2663);
nand U7666 (N_7666,N_3325,N_425);
or U7667 (N_7667,N_3374,N_369);
and U7668 (N_7668,N_1188,N_183);
and U7669 (N_7669,N_1270,N_1783);
or U7670 (N_7670,N_1947,N_1762);
nor U7671 (N_7671,N_1566,N_2682);
or U7672 (N_7672,N_591,N_2726);
nand U7673 (N_7673,N_1308,N_2901);
nand U7674 (N_7674,N_3228,N_2525);
and U7675 (N_7675,N_1362,N_940);
and U7676 (N_7676,N_419,N_2349);
or U7677 (N_7677,N_1918,N_2730);
or U7678 (N_7678,N_2747,N_1809);
or U7679 (N_7679,N_889,N_865);
and U7680 (N_7680,N_618,N_758);
nand U7681 (N_7681,N_1836,N_601);
and U7682 (N_7682,N_2774,N_2372);
and U7683 (N_7683,N_3363,N_1813);
nor U7684 (N_7684,N_1651,N_1950);
or U7685 (N_7685,N_1888,N_1295);
and U7686 (N_7686,N_2544,N_1210);
and U7687 (N_7687,N_3368,N_2876);
nand U7688 (N_7688,N_2528,N_2360);
nor U7689 (N_7689,N_1700,N_3628);
nor U7690 (N_7690,N_1182,N_2988);
and U7691 (N_7691,N_3819,N_826);
or U7692 (N_7692,N_112,N_2777);
or U7693 (N_7693,N_2119,N_32);
nor U7694 (N_7694,N_1854,N_568);
nand U7695 (N_7695,N_3709,N_1993);
or U7696 (N_7696,N_717,N_561);
nor U7697 (N_7697,N_928,N_3220);
nor U7698 (N_7698,N_3740,N_1053);
and U7699 (N_7699,N_1883,N_7);
nor U7700 (N_7700,N_2771,N_3427);
nor U7701 (N_7701,N_2032,N_3539);
nand U7702 (N_7702,N_3177,N_1898);
and U7703 (N_7703,N_2582,N_3382);
and U7704 (N_7704,N_300,N_1981);
and U7705 (N_7705,N_253,N_2958);
or U7706 (N_7706,N_1299,N_943);
nor U7707 (N_7707,N_535,N_2098);
nor U7708 (N_7708,N_930,N_3750);
nand U7709 (N_7709,N_230,N_1393);
nor U7710 (N_7710,N_2691,N_2226);
nor U7711 (N_7711,N_2043,N_2526);
or U7712 (N_7712,N_446,N_1517);
nor U7713 (N_7713,N_795,N_1332);
nand U7714 (N_7714,N_3225,N_3731);
nor U7715 (N_7715,N_3076,N_3107);
and U7716 (N_7716,N_1611,N_3691);
xnor U7717 (N_7717,N_2929,N_1536);
nor U7718 (N_7718,N_557,N_2630);
nor U7719 (N_7719,N_947,N_1702);
nand U7720 (N_7720,N_1238,N_3167);
xor U7721 (N_7721,N_594,N_1977);
or U7722 (N_7722,N_1249,N_1410);
and U7723 (N_7723,N_1510,N_3614);
and U7724 (N_7724,N_2733,N_2374);
or U7725 (N_7725,N_1340,N_57);
nand U7726 (N_7726,N_3600,N_1690);
nand U7727 (N_7727,N_398,N_2034);
and U7728 (N_7728,N_1034,N_786);
nor U7729 (N_7729,N_490,N_3202);
nor U7730 (N_7730,N_1763,N_1787);
nand U7731 (N_7731,N_1192,N_351);
nand U7732 (N_7732,N_3816,N_3668);
and U7733 (N_7733,N_256,N_3911);
nand U7734 (N_7734,N_2283,N_2134);
xnor U7735 (N_7735,N_3726,N_3028);
or U7736 (N_7736,N_2997,N_1620);
and U7737 (N_7737,N_629,N_3453);
and U7738 (N_7738,N_3495,N_1578);
or U7739 (N_7739,N_3248,N_3952);
and U7740 (N_7740,N_3289,N_2978);
nand U7741 (N_7741,N_850,N_2684);
nand U7742 (N_7742,N_3358,N_1854);
xnor U7743 (N_7743,N_3773,N_104);
and U7744 (N_7744,N_953,N_1722);
or U7745 (N_7745,N_1594,N_2012);
xor U7746 (N_7746,N_3818,N_2377);
nor U7747 (N_7747,N_2764,N_1235);
or U7748 (N_7748,N_1881,N_451);
nand U7749 (N_7749,N_885,N_3987);
nor U7750 (N_7750,N_909,N_427);
or U7751 (N_7751,N_3384,N_1988);
nand U7752 (N_7752,N_2438,N_3756);
and U7753 (N_7753,N_3829,N_1647);
nand U7754 (N_7754,N_259,N_3341);
nor U7755 (N_7755,N_1693,N_1849);
and U7756 (N_7756,N_3175,N_3285);
nor U7757 (N_7757,N_1937,N_1511);
nand U7758 (N_7758,N_3410,N_3076);
nor U7759 (N_7759,N_3303,N_993);
nor U7760 (N_7760,N_3253,N_2651);
or U7761 (N_7761,N_1340,N_2649);
xnor U7762 (N_7762,N_586,N_2890);
or U7763 (N_7763,N_596,N_3225);
and U7764 (N_7764,N_2159,N_3674);
nor U7765 (N_7765,N_1277,N_2349);
nor U7766 (N_7766,N_2224,N_1235);
nor U7767 (N_7767,N_874,N_3319);
nand U7768 (N_7768,N_3115,N_3678);
and U7769 (N_7769,N_2302,N_3756);
nand U7770 (N_7770,N_3909,N_85);
or U7771 (N_7771,N_918,N_1111);
and U7772 (N_7772,N_188,N_1706);
or U7773 (N_7773,N_464,N_324);
and U7774 (N_7774,N_1703,N_2990);
or U7775 (N_7775,N_804,N_3735);
nand U7776 (N_7776,N_3486,N_598);
and U7777 (N_7777,N_315,N_1018);
or U7778 (N_7778,N_3725,N_2092);
and U7779 (N_7779,N_2892,N_3549);
and U7780 (N_7780,N_2501,N_2582);
nand U7781 (N_7781,N_2502,N_2320);
nand U7782 (N_7782,N_2539,N_2419);
nor U7783 (N_7783,N_3745,N_804);
xnor U7784 (N_7784,N_2166,N_3838);
and U7785 (N_7785,N_2841,N_1537);
nand U7786 (N_7786,N_2926,N_3994);
and U7787 (N_7787,N_3179,N_3032);
or U7788 (N_7788,N_2420,N_3653);
or U7789 (N_7789,N_1381,N_3771);
and U7790 (N_7790,N_1460,N_1074);
and U7791 (N_7791,N_952,N_898);
nor U7792 (N_7792,N_1878,N_3353);
and U7793 (N_7793,N_3460,N_2546);
nand U7794 (N_7794,N_1161,N_594);
nand U7795 (N_7795,N_1019,N_1650);
and U7796 (N_7796,N_219,N_3345);
nor U7797 (N_7797,N_1644,N_1863);
nor U7798 (N_7798,N_245,N_524);
xnor U7799 (N_7799,N_3399,N_1126);
nor U7800 (N_7800,N_829,N_2946);
and U7801 (N_7801,N_2824,N_2407);
or U7802 (N_7802,N_72,N_847);
or U7803 (N_7803,N_3919,N_1076);
nor U7804 (N_7804,N_657,N_1748);
nand U7805 (N_7805,N_2261,N_1045);
and U7806 (N_7806,N_1802,N_1890);
nand U7807 (N_7807,N_2168,N_492);
and U7808 (N_7808,N_1797,N_3824);
and U7809 (N_7809,N_1416,N_851);
nor U7810 (N_7810,N_1319,N_3269);
nor U7811 (N_7811,N_2143,N_566);
nor U7812 (N_7812,N_3358,N_2924);
or U7813 (N_7813,N_541,N_974);
nor U7814 (N_7814,N_2950,N_521);
or U7815 (N_7815,N_542,N_3016);
and U7816 (N_7816,N_3268,N_930);
and U7817 (N_7817,N_3343,N_1880);
or U7818 (N_7818,N_3460,N_1377);
nand U7819 (N_7819,N_3928,N_3440);
nor U7820 (N_7820,N_3000,N_3540);
or U7821 (N_7821,N_2782,N_3394);
nor U7822 (N_7822,N_742,N_1778);
nor U7823 (N_7823,N_1771,N_638);
nor U7824 (N_7824,N_3691,N_2065);
and U7825 (N_7825,N_1819,N_2860);
or U7826 (N_7826,N_498,N_2002);
or U7827 (N_7827,N_1994,N_2558);
nor U7828 (N_7828,N_240,N_3155);
nor U7829 (N_7829,N_1676,N_1415);
and U7830 (N_7830,N_1139,N_1116);
nor U7831 (N_7831,N_272,N_3492);
and U7832 (N_7832,N_3074,N_1951);
or U7833 (N_7833,N_2217,N_2648);
nand U7834 (N_7834,N_3189,N_1638);
and U7835 (N_7835,N_3058,N_509);
or U7836 (N_7836,N_1249,N_2550);
xnor U7837 (N_7837,N_861,N_33);
nor U7838 (N_7838,N_2519,N_2446);
and U7839 (N_7839,N_2458,N_2307);
xnor U7840 (N_7840,N_2959,N_1298);
xnor U7841 (N_7841,N_3890,N_641);
nand U7842 (N_7842,N_2098,N_2607);
nand U7843 (N_7843,N_1285,N_2491);
nor U7844 (N_7844,N_77,N_1489);
nor U7845 (N_7845,N_3444,N_772);
nand U7846 (N_7846,N_1453,N_2688);
nor U7847 (N_7847,N_1372,N_3224);
and U7848 (N_7848,N_3253,N_2273);
and U7849 (N_7849,N_967,N_1182);
xnor U7850 (N_7850,N_2634,N_1229);
and U7851 (N_7851,N_1315,N_226);
or U7852 (N_7852,N_1123,N_3403);
nand U7853 (N_7853,N_3834,N_1674);
nand U7854 (N_7854,N_1662,N_922);
nand U7855 (N_7855,N_2918,N_1201);
nor U7856 (N_7856,N_2917,N_15);
nand U7857 (N_7857,N_3283,N_908);
nand U7858 (N_7858,N_1566,N_569);
and U7859 (N_7859,N_1605,N_2236);
nor U7860 (N_7860,N_1915,N_1096);
and U7861 (N_7861,N_3219,N_1046);
and U7862 (N_7862,N_1054,N_2106);
and U7863 (N_7863,N_1030,N_1458);
or U7864 (N_7864,N_1321,N_1448);
nand U7865 (N_7865,N_2119,N_1990);
and U7866 (N_7866,N_1537,N_765);
nor U7867 (N_7867,N_2388,N_2287);
and U7868 (N_7868,N_1648,N_1912);
nor U7869 (N_7869,N_3964,N_1084);
nor U7870 (N_7870,N_2794,N_2861);
and U7871 (N_7871,N_3823,N_2482);
nor U7872 (N_7872,N_102,N_1051);
or U7873 (N_7873,N_1100,N_2960);
nor U7874 (N_7874,N_2491,N_1888);
and U7875 (N_7875,N_2125,N_2061);
nand U7876 (N_7876,N_2294,N_2225);
or U7877 (N_7877,N_846,N_2283);
and U7878 (N_7878,N_3089,N_3863);
or U7879 (N_7879,N_167,N_1952);
nor U7880 (N_7880,N_3935,N_1136);
nand U7881 (N_7881,N_3106,N_2775);
nand U7882 (N_7882,N_3825,N_879);
or U7883 (N_7883,N_2020,N_3245);
nand U7884 (N_7884,N_3995,N_1681);
nor U7885 (N_7885,N_3977,N_2508);
and U7886 (N_7886,N_3315,N_2121);
nand U7887 (N_7887,N_1443,N_3524);
nor U7888 (N_7888,N_2895,N_3002);
xor U7889 (N_7889,N_2840,N_491);
xnor U7890 (N_7890,N_2022,N_353);
nor U7891 (N_7891,N_181,N_3585);
or U7892 (N_7892,N_2737,N_3360);
nand U7893 (N_7893,N_2406,N_2973);
nor U7894 (N_7894,N_2087,N_3744);
nand U7895 (N_7895,N_3407,N_2293);
or U7896 (N_7896,N_3567,N_457);
and U7897 (N_7897,N_3420,N_3384);
nand U7898 (N_7898,N_175,N_771);
nand U7899 (N_7899,N_1199,N_3437);
or U7900 (N_7900,N_3297,N_2912);
nor U7901 (N_7901,N_735,N_3127);
nand U7902 (N_7902,N_3378,N_582);
and U7903 (N_7903,N_2694,N_2700);
nor U7904 (N_7904,N_3969,N_768);
nand U7905 (N_7905,N_2168,N_2678);
or U7906 (N_7906,N_3489,N_3479);
or U7907 (N_7907,N_1428,N_1249);
nand U7908 (N_7908,N_2789,N_1848);
nor U7909 (N_7909,N_1120,N_1334);
nand U7910 (N_7910,N_790,N_1108);
or U7911 (N_7911,N_2333,N_3914);
nand U7912 (N_7912,N_1075,N_572);
nand U7913 (N_7913,N_433,N_2815);
and U7914 (N_7914,N_1502,N_863);
and U7915 (N_7915,N_1446,N_414);
nand U7916 (N_7916,N_2496,N_120);
nand U7917 (N_7917,N_3231,N_2077);
nor U7918 (N_7918,N_1779,N_1035);
nor U7919 (N_7919,N_2836,N_3706);
nand U7920 (N_7920,N_2397,N_1523);
xnor U7921 (N_7921,N_2176,N_1492);
and U7922 (N_7922,N_1657,N_3515);
or U7923 (N_7923,N_3321,N_3627);
nor U7924 (N_7924,N_2106,N_2897);
and U7925 (N_7925,N_3781,N_3364);
and U7926 (N_7926,N_819,N_3779);
nand U7927 (N_7927,N_316,N_1315);
and U7928 (N_7928,N_1423,N_644);
and U7929 (N_7929,N_3470,N_2068);
nor U7930 (N_7930,N_1000,N_2501);
and U7931 (N_7931,N_3334,N_2278);
and U7932 (N_7932,N_571,N_2370);
xnor U7933 (N_7933,N_2961,N_338);
or U7934 (N_7934,N_2071,N_2934);
nand U7935 (N_7935,N_566,N_65);
and U7936 (N_7936,N_524,N_2325);
and U7937 (N_7937,N_3074,N_522);
nand U7938 (N_7938,N_3604,N_2732);
or U7939 (N_7939,N_2713,N_960);
xnor U7940 (N_7940,N_2888,N_1468);
or U7941 (N_7941,N_299,N_1658);
nor U7942 (N_7942,N_3575,N_1511);
and U7943 (N_7943,N_1600,N_1040);
xnor U7944 (N_7944,N_3624,N_3186);
nor U7945 (N_7945,N_2447,N_2581);
nand U7946 (N_7946,N_3301,N_3390);
xor U7947 (N_7947,N_1733,N_2500);
nor U7948 (N_7948,N_1489,N_324);
nor U7949 (N_7949,N_1074,N_1904);
and U7950 (N_7950,N_1616,N_1539);
nor U7951 (N_7951,N_3258,N_576);
nand U7952 (N_7952,N_2777,N_1240);
xor U7953 (N_7953,N_3127,N_1205);
nor U7954 (N_7954,N_1287,N_1627);
nand U7955 (N_7955,N_1748,N_2386);
nand U7956 (N_7956,N_1872,N_2559);
and U7957 (N_7957,N_2507,N_2645);
and U7958 (N_7958,N_3613,N_2758);
or U7959 (N_7959,N_550,N_3033);
or U7960 (N_7960,N_2510,N_2311);
nor U7961 (N_7961,N_582,N_3133);
or U7962 (N_7962,N_2000,N_1561);
or U7963 (N_7963,N_1919,N_1877);
nand U7964 (N_7964,N_3843,N_3207);
xor U7965 (N_7965,N_1426,N_1935);
xor U7966 (N_7966,N_3258,N_176);
and U7967 (N_7967,N_2570,N_3375);
or U7968 (N_7968,N_3647,N_1229);
and U7969 (N_7969,N_3617,N_3547);
nand U7970 (N_7970,N_989,N_3266);
xor U7971 (N_7971,N_2842,N_10);
nor U7972 (N_7972,N_1633,N_1596);
nor U7973 (N_7973,N_1360,N_683);
or U7974 (N_7974,N_2817,N_2032);
nand U7975 (N_7975,N_653,N_584);
xor U7976 (N_7976,N_1210,N_672);
xnor U7977 (N_7977,N_194,N_1171);
and U7978 (N_7978,N_3589,N_376);
and U7979 (N_7979,N_1744,N_3854);
nand U7980 (N_7980,N_1133,N_1687);
nand U7981 (N_7981,N_3441,N_1759);
or U7982 (N_7982,N_1437,N_2638);
nand U7983 (N_7983,N_2983,N_1979);
xor U7984 (N_7984,N_289,N_1030);
and U7985 (N_7985,N_2365,N_912);
nand U7986 (N_7986,N_3832,N_2591);
nor U7987 (N_7987,N_2885,N_3271);
or U7988 (N_7988,N_1984,N_1955);
or U7989 (N_7989,N_3715,N_1262);
nor U7990 (N_7990,N_1841,N_3247);
or U7991 (N_7991,N_374,N_2957);
nand U7992 (N_7992,N_1660,N_3241);
and U7993 (N_7993,N_2831,N_2864);
or U7994 (N_7994,N_1772,N_791);
nor U7995 (N_7995,N_2926,N_2610);
nor U7996 (N_7996,N_3484,N_623);
nor U7997 (N_7997,N_511,N_506);
nand U7998 (N_7998,N_10,N_3982);
and U7999 (N_7999,N_3969,N_444);
or U8000 (N_8000,N_7351,N_5843);
nor U8001 (N_8001,N_7622,N_6340);
and U8002 (N_8002,N_4347,N_4740);
and U8003 (N_8003,N_7807,N_7638);
nor U8004 (N_8004,N_6518,N_4732);
and U8005 (N_8005,N_4768,N_5337);
nor U8006 (N_8006,N_5844,N_4437);
nor U8007 (N_8007,N_7291,N_4366);
nor U8008 (N_8008,N_7481,N_7444);
xor U8009 (N_8009,N_6549,N_5117);
nor U8010 (N_8010,N_5663,N_4622);
nor U8011 (N_8011,N_4502,N_6500);
and U8012 (N_8012,N_5669,N_5195);
nor U8013 (N_8013,N_7720,N_7657);
or U8014 (N_8014,N_4482,N_5688);
xor U8015 (N_8015,N_4526,N_5760);
and U8016 (N_8016,N_5953,N_7120);
nand U8017 (N_8017,N_5012,N_5106);
xor U8018 (N_8018,N_7978,N_4821);
and U8019 (N_8019,N_5249,N_7175);
nor U8020 (N_8020,N_5177,N_7428);
or U8021 (N_8021,N_5320,N_4422);
nand U8022 (N_8022,N_6121,N_6243);
nor U8023 (N_8023,N_4510,N_4551);
or U8024 (N_8024,N_6788,N_6111);
and U8025 (N_8025,N_5399,N_5894);
nor U8026 (N_8026,N_7031,N_4774);
and U8027 (N_8027,N_6326,N_7914);
and U8028 (N_8028,N_5707,N_5873);
xor U8029 (N_8029,N_5982,N_4518);
and U8030 (N_8030,N_4773,N_6961);
nand U8031 (N_8031,N_7061,N_7595);
nand U8032 (N_8032,N_6071,N_5803);
nand U8033 (N_8033,N_4964,N_5412);
nand U8034 (N_8034,N_7506,N_7293);
or U8035 (N_8035,N_7779,N_7688);
and U8036 (N_8036,N_6291,N_5121);
nor U8037 (N_8037,N_7078,N_7212);
nor U8038 (N_8038,N_4706,N_4573);
and U8039 (N_8039,N_7821,N_5018);
nand U8040 (N_8040,N_4642,N_5666);
or U8041 (N_8041,N_5573,N_4981);
or U8042 (N_8042,N_7517,N_7278);
nor U8043 (N_8043,N_7177,N_5950);
nor U8044 (N_8044,N_6297,N_4177);
xnor U8045 (N_8045,N_5991,N_4125);
nand U8046 (N_8046,N_4245,N_4661);
nor U8047 (N_8047,N_4084,N_4472);
nor U8048 (N_8048,N_4111,N_4559);
and U8049 (N_8049,N_5002,N_7475);
nor U8050 (N_8050,N_7183,N_4698);
or U8051 (N_8051,N_5900,N_4765);
nand U8052 (N_8052,N_5074,N_5589);
nand U8053 (N_8053,N_5271,N_7877);
or U8054 (N_8054,N_7254,N_4352);
and U8055 (N_8055,N_7512,N_4802);
nor U8056 (N_8056,N_5716,N_6379);
or U8057 (N_8057,N_4001,N_6913);
nand U8058 (N_8058,N_6919,N_6522);
nand U8059 (N_8059,N_6315,N_4763);
nor U8060 (N_8060,N_4879,N_4447);
nor U8061 (N_8061,N_5626,N_4042);
or U8062 (N_8062,N_4055,N_5442);
nor U8063 (N_8063,N_4572,N_4693);
and U8064 (N_8064,N_4299,N_7124);
or U8065 (N_8065,N_4483,N_6520);
nor U8066 (N_8066,N_5665,N_7681);
nor U8067 (N_8067,N_5777,N_6208);
nand U8068 (N_8068,N_5093,N_5618);
or U8069 (N_8069,N_6333,N_7948);
and U8070 (N_8070,N_6953,N_5565);
or U8071 (N_8071,N_5204,N_7667);
nor U8072 (N_8072,N_7007,N_7991);
nand U8073 (N_8073,N_5205,N_6877);
nor U8074 (N_8074,N_7129,N_6452);
and U8075 (N_8075,N_5785,N_4090);
and U8076 (N_8076,N_7251,N_4575);
nor U8077 (N_8077,N_5279,N_7330);
nand U8078 (N_8078,N_4527,N_6565);
xor U8079 (N_8079,N_4546,N_5741);
or U8080 (N_8080,N_7499,N_4013);
xor U8081 (N_8081,N_7787,N_6363);
and U8082 (N_8082,N_6244,N_6373);
nand U8083 (N_8083,N_6330,N_4272);
or U8084 (N_8084,N_6055,N_4373);
nor U8085 (N_8085,N_6930,N_7876);
nand U8086 (N_8086,N_7922,N_6865);
nor U8087 (N_8087,N_6677,N_6767);
nand U8088 (N_8088,N_4052,N_6424);
nand U8089 (N_8089,N_4711,N_6195);
or U8090 (N_8090,N_7326,N_4009);
and U8091 (N_8091,N_7549,N_7270);
nor U8092 (N_8092,N_6869,N_7314);
nand U8093 (N_8093,N_6741,N_5092);
or U8094 (N_8094,N_6052,N_6286);
or U8095 (N_8095,N_4249,N_7179);
nor U8096 (N_8096,N_7365,N_5221);
and U8097 (N_8097,N_4259,N_7185);
nand U8098 (N_8098,N_7013,N_5768);
and U8099 (N_8099,N_6794,N_4993);
nor U8100 (N_8100,N_4686,N_5918);
and U8101 (N_8101,N_4775,N_5465);
xnor U8102 (N_8102,N_4047,N_6868);
xor U8103 (N_8103,N_7361,N_6866);
xor U8104 (N_8104,N_5022,N_4411);
nand U8105 (N_8105,N_4105,N_4394);
or U8106 (N_8106,N_6122,N_5167);
nand U8107 (N_8107,N_5622,N_6712);
and U8108 (N_8108,N_6528,N_6893);
nand U8109 (N_8109,N_5682,N_5490);
and U8110 (N_8110,N_7508,N_7346);
nand U8111 (N_8111,N_7420,N_5076);
or U8112 (N_8112,N_5522,N_6867);
or U8113 (N_8113,N_7906,N_6150);
nand U8114 (N_8114,N_4446,N_4266);
and U8115 (N_8115,N_7846,N_5549);
or U8116 (N_8116,N_7611,N_7279);
xnor U8117 (N_8117,N_6700,N_6765);
xnor U8118 (N_8118,N_5429,N_4193);
nand U8119 (N_8119,N_6045,N_4689);
nor U8120 (N_8120,N_7718,N_6753);
nor U8121 (N_8121,N_6422,N_7114);
xnor U8122 (N_8122,N_7302,N_6447);
or U8123 (N_8123,N_5409,N_7285);
or U8124 (N_8124,N_7737,N_5331);
nand U8125 (N_8125,N_5088,N_5939);
or U8126 (N_8126,N_6364,N_7852);
and U8127 (N_8127,N_4841,N_4595);
or U8128 (N_8128,N_6415,N_6662);
and U8129 (N_8129,N_6319,N_5324);
or U8130 (N_8130,N_5096,N_4590);
and U8131 (N_8131,N_6783,N_7913);
or U8132 (N_8132,N_6858,N_5798);
nand U8133 (N_8133,N_4370,N_5747);
or U8134 (N_8134,N_7607,N_7550);
or U8135 (N_8135,N_6989,N_6745);
xor U8136 (N_8136,N_5390,N_7985);
nand U8137 (N_8137,N_5675,N_5964);
and U8138 (N_8138,N_6000,N_7648);
or U8139 (N_8139,N_6515,N_4399);
nand U8140 (N_8140,N_5788,N_4149);
nor U8141 (N_8141,N_4557,N_6095);
or U8142 (N_8142,N_5461,N_5552);
nor U8143 (N_8143,N_4852,N_6430);
nand U8144 (N_8144,N_4371,N_6709);
nand U8145 (N_8145,N_5763,N_7003);
nand U8146 (N_8146,N_7599,N_6168);
nor U8147 (N_8147,N_6604,N_4381);
or U8148 (N_8148,N_7182,N_6573);
or U8149 (N_8149,N_4623,N_7940);
and U8150 (N_8150,N_6310,N_7460);
or U8151 (N_8151,N_6671,N_7678);
nand U8152 (N_8152,N_6701,N_7992);
xor U8153 (N_8153,N_6030,N_6025);
and U8154 (N_8154,N_4761,N_6726);
or U8155 (N_8155,N_4611,N_4237);
or U8156 (N_8156,N_6349,N_4385);
and U8157 (N_8157,N_6007,N_6807);
xnor U8158 (N_8158,N_7441,N_7045);
nor U8159 (N_8159,N_6899,N_5576);
nor U8160 (N_8160,N_6497,N_5309);
nand U8161 (N_8161,N_6439,N_5598);
nand U8162 (N_8162,N_4613,N_5611);
and U8163 (N_8163,N_5828,N_5349);
nor U8164 (N_8164,N_6616,N_4662);
nor U8165 (N_8165,N_6688,N_7021);
or U8166 (N_8166,N_4577,N_7637);
nor U8167 (N_8167,N_6928,N_7433);
nor U8168 (N_8168,N_4878,N_4186);
or U8169 (N_8169,N_5888,N_6769);
nand U8170 (N_8170,N_5325,N_5445);
nand U8171 (N_8171,N_4545,N_5198);
and U8172 (N_8172,N_6203,N_5752);
or U8173 (N_8173,N_5212,N_5600);
or U8174 (N_8174,N_5045,N_7329);
nand U8175 (N_8175,N_4766,N_7315);
nor U8176 (N_8176,N_7649,N_7354);
and U8177 (N_8177,N_6336,N_4121);
nor U8178 (N_8178,N_4202,N_7818);
and U8179 (N_8179,N_7988,N_7536);
and U8180 (N_8180,N_4497,N_6747);
nor U8181 (N_8181,N_4922,N_7650);
nand U8182 (N_8182,N_6137,N_6233);
or U8183 (N_8183,N_5275,N_4585);
nand U8184 (N_8184,N_6622,N_4589);
nor U8185 (N_8185,N_5511,N_7915);
nor U8186 (N_8186,N_6394,N_5368);
or U8187 (N_8187,N_5751,N_7619);
or U8188 (N_8188,N_5898,N_4612);
nor U8189 (N_8189,N_5903,N_4669);
or U8190 (N_8190,N_5027,N_4817);
and U8191 (N_8191,N_5868,N_5266);
or U8192 (N_8192,N_6246,N_4435);
and U8193 (N_8193,N_7216,N_4428);
xor U8194 (N_8194,N_5243,N_7503);
and U8195 (N_8195,N_6482,N_5201);
nand U8196 (N_8196,N_4885,N_5234);
xnor U8197 (N_8197,N_6419,N_7799);
and U8198 (N_8198,N_7465,N_6048);
nand U8199 (N_8199,N_7792,N_4828);
or U8200 (N_8200,N_6544,N_7132);
nor U8201 (N_8201,N_7198,N_7051);
nor U8202 (N_8202,N_5263,N_5466);
nand U8203 (N_8203,N_4040,N_5211);
and U8204 (N_8204,N_6743,N_7210);
or U8205 (N_8205,N_7810,N_6925);
or U8206 (N_8206,N_6513,N_5035);
nand U8207 (N_8207,N_5531,N_6440);
nand U8208 (N_8208,N_7498,N_7248);
xor U8209 (N_8209,N_4312,N_4566);
or U8210 (N_8210,N_7079,N_5693);
nand U8211 (N_8211,N_7386,N_4273);
nand U8212 (N_8212,N_5190,N_7395);
nor U8213 (N_8213,N_6856,N_5561);
or U8214 (N_8214,N_5672,N_6230);
and U8215 (N_8215,N_6655,N_6063);
nand U8216 (N_8216,N_4891,N_7653);
nor U8217 (N_8217,N_4889,N_6385);
or U8218 (N_8218,N_7464,N_6459);
and U8219 (N_8219,N_7062,N_5515);
nand U8220 (N_8220,N_5487,N_6181);
or U8221 (N_8221,N_5543,N_7316);
nor U8222 (N_8222,N_7813,N_5638);
and U8223 (N_8223,N_5330,N_4191);
nor U8224 (N_8224,N_6713,N_6227);
nand U8225 (N_8225,N_4757,N_5793);
nor U8226 (N_8226,N_6703,N_4296);
nor U8227 (N_8227,N_6343,N_5755);
nand U8228 (N_8228,N_6200,N_6037);
or U8229 (N_8229,N_7686,N_4226);
or U8230 (N_8230,N_4951,N_5013);
nor U8231 (N_8231,N_7141,N_7770);
nand U8232 (N_8232,N_6799,N_6220);
nand U8233 (N_8233,N_7231,N_5975);
nand U8234 (N_8234,N_5459,N_5061);
and U8235 (N_8235,N_5229,N_5463);
or U8236 (N_8236,N_6977,N_4673);
nor U8237 (N_8237,N_4976,N_7245);
nor U8238 (N_8238,N_5259,N_5202);
or U8239 (N_8239,N_7029,N_5668);
nand U8240 (N_8240,N_4234,N_5696);
or U8241 (N_8241,N_6486,N_7064);
nand U8242 (N_8242,N_6884,N_7343);
or U8243 (N_8243,N_5360,N_5289);
nand U8244 (N_8244,N_7661,N_7471);
nor U8245 (N_8245,N_4323,N_7788);
nand U8246 (N_8246,N_5628,N_6069);
or U8247 (N_8247,N_5434,N_5359);
nor U8248 (N_8248,N_6076,N_5575);
or U8249 (N_8249,N_7714,N_5016);
nand U8250 (N_8250,N_5428,N_4219);
xor U8251 (N_8251,N_6491,N_4996);
nand U8252 (N_8252,N_4695,N_6873);
xor U8253 (N_8253,N_7875,N_5374);
or U8254 (N_8254,N_4342,N_4912);
nor U8255 (N_8255,N_6106,N_7783);
and U8256 (N_8256,N_4815,N_5416);
and U8257 (N_8257,N_7004,N_7998);
xor U8258 (N_8258,N_4151,N_5477);
and U8259 (N_8259,N_6320,N_4117);
nor U8260 (N_8260,N_4375,N_4178);
xnor U8261 (N_8261,N_5652,N_6940);
and U8262 (N_8262,N_7625,N_5529);
xor U8263 (N_8263,N_4128,N_7160);
and U8264 (N_8264,N_5142,N_5771);
or U8265 (N_8265,N_7771,N_4292);
nor U8266 (N_8266,N_6773,N_7037);
nor U8267 (N_8267,N_5393,N_5550);
or U8268 (N_8268,N_4911,N_4833);
and U8269 (N_8269,N_5223,N_5065);
nand U8270 (N_8270,N_5833,N_6761);
and U8271 (N_8271,N_4950,N_5339);
or U8272 (N_8272,N_6074,N_7626);
or U8273 (N_8273,N_5099,N_7096);
nand U8274 (N_8274,N_5523,N_5342);
nand U8275 (N_8275,N_7636,N_6908);
xor U8276 (N_8276,N_4604,N_4364);
nor U8277 (N_8277,N_5116,N_7387);
or U8278 (N_8278,N_6478,N_7640);
and U8279 (N_8279,N_7443,N_5871);
and U8280 (N_8280,N_4792,N_6781);
or U8281 (N_8281,N_5187,N_4239);
xor U8282 (N_8282,N_5150,N_4062);
nor U8283 (N_8283,N_4407,N_5043);
nor U8284 (N_8284,N_4903,N_4017);
or U8285 (N_8285,N_7469,N_4269);
nand U8286 (N_8286,N_6540,N_5988);
or U8287 (N_8287,N_5344,N_4894);
or U8288 (N_8288,N_7744,N_7518);
nand U8289 (N_8289,N_6169,N_5336);
nor U8290 (N_8290,N_4469,N_5674);
and U8291 (N_8291,N_7213,N_6339);
nor U8292 (N_8292,N_6141,N_6460);
nand U8293 (N_8293,N_7421,N_5458);
or U8294 (N_8294,N_7935,N_5959);
or U8295 (N_8295,N_7188,N_7946);
nor U8296 (N_8296,N_7197,N_5866);
nand U8297 (N_8297,N_7164,N_6832);
and U8298 (N_8298,N_6907,N_6876);
nand U8299 (N_8299,N_6787,N_4665);
nand U8300 (N_8300,N_6462,N_6561);
nand U8301 (N_8301,N_6724,N_5256);
nor U8302 (N_8302,N_7983,N_7271);
nand U8303 (N_8303,N_4046,N_4036);
nand U8304 (N_8304,N_6857,N_4846);
xor U8305 (N_8305,N_6635,N_6360);
nand U8306 (N_8306,N_4061,N_4890);
and U8307 (N_8307,N_7809,N_7191);
nand U8308 (N_8308,N_5799,N_5038);
nor U8309 (N_8309,N_5508,N_4944);
nand U8310 (N_8310,N_5736,N_7209);
or U8311 (N_8311,N_7313,N_6538);
nand U8312 (N_8312,N_5175,N_6646);
and U8313 (N_8313,N_4173,N_7372);
and U8314 (N_8314,N_7331,N_7423);
nand U8315 (N_8315,N_4564,N_6467);
xor U8316 (N_8316,N_7567,N_4449);
nand U8317 (N_8317,N_5354,N_4295);
or U8318 (N_8318,N_5753,N_6275);
nand U8319 (N_8319,N_5756,N_7581);
or U8320 (N_8320,N_7500,N_6372);
or U8321 (N_8321,N_5677,N_5011);
nor U8322 (N_8322,N_5502,N_6217);
nand U8323 (N_8323,N_6707,N_4560);
xor U8324 (N_8324,N_6710,N_7435);
nand U8325 (N_8325,N_6812,N_7731);
nand U8326 (N_8326,N_5946,N_5855);
nand U8327 (N_8327,N_7735,N_6389);
nand U8328 (N_8328,N_4459,N_7467);
or U8329 (N_8329,N_5955,N_7307);
nor U8330 (N_8330,N_7698,N_5456);
nor U8331 (N_8331,N_5424,N_6811);
nand U8332 (N_8332,N_6779,N_6810);
or U8333 (N_8333,N_5867,N_4132);
and U8334 (N_8334,N_6471,N_4075);
nand U8335 (N_8335,N_5494,N_6621);
and U8336 (N_8336,N_6342,N_6351);
nor U8337 (N_8337,N_7520,N_6305);
nor U8338 (N_8338,N_5154,N_6827);
or U8339 (N_8339,N_5792,N_7319);
nor U8340 (N_8340,N_6322,N_7126);
or U8341 (N_8341,N_4341,N_4087);
nand U8342 (N_8342,N_7964,N_6406);
or U8343 (N_8343,N_6772,N_7140);
or U8344 (N_8344,N_7095,N_7450);
xnor U8345 (N_8345,N_7115,N_4521);
or U8346 (N_8346,N_7038,N_7982);
or U8347 (N_8347,N_4650,N_6051);
nor U8348 (N_8348,N_4729,N_4496);
nand U8349 (N_8349,N_7349,N_7128);
and U8350 (N_8350,N_4592,N_6590);
or U8351 (N_8351,N_5037,N_5727);
and U8352 (N_8352,N_5761,N_4788);
nand U8353 (N_8353,N_4862,N_5906);
and U8354 (N_8354,N_4741,N_5094);
nand U8355 (N_8355,N_6880,N_6028);
and U8356 (N_8356,N_6681,N_5897);
or U8357 (N_8357,N_4904,N_4855);
or U8358 (N_8358,N_6979,N_5814);
nor U8359 (N_8359,N_4547,N_6759);
or U8360 (N_8360,N_6664,N_6918);
nor U8361 (N_8361,N_4576,N_6881);
nor U8362 (N_8362,N_4931,N_5968);
nand U8363 (N_8363,N_5444,N_6353);
or U8364 (N_8364,N_6417,N_5933);
nand U8365 (N_8365,N_6253,N_7000);
xor U8366 (N_8366,N_5782,N_6721);
or U8367 (N_8367,N_7939,N_7287);
nor U8368 (N_8368,N_6105,N_4637);
and U8369 (N_8369,N_4071,N_5218);
and U8370 (N_8370,N_4811,N_6526);
nand U8371 (N_8371,N_6568,N_4135);
xnor U8372 (N_8372,N_5188,N_4044);
nor U8373 (N_8373,N_6718,N_6829);
nor U8374 (N_8374,N_7963,N_5206);
nor U8375 (N_8375,N_4208,N_4384);
nand U8376 (N_8376,N_7839,N_6946);
and U8377 (N_8377,N_5007,N_5840);
nand U8378 (N_8378,N_6800,N_6805);
nor U8379 (N_8379,N_7060,N_7659);
nor U8380 (N_8380,N_5010,N_5578);
nor U8381 (N_8381,N_7170,N_4808);
and U8382 (N_8382,N_7815,N_4795);
nor U8383 (N_8383,N_6864,N_5262);
or U8384 (N_8384,N_5115,N_7082);
nand U8385 (N_8385,N_6024,N_4287);
xor U8386 (N_8386,N_6820,N_7750);
nand U8387 (N_8387,N_7620,N_4006);
nand U8388 (N_8388,N_7748,N_7259);
nand U8389 (N_8389,N_4914,N_4508);
and U8390 (N_8390,N_4721,N_5213);
xnor U8391 (N_8391,N_4909,N_7255);
nand U8392 (N_8392,N_6044,N_6241);
xor U8393 (N_8393,N_4334,N_6004);
or U8394 (N_8394,N_6601,N_4000);
nor U8395 (N_8395,N_4353,N_6149);
and U8396 (N_8396,N_5302,N_5613);
and U8397 (N_8397,N_5930,N_5836);
nor U8398 (N_8398,N_4133,N_6642);
nand U8399 (N_8399,N_6103,N_6120);
or U8400 (N_8400,N_6252,N_5895);
or U8401 (N_8401,N_6516,N_6087);
or U8402 (N_8402,N_6388,N_4785);
nor U8403 (N_8403,N_6886,N_7849);
or U8404 (N_8404,N_6553,N_7453);
nand U8405 (N_8405,N_7401,N_7122);
xor U8406 (N_8406,N_6098,N_4728);
or U8407 (N_8407,N_7778,N_7893);
and U8408 (N_8408,N_7389,N_7378);
or U8409 (N_8409,N_7702,N_6421);
or U8410 (N_8410,N_7083,N_5704);
nor U8411 (N_8411,N_5014,N_4854);
nand U8412 (N_8412,N_5264,N_6509);
and U8413 (N_8413,N_6316,N_4587);
and U8414 (N_8414,N_4355,N_5242);
or U8415 (N_8415,N_4666,N_4882);
nand U8416 (N_8416,N_6212,N_5783);
nand U8417 (N_8417,N_4454,N_6670);
or U8418 (N_8418,N_6821,N_6299);
nor U8419 (N_8419,N_7215,N_6558);
nand U8420 (N_8420,N_5199,N_5679);
and U8421 (N_8421,N_4959,N_6453);
and U8422 (N_8422,N_6112,N_5983);
and U8423 (N_8423,N_5124,N_7118);
or U8424 (N_8424,N_6454,N_4630);
or U8425 (N_8425,N_7894,N_6059);
nand U8426 (N_8426,N_6091,N_6852);
and U8427 (N_8427,N_7531,N_5270);
or U8428 (N_8428,N_6530,N_4349);
nor U8429 (N_8429,N_7406,N_5468);
nor U8430 (N_8430,N_7538,N_7711);
nor U8431 (N_8431,N_7049,N_7305);
nand U8432 (N_8432,N_7924,N_6755);
nand U8433 (N_8433,N_7033,N_6125);
or U8434 (N_8434,N_6038,N_4141);
nor U8435 (N_8435,N_6559,N_4322);
xor U8436 (N_8436,N_5128,N_4984);
nor U8437 (N_8437,N_5457,N_7050);
nor U8438 (N_8438,N_7949,N_6173);
xor U8439 (N_8439,N_5452,N_6383);
or U8440 (N_8440,N_4054,N_5352);
or U8441 (N_8441,N_4308,N_7859);
nor U8442 (N_8442,N_5499,N_5241);
xnor U8443 (N_8443,N_7655,N_4119);
or U8444 (N_8444,N_7260,N_5766);
nor U8445 (N_8445,N_7864,N_4517);
nor U8446 (N_8446,N_5881,N_5066);
and U8447 (N_8447,N_4679,N_6790);
or U8448 (N_8448,N_7135,N_4316);
and U8449 (N_8449,N_7071,N_7780);
or U8450 (N_8450,N_4632,N_6387);
nor U8451 (N_8451,N_7746,N_6944);
and U8452 (N_8452,N_6816,N_7138);
nand U8453 (N_8453,N_5322,N_5227);
nand U8454 (N_8454,N_7865,N_7828);
nor U8455 (N_8455,N_6898,N_7407);
and U8456 (N_8456,N_4973,N_6862);
and U8457 (N_8457,N_4250,N_6802);
xor U8458 (N_8458,N_4004,N_6107);
and U8459 (N_8459,N_4329,N_6554);
nand U8460 (N_8460,N_6536,N_5478);
and U8461 (N_8461,N_5535,N_5931);
or U8462 (N_8462,N_5451,N_4291);
and U8463 (N_8463,N_5729,N_7159);
nand U8464 (N_8464,N_6999,N_7579);
or U8465 (N_8465,N_4254,N_5521);
nand U8466 (N_8466,N_7505,N_5389);
and U8467 (N_8467,N_7529,N_5453);
or U8468 (N_8468,N_4015,N_6719);
nand U8469 (N_8469,N_4516,N_5048);
and U8470 (N_8470,N_7546,N_7338);
or U8471 (N_8471,N_5274,N_4391);
nor U8472 (N_8472,N_5496,N_6481);
nand U8473 (N_8473,N_5513,N_4379);
nand U8474 (N_8474,N_5113,N_5176);
xor U8475 (N_8475,N_4596,N_7396);
and U8476 (N_8476,N_4201,N_5423);
nor U8477 (N_8477,N_4888,N_5417);
or U8478 (N_8478,N_6784,N_7997);
nor U8479 (N_8479,N_6978,N_7162);
and U8480 (N_8480,N_5963,N_6611);
nand U8481 (N_8481,N_5036,N_6472);
nand U8482 (N_8482,N_6049,N_5422);
xnor U8483 (N_8483,N_7726,N_4190);
and U8484 (N_8484,N_6429,N_5922);
xnor U8485 (N_8485,N_4809,N_5790);
nand U8486 (N_8486,N_7721,N_7207);
or U8487 (N_8487,N_5643,N_6752);
nor U8488 (N_8488,N_6644,N_7928);
nor U8489 (N_8489,N_4660,N_5915);
xor U8490 (N_8490,N_6041,N_7186);
or U8491 (N_8491,N_4212,N_6947);
and U8492 (N_8492,N_7110,N_7723);
nor U8493 (N_8493,N_6182,N_4382);
nand U8494 (N_8494,N_6650,N_5411);
or U8495 (N_8495,N_4324,N_7816);
or U8496 (N_8496,N_5363,N_5607);
nor U8497 (N_8497,N_4305,N_6223);
nand U8498 (N_8498,N_6791,N_4485);
nand U8499 (N_8499,N_7006,N_4712);
and U8500 (N_8500,N_6093,N_4842);
nor U8501 (N_8501,N_4430,N_5724);
nand U8502 (N_8502,N_6465,N_6014);
xor U8503 (N_8503,N_4220,N_4387);
and U8504 (N_8504,N_5313,N_5355);
nor U8505 (N_8505,N_5372,N_5152);
and U8506 (N_8506,N_4335,N_4488);
nand U8507 (N_8507,N_4725,N_6610);
nand U8508 (N_8508,N_4672,N_5246);
nand U8509 (N_8509,N_7397,N_5657);
nor U8510 (N_8510,N_7280,N_5080);
xnor U8511 (N_8511,N_4158,N_4131);
nor U8512 (N_8512,N_7853,N_7901);
or U8513 (N_8513,N_4473,N_7556);
and U8514 (N_8514,N_5605,N_5194);
xnor U8515 (N_8515,N_7429,N_7008);
or U8516 (N_8516,N_5820,N_6404);
or U8517 (N_8517,N_4408,N_5853);
or U8518 (N_8518,N_6190,N_6945);
and U8519 (N_8519,N_4311,N_6643);
and U8520 (N_8520,N_6840,N_4197);
or U8521 (N_8521,N_4456,N_6975);
or U8522 (N_8522,N_7218,N_4812);
nor U8523 (N_8523,N_5765,N_4300);
and U8524 (N_8524,N_6434,N_7895);
xnor U8525 (N_8525,N_7320,N_4823);
nor U8526 (N_8526,N_5641,N_5020);
and U8527 (N_8527,N_4747,N_5070);
nand U8528 (N_8528,N_6186,N_4155);
xnor U8529 (N_8529,N_7918,N_5810);
nand U8530 (N_8530,N_4769,N_4876);
xnor U8531 (N_8531,N_5122,N_5911);
and U8532 (N_8532,N_7800,N_4122);
nand U8533 (N_8533,N_6665,N_7916);
and U8534 (N_8534,N_6853,N_5890);
nor U8535 (N_8535,N_7371,N_4568);
nor U8536 (N_8536,N_4525,N_6034);
nand U8537 (N_8537,N_4584,N_6010);
or U8538 (N_8538,N_7180,N_6172);
nand U8539 (N_8539,N_6312,N_5594);
or U8540 (N_8540,N_5052,N_5056);
xnor U8541 (N_8541,N_5951,N_5017);
or U8542 (N_8542,N_5558,N_5732);
nand U8543 (N_8543,N_7602,N_5003);
or U8544 (N_8544,N_5583,N_7932);
and U8545 (N_8545,N_4067,N_7616);
xnor U8546 (N_8546,N_7167,N_4362);
nor U8547 (N_8547,N_7142,N_4051);
nor U8548 (N_8548,N_4203,N_5298);
nor U8549 (N_8549,N_6020,N_5920);
and U8550 (N_8550,N_5338,N_5403);
nand U8551 (N_8551,N_7028,N_4570);
and U8552 (N_8552,N_5957,N_7094);
nor U8553 (N_8553,N_5488,N_5567);
nand U8554 (N_8554,N_7012,N_7025);
nand U8555 (N_8555,N_5388,N_5837);
xor U8556 (N_8556,N_5138,N_4089);
and U8557 (N_8557,N_4425,N_6539);
nand U8558 (N_8558,N_7919,N_7530);
xnor U8559 (N_8559,N_5284,N_4406);
or U8560 (N_8560,N_5203,N_4257);
nand U8561 (N_8561,N_6706,N_6731);
nor U8562 (N_8562,N_7570,N_4476);
nand U8563 (N_8563,N_5455,N_7009);
or U8564 (N_8564,N_7559,N_5064);
nand U8565 (N_8565,N_5267,N_4256);
nand U8566 (N_8566,N_5525,N_6796);
and U8567 (N_8567,N_4065,N_5318);
nor U8568 (N_8568,N_5288,N_6714);
nand U8569 (N_8569,N_4444,N_7763);
and U8570 (N_8570,N_7573,N_4799);
nor U8571 (N_8571,N_4176,N_6242);
nand U8572 (N_8572,N_4825,N_7297);
nand U8573 (N_8573,N_4682,N_5597);
and U8574 (N_8574,N_4389,N_6064);
and U8575 (N_8575,N_4783,N_5432);
and U8576 (N_8576,N_6261,N_4731);
nor U8577 (N_8577,N_7116,N_6205);
and U8578 (N_8578,N_5538,N_5700);
and U8579 (N_8579,N_4429,N_7829);
nand U8580 (N_8580,N_7677,N_4887);
or U8581 (N_8581,N_6119,N_6157);
nand U8582 (N_8582,N_4434,N_5956);
nand U8583 (N_8583,N_6347,N_7605);
nand U8584 (N_8584,N_5750,N_4431);
nor U8585 (N_8585,N_7225,N_6102);
or U8586 (N_8586,N_7740,N_6357);
and U8587 (N_8587,N_4232,N_7930);
nor U8588 (N_8588,N_5300,N_6889);
nand U8589 (N_8589,N_7063,N_6929);
nand U8590 (N_8590,N_6255,N_4123);
and U8591 (N_8591,N_7459,N_5644);
or U8592 (N_8592,N_4405,N_4258);
nand U8593 (N_8593,N_4869,N_4263);
nor U8594 (N_8594,N_7641,N_5207);
nor U8595 (N_8595,N_7463,N_7755);
nor U8596 (N_8596,N_7627,N_5941);
nor U8597 (N_8597,N_7540,N_6189);
nor U8598 (N_8598,N_5671,N_4625);
and U8599 (N_8599,N_6591,N_5891);
nand U8600 (N_8600,N_6123,N_4081);
nand U8601 (N_8601,N_4657,N_5006);
and U8602 (N_8602,N_6427,N_5872);
nand U8603 (N_8603,N_6042,N_5742);
nand U8604 (N_8604,N_6016,N_4990);
and U8605 (N_8605,N_7281,N_4204);
nor U8606 (N_8606,N_6211,N_5609);
nand U8607 (N_8607,N_5662,N_4819);
nand U8608 (N_8608,N_4742,N_4915);
and U8609 (N_8609,N_7490,N_4543);
nor U8610 (N_8610,N_4586,N_6717);
nand U8611 (N_8611,N_7477,N_5058);
or U8612 (N_8612,N_4106,N_6492);
nand U8613 (N_8613,N_6162,N_6689);
or U8614 (N_8614,N_5973,N_5591);
nor U8615 (N_8615,N_6966,N_4901);
and U8616 (N_8616,N_4954,N_4925);
xnor U8617 (N_8617,N_6586,N_5171);
and U8618 (N_8618,N_6113,N_7592);
xnor U8619 (N_8619,N_6872,N_4031);
xnor U8620 (N_8620,N_4424,N_7480);
nand U8621 (N_8621,N_4318,N_6307);
and U8622 (N_8622,N_5078,N_7989);
nor U8623 (N_8623,N_6514,N_7303);
nand U8624 (N_8624,N_6133,N_4754);
nand U8625 (N_8625,N_4319,N_4533);
and U8626 (N_8626,N_4302,N_5441);
nand U8627 (N_8627,N_6542,N_6057);
nor U8628 (N_8628,N_6185,N_7557);
and U8629 (N_8629,N_4986,N_6215);
nor U8630 (N_8630,N_4492,N_5801);
nand U8631 (N_8631,N_6792,N_4663);
nor U8632 (N_8632,N_4410,N_6304);
nand U8633 (N_8633,N_5829,N_5586);
and U8634 (N_8634,N_6159,N_4816);
nand U8635 (N_8635,N_6669,N_5634);
nor U8636 (N_8636,N_5307,N_7058);
nor U8637 (N_8637,N_5273,N_4494);
or U8638 (N_8638,N_4433,N_7604);
and U8639 (N_8639,N_7416,N_5410);
nor U8640 (N_8640,N_4668,N_6174);
and U8641 (N_8641,N_7200,N_5625);
and U8642 (N_8642,N_4539,N_7409);
and U8643 (N_8643,N_7385,N_7472);
or U8644 (N_8644,N_6803,N_6061);
or U8645 (N_8645,N_5215,N_5970);
or U8646 (N_8646,N_7173,N_5925);
and U8647 (N_8647,N_7087,N_7131);
nand U8648 (N_8648,N_5929,N_4978);
nand U8649 (N_8649,N_7817,N_5049);
and U8650 (N_8650,N_4466,N_6609);
nand U8651 (N_8651,N_6506,N_7668);
and U8652 (N_8652,N_7097,N_6894);
nor U8653 (N_8653,N_6960,N_4450);
and U8654 (N_8654,N_4917,N_7631);
and U8655 (N_8655,N_6626,N_6356);
nor U8656 (N_8656,N_6017,N_4077);
or U8657 (N_8657,N_4961,N_4486);
and U8658 (N_8658,N_7854,N_5436);
or U8659 (N_8659,N_5562,N_7026);
or U8660 (N_8660,N_4160,N_5068);
xor U8661 (N_8661,N_4304,N_6686);
nand U8662 (N_8662,N_4222,N_7080);
and U8663 (N_8663,N_4074,N_6390);
or U8664 (N_8664,N_5536,N_7325);
and U8665 (N_8665,N_7434,N_5965);
nand U8666 (N_8666,N_5648,N_4958);
xor U8667 (N_8667,N_6660,N_5306);
and U8668 (N_8668,N_7869,N_6942);
nand U8669 (N_8669,N_5340,N_7375);
nand U8670 (N_8670,N_7976,N_5105);
nand U8671 (N_8671,N_7340,N_7886);
or U8672 (N_8672,N_6485,N_6924);
and U8673 (N_8673,N_5353,N_5661);
and U8674 (N_8674,N_7552,N_4039);
or U8675 (N_8675,N_7724,N_6270);
nor U8676 (N_8676,N_4933,N_7310);
xor U8677 (N_8677,N_6262,N_6923);
or U8678 (N_8678,N_4134,N_4248);
or U8679 (N_8679,N_6216,N_7077);
and U8680 (N_8680,N_7455,N_4357);
or U8681 (N_8681,N_5136,N_6129);
and U8682 (N_8682,N_6104,N_5057);
nand U8683 (N_8683,N_7868,N_6289);
nor U8684 (N_8684,N_6284,N_4696);
nor U8685 (N_8685,N_6272,N_7654);
xor U8686 (N_8686,N_7885,N_6912);
and U8687 (N_8687,N_4468,N_6029);
nand U8688 (N_8688,N_7577,N_6483);
or U8689 (N_8689,N_4602,N_4095);
nand U8690 (N_8690,N_6043,N_4276);
and U8691 (N_8691,N_6570,N_4301);
or U8692 (N_8692,N_7646,N_4620);
nand U8693 (N_8693,N_7193,N_4268);
nor U8694 (N_8694,N_5237,N_4992);
and U8695 (N_8695,N_6764,N_6535);
nand U8696 (N_8696,N_6498,N_7432);
nand U8697 (N_8697,N_7634,N_5681);
or U8698 (N_8698,N_7743,N_6982);
and U8699 (N_8699,N_4899,N_7440);
and U8700 (N_8700,N_6175,N_7844);
nand U8701 (N_8701,N_7355,N_4253);
nand U8702 (N_8702,N_5908,N_6901);
and U8703 (N_8703,N_7861,N_4206);
nand U8704 (N_8704,N_4080,N_7263);
and U8705 (N_8705,N_5992,N_4946);
nor U8706 (N_8706,N_4640,N_4687);
or U8707 (N_8707,N_7911,N_7822);
nand U8708 (N_8708,N_5850,N_6450);
nand U8709 (N_8709,N_4251,N_5916);
and U8710 (N_8710,N_7156,N_4998);
nand U8711 (N_8711,N_5772,N_5329);
or U8712 (N_8712,N_4553,N_6763);
or U8713 (N_8713,N_5040,N_7838);
and U8714 (N_8714,N_6981,N_4717);
and U8715 (N_8715,N_6245,N_5725);
and U8716 (N_8716,N_5366,N_7341);
or U8717 (N_8717,N_4975,N_7522);
nand U8718 (N_8718,N_7757,N_4265);
or U8719 (N_8719,N_7760,N_4982);
and U8720 (N_8720,N_5333,N_5294);
or U8721 (N_8721,N_5553,N_7727);
xnor U8722 (N_8722,N_4606,N_4452);
and U8723 (N_8723,N_5133,N_5217);
nand U8724 (N_8724,N_5614,N_4618);
or U8725 (N_8725,N_6921,N_5371);
nor U8726 (N_8726,N_6905,N_7601);
and U8727 (N_8727,N_4070,N_4495);
nor U8728 (N_8728,N_7357,N_5153);
or U8729 (N_8729,N_6804,N_4286);
or U8730 (N_8730,N_4505,N_5210);
and U8731 (N_8731,N_7473,N_7543);
and U8732 (N_8732,N_6888,N_7937);
and U8733 (N_8733,N_4172,N_7860);
and U8734 (N_8734,N_6986,N_7461);
or U8735 (N_8735,N_4038,N_7956);
xor U8736 (N_8736,N_5846,N_5697);
and U8737 (N_8737,N_5396,N_6161);
and U8738 (N_8738,N_4534,N_4088);
nor U8739 (N_8739,N_4367,N_7912);
xnor U8740 (N_8740,N_4116,N_6762);
nor U8741 (N_8741,N_7020,N_6209);
nor U8742 (N_8742,N_4395,N_5091);
or U8743 (N_8743,N_4005,N_4048);
nand U8744 (N_8744,N_6596,N_6897);
and U8745 (N_8745,N_5492,N_6956);
or U8746 (N_8746,N_5841,N_5269);
nor U8747 (N_8747,N_5758,N_4624);
nand U8748 (N_8748,N_7442,N_4058);
or U8749 (N_8749,N_7774,N_6493);
nor U8750 (N_8750,N_7571,N_7476);
nor U8751 (N_8751,N_7588,N_5386);
or U8752 (N_8752,N_5587,N_6473);
nor U8753 (N_8753,N_4079,N_5875);
xor U8754 (N_8754,N_6006,N_4361);
nand U8755 (N_8755,N_5244,N_7165);
nand U8756 (N_8756,N_5182,N_6690);
nor U8757 (N_8757,N_6841,N_7835);
or U8758 (N_8758,N_6033,N_4196);
nor U8759 (N_8759,N_7513,N_4818);
xnor U8760 (N_8760,N_4549,N_5383);
xnor U8761 (N_8761,N_6411,N_7883);
nor U8762 (N_8762,N_7541,N_5664);
nor U8763 (N_8763,N_6580,N_6086);
and U8764 (N_8764,N_4798,N_4441);
or U8765 (N_8765,N_4810,N_5413);
nand U8766 (N_8766,N_6503,N_7719);
nand U8767 (N_8767,N_6629,N_4096);
nand U8768 (N_8768,N_7519,N_6437);
nor U8769 (N_8769,N_4779,N_6035);
nand U8770 (N_8770,N_7572,N_6331);
nor U8771 (N_8771,N_5517,N_5673);
and U8772 (N_8772,N_4949,N_5415);
xor U8773 (N_8773,N_6746,N_7786);
xor U8774 (N_8774,N_4439,N_4188);
nor U8775 (N_8775,N_7872,N_5905);
nor U8776 (N_8776,N_4014,N_6729);
and U8777 (N_8777,N_5378,N_5438);
nand U8778 (N_8778,N_4448,N_4822);
nor U8779 (N_8779,N_6578,N_5077);
nor U8780 (N_8780,N_7826,N_5582);
nand U8781 (N_8781,N_4571,N_4800);
nand U8782 (N_8782,N_6968,N_7452);
or U8783 (N_8783,N_7554,N_4556);
or U8784 (N_8784,N_7593,N_5281);
nor U8785 (N_8785,N_5647,N_4743);
nor U8786 (N_8786,N_7024,N_6969);
nand U8787 (N_8787,N_4884,N_7067);
nor U8788 (N_8788,N_5734,N_6066);
and U8789 (N_8789,N_6446,N_4491);
nand U8790 (N_8790,N_5995,N_6903);
nor U8791 (N_8791,N_4478,N_6958);
nand U8792 (N_8792,N_6381,N_6725);
nor U8793 (N_8793,N_5251,N_4776);
and U8794 (N_8794,N_7811,N_6603);
or U8795 (N_8795,N_7752,N_6595);
or U8796 (N_8796,N_6282,N_5071);
and U8797 (N_8797,N_4676,N_6597);
and U8798 (N_8798,N_7671,N_6973);
or U8799 (N_8799,N_6067,N_5042);
and U8800 (N_8800,N_6715,N_7551);
nor U8801 (N_8801,N_5539,N_4159);
nor U8802 (N_8802,N_5110,N_5633);
or U8803 (N_8803,N_6314,N_7292);
and U8804 (N_8804,N_4619,N_4956);
nand U8805 (N_8805,N_4519,N_7971);
and U8806 (N_8806,N_5404,N_6350);
nor U8807 (N_8807,N_4897,N_5512);
and U8808 (N_8808,N_5708,N_7722);
or U8809 (N_8809,N_4378,N_6202);
and U8810 (N_8810,N_7208,N_5225);
nand U8811 (N_8811,N_6692,N_4770);
or U8812 (N_8812,N_4288,N_5544);
nor U8813 (N_8813,N_4479,N_5807);
and U8814 (N_8814,N_4834,N_6623);
and U8815 (N_8815,N_6201,N_7090);
xor U8816 (N_8816,N_7534,N_6663);
or U8817 (N_8817,N_5031,N_4635);
or U8818 (N_8818,N_7134,N_6134);
nand U8819 (N_8819,N_4849,N_4236);
nand U8820 (N_8820,N_7262,N_7952);
nor U8821 (N_8821,N_4289,N_5542);
or U8822 (N_8822,N_4910,N_7585);
nand U8823 (N_8823,N_7900,N_6952);
or U8824 (N_8824,N_4678,N_4094);
nand U8825 (N_8825,N_7119,N_4943);
nand U8826 (N_8826,N_7234,N_5952);
and U8827 (N_8827,N_6116,N_5369);
xnor U8828 (N_8828,N_5402,N_7580);
nand U8829 (N_8829,N_7237,N_4401);
nor U8830 (N_8830,N_4328,N_4474);
or U8831 (N_8831,N_5316,N_5845);
or U8832 (N_8832,N_5559,N_4962);
and U8833 (N_8833,N_5852,N_7701);
and U8834 (N_8834,N_7510,N_5812);
or U8835 (N_8835,N_4118,N_5718);
and U8836 (N_8836,N_4380,N_5621);
nor U8837 (N_8837,N_6391,N_4690);
xor U8838 (N_8838,N_4597,N_4198);
nor U8839 (N_8839,N_6996,N_4908);
nor U8840 (N_8840,N_4649,N_6184);
nand U8841 (N_8841,N_5214,N_6436);
or U8842 (N_8842,N_7391,N_6524);
nor U8843 (N_8843,N_6073,N_4432);
or U8844 (N_8844,N_4514,N_7548);
and U8845 (N_8845,N_5087,N_7011);
nor U8846 (N_8846,N_7697,N_5636);
or U8847 (N_8847,N_6537,N_5147);
nand U8848 (N_8848,N_4683,N_6444);
nand U8849 (N_8849,N_5887,N_6131);
xor U8850 (N_8850,N_4164,N_7990);
and U8851 (N_8851,N_7754,N_7767);
xor U8852 (N_8852,N_5645,N_6079);
and U8853 (N_8853,N_6136,N_6728);
or U8854 (N_8854,N_7290,N_6737);
and U8855 (N_8855,N_6489,N_4820);
and U8856 (N_8856,N_4043,N_4033);
and U8857 (N_8857,N_4609,N_6099);
or U8858 (N_8858,N_4704,N_7076);
nand U8859 (N_8859,N_6891,N_4616);
nor U8860 (N_8860,N_4343,N_6012);
and U8861 (N_8861,N_7112,N_7497);
or U8862 (N_8862,N_7382,N_6587);
or U8863 (N_8863,N_7729,N_7161);
and U8864 (N_8864,N_6967,N_7187);
nand U8865 (N_8865,N_6132,N_4748);
or U8866 (N_8866,N_6734,N_4872);
or U8867 (N_8867,N_4756,N_7749);
and U8868 (N_8868,N_6566,N_4738);
nand U8869 (N_8869,N_5720,N_6126);
nand U8870 (N_8870,N_5095,N_5754);
nor U8871 (N_8871,N_4114,N_7436);
and U8872 (N_8872,N_4152,N_5776);
nand U8873 (N_8873,N_6271,N_7629);
xnor U8874 (N_8874,N_5067,N_6749);
and U8875 (N_8875,N_4610,N_7311);
and U8876 (N_8876,N_4541,N_5401);
or U8877 (N_8877,N_5842,N_6649);
or U8878 (N_8878,N_4726,N_7947);
nand U8879 (N_8879,N_5779,N_6909);
and U8880 (N_8880,N_6631,N_6420);
or U8881 (N_8881,N_5341,N_5173);
xnor U8882 (N_8882,N_6641,N_5073);
and U8883 (N_8883,N_7486,N_7765);
and U8884 (N_8884,N_7367,N_6576);
nand U8885 (N_8885,N_5362,N_6531);
or U8886 (N_8886,N_7784,N_7564);
xor U8887 (N_8887,N_4797,N_4064);
or U8888 (N_8888,N_4656,N_5893);
nand U8889 (N_8889,N_5419,N_4653);
or U8890 (N_8890,N_5857,N_5858);
xor U8891 (N_8891,N_5392,N_6490);
nor U8892 (N_8892,N_6517,N_7176);
nand U8893 (N_8893,N_6674,N_4558);
and U8894 (N_8894,N_5156,N_7715);
or U8895 (N_8895,N_5526,N_6441);
and U8896 (N_8896,N_6720,N_6825);
or U8897 (N_8897,N_6890,N_6237);
and U8898 (N_8898,N_4520,N_7241);
nor U8899 (N_8899,N_6477,N_5596);
and U8900 (N_8900,N_7252,N_6247);
or U8901 (N_8901,N_6263,N_4591);
and U8902 (N_8902,N_7703,N_5450);
nand U8903 (N_8903,N_5498,N_4414);
nor U8904 (N_8904,N_4837,N_6955);
or U8905 (N_8905,N_6954,N_7583);
or U8906 (N_8906,N_4194,N_5996);
or U8907 (N_8907,N_5961,N_6854);
nor U8908 (N_8908,N_6386,N_4297);
and U8909 (N_8909,N_4920,N_7747);
or U8910 (N_8910,N_6068,N_6684);
nor U8911 (N_8911,N_6092,N_7092);
nand U8912 (N_8912,N_4900,N_7363);
and U8913 (N_8913,N_4221,N_7873);
and U8914 (N_8914,N_7479,N_6265);
or U8915 (N_8915,N_4898,N_7273);
nor U8916 (N_8916,N_5886,N_4363);
and U8917 (N_8917,N_5437,N_6329);
and U8918 (N_8918,N_4499,N_6957);
nand U8919 (N_8919,N_4278,N_7682);
or U8920 (N_8920,N_4594,N_6256);
and U8921 (N_8921,N_6983,N_6900);
nand U8922 (N_8922,N_5985,N_6675);
nor U8923 (N_8923,N_5518,N_7938);
nand U8924 (N_8924,N_5770,N_4952);
xor U8925 (N_8925,N_4777,N_6965);
nor U8926 (N_8926,N_7692,N_6040);
nand U8927 (N_8927,N_7192,N_7908);
or U8928 (N_8928,N_7108,N_5945);
nor U8929 (N_8929,N_4063,N_6708);
xor U8930 (N_8930,N_4893,N_6412);
nand U8931 (N_8931,N_5209,N_4880);
or U8932 (N_8932,N_4332,N_6228);
or U8933 (N_8933,N_7615,N_4294);
or U8934 (N_8934,N_6366,N_4493);
and U8935 (N_8935,N_6995,N_5145);
and U8936 (N_8936,N_5365,N_7493);
and U8937 (N_8937,N_5197,N_7070);
and U8938 (N_8938,N_4814,N_5219);
nor U8939 (N_8939,N_7247,N_7137);
or U8940 (N_8940,N_7954,N_7863);
and U8941 (N_8941,N_7862,N_5889);
or U8942 (N_8942,N_6750,N_7398);
nor U8943 (N_8943,N_6118,N_4185);
nor U8944 (N_8944,N_7230,N_6831);
nor U8945 (N_8945,N_4997,N_6413);
xor U8946 (N_8946,N_5443,N_6378);
or U8947 (N_8947,N_5631,N_5702);
nand U8948 (N_8948,N_7035,N_5610);
xor U8949 (N_8949,N_5069,N_5314);
nor U8950 (N_8950,N_7411,N_4298);
xor U8951 (N_8951,N_4542,N_7793);
nor U8952 (N_8952,N_5885,N_6254);
or U8953 (N_8953,N_4786,N_4739);
or U8954 (N_8954,N_4804,N_7674);
xnor U8955 (N_8955,N_5044,N_4358);
or U8956 (N_8956,N_4252,N_7308);
nor U8957 (N_8957,N_7965,N_5160);
nand U8958 (N_8958,N_5912,N_4720);
and U8959 (N_8959,N_6620,N_5280);
nor U8960 (N_8960,N_5454,N_4563);
or U8961 (N_8961,N_7239,N_7056);
and U8962 (N_8962,N_4919,N_6985);
nand U8963 (N_8963,N_7624,N_7521);
nor U8964 (N_8964,N_4692,N_7235);
nand U8965 (N_8965,N_6056,N_5435);
nor U8966 (N_8966,N_5545,N_6934);
or U8967 (N_8967,N_7168,N_7773);
nand U8968 (N_8968,N_6705,N_7055);
nand U8969 (N_8969,N_5100,N_7484);
nor U8970 (N_8970,N_5268,N_6795);
nand U8971 (N_8971,N_6915,N_7404);
and U8972 (N_8972,N_4166,N_7902);
or U8973 (N_8973,N_7742,N_6502);
and U8974 (N_8974,N_5183,N_6797);
nor U8975 (N_8975,N_5184,N_5260);
or U8976 (N_8976,N_6479,N_6808);
and U8977 (N_8977,N_5819,N_4873);
xnor U8978 (N_8978,N_5571,N_5966);
or U8979 (N_8979,N_6896,N_4264);
nor U8980 (N_8980,N_5377,N_6801);
and U8981 (N_8981,N_5046,N_6060);
and U8982 (N_8982,N_5021,N_6138);
nor U8983 (N_8983,N_4246,N_6021);
or U8984 (N_8984,N_6870,N_5394);
xor U8985 (N_8985,N_4716,N_5714);
nand U8986 (N_8986,N_7905,N_6249);
or U8987 (N_8987,N_7337,N_4845);
nand U8988 (N_8988,N_7482,N_5149);
or U8989 (N_8989,N_4544,N_5250);
nand U8990 (N_8990,N_7258,N_4719);
xor U8991 (N_8991,N_7987,N_6606);
or U8992 (N_8992,N_5084,N_6768);
and U8993 (N_8993,N_7462,N_6736);
nand U8994 (N_8994,N_4644,N_5025);
or U8995 (N_8995,N_5381,N_7758);
or U8996 (N_8996,N_4238,N_7597);
xor U8997 (N_8997,N_4918,N_7491);
nor U8998 (N_8998,N_6593,N_6552);
nand U8999 (N_8999,N_6308,N_4670);
nor U9000 (N_9000,N_5034,N_6183);
nor U9001 (N_9001,N_5555,N_4010);
nor U9002 (N_9002,N_7145,N_4838);
and U9003 (N_9003,N_6949,N_7422);
nand U9004 (N_9004,N_4145,N_5584);
or U9005 (N_9005,N_6926,N_5179);
and U9006 (N_9006,N_4409,N_6139);
and U9007 (N_9007,N_6628,N_4913);
or U9008 (N_9008,N_4926,N_5838);
nand U9009 (N_9009,N_6602,N_7454);
or U9010 (N_9010,N_6592,N_6148);
nand U9011 (N_9011,N_7043,N_6571);
nand U9012 (N_9012,N_7348,N_7379);
or U9013 (N_9013,N_7889,N_7878);
or U9014 (N_9014,N_4813,N_7553);
and U9015 (N_9015,N_4643,N_6250);
and U9016 (N_9016,N_6678,N_5484);
xor U9017 (N_9017,N_5155,N_6855);
and U9018 (N_9018,N_5581,N_6582);
and U9019 (N_9019,N_5728,N_4144);
nor U9020 (N_9020,N_4465,N_5859);
nand U9021 (N_9021,N_7431,N_5731);
and U9022 (N_9022,N_7392,N_7250);
xor U9023 (N_9023,N_4780,N_5224);
nand U9024 (N_9024,N_7249,N_4641);
nand U9025 (N_9025,N_4645,N_5072);
and U9026 (N_9026,N_6585,N_4315);
or U9027 (N_9027,N_4377,N_5114);
xnor U9028 (N_9028,N_5408,N_6013);
xor U9029 (N_9029,N_5592,N_4601);
nor U9030 (N_9030,N_6474,N_6951);
or U9031 (N_9031,N_5258,N_4902);
and U9032 (N_9032,N_4458,N_5028);
nor U9033 (N_9033,N_7017,N_7904);
or U9034 (N_9034,N_7393,N_7644);
and U9035 (N_9035,N_7591,N_5579);
nand U9036 (N_9036,N_4883,N_5143);
xor U9037 (N_9037,N_6165,N_4402);
nand U9038 (N_9038,N_6382,N_7074);
and U9039 (N_9039,N_6950,N_5308);
and U9040 (N_9040,N_7733,N_4354);
nor U9041 (N_9041,N_5809,N_7494);
nor U9042 (N_9042,N_4445,N_6455);
and U9043 (N_9043,N_5619,N_5530);
xnor U9044 (N_9044,N_6974,N_4306);
nand U9045 (N_9045,N_5627,N_4346);
and U9046 (N_9046,N_6423,N_4303);
nand U9047 (N_9047,N_5504,N_4290);
nand U9048 (N_9048,N_7057,N_6815);
and U9049 (N_9049,N_4073,N_5196);
nand U9050 (N_9050,N_4209,N_7144);
nor U9051 (N_9051,N_5654,N_6475);
or U9052 (N_9052,N_4207,N_7857);
nor U9053 (N_9053,N_5311,N_5684);
nor U9054 (N_9054,N_5909,N_5132);
and U9055 (N_9055,N_4847,N_4213);
or U9056 (N_9056,N_4659,N_5705);
and U9057 (N_9057,N_5769,N_4032);
nand U9058 (N_9058,N_5162,N_4462);
or U9059 (N_9059,N_5146,N_7562);
nor U9060 (N_9060,N_7635,N_5949);
xnor U9061 (N_9061,N_5297,N_5534);
nand U9062 (N_9062,N_6187,N_5856);
nor U9063 (N_9063,N_4383,N_6433);
nand U9064 (N_9064,N_7511,N_7103);
nand U9065 (N_9065,N_6003,N_7621);
nor U9066 (N_9066,N_5447,N_4840);
nand U9067 (N_9067,N_7950,N_4137);
nand U9068 (N_9068,N_6698,N_5910);
and U9069 (N_9069,N_6218,N_4937);
and U9070 (N_9070,N_5089,N_6022);
and U9071 (N_9071,N_6337,N_4210);
or U9072 (N_9072,N_7931,N_5791);
and U9073 (N_9073,N_7856,N_5774);
or U9074 (N_9074,N_6771,N_4791);
and U9075 (N_9075,N_5551,N_6847);
and U9076 (N_9076,N_7921,N_4529);
and U9077 (N_9077,N_4865,N_4871);
nand U9078 (N_9078,N_6309,N_4848);
or U9079 (N_9079,N_6396,N_4148);
nor U9080 (N_9080,N_4803,N_7613);
nor U9081 (N_9081,N_6236,N_6115);
or U9082 (N_9082,N_5685,N_6600);
nor U9083 (N_9083,N_5879,N_5236);
nand U9084 (N_9084,N_4942,N_7111);
and U9085 (N_9085,N_5737,N_7693);
nor U9086 (N_9086,N_5319,N_4027);
nand U9087 (N_9087,N_7229,N_6939);
nor U9088 (N_9088,N_6327,N_7286);
and U9089 (N_9089,N_4707,N_5391);
nor U9090 (N_9090,N_7069,N_6176);
nor U9091 (N_9091,N_5053,N_7336);
or U9092 (N_9092,N_6697,N_5462);
nor U9093 (N_9093,N_4758,N_6480);
and U9094 (N_9094,N_7639,N_7827);
nor U9095 (N_9095,N_7576,N_7148);
and U9096 (N_9096,N_5039,N_4168);
nand U9097 (N_9097,N_6301,N_6377);
nor U9098 (N_9098,N_7015,N_5546);
and U9099 (N_9099,N_6036,N_4605);
nand U9100 (N_9100,N_7526,N_6997);
or U9101 (N_9101,N_5430,N_7417);
and U9102 (N_9102,N_4658,N_7048);
or U9103 (N_9103,N_6523,N_5024);
or U9104 (N_9104,N_6128,N_4896);
nor U9105 (N_9105,N_6178,N_7687);
or U9106 (N_9106,N_6702,N_7376);
xor U9107 (N_9107,N_5240,N_6819);
xor U9108 (N_9108,N_6744,N_4199);
nor U9109 (N_9109,N_7437,N_6188);
nand U9110 (N_9110,N_7284,N_6775);
nor U9111 (N_9111,N_7101,N_5335);
nand U9112 (N_9112,N_6487,N_4271);
and U9113 (N_9113,N_6704,N_5826);
and U9114 (N_9114,N_7542,N_7804);
and U9115 (N_9115,N_4522,N_5960);
or U9116 (N_9116,N_4076,N_5373);
and U9117 (N_9117,N_6008,N_4331);
nand U9118 (N_9118,N_7936,N_7656);
nand U9119 (N_9119,N_4501,N_7660);
xnor U9120 (N_9120,N_6980,N_7242);
and U9121 (N_9121,N_6575,N_5997);
and U9122 (N_9122,N_5827,N_5159);
nand U9123 (N_9123,N_4274,N_5050);
and U9124 (N_9124,N_5317,N_5144);
or U9125 (N_9125,N_5379,N_4868);
or U9126 (N_9126,N_4215,N_7672);
xnor U9127 (N_9127,N_7424,N_4599);
and U9128 (N_9128,N_4755,N_7085);
nand U9129 (N_9129,N_5863,N_6612);
nor U9130 (N_9130,N_7068,N_7776);
nand U9131 (N_9131,N_4293,N_4500);
and U9132 (N_9132,N_6550,N_4099);
nand U9133 (N_9133,N_7158,N_4593);
nand U9134 (N_9134,N_6555,N_4338);
or U9135 (N_9135,N_4326,N_5367);
or U9136 (N_9136,N_5334,N_5427);
or U9137 (N_9137,N_6438,N_7364);
or U9138 (N_9138,N_5713,N_6398);
and U9139 (N_9139,N_5232,N_4680);
nand U9140 (N_9140,N_5285,N_7970);
nor U9141 (N_9141,N_5924,N_6365);
nor U9142 (N_9142,N_4098,N_6685);
or U9143 (N_9143,N_5678,N_4700);
or U9144 (N_9144,N_7366,N_6325);
nand U9145 (N_9145,N_5940,N_4627);
nor U9146 (N_9146,N_4538,N_4484);
nor U9147 (N_9147,N_6843,N_5376);
or U9148 (N_9148,N_4218,N_4227);
or U9149 (N_9149,N_6495,N_6050);
nand U9150 (N_9150,N_7679,N_5485);
and U9151 (N_9151,N_5870,N_4113);
nor U9152 (N_9152,N_7532,N_4939);
xor U9153 (N_9153,N_5139,N_4948);
or U9154 (N_9154,N_6408,N_6235);
xor U9155 (N_9155,N_7907,N_6822);
nor U9156 (N_9156,N_6397,N_5884);
nor U9157 (N_9157,N_5998,N_6153);
or U9158 (N_9158,N_5233,N_6823);
and U9159 (N_9159,N_4651,N_5778);
nand U9160 (N_9160,N_4671,N_4535);
or U9161 (N_9161,N_7403,N_5806);
nand U9162 (N_9162,N_5590,N_5615);
or U9163 (N_9163,N_5706,N_4400);
and U9164 (N_9164,N_5656,N_7874);
nand U9165 (N_9165,N_7967,N_7150);
or U9166 (N_9166,N_7836,N_5346);
or U9167 (N_9167,N_6917,N_6192);
or U9168 (N_9168,N_7091,N_4345);
xor U9169 (N_9169,N_5676,N_6911);
and U9170 (N_9170,N_7782,N_5520);
nor U9171 (N_9171,N_4506,N_4041);
or U9172 (N_9172,N_7880,N_4285);
or U9173 (N_9173,N_4279,N_6920);
or U9174 (N_9174,N_7402,N_6144);
or U9175 (N_9175,N_7994,N_6758);
nor U9176 (N_9176,N_4277,N_6793);
nand U9177 (N_9177,N_7184,N_6716);
nor U9178 (N_9178,N_5902,N_6358);
or U9179 (N_9179,N_7053,N_4701);
nor U9180 (N_9180,N_6878,N_6835);
xnor U9181 (N_9181,N_5348,N_4337);
or U9182 (N_9182,N_7468,N_6927);
nor U9183 (N_9183,N_6367,N_6348);
nand U9184 (N_9184,N_6499,N_6084);
xnor U9185 (N_9185,N_4581,N_6594);
nand U9186 (N_9186,N_4457,N_5595);
or U9187 (N_9187,N_5570,N_6088);
nand U9188 (N_9188,N_7339,N_7708);
nand U9189 (N_9189,N_5880,N_6058);
nor U9190 (N_9190,N_6994,N_5439);
and U9191 (N_9191,N_5304,N_6931);
nor U9192 (N_9192,N_7041,N_4793);
and U9193 (N_9193,N_7466,N_6987);
or U9194 (N_9194,N_4515,N_4115);
or U9195 (N_9195,N_4053,N_5616);
xor U9196 (N_9196,N_6401,N_7563);
nor U9197 (N_9197,N_5245,N_6197);
or U9198 (N_9198,N_6543,N_6605);
or U9199 (N_9199,N_7658,N_6362);
and U9200 (N_9200,N_7651,N_7745);
nor U9201 (N_9201,N_4327,N_6395);
and U9202 (N_9202,N_6449,N_4523);
or U9203 (N_9203,N_7345,N_5361);
or U9204 (N_9204,N_7858,N_4283);
and U9205 (N_9205,N_4049,N_6680);
nand U9206 (N_9206,N_4639,N_5479);
or U9207 (N_9207,N_4735,N_7276);
nor U9208 (N_9208,N_7065,N_6837);
xor U9209 (N_9209,N_7841,N_6418);
nor U9210 (N_9210,N_7761,N_7483);
or U9211 (N_9211,N_5047,N_6277);
nor U9212 (N_9212,N_6458,N_4626);
xnor U9213 (N_9213,N_6096,N_4060);
nand U9214 (N_9214,N_4393,N_5937);
or U9215 (N_9215,N_7105,N_4022);
nand U9216 (N_9216,N_7848,N_7448);
or U9217 (N_9217,N_7923,N_5189);
nand U9218 (N_9218,N_7368,N_4309);
nor U9219 (N_9219,N_7488,N_6501);
or U9220 (N_9220,N_4436,N_5231);
nor U9221 (N_9221,N_5762,N_6916);
or U9222 (N_9222,N_7899,N_7265);
or U9223 (N_9223,N_5541,N_6280);
nand U9224 (N_9224,N_4072,N_6833);
or U9225 (N_9225,N_7516,N_5789);
or U9226 (N_9226,N_5103,N_6618);
nand U9227 (N_9227,N_4229,N_6300);
or U9228 (N_9228,N_4746,N_7334);
xor U9229 (N_9229,N_6368,N_6730);
or U9230 (N_9230,N_6167,N_5524);
nor U9231 (N_9231,N_7139,N_6266);
and U9232 (N_9232,N_7665,N_5817);
or U9233 (N_9233,N_4507,N_6990);
nand U9234 (N_9234,N_5420,N_4415);
nor U9235 (N_9235,N_5568,N_7753);
nand U9236 (N_9236,N_6194,N_6936);
and U9237 (N_9237,N_6733,N_4966);
nand U9238 (N_9238,N_5328,N_4037);
and U9239 (N_9239,N_4562,N_6222);
nor U9240 (N_9240,N_4580,N_4866);
nand U9241 (N_9241,N_5865,N_5715);
nand U9242 (N_9242,N_4412,N_7589);
nand U9243 (N_9243,N_4598,N_7953);
or U9244 (N_9244,N_6695,N_5557);
or U9245 (N_9245,N_7324,N_5148);
nand U9246 (N_9246,N_6070,N_7152);
nand U9247 (N_9247,N_6410,N_7309);
nand U9248 (N_9248,N_6824,N_6569);
xnor U9249 (N_9249,N_5295,N_5343);
or U9250 (N_9250,N_5585,N_5299);
nand U9251 (N_9251,N_6959,N_7958);
nand U9252 (N_9252,N_6124,N_7223);
or U9253 (N_9253,N_7147,N_5726);
nand U9254 (N_9254,N_7555,N_5934);
and U9255 (N_9255,N_5085,N_7974);
nand U9256 (N_9256,N_7524,N_5483);
or U9257 (N_9257,N_5687,N_6906);
nor U9258 (N_9258,N_7528,N_6130);
nor U9259 (N_9259,N_7847,N_6442);
nor U9260 (N_9260,N_7955,N_6676);
and U9261 (N_9261,N_4806,N_7896);
nor U9262 (N_9262,N_4875,N_5712);
or U9263 (N_9263,N_7294,N_4824);
or U9264 (N_9264,N_6679,N_6081);
nor U9265 (N_9265,N_5972,N_7130);
nor U9266 (N_9266,N_7027,N_5178);
and U9267 (N_9267,N_6075,N_4767);
nor U9268 (N_9268,N_5606,N_7430);
and U9269 (N_9269,N_6160,N_6047);
nand U9270 (N_9270,N_5111,N_6826);
nand U9271 (N_9271,N_6774,N_6581);
and U9272 (N_9272,N_4225,N_4314);
and U9273 (N_9273,N_5510,N_6563);
or U9274 (N_9274,N_6204,N_4127);
nor U9275 (N_9275,N_6392,N_6163);
or U9276 (N_9276,N_6294,N_4086);
or U9277 (N_9277,N_5474,N_7647);
nor U9278 (N_9278,N_4995,N_5350);
xnor U9279 (N_9279,N_7405,N_5475);
and U9280 (N_9280,N_6154,N_7683);
and U9281 (N_9281,N_5293,N_6375);
and U9282 (N_9282,N_7569,N_5748);
nand U9283 (N_9283,N_7019,N_5794);
nand U9284 (N_9284,N_4718,N_6682);
and U9285 (N_9285,N_4980,N_5834);
nor U9286 (N_9286,N_5385,N_4018);
nor U9287 (N_9287,N_6932,N_4983);
xnor U9288 (N_9288,N_4109,N_6206);
xor U9289 (N_9289,N_5569,N_4905);
nand U9290 (N_9290,N_6089,N_4930);
or U9291 (N_9291,N_7525,N_6748);
nand U9292 (N_9292,N_7690,N_4667);
and U9293 (N_9293,N_7705,N_7211);
or U9294 (N_9294,N_7321,N_7834);
or U9295 (N_9295,N_7673,N_6904);
nand U9296 (N_9296,N_5440,N_7584);
or U9297 (N_9297,N_4760,N_4947);
and U9298 (N_9298,N_5745,N_4530);
nor U9299 (N_9299,N_5009,N_6971);
xnor U9300 (N_9300,N_5257,N_6083);
nand U9301 (N_9301,N_7820,N_7790);
nand U9302 (N_9302,N_6636,N_4843);
xnor U9303 (N_9303,N_7734,N_5564);
or U9304 (N_9304,N_7040,N_4934);
nor U9305 (N_9305,N_4029,N_4351);
or U9306 (N_9306,N_4056,N_5174);
nor U9307 (N_9307,N_7451,N_5987);
xnor U9308 (N_9308,N_7109,N_4762);
nor U9309 (N_9309,N_7312,N_6993);
nand U9310 (N_9310,N_6416,N_7533);
nor U9311 (N_9311,N_7879,N_6177);
nand U9312 (N_9312,N_4861,N_4588);
xor U9313 (N_9313,N_7691,N_6828);
nand U9314 (N_9314,N_7030,N_5971);
xor U9315 (N_9315,N_4165,N_7996);
xnor U9316 (N_9316,N_4026,N_7317);
nand U9317 (N_9317,N_7881,N_5400);
nand U9318 (N_9318,N_5692,N_7333);
nor U9319 (N_9319,N_4867,N_6108);
nor U9320 (N_9320,N_5405,N_7155);
and U9321 (N_9321,N_5356,N_5540);
nand U9322 (N_9322,N_4214,N_5448);
nor U9323 (N_9323,N_5899,N_7054);
nor U9324 (N_9324,N_4652,N_5131);
and U9325 (N_9325,N_4957,N_4548);
nor U9326 (N_9326,N_6613,N_6374);
and U9327 (N_9327,N_4490,N_7814);
or U9328 (N_9328,N_4555,N_5426);
and U9329 (N_9329,N_7032,N_4614);
and U9330 (N_9330,N_5090,N_7775);
nand U9331 (N_9331,N_5800,N_5108);
nor U9332 (N_9332,N_7390,N_6584);
nor U9333 (N_9333,N_6809,N_7606);
nand U9334 (N_9334,N_7380,N_7275);
nor U9335 (N_9335,N_6938,N_7823);
or U9336 (N_9336,N_5172,N_7764);
nor U9337 (N_9337,N_7608,N_6062);
xor U9338 (N_9338,N_5332,N_4217);
nor U9339 (N_9339,N_7973,N_4540);
nor U9340 (N_9340,N_7676,N_4475);
nand U9341 (N_9341,N_7014,N_5493);
nand U9342 (N_9342,N_5680,N_5969);
or U9343 (N_9343,N_4724,N_5709);
or U9344 (N_9344,N_7898,N_4224);
xnor U9345 (N_9345,N_5944,N_5533);
or U9346 (N_9346,N_7098,N_6344);
or U9347 (N_9347,N_4730,N_5764);
nand U9348 (N_9348,N_7172,N_6711);
nor U9349 (N_9349,N_4156,N_7227);
nand U9350 (N_9350,N_4418,N_4333);
or U9351 (N_9351,N_4050,N_6231);
or U9352 (N_9352,N_7643,N_7022);
nor U9353 (N_9353,N_7492,N_4751);
nand U9354 (N_9354,N_4675,N_6668);
nand U9355 (N_9355,N_6529,N_4703);
nor U9356 (N_9356,N_5506,N_6984);
or U9357 (N_9357,N_6288,N_5851);
nor U9358 (N_9358,N_4398,N_6110);
or U9359 (N_9359,N_4831,N_5759);
nand U9360 (N_9360,N_6504,N_5473);
nand U9361 (N_9361,N_4967,N_4421);
nand U9362 (N_9362,N_5839,N_4782);
nand U9363 (N_9363,N_7845,N_5563);
nand U9364 (N_9364,N_7002,N_6461);
or U9365 (N_9365,N_5882,N_4317);
nand U9366 (N_9366,N_7427,N_4654);
and U9367 (N_9367,N_5026,N_7957);
and U9368 (N_9368,N_7146,N_5816);
and U9369 (N_9369,N_6782,N_6496);
nand U9370 (N_9370,N_4531,N_5860);
and U9371 (N_9371,N_5749,N_5686);
nand U9372 (N_9372,N_6488,N_7802);
and U9373 (N_9373,N_4138,N_6651);
nand U9374 (N_9374,N_7496,N_5980);
or U9375 (N_9375,N_7596,N_4440);
nor U9376 (N_9376,N_5818,N_6296);
nor U9377 (N_9377,N_4129,N_7781);
xnor U9378 (N_9378,N_5560,N_7943);
nor U9379 (N_9379,N_5876,N_6240);
and U9380 (N_9380,N_7154,N_6009);
nor U9381 (N_9381,N_7381,N_7267);
nor U9382 (N_9382,N_6756,N_5321);
xnor U9383 (N_9383,N_5928,N_7759);
nand U9384 (N_9384,N_4110,N_6914);
and U9385 (N_9385,N_6521,N_4471);
nor U9386 (N_9386,N_7016,N_4608);
xnor U9387 (N_9387,N_4705,N_4569);
and U9388 (N_9388,N_6470,N_5629);
nand U9389 (N_9389,N_7794,N_6548);
nor U9390 (N_9390,N_7151,N_5008);
xnor U9391 (N_9391,N_7707,N_6039);
and U9392 (N_9392,N_5265,N_7125);
xor U9393 (N_9393,N_7226,N_7470);
xor U9394 (N_9394,N_7328,N_7699);
or U9395 (N_9395,N_6384,N_6151);
nor U9396 (N_9396,N_7669,N_7501);
nand U9397 (N_9397,N_6871,N_7642);
or U9398 (N_9398,N_5208,N_4083);
and U9399 (N_9399,N_6100,N_6607);
nor U9400 (N_9400,N_4969,N_5907);
nand U9401 (N_9401,N_5140,N_4892);
nor U9402 (N_9402,N_4750,N_6258);
xor U9403 (N_9403,N_4100,N_5495);
or U9404 (N_9404,N_7547,N_5079);
nor U9405 (N_9405,N_4753,N_6346);
or U9406 (N_9406,N_5082,N_7073);
nor U9407 (N_9407,N_5967,N_4674);
nor U9408 (N_9408,N_6179,N_4877);
and U9409 (N_9409,N_7710,N_5120);
nand U9410 (N_9410,N_5059,N_4280);
nor U9411 (N_9411,N_6323,N_6654);
and U9412 (N_9412,N_6892,N_6508);
or U9413 (N_9413,N_5849,N_5186);
xnor U9414 (N_9414,N_5938,N_7664);
nor U9415 (N_9415,N_5464,N_7202);
and U9416 (N_9416,N_4023,N_4189);
and U9417 (N_9417,N_4167,N_4360);
or U9418 (N_9418,N_4275,N_7228);
or U9419 (N_9419,N_5815,N_6224);
nand U9420 (N_9420,N_7675,N_7933);
nand U9421 (N_9421,N_7969,N_5913);
or U9422 (N_9422,N_5927,N_6234);
and U9423 (N_9423,N_5164,N_5261);
nor U9424 (N_9424,N_6633,N_7288);
and U9425 (N_9425,N_4745,N_5062);
and U9426 (N_9426,N_4107,N_7233);
or U9427 (N_9427,N_6895,N_5635);
and U9428 (N_9428,N_4513,N_7716);
and U9429 (N_9429,N_4242,N_7181);
and U9430 (N_9430,N_6443,N_4647);
nor U9431 (N_9431,N_6156,N_4582);
nand U9432 (N_9432,N_5787,N_6403);
nand U9433 (N_9433,N_5001,N_6735);
nor U9434 (N_9434,N_5055,N_5926);
nand U9435 (N_9435,N_4112,N_4281);
nand U9436 (N_9436,N_4972,N_5414);
or U9437 (N_9437,N_7717,N_5098);
or U9438 (N_9438,N_6883,N_7785);
or U9439 (N_9439,N_7195,N_5127);
and U9440 (N_9440,N_7666,N_5347);
and U9441 (N_9441,N_5000,N_6101);
nand U9442 (N_9442,N_4989,N_6846);
nor U9443 (N_9443,N_4386,N_5808);
nand U9444 (N_9444,N_7633,N_7277);
or U9445 (N_9445,N_5602,N_6295);
xnor U9446 (N_9446,N_5301,N_4929);
and U9447 (N_9447,N_5351,N_7851);
nor U9448 (N_9448,N_5691,N_6109);
and U9449 (N_9449,N_5421,N_5612);
xnor U9450 (N_9450,N_6860,N_7903);
or U9451 (N_9451,N_4764,N_7220);
nor U9452 (N_9452,N_5222,N_5312);
and U9453 (N_9453,N_4261,N_4310);
and U9454 (N_9454,N_7136,N_4537);
or U9455 (N_9455,N_4991,N_6842);
nor U9456 (N_9456,N_5892,N_7798);
nand U9457 (N_9457,N_7410,N_7347);
or U9458 (N_9458,N_7789,N_7762);
nor U9459 (N_9459,N_6032,N_7413);
and U9460 (N_9460,N_6207,N_7527);
nor U9461 (N_9461,N_7066,N_4085);
and U9462 (N_9462,N_7236,N_5296);
nand U9463 (N_9463,N_5509,N_5646);
and U9464 (N_9464,N_6015,N_7891);
nor U9465 (N_9465,N_7036,N_6848);
xor U9466 (N_9466,N_4101,N_6078);
nand U9467 (N_9467,N_7204,N_5703);
or U9468 (N_9468,N_6180,N_5469);
xnor U9469 (N_9469,N_4567,N_6155);
or U9470 (N_9470,N_5041,N_7300);
nor U9471 (N_9471,N_4826,N_4344);
or U9472 (N_9472,N_5033,N_6225);
and U9473 (N_9473,N_5632,N_7384);
or U9474 (N_9474,N_6777,N_6572);
nand U9475 (N_9475,N_7018,N_7093);
nor U9476 (N_9476,N_4069,N_4374);
xnor U9477 (N_9477,N_6658,N_7840);
and U9478 (N_9478,N_5109,N_7425);
and U9479 (N_9479,N_5689,N_5137);
xnor U9480 (N_9480,N_4339,N_7171);
nor U9481 (N_9481,N_5649,N_7535);
or U9482 (N_9482,N_4708,N_4240);
or U9483 (N_9483,N_4963,N_5345);
nor U9484 (N_9484,N_4078,N_4835);
and U9485 (N_9485,N_4771,N_6645);
nand U9486 (N_9486,N_5287,N_7323);
xor U9487 (N_9487,N_7240,N_5193);
nor U9488 (N_9488,N_6143,N_7941);
or U9489 (N_9489,N_6278,N_6991);
nand U9490 (N_9490,N_7127,N_4524);
xor U9491 (N_9491,N_7523,N_5252);
or U9492 (N_9492,N_6560,N_4244);
nor U9493 (N_9493,N_7756,N_5746);
or U9494 (N_9494,N_7574,N_5624);
nand U9495 (N_9495,N_7700,N_5282);
nor U9496 (N_9496,N_5921,N_4142);
and U9497 (N_9497,N_4231,N_6199);
or U9498 (N_9498,N_5977,N_7206);
xor U9499 (N_9499,N_4184,N_6239);
and U9500 (N_9500,N_7449,N_6311);
nor U9501 (N_9501,N_6696,N_7196);
xnor U9502 (N_9502,N_4066,N_4426);
and U9503 (N_9503,N_7887,N_7439);
nand U9504 (N_9504,N_7509,N_4162);
nor U9505 (N_9505,N_5370,N_6615);
nor U9506 (N_9506,N_4480,N_5733);
or U9507 (N_9507,N_5694,N_6248);
nand U9508 (N_9508,N_7706,N_4985);
nand U9509 (N_9509,N_4104,N_4092);
nand U9510 (N_9510,N_5821,N_7089);
nand U9511 (N_9511,N_7890,N_7791);
nand U9512 (N_9512,N_5695,N_4699);
or U9513 (N_9513,N_6885,N_6090);
nor U9514 (N_9514,N_6127,N_4965);
nand U9515 (N_9515,N_4936,N_4108);
and U9516 (N_9516,N_4143,N_4935);
and U9517 (N_9517,N_7966,N_4727);
nand U9518 (N_9518,N_7342,N_4463);
or U9519 (N_9519,N_6341,N_7359);
xnor U9520 (N_9520,N_6519,N_7696);
nor U9521 (N_9521,N_4416,N_5740);
nor U9522 (N_9522,N_4858,N_6468);
or U9523 (N_9523,N_6451,N_5943);
xnor U9524 (N_9524,N_4336,N_6318);
nand U9525 (N_9525,N_4404,N_6998);
and U9526 (N_9526,N_6011,N_7507);
xnor U9527 (N_9527,N_6267,N_5864);
or U9528 (N_9528,N_6053,N_5588);
and U9529 (N_9529,N_7808,N_4340);
xnor U9530 (N_9530,N_4241,N_7327);
xnor U9531 (N_9531,N_7910,N_4419);
nor U9532 (N_9532,N_4617,N_6097);
xnor U9533 (N_9533,N_4216,N_7962);
and U9534 (N_9534,N_7274,N_4749);
nand U9535 (N_9535,N_5805,N_6393);
nor U9536 (N_9536,N_7610,N_7023);
nor U9537 (N_9537,N_7504,N_7219);
nand U9538 (N_9538,N_7945,N_5580);
and U9539 (N_9539,N_6533,N_4999);
nor U9540 (N_9540,N_5486,N_7059);
or U9541 (N_9541,N_7981,N_6567);
or U9542 (N_9542,N_7979,N_6948);
nor U9543 (N_9543,N_4677,N_6082);
nand U9544 (N_9544,N_7766,N_6583);
nor U9545 (N_9545,N_6399,N_5735);
nor U9546 (N_9546,N_5914,N_4968);
or U9547 (N_9547,N_6851,N_4565);
or U9548 (N_9548,N_4685,N_4262);
and U9549 (N_9549,N_7704,N_6361);
or U9550 (N_9550,N_7897,N_7072);
and U9551 (N_9551,N_5874,N_5667);
or U9552 (N_9552,N_7926,N_6238);
and U9553 (N_9553,N_5497,N_7149);
xor U9554 (N_9554,N_7968,N_4267);
or U9555 (N_9555,N_6334,N_7377);
nand U9556 (N_9556,N_5081,N_6221);
nor U9557 (N_9557,N_7732,N_4282);
nor U9558 (N_9558,N_6345,N_7617);
nand U9559 (N_9559,N_5923,N_5166);
and U9560 (N_9560,N_4057,N_7594);
and U9561 (N_9561,N_6077,N_4621);
nor U9562 (N_9562,N_5489,N_6634);
or U9563 (N_9563,N_5608,N_4455);
nor U9564 (N_9564,N_6836,N_4860);
or U9565 (N_9565,N_6754,N_5375);
nor U9566 (N_9566,N_4200,N_4906);
xnor U9567 (N_9567,N_6625,N_6818);
nand U9568 (N_9568,N_5500,N_5954);
and U9569 (N_9569,N_5784,N_5989);
or U9570 (N_9570,N_6723,N_4235);
nor U9571 (N_9571,N_4368,N_5528);
and U9572 (N_9572,N_5310,N_6166);
xor U9573 (N_9573,N_6171,N_4836);
nand U9574 (N_9574,N_6785,N_4020);
nand U9575 (N_9575,N_4124,N_4103);
nor U9576 (N_9576,N_6937,N_6639);
and U9577 (N_9577,N_5358,N_7283);
or U9578 (N_9578,N_7157,N_5015);
xnor U9579 (N_9579,N_7539,N_4955);
nand U9580 (N_9580,N_6525,N_5630);
and U9581 (N_9581,N_6534,N_6557);
and U9582 (N_9582,N_4477,N_6027);
nor U9583 (N_9583,N_6226,N_5226);
or U9584 (N_9584,N_5291,N_4631);
and U9585 (N_9585,N_4603,N_4807);
or U9586 (N_9586,N_6354,N_5869);
or U9587 (N_9587,N_6770,N_5283);
or U9588 (N_9588,N_5418,N_4150);
or U9589 (N_9589,N_4255,N_5796);
nor U9590 (N_9590,N_6435,N_5505);
and U9591 (N_9591,N_6407,N_5548);
and U9592 (N_9592,N_7544,N_5574);
or U9593 (N_9593,N_6324,N_7920);
or U9594 (N_9594,N_5051,N_7685);
or U9595 (N_9595,N_5305,N_4512);
and U9596 (N_9596,N_7999,N_4021);
and U9597 (N_9597,N_4453,N_5848);
nor U9598 (N_9598,N_5947,N_7335);
nand U9599 (N_9599,N_5157,N_5286);
or U9600 (N_9600,N_4805,N_7825);
and U9601 (N_9601,N_4180,N_5603);
nand U9602 (N_9602,N_6145,N_5254);
or U9603 (N_9603,N_6970,N_6739);
xnor U9604 (N_9604,N_7566,N_7614);
or U9605 (N_9605,N_5323,N_7796);
nor U9606 (N_9606,N_5699,N_7086);
nand U9607 (N_9607,N_5247,N_6732);
nand U9608 (N_9608,N_4895,N_7694);
and U9609 (N_9609,N_5978,N_6579);
nor U9610 (N_9610,N_5990,N_7117);
and U9611 (N_9611,N_6213,N_5192);
nand U9612 (N_9612,N_5942,N_6214);
nor U9613 (N_9613,N_7824,N_4691);
and U9614 (N_9614,N_7102,N_4307);
nor U9615 (N_9615,N_4140,N_7010);
nand U9616 (N_9616,N_7662,N_6210);
nor U9617 (N_9617,N_7568,N_5932);
nor U9618 (N_9618,N_4940,N_6306);
nand U9619 (N_9619,N_7925,N_7253);
nand U9620 (N_9620,N_6469,N_7113);
or U9621 (N_9621,N_4011,N_7034);
or U9622 (N_9622,N_4007,N_7741);
nor U9623 (N_9623,N_4853,N_6293);
nor U9624 (N_9624,N_4646,N_7426);
nand U9625 (N_9625,N_4988,N_7959);
nor U9626 (N_9626,N_6648,N_7415);
or U9627 (N_9627,N_4438,N_5601);
or U9628 (N_9628,N_4481,N_7598);
nor U9629 (N_9629,N_4970,N_7047);
and U9630 (N_9630,N_7100,N_7350);
nand U9631 (N_9631,N_5278,N_4830);
nor U9632 (N_9632,N_5986,N_4030);
or U9633 (N_9633,N_6861,N_4923);
xor U9634 (N_9634,N_6661,N_7344);
nand U9635 (N_9635,N_6510,N_7578);
nand U9636 (N_9636,N_7736,N_5357);
or U9637 (N_9637,N_5005,N_7304);
or U9638 (N_9638,N_4921,N_4928);
or U9639 (N_9639,N_6751,N_5527);
and U9640 (N_9640,N_4916,N_4451);
or U9641 (N_9641,N_5730,N_4157);
and U9642 (N_9642,N_5326,N_4714);
nand U9643 (N_9643,N_5917,N_4012);
nand U9644 (N_9644,N_4710,N_4851);
and U9645 (N_9645,N_6285,N_4839);
nand U9646 (N_9646,N_5655,N_7133);
and U9647 (N_9647,N_4024,N_5216);
nand U9648 (N_9648,N_7725,N_7243);
or U9649 (N_9649,N_6740,N_7689);
nor U9650 (N_9650,N_4781,N_7819);
and U9651 (N_9651,N_6229,N_7166);
and U9652 (N_9652,N_7153,N_5476);
and U9653 (N_9653,N_4702,N_4971);
nand U9654 (N_9654,N_6257,N_4907);
and U9655 (N_9655,N_5123,N_6964);
and U9656 (N_9656,N_7600,N_6757);
or U9657 (N_9657,N_6317,N_4146);
or U9658 (N_9658,N_7803,N_5126);
nand U9659 (N_9659,N_4977,N_5651);
or U9660 (N_9660,N_7680,N_4550);
xor U9661 (N_9661,N_5599,N_6722);
xnor U9662 (N_9662,N_7221,N_5200);
and U9663 (N_9663,N_7832,N_4827);
xor U9664 (N_9664,N_4927,N_5795);
or U9665 (N_9665,N_5653,N_4187);
nor U9666 (N_9666,N_6617,N_5822);
or U9667 (N_9667,N_6193,N_4097);
nand U9668 (N_9668,N_5228,N_7487);
nor U9669 (N_9669,N_7712,N_5030);
or U9670 (N_9670,N_6630,N_5083);
nor U9671 (N_9671,N_6448,N_6972);
or U9672 (N_9672,N_5639,N_4628);
nor U9673 (N_9673,N_7630,N_4392);
nor U9674 (N_9674,N_7370,N_6887);
and U9675 (N_9675,N_7373,N_4003);
nor U9676 (N_9676,N_5847,N_5292);
nor U9677 (N_9677,N_5101,N_5255);
or U9678 (N_9678,N_5395,N_6414);
or U9679 (N_9679,N_4126,N_4723);
or U9680 (N_9680,N_6992,N_7695);
nor U9681 (N_9681,N_5831,N_7044);
nand U9682 (N_9682,N_7190,N_5054);
or U9683 (N_9683,N_7081,N_7039);
nand U9684 (N_9684,N_6376,N_6328);
xnor U9685 (N_9685,N_6943,N_7609);
and U9686 (N_9686,N_7934,N_6276);
nand U9687 (N_9687,N_6380,N_7831);
or U9688 (N_9688,N_4759,N_6405);
and U9689 (N_9689,N_6085,N_6647);
and U9690 (N_9690,N_6332,N_6196);
nand U9691 (N_9691,N_6292,N_4139);
or U9692 (N_9692,N_5743,N_5604);
nor U9693 (N_9693,N_4403,N_5722);
nor U9694 (N_9694,N_5780,N_4461);
or U9695 (N_9695,N_5554,N_4093);
nand U9696 (N_9696,N_7458,N_4356);
nor U9697 (N_9697,N_5431,N_6789);
and U9698 (N_9698,N_6511,N_5962);
nor U9699 (N_9699,N_4369,N_6845);
nor U9700 (N_9700,N_5660,N_4684);
or U9701 (N_9701,N_4579,N_6466);
and U9702 (N_9702,N_4045,N_6798);
nor U9703 (N_9703,N_6046,N_7178);
nand U9704 (N_9704,N_4154,N_6902);
xnor U9705 (N_9705,N_5220,N_5767);
or U9706 (N_9706,N_7266,N_6402);
nor U9707 (N_9707,N_5004,N_7272);
and U9708 (N_9708,N_6018,N_5717);
nand U9709 (N_9709,N_4487,N_4396);
nor U9710 (N_9710,N_7394,N_5387);
or U9711 (N_9711,N_7203,N_6656);
or U9712 (N_9712,N_6687,N_6494);
nor U9713 (N_9713,N_5470,N_5112);
nor U9714 (N_9714,N_6545,N_6640);
nor U9715 (N_9715,N_5572,N_4420);
and U9716 (N_9716,N_6527,N_6146);
and U9717 (N_9717,N_4552,N_6142);
nor U9718 (N_9718,N_5482,N_5032);
nor U9719 (N_9719,N_4359,N_6158);
and U9720 (N_9720,N_4008,N_6551);
nand U9721 (N_9721,N_5711,N_5168);
nand U9722 (N_9722,N_4737,N_7892);
nor U9723 (N_9723,N_4648,N_5481);
nand U9724 (N_9724,N_6023,N_4664);
or U9725 (N_9725,N_6863,N_7322);
nand U9726 (N_9726,N_5690,N_6780);
or U9727 (N_9727,N_5683,N_5119);
nor U9728 (N_9728,N_6321,N_5642);
nand U9729 (N_9729,N_6140,N_4655);
and U9730 (N_9730,N_6359,N_6409);
or U9731 (N_9731,N_4365,N_4600);
nand U9732 (N_9732,N_5901,N_7174);
nor U9733 (N_9733,N_7769,N_5757);
nor U9734 (N_9734,N_4016,N_6786);
xnor U9735 (N_9735,N_7106,N_5180);
nand U9736 (N_9736,N_6532,N_6546);
nor U9737 (N_9737,N_5721,N_6776);
xnor U9738 (N_9738,N_7456,N_6264);
and U9739 (N_9739,N_7833,N_7489);
and U9740 (N_9740,N_7882,N_7052);
or U9741 (N_9741,N_5480,N_7268);
xnor U9742 (N_9742,N_4195,N_5984);
xnor U9743 (N_9743,N_5248,N_7298);
or U9744 (N_9744,N_4442,N_4233);
and U9745 (N_9745,N_5719,N_5999);
and U9746 (N_9746,N_5994,N_5877);
nor U9747 (N_9747,N_7383,N_4417);
nand U9748 (N_9748,N_4147,N_7445);
or U9749 (N_9749,N_5253,N_4713);
and U9750 (N_9750,N_4850,N_5813);
nand U9751 (N_9751,N_7850,N_7388);
and U9752 (N_9752,N_5507,N_5904);
nand U9753 (N_9753,N_6259,N_7457);
nand U9754 (N_9754,N_7993,N_4681);
xor U9755 (N_9755,N_5169,N_6164);
nor U9756 (N_9756,N_6935,N_6432);
or U9757 (N_9757,N_4709,N_7884);
nor U9758 (N_9758,N_7163,N_6335);
nor U9759 (N_9759,N_7474,N_6080);
or U9760 (N_9760,N_6673,N_4034);
nand U9761 (N_9761,N_5425,N_7478);
nor U9762 (N_9762,N_5397,N_7143);
xnor U9763 (N_9763,N_7269,N_5102);
nor U9764 (N_9764,N_7289,N_7360);
or U9765 (N_9765,N_5811,N_7399);
nand U9766 (N_9766,N_6445,N_5773);
nand U9767 (N_9767,N_4467,N_6657);
and U9768 (N_9768,N_7942,N_6505);
nand U9769 (N_9769,N_4388,N_5514);
nand U9770 (N_9770,N_5786,N_5075);
or U9771 (N_9771,N_7238,N_7485);
nand U9772 (N_9772,N_7986,N_5191);
or U9773 (N_9773,N_4778,N_6269);
xnor U9774 (N_9774,N_5181,N_4511);
or U9775 (N_9775,N_4390,N_5830);
and U9776 (N_9776,N_5019,N_7575);
and U9777 (N_9777,N_6941,N_6562);
or U9778 (N_9778,N_4960,N_6094);
nor U9779 (N_9779,N_5467,N_5993);
nand U9780 (N_9780,N_6547,N_7652);
and U9781 (N_9781,N_7088,N_7843);
or U9782 (N_9782,N_6251,N_6541);
and U9783 (N_9783,N_5547,N_6638);
nand U9784 (N_9784,N_6693,N_5698);
nand U9785 (N_9785,N_7189,N_5163);
or U9786 (N_9786,N_7565,N_4829);
xnor U9787 (N_9787,N_4886,N_6806);
and U9788 (N_9788,N_7205,N_4223);
nand U9789 (N_9789,N_6484,N_5979);
nand U9790 (N_9790,N_7888,N_5739);
xnor U9791 (N_9791,N_7618,N_4028);
or U9792 (N_9792,N_6962,N_4633);
or U9793 (N_9793,N_4789,N_7261);
or U9794 (N_9794,N_4102,N_5637);
nand U9795 (N_9795,N_5936,N_7984);
or U9796 (N_9796,N_5976,N_5744);
and U9797 (N_9797,N_4561,N_4174);
and U9798 (N_9798,N_4443,N_7587);
nand U9799 (N_9799,N_6564,N_6844);
nand U9800 (N_9800,N_5107,N_7842);
or U9801 (N_9801,N_7684,N_4068);
or U9802 (N_9802,N_7400,N_7951);
nand U9803 (N_9803,N_6976,N_4870);
nor U9804 (N_9804,N_6355,N_4413);
nor U9805 (N_9805,N_4722,N_4325);
or U9806 (N_9806,N_4260,N_7001);
xor U9807 (N_9807,N_5804,N_7214);
nand U9808 (N_9808,N_6742,N_5151);
and U9809 (N_9809,N_4574,N_4498);
nor U9810 (N_9810,N_7362,N_7412);
or U9811 (N_9811,N_5158,N_5640);
or U9812 (N_9812,N_4864,N_4170);
nor U9813 (N_9813,N_5623,N_4752);
nand U9814 (N_9814,N_4688,N_4372);
nor U9815 (N_9815,N_7084,N_6507);
or U9816 (N_9816,N_6431,N_6667);
nor U9817 (N_9817,N_7419,N_7801);
and U9818 (N_9818,N_6963,N_7927);
xnor U9819 (N_9819,N_7961,N_4397);
nand U9820 (N_9820,N_5364,N_4733);
xnor U9821 (N_9821,N_7545,N_6400);
or U9822 (N_9822,N_7515,N_4953);
nand U9823 (N_9823,N_6589,N_6778);
or U9824 (N_9824,N_7046,N_5532);
and U9825 (N_9825,N_7870,N_5710);
or U9826 (N_9826,N_4859,N_5935);
nor U9827 (N_9827,N_4801,N_6457);
nor U9828 (N_9828,N_5303,N_6859);
nor U9829 (N_9829,N_6830,N_6659);
xnor U9830 (N_9830,N_6274,N_5919);
and U9831 (N_9831,N_6281,N_5503);
nand U9832 (N_9832,N_7104,N_6875);
or U9833 (N_9833,N_5577,N_5315);
and U9834 (N_9834,N_4532,N_4423);
nand U9835 (N_9835,N_6273,N_7730);
nor U9836 (N_9836,N_4790,N_6005);
or U9837 (N_9837,N_7296,N_5823);
nor U9838 (N_9838,N_5471,N_5883);
and U9839 (N_9839,N_4002,N_7917);
xor U9840 (N_9840,N_5290,N_5825);
nor U9841 (N_9841,N_7812,N_5029);
xnor U9842 (N_9842,N_7353,N_4035);
or U9843 (N_9843,N_6219,N_7414);
nand U9844 (N_9844,N_4205,N_7867);
nand U9845 (N_9845,N_5824,N_5670);
nand U9846 (N_9846,N_4856,N_4181);
xor U9847 (N_9847,N_4161,N_5556);
or U9848 (N_9848,N_6632,N_6653);
or U9849 (N_9849,N_4321,N_6065);
nand U9850 (N_9850,N_4182,N_4284);
or U9851 (N_9851,N_6879,N_5060);
nor U9852 (N_9852,N_7199,N_7495);
xor U9853 (N_9853,N_6813,N_7257);
xnor U9854 (N_9854,N_5230,N_5384);
or U9855 (N_9855,N_4734,N_7972);
nand U9856 (N_9856,N_5519,N_6191);
or U9857 (N_9857,N_7795,N_6054);
nand U9858 (N_9858,N_4941,N_6683);
xnor U9859 (N_9859,N_5958,N_4772);
or U9860 (N_9860,N_7980,N_4974);
nor U9861 (N_9861,N_7318,N_5277);
nand U9862 (N_9862,N_4171,N_7537);
xor U9863 (N_9863,N_6598,N_6428);
nor U9864 (N_9864,N_5239,N_5650);
nor U9865 (N_9865,N_4019,N_7295);
nor U9866 (N_9866,N_5170,N_4247);
xor U9867 (N_9867,N_5135,N_4464);
and U9868 (N_9868,N_4994,N_4183);
nor U9869 (N_9869,N_4376,N_7709);
xnor U9870 (N_9870,N_5446,N_4528);
and U9871 (N_9871,N_5380,N_6817);
nand U9872 (N_9872,N_5948,N_6838);
and U9873 (N_9873,N_5797,N_6260);
xor U9874 (N_9874,N_7418,N_4489);
and U9875 (N_9875,N_5118,N_7628);
nand U9876 (N_9876,N_4427,N_7805);
nor U9877 (N_9877,N_5134,N_6850);
and U9878 (N_9878,N_7282,N_7645);
and U9879 (N_9879,N_5460,N_7738);
and U9880 (N_9880,N_6147,N_6002);
or U9881 (N_9881,N_6019,N_7713);
or U9882 (N_9882,N_4857,N_5537);
or U9883 (N_9883,N_4578,N_7332);
or U9884 (N_9884,N_6279,N_7005);
nor U9885 (N_9885,N_4697,N_7582);
or U9886 (N_9886,N_7797,N_6198);
or U9887 (N_9887,N_6512,N_4179);
or U9888 (N_9888,N_5161,N_5659);
or U9889 (N_9889,N_5832,N_5516);
nor U9890 (N_9890,N_7830,N_7502);
xnor U9891 (N_9891,N_7975,N_7960);
nor U9892 (N_9892,N_6268,N_4153);
nor U9893 (N_9893,N_7612,N_7739);
or U9894 (N_9894,N_7244,N_4243);
nand U9895 (N_9895,N_4784,N_7232);
and U9896 (N_9896,N_5165,N_4554);
nor U9897 (N_9897,N_6338,N_6988);
nand U9898 (N_9898,N_4736,N_4932);
nand U9899 (N_9899,N_4130,N_5130);
or U9900 (N_9900,N_5617,N_5449);
and U9901 (N_9901,N_5129,N_4874);
and U9902 (N_9902,N_7246,N_7369);
or U9903 (N_9903,N_6425,N_7623);
nand U9904 (N_9904,N_7121,N_7561);
nand U9905 (N_9905,N_6001,N_7909);
and U9906 (N_9906,N_4796,N_7222);
and U9907 (N_9907,N_4230,N_4082);
and U9908 (N_9908,N_7358,N_5658);
nand U9909 (N_9909,N_6839,N_4025);
xnor U9910 (N_9910,N_6287,N_4136);
and U9911 (N_9911,N_4638,N_4460);
xor U9912 (N_9912,N_5185,N_6627);
xor U9913 (N_9913,N_6849,N_4863);
nand U9914 (N_9914,N_6882,N_6476);
nor U9915 (N_9915,N_6694,N_5854);
or U9916 (N_9916,N_4270,N_5238);
nand U9917 (N_9917,N_6290,N_7929);
or U9918 (N_9918,N_6760,N_6619);
xnor U9919 (N_9919,N_6588,N_4945);
and U9920 (N_9920,N_7264,N_4320);
nor U9921 (N_9921,N_6303,N_7728);
nand U9922 (N_9922,N_7042,N_4832);
nand U9923 (N_9923,N_4192,N_5063);
nor U9924 (N_9924,N_6135,N_6371);
nand U9925 (N_9925,N_6369,N_7107);
nand U9926 (N_9926,N_6302,N_7099);
and U9927 (N_9927,N_7944,N_7356);
nand U9928 (N_9928,N_7806,N_6766);
xnor U9929 (N_9929,N_5406,N_5272);
nor U9930 (N_9930,N_7768,N_6933);
nor U9931 (N_9931,N_6072,N_4583);
nor U9932 (N_9932,N_6574,N_4211);
xor U9933 (N_9933,N_6170,N_7751);
xnor U9934 (N_9934,N_7123,N_7670);
and U9935 (N_9935,N_6738,N_6556);
xor U9936 (N_9936,N_4163,N_4938);
nor U9937 (N_9937,N_4350,N_5104);
or U9938 (N_9938,N_5501,N_5981);
nand U9939 (N_9939,N_6152,N_4694);
nand U9940 (N_9940,N_7632,N_6577);
nor U9941 (N_9941,N_5620,N_7777);
nand U9942 (N_9942,N_6727,N_6652);
nor U9943 (N_9943,N_4120,N_7299);
or U9944 (N_9944,N_5491,N_6699);
and U9945 (N_9945,N_7201,N_6874);
or U9946 (N_9946,N_5276,N_5472);
nand U9947 (N_9947,N_7075,N_4844);
nand U9948 (N_9948,N_4169,N_5701);
nor U9949 (N_9949,N_7560,N_7447);
xor U9950 (N_9950,N_4503,N_4787);
xor U9951 (N_9951,N_4794,N_5433);
and U9952 (N_9952,N_6283,N_5896);
and U9953 (N_9953,N_7995,N_5398);
or U9954 (N_9954,N_7301,N_6456);
nor U9955 (N_9955,N_6026,N_4091);
nand U9956 (N_9956,N_7977,N_5407);
nand U9957 (N_9957,N_7169,N_4313);
nand U9958 (N_9958,N_7855,N_4509);
or U9959 (N_9959,N_5023,N_4715);
or U9960 (N_9960,N_5802,N_6298);
nor U9961 (N_9961,N_7871,N_5382);
nor U9962 (N_9962,N_4979,N_5862);
nand U9963 (N_9963,N_7306,N_4881);
or U9964 (N_9964,N_6117,N_4924);
nor U9965 (N_9965,N_5566,N_6599);
xnor U9966 (N_9966,N_6691,N_7217);
nor U9967 (N_9967,N_4330,N_6834);
or U9968 (N_9968,N_7194,N_7590);
and U9969 (N_9969,N_4175,N_4615);
nor U9970 (N_9970,N_7663,N_7514);
nor U9971 (N_9971,N_4607,N_4348);
nand U9972 (N_9972,N_5235,N_7866);
nand U9973 (N_9973,N_5775,N_7837);
or U9974 (N_9974,N_4744,N_6922);
and U9975 (N_9975,N_5097,N_7256);
or U9976 (N_9976,N_6637,N_4636);
nor U9977 (N_9977,N_7446,N_7586);
and U9978 (N_9978,N_5141,N_6114);
nor U9979 (N_9979,N_7558,N_6910);
xnor U9980 (N_9980,N_5738,N_4536);
xnor U9981 (N_9981,N_6624,N_4470);
nor U9982 (N_9982,N_7438,N_4059);
or U9983 (N_9983,N_5974,N_6232);
or U9984 (N_9984,N_6608,N_6666);
and U9985 (N_9985,N_5125,N_5086);
nand U9986 (N_9986,N_5781,N_6352);
nand U9987 (N_9987,N_7603,N_6313);
and U9988 (N_9988,N_5327,N_6672);
xor U9989 (N_9989,N_4504,N_5878);
or U9990 (N_9990,N_5835,N_4629);
and U9991 (N_9991,N_5861,N_6031);
xor U9992 (N_9992,N_6370,N_5593);
nand U9993 (N_9993,N_4228,N_4987);
xor U9994 (N_9994,N_6614,N_7772);
or U9995 (N_9995,N_7352,N_7408);
or U9996 (N_9996,N_6814,N_6464);
or U9997 (N_9997,N_4634,N_5723);
or U9998 (N_9998,N_6426,N_6463);
nor U9999 (N_9999,N_7374,N_7224);
or U10000 (N_10000,N_7996,N_7781);
nor U10001 (N_10001,N_6123,N_6861);
xnor U10002 (N_10002,N_5234,N_7742);
nor U10003 (N_10003,N_5567,N_6154);
nand U10004 (N_10004,N_7921,N_7183);
nand U10005 (N_10005,N_6560,N_5894);
xnor U10006 (N_10006,N_4295,N_6796);
and U10007 (N_10007,N_6920,N_6873);
or U10008 (N_10008,N_5054,N_5373);
nand U10009 (N_10009,N_4799,N_4359);
or U10010 (N_10010,N_5585,N_6537);
nor U10011 (N_10011,N_4468,N_6730);
and U10012 (N_10012,N_6872,N_4540);
nor U10013 (N_10013,N_4354,N_4980);
or U10014 (N_10014,N_5322,N_4636);
nand U10015 (N_10015,N_7114,N_4119);
nand U10016 (N_10016,N_4502,N_4646);
and U10017 (N_10017,N_5141,N_5010);
xor U10018 (N_10018,N_6111,N_4524);
nand U10019 (N_10019,N_4592,N_6208);
or U10020 (N_10020,N_4297,N_6097);
nor U10021 (N_10021,N_4562,N_6766);
and U10022 (N_10022,N_5686,N_6192);
and U10023 (N_10023,N_7572,N_5063);
xnor U10024 (N_10024,N_5121,N_5307);
xor U10025 (N_10025,N_7038,N_6578);
or U10026 (N_10026,N_6440,N_4206);
nand U10027 (N_10027,N_4102,N_4340);
or U10028 (N_10028,N_7960,N_7832);
or U10029 (N_10029,N_7832,N_4901);
or U10030 (N_10030,N_5150,N_6854);
xnor U10031 (N_10031,N_7465,N_6956);
nor U10032 (N_10032,N_6018,N_5621);
nand U10033 (N_10033,N_6695,N_4503);
nor U10034 (N_10034,N_5993,N_5000);
nor U10035 (N_10035,N_6764,N_7634);
nand U10036 (N_10036,N_6846,N_6651);
xor U10037 (N_10037,N_4720,N_5464);
nand U10038 (N_10038,N_7886,N_5826);
or U10039 (N_10039,N_4011,N_6528);
and U10040 (N_10040,N_7178,N_5698);
nor U10041 (N_10041,N_6861,N_4345);
or U10042 (N_10042,N_7777,N_7146);
and U10043 (N_10043,N_5655,N_4574);
nand U10044 (N_10044,N_6470,N_4258);
or U10045 (N_10045,N_7217,N_5536);
nand U10046 (N_10046,N_7368,N_5535);
xor U10047 (N_10047,N_4626,N_6955);
nor U10048 (N_10048,N_5467,N_5484);
and U10049 (N_10049,N_4693,N_4057);
or U10050 (N_10050,N_6896,N_4814);
and U10051 (N_10051,N_7439,N_7511);
nor U10052 (N_10052,N_7983,N_4282);
nor U10053 (N_10053,N_5601,N_4893);
nand U10054 (N_10054,N_7055,N_6944);
xor U10055 (N_10055,N_5715,N_4199);
nor U10056 (N_10056,N_5168,N_6354);
or U10057 (N_10057,N_5417,N_7902);
and U10058 (N_10058,N_4557,N_6080);
nor U10059 (N_10059,N_7880,N_7565);
and U10060 (N_10060,N_5867,N_7072);
xor U10061 (N_10061,N_5016,N_7107);
xnor U10062 (N_10062,N_6224,N_7856);
nand U10063 (N_10063,N_4906,N_5783);
xnor U10064 (N_10064,N_7648,N_4558);
and U10065 (N_10065,N_6142,N_4259);
xnor U10066 (N_10066,N_4208,N_6321);
nand U10067 (N_10067,N_6817,N_7235);
nor U10068 (N_10068,N_7350,N_7769);
and U10069 (N_10069,N_7377,N_5743);
nor U10070 (N_10070,N_4760,N_7338);
and U10071 (N_10071,N_5207,N_6643);
nor U10072 (N_10072,N_6704,N_6092);
nand U10073 (N_10073,N_7170,N_5497);
or U10074 (N_10074,N_6546,N_5858);
and U10075 (N_10075,N_4294,N_4303);
nand U10076 (N_10076,N_4855,N_6500);
or U10077 (N_10077,N_7576,N_5562);
and U10078 (N_10078,N_7329,N_7873);
and U10079 (N_10079,N_6420,N_4504);
and U10080 (N_10080,N_6080,N_6733);
or U10081 (N_10081,N_5316,N_6069);
or U10082 (N_10082,N_7172,N_6248);
xor U10083 (N_10083,N_5576,N_6751);
and U10084 (N_10084,N_5136,N_7419);
nand U10085 (N_10085,N_4548,N_4638);
and U10086 (N_10086,N_5161,N_4225);
xor U10087 (N_10087,N_7276,N_5446);
or U10088 (N_10088,N_5814,N_4432);
or U10089 (N_10089,N_4005,N_5753);
nand U10090 (N_10090,N_4534,N_7417);
nand U10091 (N_10091,N_6066,N_6121);
nor U10092 (N_10092,N_5384,N_5727);
nor U10093 (N_10093,N_5690,N_7640);
nand U10094 (N_10094,N_4245,N_7463);
nor U10095 (N_10095,N_7657,N_5637);
nand U10096 (N_10096,N_7402,N_6260);
nand U10097 (N_10097,N_4762,N_5391);
or U10098 (N_10098,N_5685,N_6124);
and U10099 (N_10099,N_6815,N_7991);
nand U10100 (N_10100,N_7235,N_5131);
and U10101 (N_10101,N_7361,N_6605);
or U10102 (N_10102,N_7231,N_5839);
or U10103 (N_10103,N_4346,N_4947);
nor U10104 (N_10104,N_6809,N_6905);
and U10105 (N_10105,N_7160,N_5191);
or U10106 (N_10106,N_5241,N_6463);
nand U10107 (N_10107,N_4162,N_4759);
nor U10108 (N_10108,N_6946,N_7527);
nand U10109 (N_10109,N_4046,N_4754);
nand U10110 (N_10110,N_4795,N_6552);
or U10111 (N_10111,N_7468,N_6734);
or U10112 (N_10112,N_7967,N_5813);
and U10113 (N_10113,N_4803,N_5831);
and U10114 (N_10114,N_6108,N_6878);
or U10115 (N_10115,N_5374,N_7474);
xor U10116 (N_10116,N_7877,N_5033);
nor U10117 (N_10117,N_4229,N_4567);
or U10118 (N_10118,N_5012,N_4113);
nand U10119 (N_10119,N_6077,N_5227);
nor U10120 (N_10120,N_7015,N_7847);
nand U10121 (N_10121,N_4553,N_4740);
and U10122 (N_10122,N_7733,N_5970);
nor U10123 (N_10123,N_4008,N_6804);
and U10124 (N_10124,N_5041,N_7242);
and U10125 (N_10125,N_4549,N_6872);
nor U10126 (N_10126,N_5256,N_7858);
and U10127 (N_10127,N_4661,N_6999);
and U10128 (N_10128,N_7881,N_6606);
and U10129 (N_10129,N_7369,N_5563);
or U10130 (N_10130,N_7473,N_7470);
nand U10131 (N_10131,N_6704,N_5683);
nand U10132 (N_10132,N_7366,N_7549);
or U10133 (N_10133,N_6555,N_7885);
and U10134 (N_10134,N_6050,N_5309);
and U10135 (N_10135,N_4769,N_4565);
xnor U10136 (N_10136,N_5465,N_4237);
nand U10137 (N_10137,N_6594,N_4999);
and U10138 (N_10138,N_7116,N_4460);
or U10139 (N_10139,N_6211,N_6457);
and U10140 (N_10140,N_6360,N_6164);
or U10141 (N_10141,N_5383,N_5001);
and U10142 (N_10142,N_5331,N_7763);
and U10143 (N_10143,N_7094,N_7943);
nor U10144 (N_10144,N_7588,N_4246);
nor U10145 (N_10145,N_5746,N_7417);
or U10146 (N_10146,N_4066,N_4029);
nand U10147 (N_10147,N_6946,N_7958);
nor U10148 (N_10148,N_7810,N_6125);
nand U10149 (N_10149,N_4482,N_6987);
or U10150 (N_10150,N_5001,N_5560);
nand U10151 (N_10151,N_4834,N_7170);
xor U10152 (N_10152,N_6150,N_7168);
nor U10153 (N_10153,N_7352,N_7944);
or U10154 (N_10154,N_6255,N_7248);
or U10155 (N_10155,N_5351,N_4467);
nor U10156 (N_10156,N_5909,N_6131);
or U10157 (N_10157,N_4658,N_4421);
nand U10158 (N_10158,N_6881,N_6713);
nor U10159 (N_10159,N_7065,N_6234);
and U10160 (N_10160,N_7932,N_4049);
nand U10161 (N_10161,N_6922,N_4944);
nor U10162 (N_10162,N_4358,N_6043);
nor U10163 (N_10163,N_6133,N_6708);
nand U10164 (N_10164,N_7089,N_4870);
nor U10165 (N_10165,N_4709,N_4874);
nor U10166 (N_10166,N_7274,N_4133);
and U10167 (N_10167,N_6813,N_6880);
and U10168 (N_10168,N_4792,N_5058);
xnor U10169 (N_10169,N_4020,N_5336);
and U10170 (N_10170,N_6308,N_5378);
or U10171 (N_10171,N_7627,N_7293);
nor U10172 (N_10172,N_4746,N_7061);
and U10173 (N_10173,N_4618,N_5901);
nand U10174 (N_10174,N_5563,N_4497);
nor U10175 (N_10175,N_5689,N_7710);
nand U10176 (N_10176,N_6987,N_6858);
or U10177 (N_10177,N_4876,N_4341);
nand U10178 (N_10178,N_7970,N_5933);
and U10179 (N_10179,N_4080,N_7556);
nand U10180 (N_10180,N_7000,N_4107);
nor U10181 (N_10181,N_4126,N_7730);
or U10182 (N_10182,N_5692,N_4726);
and U10183 (N_10183,N_5473,N_6880);
nor U10184 (N_10184,N_7036,N_7287);
and U10185 (N_10185,N_4926,N_7545);
nand U10186 (N_10186,N_7853,N_6480);
nor U10187 (N_10187,N_6780,N_5301);
nor U10188 (N_10188,N_6818,N_7519);
and U10189 (N_10189,N_5232,N_5518);
and U10190 (N_10190,N_7741,N_7235);
nor U10191 (N_10191,N_4269,N_7368);
or U10192 (N_10192,N_7203,N_4824);
xor U10193 (N_10193,N_5439,N_4874);
or U10194 (N_10194,N_6563,N_4912);
or U10195 (N_10195,N_5617,N_4652);
xor U10196 (N_10196,N_6166,N_5077);
nor U10197 (N_10197,N_7914,N_7948);
and U10198 (N_10198,N_5650,N_5404);
or U10199 (N_10199,N_6539,N_4667);
and U10200 (N_10200,N_5687,N_5470);
nand U10201 (N_10201,N_4996,N_5253);
or U10202 (N_10202,N_5119,N_4365);
nand U10203 (N_10203,N_5894,N_5950);
nor U10204 (N_10204,N_5871,N_6455);
or U10205 (N_10205,N_5055,N_7552);
xnor U10206 (N_10206,N_6664,N_7354);
nor U10207 (N_10207,N_7449,N_6324);
nand U10208 (N_10208,N_4391,N_5368);
and U10209 (N_10209,N_4598,N_7009);
nand U10210 (N_10210,N_4150,N_6308);
or U10211 (N_10211,N_5442,N_7657);
nor U10212 (N_10212,N_7913,N_5342);
and U10213 (N_10213,N_7366,N_5276);
xnor U10214 (N_10214,N_4784,N_7808);
or U10215 (N_10215,N_5689,N_5847);
or U10216 (N_10216,N_4349,N_6761);
nand U10217 (N_10217,N_7816,N_6184);
nor U10218 (N_10218,N_5620,N_7156);
or U10219 (N_10219,N_6892,N_7246);
nor U10220 (N_10220,N_6474,N_5795);
and U10221 (N_10221,N_5835,N_5919);
and U10222 (N_10222,N_4975,N_6619);
and U10223 (N_10223,N_4311,N_6833);
nand U10224 (N_10224,N_5690,N_5080);
nand U10225 (N_10225,N_7531,N_5385);
or U10226 (N_10226,N_7084,N_5138);
and U10227 (N_10227,N_7525,N_7540);
nor U10228 (N_10228,N_5027,N_7634);
nor U10229 (N_10229,N_7023,N_7299);
nor U10230 (N_10230,N_7120,N_7921);
nand U10231 (N_10231,N_5436,N_6557);
or U10232 (N_10232,N_6241,N_7006);
nand U10233 (N_10233,N_4687,N_4249);
and U10234 (N_10234,N_6169,N_7141);
nand U10235 (N_10235,N_5671,N_7815);
nor U10236 (N_10236,N_4834,N_4152);
and U10237 (N_10237,N_6193,N_5546);
and U10238 (N_10238,N_6490,N_7733);
nor U10239 (N_10239,N_5920,N_4668);
and U10240 (N_10240,N_5475,N_6069);
and U10241 (N_10241,N_6980,N_7062);
or U10242 (N_10242,N_4247,N_5160);
and U10243 (N_10243,N_5481,N_5609);
nor U10244 (N_10244,N_5831,N_4728);
nor U10245 (N_10245,N_7053,N_5532);
and U10246 (N_10246,N_5707,N_7638);
nand U10247 (N_10247,N_5898,N_7988);
and U10248 (N_10248,N_5196,N_4365);
nor U10249 (N_10249,N_7472,N_6451);
and U10250 (N_10250,N_7789,N_5812);
or U10251 (N_10251,N_4236,N_4078);
nand U10252 (N_10252,N_6996,N_4074);
or U10253 (N_10253,N_6622,N_7323);
or U10254 (N_10254,N_5457,N_4203);
nand U10255 (N_10255,N_4933,N_6192);
nand U10256 (N_10256,N_4177,N_4510);
or U10257 (N_10257,N_6991,N_4512);
nor U10258 (N_10258,N_6050,N_7873);
or U10259 (N_10259,N_7109,N_4137);
xor U10260 (N_10260,N_7452,N_7612);
or U10261 (N_10261,N_4921,N_4262);
nand U10262 (N_10262,N_7322,N_6744);
nand U10263 (N_10263,N_6168,N_6184);
nor U10264 (N_10264,N_7725,N_4892);
or U10265 (N_10265,N_7210,N_6894);
nor U10266 (N_10266,N_7525,N_5632);
or U10267 (N_10267,N_7950,N_5500);
and U10268 (N_10268,N_7428,N_4619);
nand U10269 (N_10269,N_5647,N_5493);
nor U10270 (N_10270,N_5167,N_5085);
or U10271 (N_10271,N_7836,N_4209);
or U10272 (N_10272,N_7406,N_6954);
nor U10273 (N_10273,N_7545,N_6900);
or U10274 (N_10274,N_4453,N_6912);
nor U10275 (N_10275,N_4585,N_7916);
and U10276 (N_10276,N_5458,N_4510);
nand U10277 (N_10277,N_7215,N_7230);
nor U10278 (N_10278,N_6996,N_5452);
nand U10279 (N_10279,N_5611,N_4560);
xor U10280 (N_10280,N_6299,N_6359);
and U10281 (N_10281,N_5800,N_6804);
or U10282 (N_10282,N_5304,N_5493);
nor U10283 (N_10283,N_7820,N_6421);
and U10284 (N_10284,N_4577,N_7861);
nor U10285 (N_10285,N_6266,N_6524);
nand U10286 (N_10286,N_6040,N_4732);
and U10287 (N_10287,N_5765,N_6850);
or U10288 (N_10288,N_5227,N_4123);
nor U10289 (N_10289,N_6159,N_6430);
and U10290 (N_10290,N_4261,N_6249);
and U10291 (N_10291,N_5514,N_6428);
nand U10292 (N_10292,N_6681,N_6850);
and U10293 (N_10293,N_4365,N_4956);
and U10294 (N_10294,N_5051,N_6772);
nor U10295 (N_10295,N_6739,N_6582);
nand U10296 (N_10296,N_6621,N_5863);
nor U10297 (N_10297,N_6806,N_7337);
and U10298 (N_10298,N_7321,N_5043);
and U10299 (N_10299,N_7099,N_5489);
and U10300 (N_10300,N_6362,N_5246);
nand U10301 (N_10301,N_6224,N_5636);
nor U10302 (N_10302,N_7622,N_5629);
nand U10303 (N_10303,N_5953,N_6577);
nand U10304 (N_10304,N_4191,N_7717);
xor U10305 (N_10305,N_7017,N_4915);
or U10306 (N_10306,N_4194,N_5757);
nand U10307 (N_10307,N_5005,N_5040);
or U10308 (N_10308,N_5162,N_5031);
or U10309 (N_10309,N_5068,N_6678);
nor U10310 (N_10310,N_4666,N_4580);
nand U10311 (N_10311,N_7740,N_4384);
and U10312 (N_10312,N_5389,N_7865);
nand U10313 (N_10313,N_6585,N_6644);
nand U10314 (N_10314,N_7392,N_7264);
and U10315 (N_10315,N_7652,N_5942);
xor U10316 (N_10316,N_6429,N_6308);
or U10317 (N_10317,N_5296,N_4241);
and U10318 (N_10318,N_6781,N_7147);
nor U10319 (N_10319,N_7665,N_5460);
nor U10320 (N_10320,N_7402,N_6980);
nor U10321 (N_10321,N_4547,N_4089);
xor U10322 (N_10322,N_6892,N_7012);
xnor U10323 (N_10323,N_6313,N_6331);
and U10324 (N_10324,N_6706,N_7413);
and U10325 (N_10325,N_5200,N_7911);
and U10326 (N_10326,N_4484,N_5734);
and U10327 (N_10327,N_5742,N_5856);
or U10328 (N_10328,N_6631,N_5116);
or U10329 (N_10329,N_4773,N_6155);
or U10330 (N_10330,N_5643,N_7518);
or U10331 (N_10331,N_5670,N_7360);
nand U10332 (N_10332,N_7968,N_5215);
nand U10333 (N_10333,N_4539,N_4641);
xor U10334 (N_10334,N_5855,N_6281);
xor U10335 (N_10335,N_5330,N_5994);
nand U10336 (N_10336,N_4779,N_6147);
nor U10337 (N_10337,N_5106,N_4730);
and U10338 (N_10338,N_4055,N_6272);
and U10339 (N_10339,N_4023,N_4397);
nand U10340 (N_10340,N_5240,N_4558);
nand U10341 (N_10341,N_7658,N_7959);
nor U10342 (N_10342,N_4032,N_6547);
and U10343 (N_10343,N_5042,N_6114);
or U10344 (N_10344,N_6339,N_4927);
or U10345 (N_10345,N_7328,N_6323);
and U10346 (N_10346,N_5218,N_4124);
or U10347 (N_10347,N_5715,N_6580);
or U10348 (N_10348,N_5190,N_4302);
nor U10349 (N_10349,N_6337,N_6664);
nor U10350 (N_10350,N_5143,N_7688);
or U10351 (N_10351,N_4783,N_6288);
xor U10352 (N_10352,N_7525,N_7809);
or U10353 (N_10353,N_5149,N_6419);
and U10354 (N_10354,N_4175,N_6474);
or U10355 (N_10355,N_7543,N_4826);
and U10356 (N_10356,N_7532,N_7401);
nor U10357 (N_10357,N_5249,N_4833);
or U10358 (N_10358,N_7609,N_5161);
nand U10359 (N_10359,N_7234,N_5883);
and U10360 (N_10360,N_5047,N_6547);
or U10361 (N_10361,N_6635,N_5186);
nand U10362 (N_10362,N_4912,N_4953);
xor U10363 (N_10363,N_7119,N_7374);
nor U10364 (N_10364,N_5494,N_5636);
or U10365 (N_10365,N_6105,N_7304);
xor U10366 (N_10366,N_4634,N_6223);
nand U10367 (N_10367,N_7053,N_7969);
and U10368 (N_10368,N_5952,N_7361);
nand U10369 (N_10369,N_6157,N_7641);
nor U10370 (N_10370,N_7011,N_4086);
and U10371 (N_10371,N_6781,N_5940);
or U10372 (N_10372,N_5409,N_7102);
nor U10373 (N_10373,N_6122,N_4107);
and U10374 (N_10374,N_5873,N_7475);
or U10375 (N_10375,N_6873,N_6459);
nor U10376 (N_10376,N_4837,N_6224);
or U10377 (N_10377,N_4197,N_6446);
xnor U10378 (N_10378,N_7252,N_6036);
nand U10379 (N_10379,N_4040,N_6065);
nand U10380 (N_10380,N_5185,N_6260);
and U10381 (N_10381,N_7406,N_7599);
nor U10382 (N_10382,N_5412,N_6784);
and U10383 (N_10383,N_4483,N_7892);
nand U10384 (N_10384,N_6041,N_6343);
xnor U10385 (N_10385,N_5742,N_7599);
and U10386 (N_10386,N_4011,N_6556);
and U10387 (N_10387,N_4639,N_5342);
nand U10388 (N_10388,N_6693,N_7692);
nand U10389 (N_10389,N_4329,N_6826);
xnor U10390 (N_10390,N_6854,N_5666);
or U10391 (N_10391,N_4136,N_5658);
nor U10392 (N_10392,N_7463,N_6177);
nor U10393 (N_10393,N_4063,N_4767);
or U10394 (N_10394,N_5205,N_7552);
nand U10395 (N_10395,N_5696,N_4481);
nor U10396 (N_10396,N_6759,N_6340);
nand U10397 (N_10397,N_5753,N_5562);
nor U10398 (N_10398,N_5328,N_4793);
nor U10399 (N_10399,N_5171,N_7068);
nand U10400 (N_10400,N_7652,N_4875);
or U10401 (N_10401,N_4120,N_4227);
nor U10402 (N_10402,N_7551,N_7115);
xnor U10403 (N_10403,N_7776,N_5534);
or U10404 (N_10404,N_7244,N_5561);
nand U10405 (N_10405,N_4289,N_6964);
and U10406 (N_10406,N_6476,N_5495);
nor U10407 (N_10407,N_4973,N_6007);
nor U10408 (N_10408,N_7439,N_6728);
and U10409 (N_10409,N_5663,N_5468);
and U10410 (N_10410,N_7582,N_7469);
or U10411 (N_10411,N_5361,N_7044);
nor U10412 (N_10412,N_7785,N_5965);
nor U10413 (N_10413,N_7162,N_4406);
and U10414 (N_10414,N_4097,N_6659);
and U10415 (N_10415,N_5267,N_7844);
and U10416 (N_10416,N_4106,N_4776);
nand U10417 (N_10417,N_5088,N_4163);
nand U10418 (N_10418,N_6809,N_6708);
nand U10419 (N_10419,N_6906,N_4186);
nor U10420 (N_10420,N_5384,N_6696);
nor U10421 (N_10421,N_6235,N_4070);
and U10422 (N_10422,N_6496,N_4070);
or U10423 (N_10423,N_4434,N_4869);
and U10424 (N_10424,N_6936,N_6642);
xnor U10425 (N_10425,N_4629,N_6688);
nor U10426 (N_10426,N_5359,N_5990);
nor U10427 (N_10427,N_6879,N_5906);
and U10428 (N_10428,N_4449,N_7660);
xnor U10429 (N_10429,N_4559,N_6507);
xnor U10430 (N_10430,N_6016,N_7216);
and U10431 (N_10431,N_5873,N_5915);
or U10432 (N_10432,N_5357,N_7197);
or U10433 (N_10433,N_4273,N_7178);
and U10434 (N_10434,N_6792,N_4952);
nand U10435 (N_10435,N_4104,N_5471);
nor U10436 (N_10436,N_5985,N_4022);
nand U10437 (N_10437,N_5418,N_5446);
or U10438 (N_10438,N_5085,N_7360);
or U10439 (N_10439,N_7864,N_4764);
and U10440 (N_10440,N_7049,N_7439);
nand U10441 (N_10441,N_6800,N_6388);
nand U10442 (N_10442,N_5166,N_5354);
nand U10443 (N_10443,N_7864,N_6540);
nand U10444 (N_10444,N_7069,N_4568);
xnor U10445 (N_10445,N_6326,N_7965);
nand U10446 (N_10446,N_6311,N_5141);
nand U10447 (N_10447,N_7643,N_7239);
xnor U10448 (N_10448,N_6894,N_7888);
and U10449 (N_10449,N_7694,N_5202);
and U10450 (N_10450,N_5078,N_6076);
and U10451 (N_10451,N_6315,N_6411);
or U10452 (N_10452,N_6706,N_4337);
nor U10453 (N_10453,N_5150,N_7530);
and U10454 (N_10454,N_4147,N_5945);
nor U10455 (N_10455,N_5580,N_7148);
nand U10456 (N_10456,N_6886,N_4342);
and U10457 (N_10457,N_6253,N_6138);
nor U10458 (N_10458,N_5382,N_5488);
nor U10459 (N_10459,N_7573,N_5248);
nand U10460 (N_10460,N_5579,N_4089);
xnor U10461 (N_10461,N_6188,N_7364);
nor U10462 (N_10462,N_4226,N_6229);
nand U10463 (N_10463,N_5150,N_4773);
and U10464 (N_10464,N_7813,N_7405);
nand U10465 (N_10465,N_6010,N_7348);
or U10466 (N_10466,N_4152,N_7362);
or U10467 (N_10467,N_4165,N_5352);
and U10468 (N_10468,N_4722,N_7764);
and U10469 (N_10469,N_5917,N_7960);
nor U10470 (N_10470,N_4066,N_6223);
and U10471 (N_10471,N_6154,N_5046);
and U10472 (N_10472,N_4986,N_5925);
nor U10473 (N_10473,N_6365,N_4917);
nand U10474 (N_10474,N_5925,N_5800);
or U10475 (N_10475,N_6558,N_7599);
xnor U10476 (N_10476,N_4588,N_6960);
and U10477 (N_10477,N_7799,N_4639);
or U10478 (N_10478,N_7156,N_4962);
or U10479 (N_10479,N_7145,N_7626);
and U10480 (N_10480,N_5557,N_4069);
or U10481 (N_10481,N_5275,N_7610);
nor U10482 (N_10482,N_6853,N_7443);
or U10483 (N_10483,N_6211,N_6648);
nor U10484 (N_10484,N_5814,N_4647);
nand U10485 (N_10485,N_7341,N_4234);
or U10486 (N_10486,N_7202,N_7218);
nor U10487 (N_10487,N_7669,N_7682);
and U10488 (N_10488,N_4559,N_4632);
nand U10489 (N_10489,N_6650,N_4080);
and U10490 (N_10490,N_5084,N_4475);
nor U10491 (N_10491,N_5537,N_4507);
or U10492 (N_10492,N_4443,N_4457);
nor U10493 (N_10493,N_6889,N_4379);
or U10494 (N_10494,N_4261,N_4778);
nand U10495 (N_10495,N_5227,N_7362);
or U10496 (N_10496,N_7205,N_6313);
or U10497 (N_10497,N_6943,N_6683);
nand U10498 (N_10498,N_4760,N_4146);
or U10499 (N_10499,N_5472,N_5572);
nor U10500 (N_10500,N_4030,N_7031);
or U10501 (N_10501,N_4228,N_7430);
nand U10502 (N_10502,N_6708,N_6528);
xor U10503 (N_10503,N_4756,N_6814);
nand U10504 (N_10504,N_5987,N_6669);
xor U10505 (N_10505,N_6958,N_4795);
nor U10506 (N_10506,N_6251,N_4956);
or U10507 (N_10507,N_7424,N_6998);
nor U10508 (N_10508,N_4974,N_5229);
and U10509 (N_10509,N_4464,N_4696);
and U10510 (N_10510,N_4971,N_7348);
xnor U10511 (N_10511,N_4559,N_7098);
nor U10512 (N_10512,N_7229,N_6464);
and U10513 (N_10513,N_6107,N_6292);
nor U10514 (N_10514,N_4622,N_4071);
or U10515 (N_10515,N_7024,N_5880);
nor U10516 (N_10516,N_5425,N_5822);
and U10517 (N_10517,N_7822,N_5254);
or U10518 (N_10518,N_6864,N_4157);
nand U10519 (N_10519,N_4925,N_7825);
nor U10520 (N_10520,N_6976,N_7452);
nand U10521 (N_10521,N_4843,N_7401);
nor U10522 (N_10522,N_7322,N_4769);
nand U10523 (N_10523,N_7214,N_5827);
or U10524 (N_10524,N_6789,N_5526);
or U10525 (N_10525,N_6544,N_6522);
and U10526 (N_10526,N_4997,N_7006);
and U10527 (N_10527,N_6558,N_7778);
or U10528 (N_10528,N_6753,N_5595);
nand U10529 (N_10529,N_5951,N_4890);
nand U10530 (N_10530,N_6861,N_7745);
xnor U10531 (N_10531,N_4665,N_7385);
nor U10532 (N_10532,N_4013,N_4008);
or U10533 (N_10533,N_6178,N_6958);
or U10534 (N_10534,N_5138,N_7031);
nand U10535 (N_10535,N_4721,N_4740);
nand U10536 (N_10536,N_4163,N_6519);
xnor U10537 (N_10537,N_5564,N_4537);
nor U10538 (N_10538,N_4061,N_5499);
or U10539 (N_10539,N_4632,N_7253);
or U10540 (N_10540,N_5237,N_4922);
nand U10541 (N_10541,N_4215,N_5977);
nand U10542 (N_10542,N_6175,N_7923);
xnor U10543 (N_10543,N_5271,N_5873);
nor U10544 (N_10544,N_7587,N_4441);
or U10545 (N_10545,N_5324,N_6720);
xnor U10546 (N_10546,N_5135,N_6546);
nand U10547 (N_10547,N_5949,N_4165);
xor U10548 (N_10548,N_5871,N_4282);
nand U10549 (N_10549,N_4144,N_4909);
nand U10550 (N_10550,N_5749,N_5683);
or U10551 (N_10551,N_6218,N_5716);
or U10552 (N_10552,N_5150,N_7547);
and U10553 (N_10553,N_4021,N_7432);
nand U10554 (N_10554,N_5216,N_7102);
nand U10555 (N_10555,N_5849,N_7571);
nand U10556 (N_10556,N_7469,N_6190);
nand U10557 (N_10557,N_6527,N_7328);
nor U10558 (N_10558,N_7918,N_6939);
nand U10559 (N_10559,N_6591,N_7001);
nor U10560 (N_10560,N_7641,N_7053);
nand U10561 (N_10561,N_4706,N_6596);
nor U10562 (N_10562,N_5602,N_6845);
nand U10563 (N_10563,N_7935,N_4981);
nor U10564 (N_10564,N_7212,N_4213);
or U10565 (N_10565,N_4774,N_4304);
nor U10566 (N_10566,N_7058,N_6229);
nand U10567 (N_10567,N_5703,N_4838);
nand U10568 (N_10568,N_6219,N_5358);
or U10569 (N_10569,N_6566,N_7396);
nor U10570 (N_10570,N_5366,N_7003);
or U10571 (N_10571,N_7518,N_4467);
nand U10572 (N_10572,N_5350,N_7148);
or U10573 (N_10573,N_7751,N_6282);
or U10574 (N_10574,N_4675,N_7282);
or U10575 (N_10575,N_7144,N_5374);
or U10576 (N_10576,N_7854,N_4451);
nor U10577 (N_10577,N_4889,N_6502);
or U10578 (N_10578,N_7843,N_7668);
or U10579 (N_10579,N_4506,N_7336);
and U10580 (N_10580,N_7574,N_4782);
or U10581 (N_10581,N_5680,N_5918);
nor U10582 (N_10582,N_4756,N_5847);
and U10583 (N_10583,N_5491,N_6957);
xor U10584 (N_10584,N_4658,N_4473);
and U10585 (N_10585,N_5814,N_6045);
nor U10586 (N_10586,N_4995,N_6323);
nand U10587 (N_10587,N_4945,N_4059);
nand U10588 (N_10588,N_6822,N_6927);
nor U10589 (N_10589,N_4635,N_5587);
xnor U10590 (N_10590,N_6189,N_7528);
nor U10591 (N_10591,N_7316,N_7583);
xnor U10592 (N_10592,N_5946,N_5024);
and U10593 (N_10593,N_4654,N_6380);
nor U10594 (N_10594,N_5359,N_5781);
and U10595 (N_10595,N_4181,N_6200);
xnor U10596 (N_10596,N_7987,N_4039);
or U10597 (N_10597,N_7684,N_7425);
nor U10598 (N_10598,N_5597,N_5140);
nor U10599 (N_10599,N_7579,N_5020);
nand U10600 (N_10600,N_6403,N_5979);
and U10601 (N_10601,N_4946,N_4771);
or U10602 (N_10602,N_4460,N_4466);
or U10603 (N_10603,N_4022,N_6060);
nand U10604 (N_10604,N_5592,N_6787);
and U10605 (N_10605,N_5408,N_6734);
nor U10606 (N_10606,N_7675,N_5100);
nor U10607 (N_10607,N_5417,N_4146);
or U10608 (N_10608,N_5526,N_4915);
and U10609 (N_10609,N_7983,N_7935);
and U10610 (N_10610,N_6664,N_7239);
xnor U10611 (N_10611,N_6610,N_4548);
nor U10612 (N_10612,N_6396,N_5519);
and U10613 (N_10613,N_4139,N_5093);
or U10614 (N_10614,N_4952,N_6435);
or U10615 (N_10615,N_7795,N_4545);
or U10616 (N_10616,N_6669,N_4743);
nor U10617 (N_10617,N_5560,N_5391);
nor U10618 (N_10618,N_5650,N_7437);
or U10619 (N_10619,N_6844,N_4177);
or U10620 (N_10620,N_7287,N_5031);
and U10621 (N_10621,N_6047,N_4358);
nor U10622 (N_10622,N_4079,N_6487);
or U10623 (N_10623,N_6537,N_6391);
xor U10624 (N_10624,N_4200,N_4535);
and U10625 (N_10625,N_4341,N_4021);
and U10626 (N_10626,N_7632,N_6166);
nand U10627 (N_10627,N_4609,N_4219);
and U10628 (N_10628,N_4236,N_7831);
or U10629 (N_10629,N_5751,N_7180);
nand U10630 (N_10630,N_4292,N_7611);
and U10631 (N_10631,N_4031,N_6681);
or U10632 (N_10632,N_7764,N_5892);
nor U10633 (N_10633,N_7912,N_7894);
nand U10634 (N_10634,N_5273,N_6784);
nand U10635 (N_10635,N_6188,N_6412);
nand U10636 (N_10636,N_7531,N_4705);
or U10637 (N_10637,N_4570,N_5363);
or U10638 (N_10638,N_4585,N_6867);
nor U10639 (N_10639,N_5375,N_6258);
nand U10640 (N_10640,N_5697,N_5263);
xor U10641 (N_10641,N_4458,N_7132);
nand U10642 (N_10642,N_5418,N_7654);
xnor U10643 (N_10643,N_7109,N_4371);
and U10644 (N_10644,N_7016,N_5207);
or U10645 (N_10645,N_5084,N_5526);
or U10646 (N_10646,N_6613,N_5498);
or U10647 (N_10647,N_5795,N_6936);
xnor U10648 (N_10648,N_7173,N_7864);
nand U10649 (N_10649,N_6304,N_5291);
xor U10650 (N_10650,N_4243,N_5200);
nand U10651 (N_10651,N_6426,N_6686);
or U10652 (N_10652,N_6368,N_4182);
nand U10653 (N_10653,N_4080,N_6623);
nor U10654 (N_10654,N_6175,N_4561);
nand U10655 (N_10655,N_7937,N_4892);
nand U10656 (N_10656,N_6682,N_4861);
nand U10657 (N_10657,N_5128,N_4236);
nand U10658 (N_10658,N_4850,N_5255);
and U10659 (N_10659,N_4649,N_4900);
and U10660 (N_10660,N_6844,N_6434);
nand U10661 (N_10661,N_5701,N_7956);
nor U10662 (N_10662,N_6670,N_6248);
nor U10663 (N_10663,N_6450,N_4279);
and U10664 (N_10664,N_7204,N_6489);
and U10665 (N_10665,N_4792,N_7711);
or U10666 (N_10666,N_5723,N_5722);
nor U10667 (N_10667,N_4451,N_6713);
xnor U10668 (N_10668,N_6732,N_7750);
and U10669 (N_10669,N_7719,N_6787);
nand U10670 (N_10670,N_4091,N_7828);
xnor U10671 (N_10671,N_4042,N_7943);
nor U10672 (N_10672,N_4454,N_4604);
nor U10673 (N_10673,N_6044,N_6567);
and U10674 (N_10674,N_4721,N_5718);
and U10675 (N_10675,N_6906,N_6110);
and U10676 (N_10676,N_7511,N_6425);
nand U10677 (N_10677,N_4922,N_4348);
xnor U10678 (N_10678,N_5609,N_7532);
and U10679 (N_10679,N_5900,N_5970);
and U10680 (N_10680,N_5216,N_7257);
nor U10681 (N_10681,N_7133,N_6802);
nor U10682 (N_10682,N_7792,N_4590);
or U10683 (N_10683,N_4394,N_7366);
and U10684 (N_10684,N_5496,N_4720);
xor U10685 (N_10685,N_7691,N_7810);
nand U10686 (N_10686,N_5684,N_5667);
xor U10687 (N_10687,N_4934,N_7835);
or U10688 (N_10688,N_4751,N_5179);
nand U10689 (N_10689,N_6957,N_4335);
nor U10690 (N_10690,N_5833,N_6920);
nor U10691 (N_10691,N_4134,N_5599);
nor U10692 (N_10692,N_5234,N_6883);
or U10693 (N_10693,N_4833,N_7979);
or U10694 (N_10694,N_7857,N_5613);
nor U10695 (N_10695,N_5217,N_4490);
nand U10696 (N_10696,N_4593,N_4156);
nand U10697 (N_10697,N_5149,N_5288);
and U10698 (N_10698,N_4482,N_6630);
nand U10699 (N_10699,N_5389,N_4178);
and U10700 (N_10700,N_7469,N_7772);
xor U10701 (N_10701,N_4915,N_5875);
nand U10702 (N_10702,N_5805,N_5697);
nor U10703 (N_10703,N_7752,N_5571);
or U10704 (N_10704,N_6025,N_6667);
and U10705 (N_10705,N_5564,N_4889);
nor U10706 (N_10706,N_4159,N_6165);
xor U10707 (N_10707,N_7509,N_7470);
and U10708 (N_10708,N_7524,N_5577);
xnor U10709 (N_10709,N_6602,N_4789);
nand U10710 (N_10710,N_6324,N_6178);
or U10711 (N_10711,N_7577,N_4250);
nor U10712 (N_10712,N_7764,N_6815);
or U10713 (N_10713,N_5991,N_6875);
or U10714 (N_10714,N_4201,N_5055);
nor U10715 (N_10715,N_5670,N_7304);
nor U10716 (N_10716,N_5288,N_5699);
nand U10717 (N_10717,N_7754,N_5395);
nor U10718 (N_10718,N_7710,N_4235);
or U10719 (N_10719,N_6149,N_6057);
xor U10720 (N_10720,N_4287,N_6162);
nor U10721 (N_10721,N_7512,N_7011);
nand U10722 (N_10722,N_5460,N_6667);
nand U10723 (N_10723,N_5875,N_5226);
nor U10724 (N_10724,N_5114,N_6257);
nor U10725 (N_10725,N_6041,N_4188);
xor U10726 (N_10726,N_6077,N_6120);
nand U10727 (N_10727,N_6505,N_4710);
and U10728 (N_10728,N_7046,N_4704);
nand U10729 (N_10729,N_5944,N_4673);
nor U10730 (N_10730,N_5907,N_5377);
xnor U10731 (N_10731,N_7878,N_4451);
or U10732 (N_10732,N_6595,N_4867);
and U10733 (N_10733,N_4300,N_6164);
nor U10734 (N_10734,N_4152,N_4541);
nand U10735 (N_10735,N_4328,N_7334);
xnor U10736 (N_10736,N_5419,N_4940);
and U10737 (N_10737,N_6322,N_6045);
and U10738 (N_10738,N_7361,N_4472);
or U10739 (N_10739,N_7721,N_7492);
nand U10740 (N_10740,N_7502,N_7874);
nand U10741 (N_10741,N_6899,N_4328);
nor U10742 (N_10742,N_6784,N_6772);
xor U10743 (N_10743,N_6194,N_6802);
and U10744 (N_10744,N_7707,N_4421);
or U10745 (N_10745,N_5073,N_5024);
nand U10746 (N_10746,N_4991,N_5107);
nor U10747 (N_10747,N_6232,N_7022);
nor U10748 (N_10748,N_4151,N_7709);
nand U10749 (N_10749,N_7404,N_5594);
and U10750 (N_10750,N_5705,N_4348);
nor U10751 (N_10751,N_5907,N_7792);
and U10752 (N_10752,N_6143,N_6558);
nor U10753 (N_10753,N_4398,N_5968);
nand U10754 (N_10754,N_7205,N_6028);
nand U10755 (N_10755,N_7440,N_5943);
or U10756 (N_10756,N_5442,N_5735);
and U10757 (N_10757,N_7977,N_5766);
and U10758 (N_10758,N_5285,N_4746);
and U10759 (N_10759,N_4212,N_5688);
xor U10760 (N_10760,N_7598,N_4337);
or U10761 (N_10761,N_6195,N_5830);
xnor U10762 (N_10762,N_6738,N_4585);
or U10763 (N_10763,N_5470,N_6957);
and U10764 (N_10764,N_6137,N_5337);
and U10765 (N_10765,N_4073,N_4080);
nand U10766 (N_10766,N_4502,N_6183);
and U10767 (N_10767,N_6712,N_5223);
xor U10768 (N_10768,N_4097,N_7673);
and U10769 (N_10769,N_6435,N_6544);
and U10770 (N_10770,N_4010,N_5420);
nand U10771 (N_10771,N_7860,N_4549);
and U10772 (N_10772,N_7227,N_7731);
nand U10773 (N_10773,N_4800,N_4135);
nand U10774 (N_10774,N_7124,N_5805);
nand U10775 (N_10775,N_5635,N_5179);
nand U10776 (N_10776,N_4519,N_6371);
nand U10777 (N_10777,N_7063,N_4643);
xor U10778 (N_10778,N_5467,N_6503);
nand U10779 (N_10779,N_6268,N_6515);
nand U10780 (N_10780,N_6845,N_4448);
nand U10781 (N_10781,N_7876,N_5337);
and U10782 (N_10782,N_4409,N_7073);
and U10783 (N_10783,N_5740,N_6070);
nand U10784 (N_10784,N_7746,N_7292);
nand U10785 (N_10785,N_7099,N_7989);
or U10786 (N_10786,N_4591,N_6188);
or U10787 (N_10787,N_6322,N_4363);
nand U10788 (N_10788,N_7616,N_6236);
nand U10789 (N_10789,N_6705,N_4449);
nor U10790 (N_10790,N_6410,N_5583);
and U10791 (N_10791,N_4913,N_4786);
or U10792 (N_10792,N_6419,N_6633);
nand U10793 (N_10793,N_4610,N_7400);
nor U10794 (N_10794,N_6694,N_7994);
nand U10795 (N_10795,N_7951,N_5153);
nor U10796 (N_10796,N_6986,N_5472);
xnor U10797 (N_10797,N_5379,N_5079);
or U10798 (N_10798,N_4840,N_4410);
and U10799 (N_10799,N_6114,N_5692);
and U10800 (N_10800,N_5062,N_7630);
or U10801 (N_10801,N_6776,N_6471);
nand U10802 (N_10802,N_6958,N_6313);
nand U10803 (N_10803,N_6482,N_7079);
or U10804 (N_10804,N_7786,N_7014);
and U10805 (N_10805,N_6469,N_6932);
and U10806 (N_10806,N_4505,N_4232);
and U10807 (N_10807,N_5591,N_6322);
nand U10808 (N_10808,N_7973,N_6349);
and U10809 (N_10809,N_4677,N_5025);
nand U10810 (N_10810,N_5381,N_7712);
nand U10811 (N_10811,N_5929,N_5507);
and U10812 (N_10812,N_6518,N_4570);
nand U10813 (N_10813,N_6149,N_6616);
nand U10814 (N_10814,N_7856,N_7151);
nor U10815 (N_10815,N_4334,N_7551);
nand U10816 (N_10816,N_5307,N_4305);
and U10817 (N_10817,N_6886,N_6210);
xnor U10818 (N_10818,N_5526,N_4200);
or U10819 (N_10819,N_5928,N_5513);
nor U10820 (N_10820,N_6373,N_7787);
or U10821 (N_10821,N_5031,N_4118);
nor U10822 (N_10822,N_4343,N_5892);
and U10823 (N_10823,N_4602,N_5147);
and U10824 (N_10824,N_4377,N_4066);
nor U10825 (N_10825,N_5660,N_6512);
or U10826 (N_10826,N_4435,N_7696);
or U10827 (N_10827,N_7049,N_5555);
and U10828 (N_10828,N_4753,N_4578);
xor U10829 (N_10829,N_6473,N_5906);
or U10830 (N_10830,N_4636,N_5034);
nand U10831 (N_10831,N_7709,N_7748);
or U10832 (N_10832,N_4470,N_4607);
and U10833 (N_10833,N_7088,N_6307);
nor U10834 (N_10834,N_7848,N_7519);
nor U10835 (N_10835,N_7523,N_4833);
nor U10836 (N_10836,N_4837,N_4727);
or U10837 (N_10837,N_4101,N_7373);
nor U10838 (N_10838,N_7329,N_5030);
and U10839 (N_10839,N_4197,N_5057);
and U10840 (N_10840,N_5476,N_7068);
nor U10841 (N_10841,N_4622,N_4865);
nor U10842 (N_10842,N_6162,N_6428);
xor U10843 (N_10843,N_7374,N_6131);
xor U10844 (N_10844,N_7887,N_5826);
or U10845 (N_10845,N_7438,N_6263);
xnor U10846 (N_10846,N_6468,N_5724);
nand U10847 (N_10847,N_6225,N_5378);
nor U10848 (N_10848,N_6431,N_6065);
and U10849 (N_10849,N_6431,N_5915);
nand U10850 (N_10850,N_6580,N_7963);
nor U10851 (N_10851,N_4951,N_4424);
nand U10852 (N_10852,N_6580,N_7362);
nor U10853 (N_10853,N_5180,N_6336);
and U10854 (N_10854,N_4756,N_7012);
or U10855 (N_10855,N_5065,N_5340);
or U10856 (N_10856,N_6056,N_6768);
nand U10857 (N_10857,N_6550,N_6817);
xor U10858 (N_10858,N_5998,N_7074);
or U10859 (N_10859,N_7371,N_6652);
nand U10860 (N_10860,N_5044,N_7138);
nand U10861 (N_10861,N_7328,N_4074);
and U10862 (N_10862,N_5072,N_7798);
and U10863 (N_10863,N_4015,N_7508);
or U10864 (N_10864,N_7896,N_7618);
and U10865 (N_10865,N_7110,N_6155);
nor U10866 (N_10866,N_7875,N_7107);
or U10867 (N_10867,N_4664,N_6534);
or U10868 (N_10868,N_5505,N_7557);
nand U10869 (N_10869,N_6259,N_7125);
nor U10870 (N_10870,N_4861,N_6194);
and U10871 (N_10871,N_4960,N_4685);
nor U10872 (N_10872,N_5835,N_6759);
and U10873 (N_10873,N_5167,N_4248);
nor U10874 (N_10874,N_4237,N_7196);
and U10875 (N_10875,N_7842,N_4484);
nand U10876 (N_10876,N_4675,N_6827);
and U10877 (N_10877,N_6471,N_7161);
nand U10878 (N_10878,N_4209,N_4504);
or U10879 (N_10879,N_5863,N_6896);
and U10880 (N_10880,N_4053,N_5984);
nand U10881 (N_10881,N_4798,N_5528);
nand U10882 (N_10882,N_6958,N_7194);
nor U10883 (N_10883,N_5866,N_4233);
and U10884 (N_10884,N_4430,N_5698);
nor U10885 (N_10885,N_4316,N_5104);
nand U10886 (N_10886,N_5856,N_7918);
nand U10887 (N_10887,N_6739,N_5729);
and U10888 (N_10888,N_7893,N_7351);
nor U10889 (N_10889,N_5707,N_4252);
and U10890 (N_10890,N_5904,N_6882);
nand U10891 (N_10891,N_7357,N_7609);
nor U10892 (N_10892,N_5834,N_4357);
nand U10893 (N_10893,N_5061,N_4877);
nor U10894 (N_10894,N_7278,N_7971);
xnor U10895 (N_10895,N_4929,N_7953);
nor U10896 (N_10896,N_7971,N_5118);
xnor U10897 (N_10897,N_7617,N_4322);
and U10898 (N_10898,N_7389,N_4182);
nor U10899 (N_10899,N_7723,N_5328);
and U10900 (N_10900,N_5881,N_5357);
or U10901 (N_10901,N_5470,N_5624);
and U10902 (N_10902,N_7055,N_4087);
nand U10903 (N_10903,N_6134,N_6683);
or U10904 (N_10904,N_7274,N_7608);
or U10905 (N_10905,N_5055,N_7613);
and U10906 (N_10906,N_4876,N_6713);
or U10907 (N_10907,N_4676,N_4607);
or U10908 (N_10908,N_6129,N_4253);
nand U10909 (N_10909,N_4690,N_7048);
or U10910 (N_10910,N_4316,N_7269);
nor U10911 (N_10911,N_7747,N_6734);
and U10912 (N_10912,N_5948,N_6511);
xor U10913 (N_10913,N_4347,N_4853);
xnor U10914 (N_10914,N_4068,N_7930);
or U10915 (N_10915,N_5139,N_7810);
nand U10916 (N_10916,N_6648,N_4145);
or U10917 (N_10917,N_6598,N_4204);
and U10918 (N_10918,N_5383,N_7720);
or U10919 (N_10919,N_7385,N_7442);
nand U10920 (N_10920,N_6746,N_6612);
nor U10921 (N_10921,N_5350,N_5200);
nor U10922 (N_10922,N_7198,N_5860);
xor U10923 (N_10923,N_7589,N_5003);
nor U10924 (N_10924,N_7461,N_7121);
nand U10925 (N_10925,N_6948,N_7772);
or U10926 (N_10926,N_5562,N_6225);
xor U10927 (N_10927,N_6716,N_6356);
nand U10928 (N_10928,N_7478,N_6800);
or U10929 (N_10929,N_7169,N_6174);
xor U10930 (N_10930,N_7044,N_4092);
or U10931 (N_10931,N_5106,N_7223);
or U10932 (N_10932,N_4019,N_7477);
nand U10933 (N_10933,N_4351,N_4779);
nor U10934 (N_10934,N_5000,N_4790);
and U10935 (N_10935,N_6629,N_5114);
and U10936 (N_10936,N_7488,N_7720);
nand U10937 (N_10937,N_7256,N_6492);
nor U10938 (N_10938,N_5740,N_5261);
nor U10939 (N_10939,N_4865,N_7578);
and U10940 (N_10940,N_5314,N_7620);
and U10941 (N_10941,N_4161,N_4585);
nand U10942 (N_10942,N_6087,N_6486);
nand U10943 (N_10943,N_5555,N_4073);
xnor U10944 (N_10944,N_5002,N_6224);
nand U10945 (N_10945,N_7663,N_6258);
nand U10946 (N_10946,N_5022,N_4849);
nand U10947 (N_10947,N_5033,N_5379);
or U10948 (N_10948,N_5016,N_4583);
or U10949 (N_10949,N_7170,N_5018);
nand U10950 (N_10950,N_7267,N_4725);
and U10951 (N_10951,N_7846,N_4840);
or U10952 (N_10952,N_7178,N_7690);
nor U10953 (N_10953,N_4736,N_5208);
or U10954 (N_10954,N_4810,N_5118);
xor U10955 (N_10955,N_4543,N_4971);
and U10956 (N_10956,N_5352,N_4501);
xor U10957 (N_10957,N_4132,N_5493);
or U10958 (N_10958,N_4929,N_4821);
and U10959 (N_10959,N_6842,N_4082);
xnor U10960 (N_10960,N_7436,N_4459);
nor U10961 (N_10961,N_4240,N_4219);
nand U10962 (N_10962,N_6653,N_7319);
nor U10963 (N_10963,N_7168,N_7894);
or U10964 (N_10964,N_4690,N_7705);
and U10965 (N_10965,N_6723,N_4535);
and U10966 (N_10966,N_7488,N_6686);
and U10967 (N_10967,N_4404,N_4542);
or U10968 (N_10968,N_7635,N_4625);
xnor U10969 (N_10969,N_5349,N_4087);
nor U10970 (N_10970,N_4376,N_4785);
nand U10971 (N_10971,N_6102,N_5623);
and U10972 (N_10972,N_4860,N_5077);
xor U10973 (N_10973,N_6082,N_7226);
or U10974 (N_10974,N_7017,N_7679);
nor U10975 (N_10975,N_5121,N_5421);
and U10976 (N_10976,N_7851,N_4767);
and U10977 (N_10977,N_4628,N_4859);
and U10978 (N_10978,N_5859,N_7288);
and U10979 (N_10979,N_5885,N_5592);
or U10980 (N_10980,N_7418,N_5653);
and U10981 (N_10981,N_5603,N_5953);
nor U10982 (N_10982,N_7032,N_4325);
nand U10983 (N_10983,N_7710,N_7435);
nor U10984 (N_10984,N_4370,N_6539);
xnor U10985 (N_10985,N_5904,N_4264);
nor U10986 (N_10986,N_6966,N_7469);
nor U10987 (N_10987,N_6225,N_6420);
and U10988 (N_10988,N_4881,N_5993);
xor U10989 (N_10989,N_4335,N_4798);
nor U10990 (N_10990,N_7413,N_6806);
and U10991 (N_10991,N_4498,N_6067);
and U10992 (N_10992,N_5156,N_6489);
and U10993 (N_10993,N_5333,N_7289);
nand U10994 (N_10994,N_6415,N_4930);
and U10995 (N_10995,N_7319,N_4777);
and U10996 (N_10996,N_4458,N_4545);
nor U10997 (N_10997,N_4447,N_4222);
nor U10998 (N_10998,N_7143,N_5351);
nand U10999 (N_10999,N_4001,N_6750);
xnor U11000 (N_11000,N_4955,N_4226);
nand U11001 (N_11001,N_6903,N_4541);
or U11002 (N_11002,N_5052,N_4333);
nor U11003 (N_11003,N_7842,N_6007);
nor U11004 (N_11004,N_4191,N_5647);
and U11005 (N_11005,N_4394,N_7432);
nand U11006 (N_11006,N_7306,N_7384);
or U11007 (N_11007,N_7825,N_4887);
or U11008 (N_11008,N_6096,N_5846);
and U11009 (N_11009,N_4695,N_7402);
xnor U11010 (N_11010,N_5140,N_4090);
nor U11011 (N_11011,N_7699,N_6748);
nor U11012 (N_11012,N_7911,N_6344);
xnor U11013 (N_11013,N_5829,N_6692);
and U11014 (N_11014,N_5015,N_6029);
or U11015 (N_11015,N_6475,N_4904);
or U11016 (N_11016,N_6233,N_6498);
nand U11017 (N_11017,N_6569,N_6209);
nor U11018 (N_11018,N_5477,N_7733);
and U11019 (N_11019,N_4662,N_6726);
nand U11020 (N_11020,N_5980,N_6222);
and U11021 (N_11021,N_4288,N_4217);
xnor U11022 (N_11022,N_7817,N_6551);
or U11023 (N_11023,N_6869,N_6711);
and U11024 (N_11024,N_6030,N_7574);
nor U11025 (N_11025,N_7741,N_4489);
nand U11026 (N_11026,N_5129,N_5045);
nand U11027 (N_11027,N_7355,N_4609);
and U11028 (N_11028,N_7228,N_5834);
nand U11029 (N_11029,N_6365,N_5429);
nand U11030 (N_11030,N_5394,N_7315);
and U11031 (N_11031,N_5596,N_7790);
nor U11032 (N_11032,N_4589,N_4435);
nand U11033 (N_11033,N_7061,N_5905);
nand U11034 (N_11034,N_7073,N_7935);
and U11035 (N_11035,N_5435,N_4915);
nor U11036 (N_11036,N_6660,N_6943);
and U11037 (N_11037,N_6351,N_4066);
nand U11038 (N_11038,N_7760,N_6828);
or U11039 (N_11039,N_7808,N_7681);
and U11040 (N_11040,N_7722,N_6304);
and U11041 (N_11041,N_6056,N_7966);
or U11042 (N_11042,N_5178,N_6507);
or U11043 (N_11043,N_5620,N_6985);
nor U11044 (N_11044,N_5608,N_5057);
or U11045 (N_11045,N_5965,N_4999);
and U11046 (N_11046,N_7054,N_5509);
nor U11047 (N_11047,N_7198,N_7876);
nor U11048 (N_11048,N_6521,N_4413);
nor U11049 (N_11049,N_7606,N_5849);
nand U11050 (N_11050,N_7820,N_6672);
nand U11051 (N_11051,N_6268,N_5815);
or U11052 (N_11052,N_4345,N_5587);
nor U11053 (N_11053,N_6993,N_5924);
nand U11054 (N_11054,N_4882,N_7371);
nand U11055 (N_11055,N_5698,N_5547);
and U11056 (N_11056,N_4281,N_7118);
nor U11057 (N_11057,N_4158,N_5546);
or U11058 (N_11058,N_6076,N_5137);
and U11059 (N_11059,N_4025,N_6296);
and U11060 (N_11060,N_4097,N_4361);
and U11061 (N_11061,N_7367,N_7373);
nand U11062 (N_11062,N_5292,N_4818);
nor U11063 (N_11063,N_4813,N_5414);
or U11064 (N_11064,N_7737,N_4462);
or U11065 (N_11065,N_7410,N_7699);
nand U11066 (N_11066,N_4815,N_6812);
nand U11067 (N_11067,N_7727,N_5890);
and U11068 (N_11068,N_5435,N_5006);
nor U11069 (N_11069,N_6771,N_7566);
nor U11070 (N_11070,N_5078,N_7617);
and U11071 (N_11071,N_5601,N_4868);
nor U11072 (N_11072,N_7571,N_5390);
xnor U11073 (N_11073,N_6689,N_6272);
and U11074 (N_11074,N_6254,N_6354);
and U11075 (N_11075,N_6041,N_5372);
nand U11076 (N_11076,N_6069,N_5341);
or U11077 (N_11077,N_7619,N_4326);
xnor U11078 (N_11078,N_5904,N_6045);
nand U11079 (N_11079,N_7464,N_5826);
nand U11080 (N_11080,N_7040,N_7263);
nor U11081 (N_11081,N_6623,N_6994);
and U11082 (N_11082,N_4477,N_5326);
nand U11083 (N_11083,N_7041,N_6611);
or U11084 (N_11084,N_4437,N_5893);
or U11085 (N_11085,N_7055,N_4850);
nand U11086 (N_11086,N_7858,N_6733);
or U11087 (N_11087,N_6419,N_6399);
or U11088 (N_11088,N_6017,N_5796);
nor U11089 (N_11089,N_4479,N_4146);
and U11090 (N_11090,N_4379,N_5270);
or U11091 (N_11091,N_6545,N_5162);
nor U11092 (N_11092,N_4232,N_6730);
and U11093 (N_11093,N_6495,N_4729);
nor U11094 (N_11094,N_7194,N_7699);
nand U11095 (N_11095,N_4941,N_4643);
or U11096 (N_11096,N_4284,N_4972);
and U11097 (N_11097,N_6955,N_5518);
or U11098 (N_11098,N_5686,N_4348);
and U11099 (N_11099,N_7981,N_6320);
nand U11100 (N_11100,N_4863,N_4862);
and U11101 (N_11101,N_4709,N_5689);
nand U11102 (N_11102,N_4303,N_7708);
nor U11103 (N_11103,N_4058,N_4936);
or U11104 (N_11104,N_4189,N_7427);
and U11105 (N_11105,N_5918,N_5619);
or U11106 (N_11106,N_7505,N_4523);
nor U11107 (N_11107,N_6384,N_6707);
nand U11108 (N_11108,N_5689,N_6579);
and U11109 (N_11109,N_7919,N_6331);
nand U11110 (N_11110,N_6511,N_6314);
nand U11111 (N_11111,N_4127,N_6325);
and U11112 (N_11112,N_5890,N_5448);
nand U11113 (N_11113,N_6367,N_7355);
nand U11114 (N_11114,N_4366,N_4180);
xor U11115 (N_11115,N_6299,N_7983);
nor U11116 (N_11116,N_7668,N_4585);
or U11117 (N_11117,N_7650,N_7950);
or U11118 (N_11118,N_4255,N_7083);
or U11119 (N_11119,N_5106,N_5832);
or U11120 (N_11120,N_5458,N_7200);
or U11121 (N_11121,N_6909,N_7747);
nor U11122 (N_11122,N_6091,N_4514);
or U11123 (N_11123,N_5934,N_7198);
xnor U11124 (N_11124,N_7231,N_6266);
nand U11125 (N_11125,N_6964,N_7467);
and U11126 (N_11126,N_4964,N_6490);
nor U11127 (N_11127,N_6207,N_5465);
nor U11128 (N_11128,N_7987,N_5200);
or U11129 (N_11129,N_7304,N_4038);
and U11130 (N_11130,N_7484,N_5741);
nand U11131 (N_11131,N_7706,N_4379);
nand U11132 (N_11132,N_4817,N_7084);
and U11133 (N_11133,N_7271,N_4082);
or U11134 (N_11134,N_5649,N_7809);
or U11135 (N_11135,N_5387,N_4361);
or U11136 (N_11136,N_6614,N_5189);
nand U11137 (N_11137,N_5018,N_4065);
nor U11138 (N_11138,N_6818,N_5089);
or U11139 (N_11139,N_6472,N_7555);
xnor U11140 (N_11140,N_6083,N_5524);
nor U11141 (N_11141,N_7315,N_5424);
or U11142 (N_11142,N_7435,N_7167);
or U11143 (N_11143,N_6956,N_7082);
nand U11144 (N_11144,N_5397,N_4350);
nor U11145 (N_11145,N_7251,N_5850);
and U11146 (N_11146,N_6073,N_4784);
or U11147 (N_11147,N_7843,N_4003);
nand U11148 (N_11148,N_6030,N_5609);
and U11149 (N_11149,N_7299,N_5616);
and U11150 (N_11150,N_4637,N_7757);
or U11151 (N_11151,N_4276,N_7752);
and U11152 (N_11152,N_4775,N_5500);
nor U11153 (N_11153,N_6090,N_5613);
nor U11154 (N_11154,N_5337,N_6072);
and U11155 (N_11155,N_7275,N_6230);
nor U11156 (N_11156,N_5537,N_7525);
nor U11157 (N_11157,N_6332,N_4346);
and U11158 (N_11158,N_5031,N_7298);
nand U11159 (N_11159,N_4901,N_6594);
nor U11160 (N_11160,N_7476,N_7215);
or U11161 (N_11161,N_7800,N_4228);
nand U11162 (N_11162,N_7548,N_7104);
or U11163 (N_11163,N_5936,N_5755);
and U11164 (N_11164,N_5410,N_7161);
xor U11165 (N_11165,N_5597,N_5612);
nor U11166 (N_11166,N_5239,N_7472);
nor U11167 (N_11167,N_6126,N_7646);
or U11168 (N_11168,N_5091,N_6558);
and U11169 (N_11169,N_4144,N_5383);
nor U11170 (N_11170,N_5538,N_5748);
xnor U11171 (N_11171,N_5315,N_5105);
nor U11172 (N_11172,N_5742,N_5233);
and U11173 (N_11173,N_4257,N_5255);
or U11174 (N_11174,N_5366,N_4159);
or U11175 (N_11175,N_7755,N_4864);
nor U11176 (N_11176,N_6330,N_7926);
nor U11177 (N_11177,N_5986,N_4548);
or U11178 (N_11178,N_5576,N_7332);
nand U11179 (N_11179,N_4721,N_4675);
nand U11180 (N_11180,N_7162,N_6647);
nand U11181 (N_11181,N_5003,N_4922);
and U11182 (N_11182,N_6894,N_4996);
or U11183 (N_11183,N_7380,N_7040);
and U11184 (N_11184,N_5966,N_4310);
and U11185 (N_11185,N_6774,N_4100);
nor U11186 (N_11186,N_7718,N_6281);
and U11187 (N_11187,N_7997,N_4253);
nand U11188 (N_11188,N_7683,N_5419);
or U11189 (N_11189,N_5810,N_5055);
and U11190 (N_11190,N_4801,N_6481);
and U11191 (N_11191,N_7217,N_7608);
nor U11192 (N_11192,N_4185,N_4256);
or U11193 (N_11193,N_4546,N_5456);
and U11194 (N_11194,N_7937,N_4815);
xor U11195 (N_11195,N_6648,N_5027);
nand U11196 (N_11196,N_5661,N_6609);
xnor U11197 (N_11197,N_4249,N_4091);
and U11198 (N_11198,N_7108,N_7286);
xor U11199 (N_11199,N_7424,N_6426);
nand U11200 (N_11200,N_7432,N_7509);
nand U11201 (N_11201,N_5086,N_6639);
nand U11202 (N_11202,N_4835,N_4668);
or U11203 (N_11203,N_6438,N_6448);
and U11204 (N_11204,N_7960,N_5068);
nor U11205 (N_11205,N_7278,N_5021);
nor U11206 (N_11206,N_7227,N_4112);
and U11207 (N_11207,N_4617,N_7192);
and U11208 (N_11208,N_7070,N_6663);
nor U11209 (N_11209,N_7112,N_6804);
and U11210 (N_11210,N_5480,N_7515);
and U11211 (N_11211,N_6861,N_5503);
or U11212 (N_11212,N_7825,N_6675);
xor U11213 (N_11213,N_7277,N_5501);
or U11214 (N_11214,N_4921,N_4829);
or U11215 (N_11215,N_5383,N_6813);
nand U11216 (N_11216,N_4913,N_4802);
or U11217 (N_11217,N_4678,N_4643);
nand U11218 (N_11218,N_4377,N_7039);
nor U11219 (N_11219,N_5858,N_5436);
nand U11220 (N_11220,N_7206,N_7780);
nand U11221 (N_11221,N_5607,N_4275);
or U11222 (N_11222,N_5034,N_5057);
and U11223 (N_11223,N_5933,N_7901);
and U11224 (N_11224,N_4889,N_5609);
and U11225 (N_11225,N_7417,N_5279);
and U11226 (N_11226,N_5180,N_6404);
and U11227 (N_11227,N_5267,N_4118);
nor U11228 (N_11228,N_4960,N_6279);
nand U11229 (N_11229,N_7481,N_6418);
nand U11230 (N_11230,N_7648,N_6064);
nand U11231 (N_11231,N_5537,N_7049);
and U11232 (N_11232,N_5540,N_5937);
xor U11233 (N_11233,N_4999,N_6321);
or U11234 (N_11234,N_6269,N_6542);
or U11235 (N_11235,N_7148,N_4753);
or U11236 (N_11236,N_6454,N_4024);
nor U11237 (N_11237,N_6736,N_7499);
or U11238 (N_11238,N_7648,N_4364);
and U11239 (N_11239,N_7199,N_5696);
nor U11240 (N_11240,N_7866,N_5370);
and U11241 (N_11241,N_7447,N_5813);
nor U11242 (N_11242,N_5150,N_4429);
and U11243 (N_11243,N_6607,N_5709);
or U11244 (N_11244,N_7299,N_6596);
and U11245 (N_11245,N_5382,N_7343);
or U11246 (N_11246,N_4794,N_4944);
or U11247 (N_11247,N_6483,N_7022);
nand U11248 (N_11248,N_7292,N_7195);
and U11249 (N_11249,N_6982,N_6016);
nand U11250 (N_11250,N_6310,N_6390);
and U11251 (N_11251,N_6376,N_5660);
and U11252 (N_11252,N_6853,N_6127);
and U11253 (N_11253,N_7352,N_5640);
nand U11254 (N_11254,N_7670,N_7053);
or U11255 (N_11255,N_7312,N_7696);
nor U11256 (N_11256,N_4393,N_5863);
nand U11257 (N_11257,N_6960,N_7902);
nor U11258 (N_11258,N_5199,N_6563);
or U11259 (N_11259,N_4645,N_4245);
nand U11260 (N_11260,N_5363,N_5751);
nand U11261 (N_11261,N_6815,N_7548);
nand U11262 (N_11262,N_6400,N_4850);
nand U11263 (N_11263,N_4856,N_7050);
or U11264 (N_11264,N_5308,N_5157);
or U11265 (N_11265,N_6571,N_5625);
nand U11266 (N_11266,N_5338,N_4813);
nor U11267 (N_11267,N_6457,N_7246);
and U11268 (N_11268,N_4703,N_4327);
nor U11269 (N_11269,N_4789,N_7680);
nor U11270 (N_11270,N_7140,N_4368);
or U11271 (N_11271,N_4010,N_7888);
or U11272 (N_11272,N_5814,N_5126);
or U11273 (N_11273,N_7582,N_6611);
and U11274 (N_11274,N_6844,N_6092);
nand U11275 (N_11275,N_5102,N_4432);
and U11276 (N_11276,N_5425,N_6750);
nand U11277 (N_11277,N_6199,N_6908);
and U11278 (N_11278,N_6085,N_6733);
and U11279 (N_11279,N_6888,N_6365);
and U11280 (N_11280,N_4600,N_4787);
or U11281 (N_11281,N_5534,N_5081);
nor U11282 (N_11282,N_6184,N_6385);
nand U11283 (N_11283,N_6405,N_4598);
or U11284 (N_11284,N_5022,N_6655);
nor U11285 (N_11285,N_6396,N_4873);
nor U11286 (N_11286,N_7265,N_4235);
or U11287 (N_11287,N_7437,N_4287);
nand U11288 (N_11288,N_5445,N_7285);
nor U11289 (N_11289,N_6649,N_7318);
nand U11290 (N_11290,N_6450,N_7029);
xor U11291 (N_11291,N_7735,N_6210);
nor U11292 (N_11292,N_7556,N_5261);
and U11293 (N_11293,N_5674,N_4548);
nand U11294 (N_11294,N_5339,N_6560);
nand U11295 (N_11295,N_5269,N_7418);
xor U11296 (N_11296,N_6499,N_6071);
or U11297 (N_11297,N_4143,N_5723);
nand U11298 (N_11298,N_7957,N_4884);
and U11299 (N_11299,N_4783,N_5110);
xor U11300 (N_11300,N_6790,N_5346);
nor U11301 (N_11301,N_4456,N_6923);
and U11302 (N_11302,N_4703,N_6096);
and U11303 (N_11303,N_7773,N_4741);
nor U11304 (N_11304,N_6070,N_6525);
xnor U11305 (N_11305,N_6759,N_7784);
nand U11306 (N_11306,N_4867,N_5944);
xnor U11307 (N_11307,N_7792,N_5830);
nand U11308 (N_11308,N_6813,N_5494);
nand U11309 (N_11309,N_6340,N_5801);
nor U11310 (N_11310,N_6241,N_4588);
nor U11311 (N_11311,N_6257,N_5579);
and U11312 (N_11312,N_7507,N_4493);
nand U11313 (N_11313,N_7619,N_5412);
nor U11314 (N_11314,N_6244,N_7286);
or U11315 (N_11315,N_5118,N_6866);
nand U11316 (N_11316,N_4928,N_7590);
or U11317 (N_11317,N_7222,N_7401);
xnor U11318 (N_11318,N_6192,N_5406);
and U11319 (N_11319,N_4804,N_7203);
nand U11320 (N_11320,N_6021,N_4992);
and U11321 (N_11321,N_7768,N_7575);
and U11322 (N_11322,N_5222,N_4494);
nor U11323 (N_11323,N_7147,N_6101);
nor U11324 (N_11324,N_7497,N_5212);
nand U11325 (N_11325,N_6208,N_6643);
xnor U11326 (N_11326,N_7752,N_6274);
or U11327 (N_11327,N_5942,N_6010);
or U11328 (N_11328,N_6733,N_7511);
nor U11329 (N_11329,N_4010,N_5907);
nor U11330 (N_11330,N_6408,N_7106);
and U11331 (N_11331,N_7408,N_5807);
or U11332 (N_11332,N_4275,N_5556);
or U11333 (N_11333,N_4193,N_4342);
nor U11334 (N_11334,N_6137,N_4939);
nand U11335 (N_11335,N_7527,N_4721);
or U11336 (N_11336,N_6794,N_7394);
or U11337 (N_11337,N_7763,N_7369);
nand U11338 (N_11338,N_4668,N_4207);
and U11339 (N_11339,N_6829,N_6717);
nand U11340 (N_11340,N_5463,N_6836);
or U11341 (N_11341,N_6381,N_7903);
xnor U11342 (N_11342,N_6167,N_7744);
or U11343 (N_11343,N_6234,N_6405);
xnor U11344 (N_11344,N_6625,N_5347);
nor U11345 (N_11345,N_4347,N_6033);
and U11346 (N_11346,N_5753,N_6567);
nor U11347 (N_11347,N_4731,N_6913);
nor U11348 (N_11348,N_7511,N_7329);
nand U11349 (N_11349,N_4863,N_6519);
nand U11350 (N_11350,N_6829,N_5109);
nor U11351 (N_11351,N_7671,N_7422);
nand U11352 (N_11352,N_5138,N_6869);
and U11353 (N_11353,N_6613,N_5799);
or U11354 (N_11354,N_6994,N_4008);
and U11355 (N_11355,N_4016,N_6749);
and U11356 (N_11356,N_5517,N_6388);
nor U11357 (N_11357,N_7170,N_4876);
and U11358 (N_11358,N_7721,N_7452);
and U11359 (N_11359,N_6393,N_7519);
xor U11360 (N_11360,N_7121,N_7136);
nor U11361 (N_11361,N_4903,N_7934);
and U11362 (N_11362,N_6990,N_7269);
or U11363 (N_11363,N_6512,N_6472);
and U11364 (N_11364,N_5602,N_7312);
and U11365 (N_11365,N_5141,N_5223);
and U11366 (N_11366,N_6966,N_6538);
nand U11367 (N_11367,N_5696,N_4410);
nor U11368 (N_11368,N_7556,N_6644);
and U11369 (N_11369,N_6903,N_6034);
xnor U11370 (N_11370,N_5756,N_7143);
or U11371 (N_11371,N_7005,N_6840);
nor U11372 (N_11372,N_7862,N_5497);
nand U11373 (N_11373,N_5610,N_7576);
or U11374 (N_11374,N_4141,N_6832);
xor U11375 (N_11375,N_4357,N_5958);
and U11376 (N_11376,N_6613,N_6264);
or U11377 (N_11377,N_7854,N_5938);
nor U11378 (N_11378,N_7119,N_7521);
and U11379 (N_11379,N_4740,N_4256);
and U11380 (N_11380,N_4010,N_4339);
nand U11381 (N_11381,N_6233,N_5482);
nand U11382 (N_11382,N_6848,N_5014);
nand U11383 (N_11383,N_6356,N_5647);
nand U11384 (N_11384,N_6848,N_5429);
xor U11385 (N_11385,N_7350,N_5764);
or U11386 (N_11386,N_6481,N_7514);
and U11387 (N_11387,N_5909,N_6733);
or U11388 (N_11388,N_5271,N_4616);
xor U11389 (N_11389,N_6877,N_4092);
nand U11390 (N_11390,N_7150,N_4242);
nor U11391 (N_11391,N_6598,N_5591);
and U11392 (N_11392,N_6377,N_4172);
or U11393 (N_11393,N_4390,N_4041);
nand U11394 (N_11394,N_7334,N_6080);
or U11395 (N_11395,N_4404,N_5722);
or U11396 (N_11396,N_7215,N_4116);
nor U11397 (N_11397,N_4287,N_5882);
and U11398 (N_11398,N_7035,N_5866);
nor U11399 (N_11399,N_7991,N_4476);
and U11400 (N_11400,N_5202,N_5445);
or U11401 (N_11401,N_5962,N_4816);
nand U11402 (N_11402,N_5799,N_7524);
or U11403 (N_11403,N_5350,N_5320);
and U11404 (N_11404,N_6538,N_7664);
or U11405 (N_11405,N_4775,N_4035);
and U11406 (N_11406,N_7802,N_6557);
or U11407 (N_11407,N_6596,N_6854);
or U11408 (N_11408,N_7093,N_6257);
nor U11409 (N_11409,N_6610,N_7130);
nor U11410 (N_11410,N_7283,N_6208);
xor U11411 (N_11411,N_6267,N_4500);
nor U11412 (N_11412,N_5582,N_4166);
or U11413 (N_11413,N_6022,N_7043);
nand U11414 (N_11414,N_4016,N_7410);
nor U11415 (N_11415,N_6841,N_4934);
nor U11416 (N_11416,N_4975,N_5773);
nor U11417 (N_11417,N_6799,N_4292);
or U11418 (N_11418,N_6988,N_4688);
and U11419 (N_11419,N_6734,N_6962);
or U11420 (N_11420,N_6038,N_6496);
and U11421 (N_11421,N_7103,N_4777);
nor U11422 (N_11422,N_7716,N_4561);
nor U11423 (N_11423,N_4860,N_5470);
and U11424 (N_11424,N_7603,N_7959);
xnor U11425 (N_11425,N_5655,N_7245);
nand U11426 (N_11426,N_7417,N_6706);
xor U11427 (N_11427,N_4134,N_6712);
nand U11428 (N_11428,N_4128,N_7574);
xor U11429 (N_11429,N_4942,N_6443);
nand U11430 (N_11430,N_5225,N_4473);
nor U11431 (N_11431,N_4085,N_5911);
nand U11432 (N_11432,N_5830,N_6107);
or U11433 (N_11433,N_6230,N_6562);
nand U11434 (N_11434,N_6765,N_7559);
nor U11435 (N_11435,N_5435,N_7379);
and U11436 (N_11436,N_5908,N_5133);
or U11437 (N_11437,N_7526,N_7948);
and U11438 (N_11438,N_5942,N_6083);
nor U11439 (N_11439,N_5960,N_6448);
xor U11440 (N_11440,N_6338,N_6081);
nand U11441 (N_11441,N_6568,N_6456);
nor U11442 (N_11442,N_7715,N_4622);
or U11443 (N_11443,N_4984,N_6048);
and U11444 (N_11444,N_5681,N_7813);
and U11445 (N_11445,N_4065,N_6081);
and U11446 (N_11446,N_4860,N_5324);
or U11447 (N_11447,N_5699,N_6919);
or U11448 (N_11448,N_6220,N_5156);
or U11449 (N_11449,N_6867,N_7686);
or U11450 (N_11450,N_4790,N_6264);
nor U11451 (N_11451,N_4503,N_5166);
xor U11452 (N_11452,N_7534,N_7309);
and U11453 (N_11453,N_5292,N_5142);
xnor U11454 (N_11454,N_5105,N_7102);
and U11455 (N_11455,N_6417,N_5303);
nor U11456 (N_11456,N_6600,N_7549);
or U11457 (N_11457,N_7972,N_4045);
and U11458 (N_11458,N_6484,N_5767);
and U11459 (N_11459,N_4598,N_7947);
nand U11460 (N_11460,N_7135,N_5286);
nand U11461 (N_11461,N_4248,N_7697);
xor U11462 (N_11462,N_6972,N_4410);
or U11463 (N_11463,N_7882,N_5685);
nand U11464 (N_11464,N_7549,N_4858);
nand U11465 (N_11465,N_5647,N_4811);
nand U11466 (N_11466,N_7334,N_7207);
or U11467 (N_11467,N_7230,N_4073);
and U11468 (N_11468,N_7537,N_7447);
nor U11469 (N_11469,N_6850,N_4581);
or U11470 (N_11470,N_7751,N_7040);
and U11471 (N_11471,N_4471,N_5898);
and U11472 (N_11472,N_5781,N_7351);
nand U11473 (N_11473,N_4209,N_4505);
nand U11474 (N_11474,N_5083,N_4545);
and U11475 (N_11475,N_4694,N_6474);
nand U11476 (N_11476,N_7336,N_7752);
nand U11477 (N_11477,N_4849,N_7363);
nor U11478 (N_11478,N_4394,N_5982);
or U11479 (N_11479,N_6251,N_7454);
or U11480 (N_11480,N_7103,N_5843);
and U11481 (N_11481,N_4527,N_4496);
or U11482 (N_11482,N_7760,N_6366);
or U11483 (N_11483,N_5047,N_6693);
or U11484 (N_11484,N_6420,N_7372);
nor U11485 (N_11485,N_4630,N_4340);
and U11486 (N_11486,N_5549,N_5819);
or U11487 (N_11487,N_6906,N_6716);
nand U11488 (N_11488,N_5865,N_6291);
xor U11489 (N_11489,N_4857,N_7740);
nor U11490 (N_11490,N_5805,N_5810);
or U11491 (N_11491,N_7188,N_7076);
and U11492 (N_11492,N_6453,N_5930);
nor U11493 (N_11493,N_5759,N_5888);
or U11494 (N_11494,N_5944,N_7660);
or U11495 (N_11495,N_7613,N_7715);
nand U11496 (N_11496,N_7532,N_4314);
and U11497 (N_11497,N_5158,N_6353);
nand U11498 (N_11498,N_6605,N_4038);
nand U11499 (N_11499,N_6710,N_5524);
nand U11500 (N_11500,N_4064,N_7923);
xor U11501 (N_11501,N_4071,N_7629);
nand U11502 (N_11502,N_6620,N_4619);
or U11503 (N_11503,N_4969,N_4683);
nand U11504 (N_11504,N_4554,N_7560);
nor U11505 (N_11505,N_7603,N_6334);
nand U11506 (N_11506,N_7860,N_6302);
or U11507 (N_11507,N_4599,N_5159);
nand U11508 (N_11508,N_4411,N_6415);
nor U11509 (N_11509,N_7413,N_4910);
nor U11510 (N_11510,N_5739,N_7193);
and U11511 (N_11511,N_7223,N_4138);
nand U11512 (N_11512,N_6147,N_7784);
or U11513 (N_11513,N_4171,N_7334);
nor U11514 (N_11514,N_5001,N_6548);
and U11515 (N_11515,N_5035,N_6379);
and U11516 (N_11516,N_7216,N_7130);
or U11517 (N_11517,N_7301,N_6667);
or U11518 (N_11518,N_6129,N_6029);
nor U11519 (N_11519,N_6402,N_7725);
or U11520 (N_11520,N_7702,N_6278);
and U11521 (N_11521,N_7990,N_4759);
nand U11522 (N_11522,N_7466,N_7153);
or U11523 (N_11523,N_6517,N_5237);
nor U11524 (N_11524,N_7158,N_7900);
nand U11525 (N_11525,N_6807,N_6061);
nand U11526 (N_11526,N_7462,N_7510);
and U11527 (N_11527,N_7755,N_7153);
xor U11528 (N_11528,N_4952,N_5891);
nor U11529 (N_11529,N_7851,N_6846);
and U11530 (N_11530,N_5719,N_6222);
nand U11531 (N_11531,N_5239,N_4644);
or U11532 (N_11532,N_7707,N_6242);
and U11533 (N_11533,N_6840,N_4162);
or U11534 (N_11534,N_5137,N_6146);
and U11535 (N_11535,N_7094,N_7307);
nand U11536 (N_11536,N_5670,N_7326);
and U11537 (N_11537,N_7989,N_7900);
xor U11538 (N_11538,N_4738,N_7928);
nand U11539 (N_11539,N_5128,N_6985);
nand U11540 (N_11540,N_4702,N_5246);
or U11541 (N_11541,N_5117,N_6434);
nand U11542 (N_11542,N_6900,N_7564);
and U11543 (N_11543,N_6077,N_5791);
nor U11544 (N_11544,N_4510,N_7490);
nor U11545 (N_11545,N_7214,N_7410);
nor U11546 (N_11546,N_6461,N_6386);
and U11547 (N_11547,N_5316,N_4927);
nand U11548 (N_11548,N_5781,N_7754);
and U11549 (N_11549,N_6242,N_4792);
or U11550 (N_11550,N_6745,N_4151);
nand U11551 (N_11551,N_7824,N_5890);
and U11552 (N_11552,N_5545,N_7905);
and U11553 (N_11553,N_5016,N_5213);
nor U11554 (N_11554,N_7854,N_5975);
or U11555 (N_11555,N_7891,N_7146);
and U11556 (N_11556,N_7600,N_5176);
nor U11557 (N_11557,N_4927,N_7771);
and U11558 (N_11558,N_7337,N_7870);
and U11559 (N_11559,N_5202,N_7638);
or U11560 (N_11560,N_6986,N_4163);
nor U11561 (N_11561,N_5135,N_7581);
nor U11562 (N_11562,N_5189,N_7123);
nor U11563 (N_11563,N_4945,N_6573);
nor U11564 (N_11564,N_7291,N_7930);
and U11565 (N_11565,N_7771,N_5068);
nor U11566 (N_11566,N_7773,N_4627);
and U11567 (N_11567,N_7561,N_5404);
nor U11568 (N_11568,N_6190,N_4612);
or U11569 (N_11569,N_5048,N_5674);
or U11570 (N_11570,N_4615,N_4806);
nand U11571 (N_11571,N_7965,N_4506);
and U11572 (N_11572,N_7455,N_6261);
or U11573 (N_11573,N_6524,N_6359);
nor U11574 (N_11574,N_4091,N_4529);
and U11575 (N_11575,N_6286,N_4757);
or U11576 (N_11576,N_7926,N_5636);
and U11577 (N_11577,N_6131,N_4616);
or U11578 (N_11578,N_4368,N_5355);
or U11579 (N_11579,N_5699,N_4135);
nor U11580 (N_11580,N_5297,N_6855);
and U11581 (N_11581,N_6125,N_7964);
nor U11582 (N_11582,N_6981,N_6209);
and U11583 (N_11583,N_6964,N_7704);
or U11584 (N_11584,N_4796,N_7211);
nand U11585 (N_11585,N_4143,N_4433);
nor U11586 (N_11586,N_5237,N_4823);
and U11587 (N_11587,N_6597,N_7300);
and U11588 (N_11588,N_7986,N_5424);
xnor U11589 (N_11589,N_5232,N_4191);
nor U11590 (N_11590,N_6064,N_5661);
xnor U11591 (N_11591,N_4937,N_4328);
nor U11592 (N_11592,N_4932,N_5625);
or U11593 (N_11593,N_7974,N_5616);
or U11594 (N_11594,N_7396,N_4570);
or U11595 (N_11595,N_4704,N_6700);
nor U11596 (N_11596,N_6558,N_5068);
and U11597 (N_11597,N_5983,N_5042);
or U11598 (N_11598,N_7302,N_7508);
xor U11599 (N_11599,N_4401,N_5045);
or U11600 (N_11600,N_4272,N_7638);
or U11601 (N_11601,N_5311,N_5200);
or U11602 (N_11602,N_6312,N_7903);
and U11603 (N_11603,N_5724,N_6765);
nand U11604 (N_11604,N_7222,N_6419);
and U11605 (N_11605,N_4242,N_5077);
nand U11606 (N_11606,N_6705,N_4103);
nor U11607 (N_11607,N_6863,N_4591);
and U11608 (N_11608,N_5041,N_6547);
nor U11609 (N_11609,N_7905,N_6121);
nand U11610 (N_11610,N_4458,N_4747);
and U11611 (N_11611,N_6205,N_5790);
nand U11612 (N_11612,N_6230,N_4424);
xor U11613 (N_11613,N_7110,N_7833);
and U11614 (N_11614,N_7060,N_7805);
and U11615 (N_11615,N_6218,N_6039);
nand U11616 (N_11616,N_7457,N_7672);
nor U11617 (N_11617,N_5559,N_5541);
nand U11618 (N_11618,N_6810,N_4285);
nand U11619 (N_11619,N_6458,N_7399);
and U11620 (N_11620,N_7086,N_4014);
nand U11621 (N_11621,N_7659,N_4146);
or U11622 (N_11622,N_6486,N_7012);
and U11623 (N_11623,N_7501,N_6967);
and U11624 (N_11624,N_5486,N_7272);
nand U11625 (N_11625,N_6776,N_6834);
and U11626 (N_11626,N_4462,N_6949);
nor U11627 (N_11627,N_5416,N_4548);
nor U11628 (N_11628,N_7930,N_5722);
nor U11629 (N_11629,N_4190,N_7220);
and U11630 (N_11630,N_5693,N_5289);
or U11631 (N_11631,N_4319,N_5370);
or U11632 (N_11632,N_4387,N_4900);
nor U11633 (N_11633,N_5628,N_6151);
nand U11634 (N_11634,N_4794,N_5344);
nor U11635 (N_11635,N_6996,N_5634);
nand U11636 (N_11636,N_7812,N_7770);
or U11637 (N_11637,N_7047,N_6685);
nand U11638 (N_11638,N_4347,N_6931);
nor U11639 (N_11639,N_7714,N_4175);
nand U11640 (N_11640,N_7594,N_5633);
nand U11641 (N_11641,N_4666,N_4525);
or U11642 (N_11642,N_4937,N_5915);
nand U11643 (N_11643,N_7188,N_4822);
or U11644 (N_11644,N_5288,N_6037);
nand U11645 (N_11645,N_7955,N_7872);
nor U11646 (N_11646,N_7692,N_5278);
xor U11647 (N_11647,N_4566,N_5404);
xor U11648 (N_11648,N_6826,N_7746);
nand U11649 (N_11649,N_6226,N_7665);
nor U11650 (N_11650,N_6906,N_5375);
or U11651 (N_11651,N_6634,N_6872);
and U11652 (N_11652,N_6134,N_7336);
and U11653 (N_11653,N_4479,N_7355);
nor U11654 (N_11654,N_5266,N_5956);
nor U11655 (N_11655,N_5347,N_4591);
xor U11656 (N_11656,N_5579,N_6949);
nor U11657 (N_11657,N_7684,N_7940);
nor U11658 (N_11658,N_5814,N_4490);
or U11659 (N_11659,N_7498,N_6444);
or U11660 (N_11660,N_6942,N_6357);
and U11661 (N_11661,N_4685,N_5817);
xnor U11662 (N_11662,N_4187,N_6243);
nor U11663 (N_11663,N_7559,N_6647);
or U11664 (N_11664,N_5684,N_5875);
and U11665 (N_11665,N_5908,N_6732);
or U11666 (N_11666,N_4594,N_7318);
or U11667 (N_11667,N_4993,N_6407);
and U11668 (N_11668,N_4469,N_4251);
nand U11669 (N_11669,N_7367,N_4134);
or U11670 (N_11670,N_6726,N_6334);
or U11671 (N_11671,N_7132,N_6246);
or U11672 (N_11672,N_4906,N_4167);
and U11673 (N_11673,N_4804,N_6319);
nor U11674 (N_11674,N_7970,N_5320);
nand U11675 (N_11675,N_7049,N_6430);
or U11676 (N_11676,N_5336,N_6284);
nor U11677 (N_11677,N_4875,N_4856);
and U11678 (N_11678,N_6442,N_7198);
xnor U11679 (N_11679,N_5557,N_4298);
nor U11680 (N_11680,N_7618,N_5958);
nor U11681 (N_11681,N_7248,N_7918);
nand U11682 (N_11682,N_7481,N_6276);
and U11683 (N_11683,N_7822,N_7174);
nand U11684 (N_11684,N_5670,N_6867);
or U11685 (N_11685,N_6176,N_6646);
or U11686 (N_11686,N_7729,N_4256);
xnor U11687 (N_11687,N_6579,N_4002);
or U11688 (N_11688,N_7461,N_5143);
nor U11689 (N_11689,N_6969,N_5514);
nor U11690 (N_11690,N_7306,N_5772);
nand U11691 (N_11691,N_7878,N_5030);
or U11692 (N_11692,N_4641,N_4780);
nor U11693 (N_11693,N_7673,N_5530);
nand U11694 (N_11694,N_4318,N_4959);
nor U11695 (N_11695,N_6876,N_7520);
and U11696 (N_11696,N_7280,N_5331);
nor U11697 (N_11697,N_5284,N_4974);
nor U11698 (N_11698,N_4121,N_5080);
or U11699 (N_11699,N_6573,N_4220);
nand U11700 (N_11700,N_7852,N_4681);
or U11701 (N_11701,N_6957,N_6484);
or U11702 (N_11702,N_5338,N_6026);
xor U11703 (N_11703,N_6795,N_5456);
nor U11704 (N_11704,N_4566,N_5985);
nor U11705 (N_11705,N_5806,N_7466);
and U11706 (N_11706,N_4877,N_5901);
nand U11707 (N_11707,N_6962,N_7518);
nand U11708 (N_11708,N_6960,N_4476);
nand U11709 (N_11709,N_7748,N_7871);
xor U11710 (N_11710,N_5679,N_5720);
nand U11711 (N_11711,N_4030,N_4083);
and U11712 (N_11712,N_5032,N_7264);
nand U11713 (N_11713,N_7188,N_6485);
and U11714 (N_11714,N_5086,N_7243);
nor U11715 (N_11715,N_7846,N_4158);
nor U11716 (N_11716,N_4175,N_7817);
nand U11717 (N_11717,N_6781,N_5666);
or U11718 (N_11718,N_7280,N_6400);
and U11719 (N_11719,N_6792,N_4779);
nand U11720 (N_11720,N_5769,N_4253);
xor U11721 (N_11721,N_6298,N_5935);
and U11722 (N_11722,N_4190,N_7604);
and U11723 (N_11723,N_5016,N_6544);
nand U11724 (N_11724,N_5925,N_4985);
nand U11725 (N_11725,N_4889,N_7202);
nand U11726 (N_11726,N_4759,N_7674);
or U11727 (N_11727,N_7956,N_7413);
nor U11728 (N_11728,N_4465,N_6550);
and U11729 (N_11729,N_6484,N_7231);
nand U11730 (N_11730,N_4818,N_4481);
or U11731 (N_11731,N_7904,N_5212);
nor U11732 (N_11732,N_7566,N_5146);
or U11733 (N_11733,N_5675,N_5561);
nor U11734 (N_11734,N_6008,N_6634);
and U11735 (N_11735,N_5076,N_5276);
or U11736 (N_11736,N_4219,N_7795);
and U11737 (N_11737,N_5703,N_5757);
or U11738 (N_11738,N_5214,N_4937);
and U11739 (N_11739,N_6567,N_6966);
nor U11740 (N_11740,N_5266,N_4350);
nor U11741 (N_11741,N_6941,N_6327);
nand U11742 (N_11742,N_6960,N_4977);
and U11743 (N_11743,N_5083,N_5345);
nor U11744 (N_11744,N_7160,N_7492);
nand U11745 (N_11745,N_4615,N_6097);
nor U11746 (N_11746,N_7344,N_4857);
nor U11747 (N_11747,N_5062,N_7309);
xor U11748 (N_11748,N_7131,N_6466);
xnor U11749 (N_11749,N_4770,N_6625);
nor U11750 (N_11750,N_4542,N_5549);
xnor U11751 (N_11751,N_7632,N_6044);
and U11752 (N_11752,N_4672,N_7947);
nor U11753 (N_11753,N_6372,N_5582);
xor U11754 (N_11754,N_6421,N_7108);
nor U11755 (N_11755,N_6160,N_6582);
xnor U11756 (N_11756,N_4205,N_4707);
nor U11757 (N_11757,N_7362,N_5866);
nor U11758 (N_11758,N_6203,N_5884);
xor U11759 (N_11759,N_6673,N_7078);
nand U11760 (N_11760,N_6583,N_6797);
and U11761 (N_11761,N_5519,N_6457);
and U11762 (N_11762,N_4806,N_4957);
or U11763 (N_11763,N_7403,N_6843);
and U11764 (N_11764,N_7039,N_5894);
or U11765 (N_11765,N_4229,N_7316);
nor U11766 (N_11766,N_6144,N_5077);
nand U11767 (N_11767,N_6779,N_4404);
xnor U11768 (N_11768,N_6195,N_5321);
nand U11769 (N_11769,N_5597,N_4414);
or U11770 (N_11770,N_7464,N_6751);
xor U11771 (N_11771,N_7208,N_4285);
and U11772 (N_11772,N_6979,N_5073);
or U11773 (N_11773,N_4821,N_6259);
nand U11774 (N_11774,N_5394,N_6182);
nor U11775 (N_11775,N_5330,N_5148);
or U11776 (N_11776,N_7299,N_6830);
or U11777 (N_11777,N_7481,N_4176);
nand U11778 (N_11778,N_4207,N_6830);
nand U11779 (N_11779,N_4282,N_5122);
or U11780 (N_11780,N_5979,N_5689);
nand U11781 (N_11781,N_6149,N_6927);
nand U11782 (N_11782,N_4085,N_5946);
nand U11783 (N_11783,N_4498,N_4683);
nor U11784 (N_11784,N_5785,N_7436);
xnor U11785 (N_11785,N_7820,N_6786);
nand U11786 (N_11786,N_5217,N_4369);
xor U11787 (N_11787,N_7537,N_6454);
nor U11788 (N_11788,N_4818,N_4227);
xor U11789 (N_11789,N_7503,N_6065);
nor U11790 (N_11790,N_6433,N_4312);
or U11791 (N_11791,N_4557,N_5005);
nand U11792 (N_11792,N_7731,N_5270);
nand U11793 (N_11793,N_5532,N_7379);
or U11794 (N_11794,N_4568,N_7087);
and U11795 (N_11795,N_7359,N_6659);
xnor U11796 (N_11796,N_4450,N_4062);
nor U11797 (N_11797,N_4329,N_5070);
nor U11798 (N_11798,N_7936,N_4177);
or U11799 (N_11799,N_5415,N_6280);
or U11800 (N_11800,N_5836,N_5348);
nand U11801 (N_11801,N_4462,N_6038);
xor U11802 (N_11802,N_5980,N_6247);
nand U11803 (N_11803,N_7088,N_7279);
and U11804 (N_11804,N_5447,N_7965);
nor U11805 (N_11805,N_4853,N_4825);
or U11806 (N_11806,N_4310,N_4967);
or U11807 (N_11807,N_5865,N_4561);
and U11808 (N_11808,N_4174,N_5827);
and U11809 (N_11809,N_6286,N_5679);
xor U11810 (N_11810,N_6488,N_5594);
nor U11811 (N_11811,N_7575,N_4047);
nand U11812 (N_11812,N_4440,N_6333);
nand U11813 (N_11813,N_5997,N_6646);
and U11814 (N_11814,N_4704,N_4133);
and U11815 (N_11815,N_6351,N_6212);
or U11816 (N_11816,N_5955,N_6348);
or U11817 (N_11817,N_4785,N_4411);
and U11818 (N_11818,N_5185,N_4369);
and U11819 (N_11819,N_6057,N_4368);
nor U11820 (N_11820,N_7758,N_7537);
and U11821 (N_11821,N_7507,N_6481);
nand U11822 (N_11822,N_5017,N_5354);
nand U11823 (N_11823,N_6818,N_6366);
or U11824 (N_11824,N_4329,N_5075);
nand U11825 (N_11825,N_4496,N_6069);
xnor U11826 (N_11826,N_7519,N_5554);
nor U11827 (N_11827,N_5701,N_5000);
xor U11828 (N_11828,N_6398,N_6960);
nor U11829 (N_11829,N_6167,N_4167);
and U11830 (N_11830,N_6380,N_4967);
nor U11831 (N_11831,N_7516,N_6006);
or U11832 (N_11832,N_5644,N_5765);
or U11833 (N_11833,N_4995,N_4883);
nand U11834 (N_11834,N_6377,N_7942);
and U11835 (N_11835,N_5661,N_6266);
or U11836 (N_11836,N_6257,N_6623);
nor U11837 (N_11837,N_6936,N_7613);
or U11838 (N_11838,N_7812,N_5718);
nor U11839 (N_11839,N_7318,N_7580);
nor U11840 (N_11840,N_4674,N_5344);
or U11841 (N_11841,N_6759,N_4627);
nor U11842 (N_11842,N_5531,N_4951);
or U11843 (N_11843,N_4734,N_5498);
nor U11844 (N_11844,N_5699,N_5359);
or U11845 (N_11845,N_6643,N_5554);
or U11846 (N_11846,N_5749,N_6685);
nor U11847 (N_11847,N_5979,N_4372);
or U11848 (N_11848,N_7393,N_6079);
and U11849 (N_11849,N_7366,N_4538);
and U11850 (N_11850,N_7583,N_4535);
nand U11851 (N_11851,N_7210,N_6089);
and U11852 (N_11852,N_4535,N_4391);
or U11853 (N_11853,N_4064,N_4440);
nand U11854 (N_11854,N_6281,N_7120);
nand U11855 (N_11855,N_7039,N_6871);
nand U11856 (N_11856,N_4179,N_7191);
nor U11857 (N_11857,N_5567,N_7578);
or U11858 (N_11858,N_5166,N_6563);
nand U11859 (N_11859,N_6156,N_4253);
and U11860 (N_11860,N_4087,N_7570);
and U11861 (N_11861,N_4864,N_7714);
nor U11862 (N_11862,N_7010,N_6010);
and U11863 (N_11863,N_6113,N_4661);
nand U11864 (N_11864,N_5312,N_4516);
nor U11865 (N_11865,N_5820,N_4737);
xnor U11866 (N_11866,N_5035,N_5275);
or U11867 (N_11867,N_5780,N_4746);
and U11868 (N_11868,N_4896,N_4558);
nand U11869 (N_11869,N_7347,N_4664);
or U11870 (N_11870,N_7186,N_5429);
and U11871 (N_11871,N_6089,N_6858);
or U11872 (N_11872,N_4405,N_4940);
and U11873 (N_11873,N_6522,N_4813);
nand U11874 (N_11874,N_7477,N_4567);
or U11875 (N_11875,N_4699,N_7513);
nand U11876 (N_11876,N_4149,N_6280);
nand U11877 (N_11877,N_7606,N_6649);
or U11878 (N_11878,N_4540,N_7522);
xnor U11879 (N_11879,N_6754,N_4805);
and U11880 (N_11880,N_7591,N_6639);
nor U11881 (N_11881,N_4514,N_7183);
and U11882 (N_11882,N_7066,N_6716);
nand U11883 (N_11883,N_5656,N_5233);
nor U11884 (N_11884,N_4624,N_4875);
xor U11885 (N_11885,N_4270,N_7953);
xor U11886 (N_11886,N_4740,N_4064);
nand U11887 (N_11887,N_4749,N_6609);
nor U11888 (N_11888,N_6410,N_5892);
nand U11889 (N_11889,N_6421,N_4755);
or U11890 (N_11890,N_7340,N_6008);
nand U11891 (N_11891,N_5314,N_5967);
nor U11892 (N_11892,N_4093,N_4728);
and U11893 (N_11893,N_6858,N_5324);
nor U11894 (N_11894,N_6240,N_4381);
nand U11895 (N_11895,N_6318,N_7200);
nand U11896 (N_11896,N_7700,N_6420);
and U11897 (N_11897,N_5307,N_7474);
nand U11898 (N_11898,N_5547,N_4158);
nor U11899 (N_11899,N_4267,N_7479);
or U11900 (N_11900,N_6983,N_4382);
nor U11901 (N_11901,N_6811,N_5660);
and U11902 (N_11902,N_7798,N_4598);
nor U11903 (N_11903,N_4343,N_4544);
or U11904 (N_11904,N_6628,N_6939);
nor U11905 (N_11905,N_4483,N_5979);
or U11906 (N_11906,N_7753,N_5705);
xor U11907 (N_11907,N_5704,N_7296);
or U11908 (N_11908,N_6721,N_7688);
nand U11909 (N_11909,N_5453,N_4642);
and U11910 (N_11910,N_4950,N_7664);
or U11911 (N_11911,N_5539,N_5532);
nand U11912 (N_11912,N_6434,N_5061);
and U11913 (N_11913,N_7494,N_6210);
nor U11914 (N_11914,N_7065,N_7826);
nand U11915 (N_11915,N_6133,N_5721);
nand U11916 (N_11916,N_7905,N_7840);
nor U11917 (N_11917,N_4323,N_4290);
nor U11918 (N_11918,N_7034,N_6804);
xor U11919 (N_11919,N_5476,N_4322);
nor U11920 (N_11920,N_6977,N_6819);
or U11921 (N_11921,N_6934,N_5501);
or U11922 (N_11922,N_7686,N_4616);
and U11923 (N_11923,N_6422,N_4089);
or U11924 (N_11924,N_5242,N_6833);
nor U11925 (N_11925,N_7542,N_7315);
nand U11926 (N_11926,N_7474,N_4017);
nand U11927 (N_11927,N_6362,N_5105);
nor U11928 (N_11928,N_4303,N_7945);
or U11929 (N_11929,N_5959,N_5396);
or U11930 (N_11930,N_4845,N_6456);
or U11931 (N_11931,N_6302,N_5674);
nor U11932 (N_11932,N_6999,N_4018);
nand U11933 (N_11933,N_6597,N_6360);
or U11934 (N_11934,N_5997,N_4395);
or U11935 (N_11935,N_6454,N_5570);
or U11936 (N_11936,N_5875,N_5889);
or U11937 (N_11937,N_4867,N_4292);
xor U11938 (N_11938,N_4117,N_6775);
and U11939 (N_11939,N_5691,N_5967);
or U11940 (N_11940,N_6199,N_6851);
nor U11941 (N_11941,N_6974,N_5957);
nand U11942 (N_11942,N_6980,N_6256);
xnor U11943 (N_11943,N_6788,N_4284);
nand U11944 (N_11944,N_4417,N_6077);
nand U11945 (N_11945,N_4764,N_6820);
or U11946 (N_11946,N_6969,N_6404);
or U11947 (N_11947,N_5069,N_4652);
or U11948 (N_11948,N_6416,N_7367);
nor U11949 (N_11949,N_7898,N_7618);
nand U11950 (N_11950,N_4342,N_5181);
and U11951 (N_11951,N_7567,N_6382);
nand U11952 (N_11952,N_5367,N_7658);
xnor U11953 (N_11953,N_7288,N_6210);
nand U11954 (N_11954,N_5199,N_7931);
or U11955 (N_11955,N_6417,N_6242);
nand U11956 (N_11956,N_5738,N_6812);
and U11957 (N_11957,N_4303,N_6289);
xor U11958 (N_11958,N_4244,N_6439);
and U11959 (N_11959,N_6362,N_6406);
nor U11960 (N_11960,N_5150,N_7294);
nor U11961 (N_11961,N_4749,N_6835);
xnor U11962 (N_11962,N_6845,N_7390);
nand U11963 (N_11963,N_6281,N_6596);
or U11964 (N_11964,N_7317,N_4547);
and U11965 (N_11965,N_7024,N_5637);
and U11966 (N_11966,N_6768,N_6514);
xnor U11967 (N_11967,N_6111,N_7140);
xor U11968 (N_11968,N_7524,N_5375);
or U11969 (N_11969,N_4646,N_7998);
or U11970 (N_11970,N_5856,N_7669);
nor U11971 (N_11971,N_6783,N_4173);
or U11972 (N_11972,N_5751,N_5957);
nand U11973 (N_11973,N_5774,N_7145);
xor U11974 (N_11974,N_4148,N_7761);
nand U11975 (N_11975,N_5763,N_6959);
or U11976 (N_11976,N_7604,N_7511);
nor U11977 (N_11977,N_4091,N_5921);
xor U11978 (N_11978,N_4628,N_5208);
nand U11979 (N_11979,N_6176,N_5529);
xor U11980 (N_11980,N_4311,N_5876);
and U11981 (N_11981,N_4920,N_6440);
nor U11982 (N_11982,N_4886,N_5492);
nand U11983 (N_11983,N_4282,N_4222);
and U11984 (N_11984,N_4171,N_5092);
or U11985 (N_11985,N_5883,N_7827);
and U11986 (N_11986,N_5510,N_7989);
and U11987 (N_11987,N_7414,N_7308);
nor U11988 (N_11988,N_4755,N_4872);
nor U11989 (N_11989,N_6980,N_6429);
and U11990 (N_11990,N_5522,N_7763);
and U11991 (N_11991,N_4779,N_4013);
and U11992 (N_11992,N_5819,N_6694);
or U11993 (N_11993,N_7523,N_4096);
and U11994 (N_11994,N_7339,N_7276);
xnor U11995 (N_11995,N_7247,N_4090);
nand U11996 (N_11996,N_6087,N_4905);
nor U11997 (N_11997,N_6319,N_6121);
xor U11998 (N_11998,N_7888,N_6153);
nand U11999 (N_11999,N_7262,N_7404);
or U12000 (N_12000,N_11647,N_9011);
or U12001 (N_12001,N_8732,N_10455);
and U12002 (N_12002,N_10530,N_8713);
or U12003 (N_12003,N_10976,N_11610);
and U12004 (N_12004,N_8674,N_11532);
or U12005 (N_12005,N_10294,N_8703);
nand U12006 (N_12006,N_11227,N_8447);
and U12007 (N_12007,N_9570,N_11615);
xor U12008 (N_12008,N_9194,N_11894);
and U12009 (N_12009,N_8688,N_9975);
nand U12010 (N_12010,N_9938,N_11165);
or U12011 (N_12011,N_9572,N_8277);
nand U12012 (N_12012,N_9984,N_11793);
nor U12013 (N_12013,N_10064,N_9457);
and U12014 (N_12014,N_9400,N_11932);
or U12015 (N_12015,N_9514,N_11650);
nand U12016 (N_12016,N_10839,N_11985);
nor U12017 (N_12017,N_9836,N_11789);
or U12018 (N_12018,N_10742,N_9109);
xnor U12019 (N_12019,N_11234,N_9258);
or U12020 (N_12020,N_11867,N_10861);
xnor U12021 (N_12021,N_10424,N_11443);
and U12022 (N_12022,N_8931,N_10324);
nor U12023 (N_12023,N_9104,N_11449);
xnor U12024 (N_12024,N_9448,N_11909);
nand U12025 (N_12025,N_10554,N_11683);
nor U12026 (N_12026,N_9830,N_9227);
nor U12027 (N_12027,N_11982,N_8499);
nand U12028 (N_12028,N_11111,N_11711);
or U12029 (N_12029,N_11902,N_10737);
and U12030 (N_12030,N_10917,N_10168);
xnor U12031 (N_12031,N_9994,N_8344);
nor U12032 (N_12032,N_10415,N_11682);
nand U12033 (N_12033,N_9134,N_8342);
or U12034 (N_12034,N_9107,N_10432);
or U12035 (N_12035,N_10134,N_8837);
and U12036 (N_12036,N_9360,N_11228);
or U12037 (N_12037,N_8297,N_11336);
and U12038 (N_12038,N_9912,N_11915);
xor U12039 (N_12039,N_8336,N_8070);
nor U12040 (N_12040,N_8612,N_9822);
nand U12041 (N_12041,N_9182,N_11980);
nor U12042 (N_12042,N_9596,N_11887);
nor U12043 (N_12043,N_9166,N_10207);
or U12044 (N_12044,N_9467,N_8908);
xnor U12045 (N_12045,N_10572,N_11349);
nand U12046 (N_12046,N_8477,N_8108);
nand U12047 (N_12047,N_8268,N_9455);
nor U12048 (N_12048,N_11340,N_8259);
nand U12049 (N_12049,N_10338,N_9224);
or U12050 (N_12050,N_9831,N_9105);
or U12051 (N_12051,N_9679,N_8444);
nand U12052 (N_12052,N_8074,N_9976);
or U12053 (N_12053,N_11577,N_10582);
nand U12054 (N_12054,N_9721,N_8968);
nand U12055 (N_12055,N_11245,N_8386);
and U12056 (N_12056,N_11448,N_11596);
nand U12057 (N_12057,N_8044,N_8399);
nand U12058 (N_12058,N_9432,N_8600);
nor U12059 (N_12059,N_10702,N_9311);
xor U12060 (N_12060,N_10150,N_9066);
nor U12061 (N_12061,N_9126,N_8207);
and U12062 (N_12062,N_11490,N_10221);
xor U12063 (N_12063,N_8029,N_8003);
xnor U12064 (N_12064,N_8747,N_11465);
nor U12065 (N_12065,N_11433,N_11531);
nand U12066 (N_12066,N_11220,N_10853);
and U12067 (N_12067,N_9404,N_8952);
nand U12068 (N_12068,N_11613,N_10716);
nand U12069 (N_12069,N_8173,N_8187);
nand U12070 (N_12070,N_11566,N_9137);
nor U12071 (N_12071,N_8402,N_10195);
nand U12072 (N_12072,N_10587,N_9284);
nand U12073 (N_12073,N_11099,N_9363);
and U12074 (N_12074,N_8682,N_11046);
or U12075 (N_12075,N_11469,N_9072);
or U12076 (N_12076,N_11677,N_10916);
or U12077 (N_12077,N_8472,N_8198);
xor U12078 (N_12078,N_9700,N_9743);
nor U12079 (N_12079,N_10884,N_8991);
xor U12080 (N_12080,N_10577,N_10343);
nor U12081 (N_12081,N_8624,N_8690);
or U12082 (N_12082,N_9250,N_8239);
or U12083 (N_12083,N_9030,N_8417);
xor U12084 (N_12084,N_9565,N_11248);
nor U12085 (N_12085,N_10416,N_10192);
nand U12086 (N_12086,N_11590,N_9583);
nand U12087 (N_12087,N_9487,N_11972);
and U12088 (N_12088,N_10220,N_9320);
xnor U12089 (N_12089,N_8067,N_11146);
nor U12090 (N_12090,N_11664,N_8346);
and U12091 (N_12091,N_11246,N_9767);
nor U12092 (N_12092,N_9128,N_11749);
nand U12093 (N_12093,N_8271,N_11484);
nor U12094 (N_12094,N_8007,N_11089);
xor U12095 (N_12095,N_11928,N_10399);
nand U12096 (N_12096,N_9395,N_11178);
nand U12097 (N_12097,N_8531,N_9275);
nor U12098 (N_12098,N_9559,N_8214);
or U12099 (N_12099,N_8331,N_8588);
and U12100 (N_12100,N_11374,N_11693);
nand U12101 (N_12101,N_11212,N_11292);
nand U12102 (N_12102,N_11468,N_10512);
or U12103 (N_12103,N_11062,N_10678);
nor U12104 (N_12104,N_8670,N_10518);
nand U12105 (N_12105,N_9242,N_11203);
nor U12106 (N_12106,N_11093,N_8753);
nand U12107 (N_12107,N_10404,N_10380);
and U12108 (N_12108,N_11418,N_10820);
nand U12109 (N_12109,N_9093,N_11026);
and U12110 (N_12110,N_10546,N_11736);
and U12111 (N_12111,N_8419,N_11954);
or U12112 (N_12112,N_9452,N_10879);
or U12113 (N_12113,N_8864,N_9716);
and U12114 (N_12114,N_8653,N_9353);
or U12115 (N_12115,N_11969,N_10584);
and U12116 (N_12116,N_10501,N_8564);
nor U12117 (N_12117,N_11522,N_11463);
and U12118 (N_12118,N_9058,N_11348);
nand U12119 (N_12119,N_9887,N_8665);
or U12120 (N_12120,N_9437,N_10037);
nand U12121 (N_12121,N_10985,N_11014);
xor U12122 (N_12122,N_9842,N_10537);
nand U12123 (N_12123,N_8977,N_9903);
nand U12124 (N_12124,N_10379,N_9879);
or U12125 (N_12125,N_10001,N_8311);
nand U12126 (N_12126,N_11413,N_10472);
nor U12127 (N_12127,N_11161,N_9026);
nor U12128 (N_12128,N_8216,N_8549);
and U12129 (N_12129,N_8082,N_9946);
xnor U12130 (N_12130,N_9986,N_9053);
or U12131 (N_12131,N_8269,N_10075);
nor U12132 (N_12132,N_9874,N_11755);
and U12133 (N_12133,N_9253,N_8850);
or U12134 (N_12134,N_8159,N_8878);
and U12135 (N_12135,N_11482,N_10610);
or U12136 (N_12136,N_10034,N_9056);
or U12137 (N_12137,N_8761,N_11629);
nor U12138 (N_12138,N_8295,N_11231);
or U12139 (N_12139,N_9853,N_9422);
nor U12140 (N_12140,N_9713,N_8835);
and U12141 (N_12141,N_10239,N_9435);
and U12142 (N_12142,N_11600,N_10061);
nor U12143 (N_12143,N_9140,N_11565);
and U12144 (N_12144,N_11023,N_10315);
and U12145 (N_12145,N_11611,N_8473);
and U12146 (N_12146,N_8847,N_8806);
nand U12147 (N_12147,N_11086,N_8493);
or U12148 (N_12148,N_8022,N_8001);
nand U12149 (N_12149,N_11423,N_10918);
nand U12150 (N_12150,N_8140,N_11623);
nand U12151 (N_12151,N_10878,N_11807);
nor U12152 (N_12152,N_11095,N_8749);
nor U12153 (N_12153,N_11714,N_10848);
nand U12154 (N_12154,N_8085,N_10511);
nor U12155 (N_12155,N_11801,N_9247);
nor U12156 (N_12156,N_8411,N_10515);
nand U12157 (N_12157,N_9013,N_8695);
and U12158 (N_12158,N_10564,N_9619);
and U12159 (N_12159,N_10476,N_11656);
xor U12160 (N_12160,N_8936,N_8142);
nor U12161 (N_12161,N_9560,N_8916);
or U12162 (N_12162,N_8405,N_10965);
or U12163 (N_12163,N_8476,N_9734);
xor U12164 (N_12164,N_11335,N_8450);
or U12165 (N_12165,N_11820,N_10750);
nand U12166 (N_12166,N_10816,N_10935);
nand U12167 (N_12167,N_11857,N_10382);
and U12168 (N_12168,N_11011,N_11300);
and U12169 (N_12169,N_8481,N_10883);
nand U12170 (N_12170,N_8807,N_9699);
nand U12171 (N_12171,N_11988,N_8971);
or U12172 (N_12172,N_9664,N_11068);
nand U12173 (N_12173,N_8731,N_11944);
or U12174 (N_12174,N_8182,N_11117);
and U12175 (N_12175,N_8061,N_11122);
nor U12176 (N_12176,N_8275,N_8869);
and U12177 (N_12177,N_8894,N_8560);
nand U12178 (N_12178,N_9660,N_11655);
xnor U12179 (N_12179,N_8967,N_10639);
or U12180 (N_12180,N_11872,N_11933);
nand U12181 (N_12181,N_8743,N_9564);
nor U12182 (N_12182,N_10082,N_11038);
nor U12183 (N_12183,N_8354,N_8981);
nor U12184 (N_12184,N_11169,N_11390);
or U12185 (N_12185,N_10891,N_10200);
and U12186 (N_12186,N_8147,N_10912);
nand U12187 (N_12187,N_10780,N_10489);
and U12188 (N_12188,N_11045,N_10899);
or U12189 (N_12189,N_8721,N_10252);
or U12190 (N_12190,N_8795,N_8832);
and U12191 (N_12191,N_10233,N_9703);
or U12192 (N_12192,N_8441,N_10442);
and U12193 (N_12193,N_11271,N_11657);
and U12194 (N_12194,N_8525,N_11121);
nand U12195 (N_12195,N_10216,N_8464);
nor U12196 (N_12196,N_8597,N_10056);
nor U12197 (N_12197,N_8640,N_10579);
or U12198 (N_12198,N_9819,N_9111);
nor U12199 (N_12199,N_10967,N_11029);
or U12200 (N_12200,N_9654,N_10269);
xnor U12201 (N_12201,N_11496,N_10612);
nand U12202 (N_12202,N_10445,N_9554);
nor U12203 (N_12203,N_9313,N_8577);
or U12204 (N_12204,N_8635,N_9981);
or U12205 (N_12205,N_10766,N_10544);
nor U12206 (N_12206,N_11030,N_9955);
nor U12207 (N_12207,N_8057,N_8824);
or U12208 (N_12208,N_11471,N_11575);
nor U12209 (N_12209,N_8181,N_10251);
xor U12210 (N_12210,N_9155,N_11144);
nand U12211 (N_12211,N_9511,N_10851);
nand U12212 (N_12212,N_9201,N_11022);
nand U12213 (N_12213,N_10413,N_10684);
and U12214 (N_12214,N_10059,N_9607);
nand U12215 (N_12215,N_9945,N_9573);
nand U12216 (N_12216,N_11622,N_11659);
nand U12217 (N_12217,N_11091,N_9029);
or U12218 (N_12218,N_8118,N_9672);
or U12219 (N_12219,N_9526,N_10290);
or U12220 (N_12220,N_11183,N_11432);
and U12221 (N_12221,N_8089,N_8486);
and U12222 (N_12222,N_10295,N_11377);
xnor U12223 (N_12223,N_8491,N_8449);
nor U12224 (N_12224,N_10845,N_11997);
or U12225 (N_12225,N_10408,N_10213);
and U12226 (N_12226,N_8808,N_9826);
nor U12227 (N_12227,N_8179,N_11759);
nor U12228 (N_12228,N_9845,N_10040);
or U12229 (N_12229,N_9517,N_8265);
nor U12230 (N_12230,N_8408,N_9388);
or U12231 (N_12231,N_11900,N_8812);
xor U12232 (N_12232,N_8112,N_10648);
nand U12233 (N_12233,N_9031,N_9318);
nand U12234 (N_12234,N_8434,N_11576);
nor U12235 (N_12235,N_9054,N_8523);
nor U12236 (N_12236,N_9589,N_10519);
or U12237 (N_12237,N_9235,N_8765);
nand U12238 (N_12238,N_9894,N_11096);
nor U12239 (N_12239,N_9685,N_10688);
and U12240 (N_12240,N_9043,N_10151);
and U12241 (N_12241,N_11644,N_11703);
xnor U12242 (N_12242,N_11354,N_10398);
nand U12243 (N_12243,N_9491,N_9528);
or U12244 (N_12244,N_10254,N_10317);
and U12245 (N_12245,N_11207,N_8851);
or U12246 (N_12246,N_9369,N_10227);
xor U12247 (N_12247,N_9101,N_11937);
or U12248 (N_12248,N_9621,N_8648);
and U12249 (N_12249,N_11466,N_11055);
or U12250 (N_12250,N_9793,N_8252);
nand U12251 (N_12251,N_8905,N_11367);
or U12252 (N_12252,N_8059,N_8261);
nor U12253 (N_12253,N_9979,N_8668);
nor U12254 (N_12254,N_8006,N_9156);
and U12255 (N_12255,N_9060,N_10031);
nor U12256 (N_12256,N_8789,N_9788);
nand U12257 (N_12257,N_9091,N_11483);
nor U12258 (N_12258,N_9418,N_11572);
nand U12259 (N_12259,N_8367,N_11235);
nand U12260 (N_12260,N_9944,N_8002);
nor U12261 (N_12261,N_10854,N_11078);
nand U12262 (N_12262,N_11742,N_11306);
or U12263 (N_12263,N_8959,N_10760);
nand U12264 (N_12264,N_11559,N_9297);
nand U12265 (N_12265,N_9474,N_9714);
and U12266 (N_12266,N_9334,N_8904);
nor U12267 (N_12267,N_9493,N_11201);
nand U12268 (N_12268,N_8706,N_9186);
nand U12269 (N_12269,N_10029,N_9612);
or U12270 (N_12270,N_9886,N_8236);
or U12271 (N_12271,N_11036,N_8226);
and U12272 (N_12272,N_11239,N_8522);
nor U12273 (N_12273,N_11603,N_9658);
nand U12274 (N_12274,N_9356,N_9578);
nand U12275 (N_12275,N_8698,N_11082);
nand U12276 (N_12276,N_10671,N_11304);
or U12277 (N_12277,N_9231,N_10426);
nand U12278 (N_12278,N_9215,N_11541);
nand U12279 (N_12279,N_10656,N_10817);
nor U12280 (N_12280,N_10000,N_8361);
xor U12281 (N_12281,N_8857,N_8209);
and U12282 (N_12282,N_10348,N_11148);
nand U12283 (N_12283,N_10533,N_9648);
and U12284 (N_12284,N_10531,N_10043);
or U12285 (N_12285,N_10499,N_9266);
or U12286 (N_12286,N_10473,N_11870);
and U12287 (N_12287,N_11869,N_10521);
and U12288 (N_12288,N_8774,N_11792);
nand U12289 (N_12289,N_10253,N_8911);
nor U12290 (N_12290,N_11296,N_8117);
nor U12291 (N_12291,N_8786,N_8772);
or U12292 (N_12292,N_11607,N_8136);
nor U12293 (N_12293,N_11673,N_10764);
nor U12294 (N_12294,N_11593,N_8780);
and U12295 (N_12295,N_11560,N_8319);
and U12296 (N_12296,N_8521,N_9278);
nor U12297 (N_12297,N_8219,N_10797);
and U12298 (N_12298,N_10433,N_11511);
nand U12299 (N_12299,N_8551,N_10673);
nor U12300 (N_12300,N_8675,N_8858);
nor U12301 (N_12301,N_8170,N_10165);
nor U12302 (N_12302,N_10339,N_10858);
xor U12303 (N_12303,N_9960,N_9728);
nand U12304 (N_12304,N_11184,N_11290);
nor U12305 (N_12305,N_9846,N_10135);
or U12306 (N_12306,N_11224,N_11003);
and U12307 (N_12307,N_10312,N_11415);
or U12308 (N_12308,N_10677,N_11131);
nor U12309 (N_12309,N_8664,N_9814);
or U12310 (N_12310,N_9602,N_9744);
or U12311 (N_12311,N_8072,N_9020);
nand U12312 (N_12312,N_8567,N_9661);
nor U12313 (N_12313,N_9824,N_8188);
nor U12314 (N_12314,N_9597,N_8392);
nand U12315 (N_12315,N_8422,N_9723);
nor U12316 (N_12316,N_8679,N_9539);
nand U12317 (N_12317,N_11426,N_9791);
nor U12318 (N_12318,N_11193,N_10155);
nand U12319 (N_12319,N_10255,N_9248);
and U12320 (N_12320,N_8819,N_8393);
and U12321 (N_12321,N_9234,N_11400);
nor U12322 (N_12322,N_10388,N_10553);
nand U12323 (N_12323,N_10856,N_8502);
xor U12324 (N_12324,N_10555,N_8797);
xor U12325 (N_12325,N_10154,N_11680);
or U12326 (N_12326,N_10403,N_11083);
nand U12327 (N_12327,N_8183,N_11993);
and U12328 (N_12328,N_10145,N_8250);
nor U12329 (N_12329,N_8875,N_11343);
xnor U12330 (N_12330,N_8141,N_8056);
nor U12331 (N_12331,N_9600,N_9562);
nand U12332 (N_12332,N_8069,N_11259);
nor U12333 (N_12333,N_10423,N_10890);
xnor U12334 (N_12334,N_11355,N_11523);
and U12335 (N_12335,N_11788,N_10568);
nor U12336 (N_12336,N_8724,N_9425);
nand U12337 (N_12337,N_8933,N_11485);
nand U12338 (N_12338,N_8841,N_10328);
or U12339 (N_12339,N_11977,N_10468);
nand U12340 (N_12340,N_9323,N_11581);
nand U12341 (N_12341,N_9127,N_8253);
nand U12342 (N_12342,N_11106,N_9580);
xor U12343 (N_12343,N_8917,N_10974);
xnor U12344 (N_12344,N_8678,N_10093);
nand U12345 (N_12345,N_10514,N_11725);
or U12346 (N_12346,N_10924,N_8415);
nand U12347 (N_12347,N_9015,N_8960);
and U12348 (N_12348,N_8340,N_10488);
and U12349 (N_12349,N_11110,N_11457);
and U12350 (N_12350,N_9270,N_9471);
nand U12351 (N_12351,N_11614,N_11351);
nand U12352 (N_12352,N_9646,N_9987);
and U12353 (N_12353,N_8840,N_10050);
nand U12354 (N_12354,N_10146,N_10222);
and U12355 (N_12355,N_9629,N_11402);
xnor U12356 (N_12356,N_11830,N_8424);
and U12357 (N_12357,N_10331,N_11444);
nor U12358 (N_12358,N_8083,N_8025);
nand U12359 (N_12359,N_10602,N_11670);
or U12360 (N_12360,N_9362,N_9614);
nand U12361 (N_12361,N_10710,N_8687);
or U12362 (N_12362,N_10888,N_9964);
or U12363 (N_12363,N_9468,N_9817);
and U12364 (N_12364,N_11098,N_10769);
nand U12365 (N_12365,N_8625,N_9708);
xor U12366 (N_12366,N_8459,N_8728);
nand U12367 (N_12367,N_10560,N_10827);
nand U12368 (N_12368,N_8620,N_9176);
and U12369 (N_12369,N_11186,N_10563);
and U12370 (N_12370,N_10049,N_10318);
nand U12371 (N_12371,N_11533,N_9158);
and U12372 (N_12372,N_10263,N_9928);
or U12373 (N_12373,N_10421,N_11844);
nor U12374 (N_12374,N_11707,N_11375);
or U12375 (N_12375,N_11440,N_9704);
nor U12376 (N_12376,N_9599,N_9820);
or U12377 (N_12377,N_8037,N_8048);
nor U12378 (N_12378,N_9113,N_8049);
nand U12379 (N_12379,N_10524,N_9540);
nand U12380 (N_12380,N_11437,N_10825);
and U12381 (N_12381,N_10798,N_9782);
xnor U12382 (N_12382,N_10391,N_11925);
or U12383 (N_12383,N_8194,N_10900);
and U12384 (N_12384,N_8719,N_10559);
nand U12385 (N_12385,N_11505,N_8536);
nor U12386 (N_12386,N_11967,N_9315);
nor U12387 (N_12387,N_11316,N_11585);
xnor U12388 (N_12388,N_8184,N_11976);
nor U12389 (N_12389,N_9106,N_8763);
nor U12390 (N_12390,N_8337,N_9933);
nand U12391 (N_12391,N_11453,N_8384);
or U12392 (N_12392,N_8264,N_11164);
nor U12393 (N_12393,N_11174,N_9386);
and U12394 (N_12394,N_8145,N_10870);
and U12395 (N_12395,N_8902,N_9390);
or U12396 (N_12396,N_9193,N_10680);
or U12397 (N_12397,N_10614,N_8714);
or U12398 (N_12398,N_10006,N_11251);
nand U12399 (N_12399,N_8152,N_11591);
xnor U12400 (N_12400,N_9399,N_8185);
and U12401 (N_12401,N_10007,N_8529);
or U12402 (N_12402,N_11574,N_11200);
or U12403 (N_12403,N_8106,N_8762);
nor U12404 (N_12404,N_8920,N_10536);
and U12405 (N_12405,N_10545,N_8873);
or U12406 (N_12406,N_9022,N_8128);
xnor U12407 (N_12407,N_9119,N_11851);
nor U12408 (N_12408,N_8518,N_10457);
nand U12409 (N_12409,N_11092,N_9898);
or U12410 (N_12410,N_11425,N_9497);
and U12411 (N_12411,N_11424,N_9032);
nor U12412 (N_12412,N_8613,N_10789);
nand U12413 (N_12413,N_9384,N_8669);
and U12414 (N_12414,N_10152,N_10204);
nor U12415 (N_12415,N_9908,N_9913);
or U12416 (N_12416,N_8487,N_8626);
xnor U12417 (N_12417,N_8132,N_11477);
nand U12418 (N_12418,N_10458,N_9882);
nor U12419 (N_12419,N_10142,N_11602);
nor U12420 (N_12420,N_9576,N_10359);
nand U12421 (N_12421,N_9325,N_8407);
xor U12422 (N_12422,N_8376,N_10989);
nor U12423 (N_12423,N_8889,N_8144);
or U12424 (N_12424,N_10625,N_10068);
nand U12425 (N_12425,N_9725,N_8978);
and U12426 (N_12426,N_9816,N_11139);
nor U12427 (N_12427,N_9283,N_9477);
xor U12428 (N_12428,N_10660,N_8178);
or U12429 (N_12429,N_10663,N_8323);
nor U12430 (N_12430,N_9379,N_10073);
or U12431 (N_12431,N_11518,N_9959);
nand U12432 (N_12432,N_10025,N_9790);
and U12433 (N_12433,N_10908,N_8125);
or U12434 (N_12434,N_8333,N_9929);
or U12435 (N_12435,N_10212,N_8026);
nand U12436 (N_12436,N_10689,N_11978);
xor U12437 (N_12437,N_10450,N_10492);
or U12438 (N_12438,N_10837,N_9593);
or U12439 (N_12439,N_10032,N_10232);
xor U12440 (N_12440,N_10709,N_11070);
nand U12441 (N_12441,N_8364,N_9655);
nor U12442 (N_12442,N_11893,N_9496);
nor U12443 (N_12443,N_9133,N_9584);
xor U12444 (N_12444,N_10011,N_9044);
nand U12445 (N_12445,N_9067,N_10451);
nor U12446 (N_12446,N_8439,N_11478);
and U12447 (N_12447,N_10988,N_11347);
xnor U12448 (N_12448,N_11039,N_8833);
nand U12449 (N_12449,N_10358,N_9008);
or U12450 (N_12450,N_9883,N_9623);
or U12451 (N_12451,N_8595,N_10199);
and U12452 (N_12452,N_8834,N_8621);
and U12453 (N_12453,N_8005,N_8148);
and U12454 (N_12454,N_11476,N_11504);
or U12455 (N_12455,N_8896,N_8677);
or U12456 (N_12456,N_8579,N_8707);
and U12457 (N_12457,N_11984,N_8543);
or U12458 (N_12458,N_11860,N_8230);
and U12459 (N_12459,N_9052,N_9818);
xnor U12460 (N_12460,N_8629,N_9701);
nand U12461 (N_12461,N_11959,N_10360);
and U12462 (N_12462,N_10306,N_10024);
or U12463 (N_12463,N_11364,N_10840);
and U12464 (N_12464,N_11685,N_9557);
or U12465 (N_12465,N_8532,N_10783);
xor U12466 (N_12466,N_9717,N_8658);
nand U12467 (N_12467,N_8313,N_10504);
or U12468 (N_12468,N_8042,N_11927);
nor U12469 (N_12469,N_8614,N_8235);
nand U12470 (N_12470,N_8590,N_11243);
or U12471 (N_12471,N_11315,N_11053);
or U12472 (N_12472,N_8782,N_8995);
and U12473 (N_12473,N_8113,N_11743);
and U12474 (N_12474,N_8350,N_8652);
and U12475 (N_12475,N_8501,N_9922);
nand U12476 (N_12476,N_9291,N_8222);
nor U12477 (N_12477,N_10513,N_9049);
and U12478 (N_12478,N_11502,N_8647);
or U12479 (N_12479,N_11689,N_9951);
nand U12480 (N_12480,N_10217,N_11542);
xnor U12481 (N_12481,N_8339,N_8517);
nand U12482 (N_12482,N_11419,N_10727);
xnor U12483 (N_12483,N_10397,N_9191);
nand U12484 (N_12484,N_11077,N_8086);
nand U12485 (N_12485,N_9983,N_11420);
or U12486 (N_12486,N_10196,N_9358);
and U12487 (N_12487,N_9890,N_10051);
or U12488 (N_12488,N_9825,N_8802);
nor U12489 (N_12489,N_8305,N_11346);
nor U12490 (N_12490,N_8195,N_8394);
nand U12491 (N_12491,N_11834,N_10116);
xnor U12492 (N_12492,N_9147,N_9500);
xor U12493 (N_12493,N_8512,N_10431);
and U12494 (N_12494,N_11744,N_11561);
nor U12495 (N_12495,N_11217,N_8711);
or U12496 (N_12496,N_10378,N_10268);
nand U12497 (N_12497,N_8910,N_11731);
nand U12498 (N_12498,N_11878,N_8615);
nand U12499 (N_12499,N_10087,N_10608);
and U12500 (N_12500,N_8701,N_11587);
nand U12501 (N_12501,N_8803,N_10721);
nand U12502 (N_12502,N_11580,N_11962);
nor U12503 (N_12503,N_10757,N_9018);
nor U12504 (N_12504,N_9472,N_9281);
nand U12505 (N_12505,N_10836,N_8330);
nand U12506 (N_12506,N_9985,N_10149);
xnor U12507 (N_12507,N_10466,N_8204);
and U12508 (N_12508,N_9401,N_8606);
nand U12509 (N_12509,N_11999,N_9843);
or U12510 (N_12510,N_10021,N_10387);
or U12511 (N_12511,N_10009,N_9163);
and U12512 (N_12512,N_10443,N_10079);
or U12513 (N_12513,N_10647,N_10903);
xnor U12514 (N_12514,N_10548,N_11264);
or U12515 (N_12515,N_9398,N_9915);
nor U12516 (N_12516,N_10479,N_11185);
and U12517 (N_12517,N_8189,N_9064);
or U12518 (N_12518,N_10676,N_9544);
nand U12519 (N_12519,N_10735,N_11642);
or U12520 (N_12520,N_8369,N_10482);
or U12521 (N_12521,N_9792,N_10249);
nand U12522 (N_12522,N_10161,N_8237);
and U12523 (N_12523,N_10897,N_11267);
nand U12524 (N_12524,N_10215,N_11599);
nand U12525 (N_12525,N_10230,N_8166);
nor U12526 (N_12526,N_9162,N_11983);
and U12527 (N_12527,N_11639,N_10223);
xnor U12528 (N_12528,N_9310,N_10118);
xnor U12529 (N_12529,N_8455,N_11612);
nand U12530 (N_12530,N_8510,N_9293);
nor U12531 (N_12531,N_9068,N_10998);
or U12532 (N_12532,N_8874,N_8467);
nand U12533 (N_12533,N_10860,N_11621);
and U12534 (N_12534,N_8463,N_11880);
nor U12535 (N_12535,N_11798,N_10613);
nand U12536 (N_12536,N_11028,N_9850);
nor U12537 (N_12537,N_11665,N_11886);
or U12538 (N_12538,N_10475,N_9001);
nand U12539 (N_12539,N_10892,N_8167);
xnor U12540 (N_12540,N_11708,N_9004);
nand U12541 (N_12541,N_10952,N_11582);
and U12542 (N_12542,N_11392,N_9902);
and U12543 (N_12543,N_10951,N_9178);
nor U12544 (N_12544,N_9918,N_11137);
and U12545 (N_12545,N_9694,N_11263);
nand U12546 (N_12546,N_8201,N_9622);
nor U12547 (N_12547,N_10367,N_11479);
and U12548 (N_12548,N_11408,N_9375);
nor U12549 (N_12549,N_8627,N_9131);
nand U12550 (N_12550,N_8796,N_11911);
xnor U12551 (N_12551,N_8068,N_11538);
nor U12552 (N_12552,N_11536,N_8483);
or U12553 (N_12553,N_10543,N_11679);
nand U12554 (N_12554,N_8771,N_9865);
nor U12555 (N_12555,N_9424,N_8143);
and U12556 (N_12556,N_8836,N_10753);
nand U12557 (N_12557,N_8058,N_10463);
and U12558 (N_12558,N_10734,N_11626);
nor U12559 (N_12559,N_11778,N_11240);
or U12560 (N_12560,N_9747,N_10356);
nand U12561 (N_12561,N_9301,N_10163);
nand U12562 (N_12562,N_8047,N_10325);
xnor U12563 (N_12563,N_11594,N_10157);
nor U12564 (N_12564,N_9169,N_9777);
nor U12565 (N_12565,N_9862,N_11385);
or U12566 (N_12566,N_9385,N_11741);
and U12567 (N_12567,N_8471,N_9549);
nand U12568 (N_12568,N_10203,N_11919);
xor U12569 (N_12569,N_10552,N_10366);
nand U12570 (N_12570,N_11196,N_9802);
nor U12571 (N_12571,N_11784,N_10975);
or U12572 (N_12572,N_11627,N_9916);
nand U12573 (N_12573,N_9548,N_10386);
nor U12574 (N_12574,N_9330,N_10626);
xor U12575 (N_12575,N_9712,N_9336);
or U12576 (N_12576,N_9932,N_11586);
nand U12577 (N_12577,N_8038,N_9719);
and U12578 (N_12578,N_11396,N_8254);
and U12579 (N_12579,N_8561,N_9442);
xor U12580 (N_12580,N_9770,N_10937);
or U12581 (N_12581,N_8944,N_10088);
or U12582 (N_12582,N_9624,N_11314);
or U12583 (N_12583,N_11080,N_8465);
nand U12584 (N_12584,N_9139,N_11190);
or U12585 (N_12585,N_9998,N_8604);
nor U12586 (N_12586,N_8322,N_11008);
xor U12587 (N_12587,N_8898,N_10767);
nor U12588 (N_12588,N_11970,N_8197);
or U12589 (N_12589,N_9531,N_10730);
or U12590 (N_12590,N_10119,N_11812);
and U12591 (N_12591,N_10407,N_11088);
nor U12592 (N_12592,N_8733,N_10969);
or U12593 (N_12593,N_9436,N_11633);
nand U12594 (N_12594,N_9335,N_9365);
nand U12595 (N_12595,N_10506,N_8958);
and U12596 (N_12596,N_8014,N_8084);
nor U12597 (N_12597,N_8395,N_11929);
or U12598 (N_12598,N_8371,N_10201);
and U12599 (N_12599,N_8586,N_10785);
nand U12600 (N_12600,N_8700,N_9804);
nor U12601 (N_12601,N_11732,N_9848);
nor U12602 (N_12602,N_8645,N_10934);
or U12603 (N_12603,N_9668,N_11333);
nor U12604 (N_12604,N_9216,N_11339);
nor U12605 (N_12605,N_10540,N_8500);
xor U12606 (N_12606,N_11059,N_11156);
and U12607 (N_12607,N_11279,N_11728);
or U12608 (N_12608,N_9567,N_8783);
and U12609 (N_12609,N_10427,N_9420);
nand U12610 (N_12610,N_9486,N_11473);
or U12611 (N_12611,N_11142,N_11775);
nand U12612 (N_12612,N_10907,N_10630);
nor U12613 (N_12613,N_8373,N_10715);
and U12614 (N_12614,N_9763,N_9996);
and U12615 (N_12615,N_9110,N_9316);
and U12616 (N_12616,N_10052,N_8770);
and U12617 (N_12617,N_9992,N_9821);
nor U12618 (N_12618,N_11794,N_10419);
nor U12619 (N_12619,N_8480,N_11353);
or U12620 (N_12620,N_10640,N_10526);
and U12621 (N_12621,N_10635,N_11064);
or U12622 (N_12622,N_10500,N_9604);
or U12623 (N_12623,N_8726,N_10089);
xor U12624 (N_12624,N_8232,N_11712);
xor U12625 (N_12625,N_9051,N_8895);
nand U12626 (N_12626,N_11103,N_9534);
nand U12627 (N_12627,N_11105,N_11724);
or U12628 (N_12628,N_8565,N_9189);
nor U12629 (N_12629,N_10235,N_8537);
or U12630 (N_12630,N_8080,N_9461);
or U12631 (N_12631,N_11868,N_11108);
and U12632 (N_12632,N_8224,N_9366);
xor U12633 (N_12633,N_10130,N_9125);
or U12634 (N_12634,N_9263,N_8868);
and U12635 (N_12635,N_8206,N_9207);
nand U12636 (N_12636,N_11172,N_11589);
nand U12637 (N_12637,N_11802,N_8720);
xor U12638 (N_12638,N_9729,N_8973);
nand U12639 (N_12639,N_10523,N_10405);
nand U12640 (N_12640,N_9633,N_11964);
and U12641 (N_12641,N_10095,N_9801);
nor U12642 (N_12642,N_10705,N_11363);
and U12643 (N_12643,N_11018,N_11035);
nand U12644 (N_12644,N_9784,N_11843);
nand U12645 (N_12645,N_11720,N_11133);
xor U12646 (N_12646,N_9023,N_9115);
xor U12647 (N_12647,N_10847,N_11226);
nor U12648 (N_12648,N_10866,N_9710);
nand U12649 (N_12649,N_9598,N_11150);
or U12650 (N_12650,N_8256,N_9080);
or U12651 (N_12651,N_8571,N_8799);
and U12652 (N_12652,N_10874,N_11813);
nor U12653 (N_12653,N_8199,N_10502);
xor U12654 (N_12654,N_10452,N_9381);
xor U12655 (N_12655,N_10172,N_10147);
nand U12656 (N_12656,N_10982,N_9656);
nand U12657 (N_12657,N_8693,N_10234);
nor U12658 (N_12658,N_10373,N_9100);
nor U12659 (N_12659,N_11252,N_8545);
nor U12660 (N_12660,N_8137,N_8742);
and U12661 (N_12661,N_9416,N_8641);
or U12662 (N_12662,N_8541,N_10417);
nor U12663 (N_12663,N_11740,N_11330);
and U12664 (N_12664,N_11949,N_9075);
nor U12665 (N_12665,N_10842,N_9426);
xnor U12666 (N_12666,N_11393,N_8215);
nor U12667 (N_12667,N_8282,N_8338);
nand U12668 (N_12668,N_11715,N_9601);
nand U12669 (N_12669,N_10193,N_11645);
and U12670 (N_12670,N_10341,N_11753);
nor U12671 (N_12671,N_11620,N_11609);
xor U12672 (N_12672,N_11898,N_9741);
or U12673 (N_12673,N_11848,N_9896);
nand U12674 (N_12674,N_10381,N_11302);
and U12675 (N_12675,N_8285,N_11056);
or U12676 (N_12676,N_9610,N_9515);
nor U12677 (N_12677,N_10401,N_11492);
and U12678 (N_12678,N_8396,N_11810);
nand U12679 (N_12679,N_8831,N_8129);
nand U12680 (N_12680,N_11303,N_11604);
nand U12681 (N_12681,N_8023,N_11563);
nand U12682 (N_12682,N_11950,N_8856);
or U12683 (N_12683,N_9282,N_11311);
xnor U12684 (N_12684,N_9209,N_9521);
and U12685 (N_12685,N_9454,N_8095);
or U12686 (N_12686,N_11781,N_9556);
and U12687 (N_12687,N_8897,N_11669);
xnor U12688 (N_12688,N_9261,N_11829);
and U12689 (N_12689,N_9447,N_9005);
or U12690 (N_12690,N_11294,N_9303);
or U12691 (N_12691,N_9393,N_11947);
or U12692 (N_12692,N_10628,N_9608);
nor U12693 (N_12693,N_10801,N_8918);
xnor U12694 (N_12694,N_11170,N_10733);
or U12695 (N_12695,N_9084,N_9632);
and U12696 (N_12696,N_11904,N_9343);
or U12697 (N_12697,N_10330,N_10180);
nand U12698 (N_12698,N_9724,N_11265);
nand U12699 (N_12699,N_10708,N_10287);
or U12700 (N_12700,N_10357,N_10036);
nor U12701 (N_12701,N_10375,N_8410);
nand U12702 (N_12702,N_10102,N_10002);
xor U12703 (N_12703,N_9259,N_9295);
and U12704 (N_12704,N_11276,N_10541);
nor U12705 (N_12705,N_9214,N_10624);
nand U12706 (N_12706,N_10184,N_11266);
or U12707 (N_12707,N_8318,N_8787);
nor U12708 (N_12708,N_8659,N_9835);
and U12709 (N_12709,N_8976,N_8655);
or U12710 (N_12710,N_9732,N_11651);
xor U12711 (N_12711,N_10616,N_11350);
nand U12712 (N_12712,N_10074,N_10669);
nand U12713 (N_12713,N_9581,N_9606);
or U12714 (N_12714,N_8734,N_11373);
nor U12715 (N_12715,N_8838,N_10813);
or U12716 (N_12716,N_8397,N_9662);
xor U12717 (N_12717,N_11750,N_8846);
nand U12718 (N_12718,N_9383,N_8775);
and U12719 (N_12719,N_8102,N_9768);
nand U12720 (N_12720,N_11114,N_10107);
or U12721 (N_12721,N_10867,N_11500);
and U12722 (N_12722,N_11635,N_9144);
or U12723 (N_12723,N_9351,N_9839);
xor U12724 (N_12724,N_9480,N_11646);
nor U12725 (N_12725,N_8028,N_11113);
xnor U12726 (N_12726,N_11435,N_8651);
nand U12727 (N_12727,N_11166,N_10469);
and U12728 (N_12728,N_9161,N_8359);
or U12729 (N_12729,N_11855,N_11837);
xnor U12730 (N_12730,N_9050,N_9884);
nand U12731 (N_12731,N_8923,N_8962);
nor U12732 (N_12732,N_11628,N_11237);
nor U12733 (N_12733,N_10335,N_9751);
or U12734 (N_12734,N_8097,N_10665);
and U12735 (N_12735,N_8622,N_9221);
nor U12736 (N_12736,N_10674,N_10583);
and U12737 (N_12737,N_8120,N_10126);
or U12738 (N_12738,N_10448,N_9002);
nand U12739 (N_12739,N_8891,N_9332);
nand U12740 (N_12740,N_11624,N_10332);
nand U12741 (N_12741,N_10363,N_11097);
or U12742 (N_12742,N_9095,N_9618);
and U12743 (N_12743,N_8245,N_8696);
xor U12744 (N_12744,N_11280,N_10441);
nand U12745 (N_12745,N_8009,N_10601);
nand U12746 (N_12746,N_11871,N_11852);
nand U12747 (N_12747,N_9153,N_11549);
and U12748 (N_12748,N_9079,N_9575);
nand U12749 (N_12749,N_10278,N_8094);
nor U12750 (N_12750,N_8306,N_9641);
nor U12751 (N_12751,N_11838,N_8725);
xnor U12752 (N_12752,N_8485,N_8150);
and U12753 (N_12753,N_10020,N_8723);
and U12754 (N_12754,N_9120,N_10898);
or U12755 (N_12755,N_8283,N_11357);
nor U12756 (N_12756,N_8470,N_10376);
nor U12757 (N_12757,N_10270,N_8888);
nand U12758 (N_12758,N_9164,N_8555);
and U12759 (N_12759,N_11019,N_8764);
nand U12760 (N_12760,N_11427,N_9484);
and U12761 (N_12761,N_9047,N_11312);
nand U12762 (N_12762,N_8666,N_8535);
and U12763 (N_12763,N_8854,N_11571);
nor U12764 (N_12764,N_11049,N_11205);
nand U12765 (N_12765,N_11051,N_9785);
or U12766 (N_12766,N_11487,N_11818);
nand U12767 (N_12767,N_10700,N_9752);
or U12768 (N_12768,N_9543,N_8524);
xnor U12769 (N_12769,N_11643,N_10759);
or U12770 (N_12770,N_9327,N_10078);
xor U12771 (N_12771,N_9225,N_9635);
nor U12772 (N_12772,N_9594,N_8746);
xnor U12773 (N_12773,N_8526,N_9634);
xor U12774 (N_12774,N_8168,N_9273);
nand U12775 (N_12775,N_8506,N_8801);
and U12776 (N_12776,N_11671,N_8383);
or U12777 (N_12777,N_11617,N_9208);
nand U12778 (N_12778,N_9529,N_11562);
and U12779 (N_12779,N_11699,N_8377);
nand U12780 (N_12780,N_11552,N_8759);
and U12781 (N_12781,N_10751,N_9232);
and U12782 (N_12782,N_11254,N_10586);
or U12783 (N_12783,N_9308,N_9413);
nand U12784 (N_12784,N_10496,N_8303);
and U12785 (N_12785,N_8110,N_8816);
nor U12786 (N_12786,N_8716,N_8709);
and U12787 (N_12787,N_9445,N_9433);
and U12788 (N_12788,N_11158,N_9089);
nor U12789 (N_12789,N_11134,N_10527);
xor U12790 (N_12790,N_10773,N_11652);
nand U12791 (N_12791,N_8871,N_8414);
or U12792 (N_12792,N_8900,N_9349);
and U12793 (N_12793,N_9149,N_11138);
xor U12794 (N_12794,N_9972,N_9458);
and U12795 (N_12795,N_8327,N_11795);
nor U12796 (N_12796,N_11509,N_8010);
or U12797 (N_12797,N_10323,N_9010);
nand U12798 (N_12798,N_10570,N_11145);
xnor U12799 (N_12799,N_11155,N_8123);
xor U12800 (N_12800,N_9995,N_8018);
nor U12801 (N_12801,N_10922,N_10776);
and U12802 (N_12802,N_11592,N_8814);
or U12803 (N_12803,N_11762,N_8752);
or U12804 (N_12804,N_10926,N_11508);
nor U12805 (N_12805,N_10516,N_9649);
or U12806 (N_12806,N_8903,N_8941);
and U12807 (N_12807,N_9762,N_11821);
nand U12808 (N_12808,N_10670,N_10296);
or U12809 (N_12809,N_11748,N_10679);
and U12810 (N_12810,N_9145,N_8479);
nor U12811 (N_12811,N_10175,N_8671);
and U12812 (N_12812,N_11735,N_11460);
nand U12813 (N_12813,N_9905,N_11202);
and U12814 (N_12814,N_11406,N_9483);
nor U12815 (N_12815,N_9346,N_8334);
nand U12816 (N_12816,N_9997,N_11684);
or U12817 (N_12817,N_11700,N_10444);
and U12818 (N_12818,N_9591,N_9233);
and U12819 (N_12819,N_10420,N_10098);
or U12820 (N_12820,N_11175,N_8452);
or U12821 (N_12821,N_8618,N_8064);
nor U12822 (N_12822,N_9244,N_9441);
or U12823 (N_12823,N_11981,N_9071);
nor U12824 (N_12824,N_8328,N_9482);
xor U12825 (N_12825,N_10247,N_8530);
nand U12826 (N_12826,N_11273,N_10174);
nand U12827 (N_12827,N_11079,N_8073);
nor U12828 (N_12828,N_8119,N_10422);
and U12829 (N_12829,N_10865,N_9187);
xor U12830 (N_12830,N_11814,N_10578);
xor U12831 (N_12831,N_9666,N_10873);
or U12832 (N_12832,N_11926,N_11547);
nor U12833 (N_12833,N_9759,N_8997);
and U12834 (N_12834,N_10606,N_9677);
or U12835 (N_12835,N_9469,N_10919);
and U12836 (N_12836,N_9891,N_10494);
and U12837 (N_12837,N_10094,N_8175);
nor U12838 (N_12838,N_11945,N_9737);
nor U12839 (N_12839,N_9083,N_10377);
nor U12840 (N_12840,N_8839,N_11071);
and U12841 (N_12841,N_10995,N_11494);
nand U12842 (N_12842,N_9558,N_8913);
nor U12843 (N_12843,N_11034,N_8041);
nor U12844 (N_12844,N_10909,N_10085);
or U12845 (N_12845,N_8504,N_8093);
nand U12846 (N_12846,N_10862,N_8220);
xor U12847 (N_12847,N_11941,N_8079);
xor U12848 (N_12848,N_10293,N_9309);
nor U12849 (N_12849,N_11278,N_9279);
or U12850 (N_12850,N_10505,N_8398);
and U12851 (N_12851,N_8637,N_10593);
nand U12852 (N_12852,N_9639,N_8172);
nor U12853 (N_12853,N_9337,N_9154);
nand U12854 (N_12854,N_10008,N_8375);
or U12855 (N_12855,N_8013,N_10720);
xnor U12856 (N_12856,N_10176,N_9367);
or U12857 (N_12857,N_10105,N_10979);
nor U12858 (N_12858,N_11301,N_11955);
and U12859 (N_12859,N_8050,N_8077);
or U12860 (N_12860,N_11567,N_11177);
or U12861 (N_12861,N_8289,N_9451);
nand U12862 (N_12862,N_11632,N_9298);
nand U12863 (N_12863,N_8912,N_8278);
or U12864 (N_12864,N_11579,N_10242);
nor U12865 (N_12865,N_8234,N_9667);
xor U12866 (N_12866,N_8286,N_9970);
or U12867 (N_12867,N_9136,N_10698);
or U12868 (N_12868,N_11409,N_11569);
xnor U12869 (N_12869,N_11006,N_8248);
xor U12870 (N_12870,N_8527,N_11923);
nor U12871 (N_12871,N_10462,N_11992);
nand U12872 (N_12872,N_8957,N_9706);
nand U12873 (N_12873,N_11811,N_10055);
nor U12874 (N_12874,N_10258,N_10652);
or U12875 (N_12875,N_10402,N_9355);
or U12876 (N_12876,N_9460,N_8109);
nor U12877 (N_12877,N_11882,N_11666);
or U12878 (N_12878,N_10528,N_10885);
nor U12879 (N_12879,N_9212,N_9368);
and U12880 (N_12880,N_8569,N_11548);
xnor U12881 (N_12881,N_8329,N_10931);
and U12882 (N_12882,N_11397,N_8310);
xnor U12883 (N_12883,N_8815,N_11027);
and U12884 (N_12884,N_8272,N_9081);
and U12885 (N_12885,N_8926,N_11445);
nand U12886 (N_12886,N_9698,N_11823);
nor U12887 (N_12887,N_11935,N_10534);
nor U12888 (N_12888,N_10929,N_11386);
and U12889 (N_12889,N_9627,N_9143);
nand U12890 (N_12890,N_9190,N_8691);
or U12891 (N_12891,N_9855,N_11358);
and U12892 (N_12892,N_9076,N_8063);
or U12893 (N_12893,N_8458,N_8562);
or U12894 (N_12894,N_9948,N_9198);
nand U12895 (N_12895,N_8639,N_8497);
and U12896 (N_12896,N_11716,N_9512);
and U12897 (N_12897,N_11678,N_11564);
nor U12898 (N_12898,N_10877,N_8929);
nor U12899 (N_12899,N_8538,N_11157);
nor U12900 (N_12900,N_10225,N_9170);
nand U12901 (N_12901,N_10831,N_9806);
or U12902 (N_12902,N_10609,N_8391);
nor U12903 (N_12903,N_11737,N_10571);
or U12904 (N_12904,N_11636,N_11236);
xnor U12905 (N_12905,N_10259,N_9062);
nor U12906 (N_12906,N_10749,N_9899);
nand U12907 (N_12907,N_8060,N_9434);
nor U12908 (N_12908,N_8091,N_10231);
or U12909 (N_12909,N_9934,N_10902);
nor U12910 (N_12910,N_8078,N_9440);
or U12911 (N_12911,N_8345,N_11282);
xor U12912 (N_12912,N_8580,N_10246);
nand U12913 (N_12913,N_10592,N_10744);
nor U12914 (N_12914,N_9682,N_11662);
nand U12915 (N_12915,N_8611,N_11786);
and U12916 (N_12916,N_10623,N_11881);
or U12917 (N_12917,N_9742,N_11771);
and U12918 (N_12918,N_9150,N_11331);
nor U12919 (N_12919,N_9344,N_9302);
nand U12920 (N_12920,N_9495,N_9756);
nand U12921 (N_12921,N_9595,N_8162);
nand U12922 (N_12922,N_10438,N_8712);
nor U12923 (N_12923,N_11833,N_9781);
nand U12924 (N_12924,N_9129,N_9446);
nand U12925 (N_12925,N_8566,N_9459);
nand U12926 (N_12926,N_10643,N_9502);
nor U12927 (N_12927,N_8552,N_11951);
or U12928 (N_12928,N_8676,N_11163);
and U12929 (N_12929,N_8435,N_11751);
or U12930 (N_12930,N_11456,N_9566);
nand U12931 (N_12931,N_11160,N_9396);
nand U12932 (N_12932,N_11261,N_8071);
or U12933 (N_12933,N_8956,N_9536);
and U12934 (N_12934,N_8429,N_9088);
nand U12935 (N_12935,N_8428,N_9319);
or U12936 (N_12936,N_8008,N_10198);
or U12937 (N_12937,N_11584,N_9338);
nor U12938 (N_12938,N_11746,N_9000);
and U12939 (N_12939,N_8630,N_8382);
or U12940 (N_12940,N_10281,N_8950);
and U12941 (N_12941,N_11876,N_10301);
xor U12942 (N_12942,N_11913,N_11429);
and U12943 (N_12943,N_8975,N_9427);
and U12944 (N_12944,N_10600,N_9776);
nor U12945 (N_12945,N_8591,N_11211);
or U12946 (N_12946,N_10886,N_8758);
nand U12947 (N_12947,N_9142,N_11835);
or U12948 (N_12948,N_11120,N_10316);
and U12949 (N_12949,N_9226,N_10045);
or U12950 (N_12950,N_11293,N_11595);
or U12951 (N_12951,N_9415,N_11329);
nand U12952 (N_12952,N_8433,N_8349);
nand U12953 (N_12953,N_8938,N_9718);
nand U12954 (N_12954,N_10517,N_10291);
nand U12955 (N_12955,N_8290,N_10264);
nor U12956 (N_12956,N_10765,N_10160);
xor U12957 (N_12957,N_11777,N_11727);
xnor U12958 (N_12958,N_8461,N_8879);
or U12959 (N_12959,N_10955,N_10190);
xor U12960 (N_12960,N_10046,N_10997);
nor U12961 (N_12961,N_10015,N_11758);
xor U12962 (N_12962,N_11858,N_9823);
and U12963 (N_12963,N_8514,N_10950);
nor U12964 (N_12964,N_10693,N_8017);
or U12965 (N_12965,N_9935,N_10990);
and U12966 (N_12966,N_11756,N_9827);
nor U12967 (N_12967,N_10226,N_11428);
or U12968 (N_12968,N_8951,N_9274);
or U12969 (N_12969,N_10770,N_11125);
nor U12970 (N_12970,N_11815,N_9324);
or U12971 (N_12971,N_8488,N_11570);
nand U12972 (N_12972,N_9146,N_9730);
xnor U12973 (N_12973,N_9276,N_10012);
or U12974 (N_12974,N_11663,N_9251);
nor U12975 (N_12975,N_11001,N_11274);
xnor U12976 (N_12976,N_10022,N_8934);
and U12977 (N_12977,N_9523,N_8948);
and U12978 (N_12978,N_9693,N_8955);
or U12979 (N_12979,N_8190,N_9684);
nand U12980 (N_12980,N_8784,N_11167);
nand U12981 (N_12981,N_10266,N_8255);
xor U12982 (N_12982,N_11757,N_10607);
and U12983 (N_12983,N_10162,N_9690);
and U12984 (N_12984,N_10454,N_10725);
nor U12985 (N_12985,N_8031,N_8609);
and U12986 (N_12986,N_10632,N_10802);
and U12987 (N_12987,N_10646,N_11529);
or U12988 (N_12988,N_8791,N_9738);
nand U12989 (N_12989,N_9456,N_9307);
or U12990 (N_12990,N_8210,N_10971);
nand U12991 (N_12991,N_11462,N_11634);
nand U12992 (N_12992,N_8016,N_8100);
and U12993 (N_12993,N_10211,N_8638);
and U12994 (N_12994,N_9289,N_11387);
and U12995 (N_12995,N_8478,N_8004);
and U12996 (N_12996,N_9430,N_8755);
or U12997 (N_12997,N_9947,N_11065);
or U12998 (N_12998,N_11395,N_11686);
nor U12999 (N_12999,N_11495,N_11975);
xnor U13000 (N_13000,N_10804,N_11376);
nor U13001 (N_13001,N_10272,N_9326);
nand U13002 (N_13002,N_9092,N_8213);
xnor U13003 (N_13003,N_9809,N_10539);
and U13004 (N_13004,N_8200,N_10793);
nor U13005 (N_13005,N_8174,N_10594);
nor U13006 (N_13006,N_10591,N_10224);
nor U13007 (N_13007,N_8680,N_11768);
nor U13008 (N_13008,N_10307,N_11206);
or U13009 (N_13009,N_10761,N_8228);
xor U13010 (N_13010,N_11826,N_9609);
nand U13011 (N_13011,N_10940,N_9165);
nor U13012 (N_13012,N_11767,N_11042);
or U13013 (N_13013,N_8218,N_10308);
or U13014 (N_13014,N_10300,N_10739);
and U13015 (N_13015,N_11232,N_9267);
nor U13016 (N_13016,N_9605,N_9888);
nor U13017 (N_13017,N_9397,N_8681);
nand U13018 (N_13018,N_9518,N_8280);
xor U13019 (N_13019,N_10137,N_10731);
nand U13020 (N_13020,N_9625,N_11747);
nand U13021 (N_13021,N_11075,N_11480);
or U13022 (N_13022,N_9342,N_9881);
xor U13023 (N_13023,N_8462,N_9588);
and U13024 (N_13024,N_8296,N_8427);
and U13025 (N_13025,N_11281,N_8133);
or U13026 (N_13026,N_9731,N_10945);
and U13027 (N_13027,N_11776,N_11401);
nor U13028 (N_13028,N_8300,N_10992);
and U13029 (N_13029,N_10013,N_8852);
and U13030 (N_13030,N_11825,N_11499);
nor U13031 (N_13031,N_8164,N_11021);
and U13032 (N_13032,N_10241,N_8308);
or U13033 (N_13033,N_11284,N_8288);
or U13034 (N_13034,N_11850,N_9408);
or U13035 (N_13035,N_10510,N_8312);
nand U13036 (N_13036,N_8494,N_10334);
and U13037 (N_13037,N_10695,N_11806);
or U13038 (N_13038,N_10352,N_9063);
or U13039 (N_13039,N_10275,N_10771);
nor U13040 (N_13040,N_8372,N_11979);
xor U13041 (N_13041,N_9159,N_9620);
or U13042 (N_13042,N_8736,N_11140);
xor U13043 (N_13043,N_9389,N_11112);
or U13044 (N_13044,N_11832,N_9873);
and U13045 (N_13045,N_8605,N_8015);
and U13046 (N_13046,N_9761,N_9213);
nand U13047 (N_13047,N_10065,N_10177);
nand U13048 (N_13048,N_11896,N_10097);
and U13049 (N_13049,N_10123,N_10752);
nor U13050 (N_13050,N_11824,N_8985);
nand U13051 (N_13051,N_11277,N_11043);
nor U13052 (N_13052,N_8482,N_11345);
xor U13053 (N_13053,N_10826,N_8474);
nor U13054 (N_13054,N_9859,N_8291);
xor U13055 (N_13055,N_8739,N_10305);
and U13056 (N_13056,N_10828,N_10311);
and U13057 (N_13057,N_10895,N_8735);
nor U13058 (N_13058,N_9926,N_8315);
nand U13059 (N_13059,N_10964,N_10329);
or U13060 (N_13060,N_11526,N_10250);
nor U13061 (N_13061,N_11439,N_8196);
nor U13062 (N_13062,N_10171,N_8343);
nor U13063 (N_13063,N_9288,N_11101);
xnor U13064 (N_13064,N_11102,N_11151);
nor U13065 (N_13065,N_11149,N_9858);
or U13066 (N_13066,N_9069,N_8208);
nand U13067 (N_13067,N_10942,N_10687);
or U13068 (N_13068,N_11884,N_10342);
and U13069 (N_13069,N_9464,N_10799);
xor U13070 (N_13070,N_11116,N_10968);
nor U13071 (N_13071,N_11761,N_9160);
nor U13072 (N_13072,N_11897,N_9021);
or U13073 (N_13073,N_10181,N_9470);
and U13074 (N_13074,N_10525,N_8684);
nand U13075 (N_13075,N_11847,N_9012);
and U13076 (N_13076,N_11694,N_11288);
nor U13077 (N_13077,N_11554,N_11917);
or U13078 (N_13078,N_9524,N_10713);
nor U13079 (N_13079,N_11176,N_8107);
or U13080 (N_13080,N_11903,N_8643);
and U13081 (N_13081,N_10465,N_9220);
or U13082 (N_13082,N_10661,N_11272);
nor U13083 (N_13083,N_8240,N_8363);
nand U13084 (N_13084,N_11258,N_11940);
and U13085 (N_13085,N_8964,N_11084);
nand U13086 (N_13086,N_8243,N_10120);
xnor U13087 (N_13087,N_11920,N_11322);
and U13088 (N_13088,N_10128,N_10077);
nor U13089 (N_13089,N_11905,N_9665);
nor U13090 (N_13090,N_8827,N_9851);
nand U13091 (N_13091,N_8032,N_8539);
xor U13092 (N_13092,N_9727,N_11734);
and U13093 (N_13093,N_11931,N_11352);
nor U13094 (N_13094,N_11464,N_8161);
or U13095 (N_13095,N_11054,N_8921);
or U13096 (N_13096,N_11063,N_11991);
nand U13097 (N_13097,N_11924,N_11317);
xnor U13098 (N_13098,N_8818,N_9364);
nand U13099 (N_13099,N_10574,N_10111);
nor U13100 (N_13100,N_8689,N_11551);
nor U13101 (N_13101,N_8777,N_11998);
nor U13102 (N_13102,N_8416,N_9138);
or U13103 (N_13103,N_10276,N_9642);
xor U13104 (N_13104,N_8557,N_10484);
nor U13105 (N_13105,N_11631,N_8919);
and U13106 (N_13106,N_11342,N_9921);
nand U13107 (N_13107,N_10963,N_8304);
or U13108 (N_13108,N_8654,N_8792);
or U13109 (N_13109,N_11960,N_9880);
xor U13110 (N_13110,N_11558,N_11458);
and U13111 (N_13111,N_10136,N_8883);
or U13112 (N_13112,N_9376,N_9025);
nor U13113 (N_13113,N_10561,N_11060);
and U13114 (N_13114,N_8307,N_9692);
nand U13115 (N_13115,N_8438,N_11891);
or U13116 (N_13116,N_8131,N_9705);
nor U13117 (N_13117,N_10875,N_10114);
and U13118 (N_13118,N_10724,N_11859);
or U13119 (N_13119,N_8317,N_8055);
or U13120 (N_13120,N_8368,N_8126);
nand U13121 (N_13121,N_10993,N_10808);
xor U13122 (N_13122,N_10852,N_8251);
nor U13123 (N_13123,N_10158,N_9778);
nand U13124 (N_13124,N_8632,N_10132);
and U13125 (N_13125,N_10283,N_11005);
or U13126 (N_13126,N_9406,N_9492);
nor U13127 (N_13127,N_8697,N_11963);
nand U13128 (N_13128,N_11512,N_8374);
xnor U13129 (N_13129,N_11422,N_9210);
nand U13130 (N_13130,N_10581,N_11760);
nor U13131 (N_13131,N_8924,N_8238);
nand U13132 (N_13132,N_11147,N_8859);
or U13133 (N_13133,N_11040,N_11828);
nand U13134 (N_13134,N_11472,N_8880);
nor U13135 (N_13135,N_11275,N_8660);
and U13136 (N_13136,N_10014,N_11488);
nand U13137 (N_13137,N_9991,N_10456);
xnor U13138 (N_13138,N_11389,N_8996);
nand U13139 (N_13139,N_10706,N_8274);
and U13140 (N_13140,N_10298,N_11384);
or U13141 (N_13141,N_11126,N_9329);
and U13142 (N_13142,N_9695,N_10245);
nand U13143 (N_13143,N_11135,N_11404);
nor U13144 (N_13144,N_11199,N_9711);
or U13145 (N_13145,N_10650,N_11256);
nand U13146 (N_13146,N_10092,N_10238);
nand U13147 (N_13147,N_9055,N_8103);
and U13148 (N_13148,N_10058,N_11939);
or U13149 (N_13149,N_8509,N_8662);
nor U13150 (N_13150,N_9269,N_8906);
or U13151 (N_13151,N_11090,N_8617);
and U13152 (N_13152,N_11050,N_8165);
and U13153 (N_13153,N_11359,N_11698);
nor U13154 (N_13154,N_8503,N_11475);
nand U13155 (N_13155,N_9255,N_10745);
nand U13156 (N_13156,N_8065,N_8519);
or U13157 (N_13157,N_11723,N_10071);
nand U13158 (N_13158,N_10507,N_8380);
and U13159 (N_13159,N_8610,N_8127);
nand U13160 (N_13160,N_9239,N_10351);
nand U13161 (N_13161,N_10598,N_8421);
nand U13162 (N_13162,N_11654,N_10717);
xnor U13163 (N_13163,N_9613,N_10038);
nand U13164 (N_13164,N_8794,N_8937);
nand U13165 (N_13165,N_10467,N_9354);
xnor U13166 (N_13166,N_9962,N_11953);
nor U13167 (N_13167,N_9003,N_9314);
or U13168 (N_13168,N_8299,N_10787);
xor U13169 (N_13169,N_9371,N_10535);
and U13170 (N_13170,N_8578,N_10946);
nand U13171 (N_13171,N_10214,N_8842);
nor U13172 (N_13172,N_8704,N_8940);
and U13173 (N_13173,N_11230,N_8432);
nor U13174 (N_13174,N_9854,N_11291);
or U13175 (N_13175,N_9828,N_10729);
xor U13176 (N_13176,N_9179,N_10863);
nor U13177 (N_13177,N_10649,N_11875);
and U13178 (N_13178,N_8528,N_10478);
nand U13179 (N_13179,N_10354,N_8425);
nor U13180 (N_13180,N_10228,N_10986);
nor U13181 (N_13181,N_9317,N_9102);
and U13182 (N_13182,N_9800,N_9958);
or U13183 (N_13183,N_11936,N_10449);
and U13184 (N_13184,N_11785,N_8585);
nor U13185 (N_13185,N_8729,N_9740);
and U13186 (N_13186,N_8341,N_9294);
xnor U13187 (N_13187,N_10447,N_9038);
or U13188 (N_13188,N_10562,N_10796);
or U13189 (N_13189,N_11430,N_10617);
nor U13190 (N_13190,N_10807,N_11958);
nor U13191 (N_13191,N_9230,N_10310);
or U13192 (N_13192,N_11058,N_11209);
xor U13193 (N_13193,N_11764,N_8988);
and U13194 (N_13194,N_8456,N_11706);
and U13195 (N_13195,N_11242,N_8656);
or U13196 (N_13196,N_11037,N_9636);
nor U13197 (N_13197,N_8813,N_9222);
or U13198 (N_13198,N_8939,N_9953);
and U13199 (N_13199,N_11630,N_9561);
and U13200 (N_13200,N_11044,N_9670);
nor U13201 (N_13201,N_9019,N_8221);
nand U13202 (N_13202,N_11233,N_9735);
or U13203 (N_13203,N_10683,N_9402);
nand U13204 (N_13204,N_8515,N_11618);
nor U13205 (N_13205,N_8992,N_11136);
nand U13206 (N_13206,N_11840,N_11921);
nand U13207 (N_13207,N_9114,N_8225);
and U13208 (N_13208,N_8804,N_9769);
and U13209 (N_13209,N_8845,N_8877);
and U13210 (N_13210,N_11539,N_9192);
and U13211 (N_13211,N_11067,N_11800);
nor U13212 (N_13212,N_11696,N_8052);
or U13213 (N_13213,N_10758,N_8105);
nor U13214 (N_13214,N_8114,N_11995);
xor U13215 (N_13215,N_10314,N_9321);
nand U13216 (N_13216,N_9505,N_8544);
nand U13217 (N_13217,N_10740,N_9669);
or U13218 (N_13218,N_8649,N_9265);
xnor U13219 (N_13219,N_8558,N_8045);
and U13220 (N_13220,N_10429,N_10297);
nor U13221 (N_13221,N_8882,N_10621);
and U13222 (N_13222,N_11517,N_9966);
nand U13223 (N_13223,N_10915,N_10815);
and U13224 (N_13224,N_9438,N_10970);
or U13225 (N_13225,N_8388,N_10538);
and U13226 (N_13226,N_8358,N_10823);
and U13227 (N_13227,N_8293,N_11269);
xor U13228 (N_13228,N_8451,N_8779);
xnor U13229 (N_13229,N_8863,N_11344);
nor U13230 (N_13230,N_10353,N_10490);
or U13231 (N_13231,N_10090,N_11327);
xnor U13232 (N_13232,N_9174,N_11031);
or U13233 (N_13233,N_11968,N_11041);
and U13234 (N_13234,N_11779,N_10704);
or U13235 (N_13235,N_8298,N_9123);
or U13236 (N_13236,N_11371,N_10430);
nand U13237 (N_13237,N_11299,N_10775);
and U13238 (N_13238,N_10299,N_8088);
xor U13239 (N_13239,N_8385,N_10711);
nand U13240 (N_13240,N_9982,N_11908);
xor U13241 (N_13241,N_11763,N_8362);
or U13242 (N_13242,N_9040,N_9009);
nand U13243 (N_13243,N_10682,N_10368);
or U13244 (N_13244,N_10205,N_8608);
and U13245 (N_13245,N_11942,N_11009);
xor U13246 (N_13246,N_9204,N_9925);
nand U13247 (N_13247,N_8335,N_8266);
nor U13248 (N_13248,N_8158,N_9967);
nand U13249 (N_13249,N_8881,N_8087);
or U13250 (N_13250,N_9405,N_10041);
and U13251 (N_13251,N_10696,N_10850);
and U13252 (N_13252,N_11853,N_11123);
or U13253 (N_13253,N_11307,N_9637);
or U13254 (N_13254,N_9841,N_9659);
nor U13255 (N_13255,N_9241,N_8694);
nor U13256 (N_13256,N_8984,N_9361);
nand U13257 (N_13257,N_9537,N_9195);
nand U13258 (N_13258,N_8492,N_11892);
nand U13259 (N_13259,N_10782,N_9653);
or U13260 (N_13260,N_9755,N_8054);
and U13261 (N_13261,N_9391,N_10115);
nor U13262 (N_13262,N_10887,N_8231);
xor U13263 (N_13263,N_8420,N_11337);
nor U13264 (N_13264,N_11966,N_8460);
xnor U13265 (N_13265,N_8672,N_10194);
and U13266 (N_13266,N_11087,N_8547);
or U13267 (N_13267,N_8203,N_8636);
nand U13268 (N_13268,N_10958,N_9942);
nand U13269 (N_13269,N_10100,N_8134);
or U13270 (N_13270,N_10746,N_9228);
and U13271 (N_13271,N_10547,N_9774);
xor U13272 (N_13272,N_9552,N_8599);
and U13273 (N_13273,N_11710,N_9331);
xor U13274 (N_13274,N_8744,N_10911);
and U13275 (N_13275,N_11370,N_8027);
nand U13276 (N_13276,N_8096,N_10786);
nor U13277 (N_13277,N_10117,N_8418);
or U13278 (N_13278,N_9577,N_10636);
xor U13279 (N_13279,N_8966,N_11238);
nor U13280 (N_13280,N_8644,N_8294);
nor U13281 (N_13281,N_9787,N_11660);
nand U13282 (N_13282,N_9815,N_8589);
nand U13283 (N_13283,N_10362,N_11520);
or U13284 (N_13284,N_8507,N_8276);
nand U13285 (N_13285,N_8570,N_10961);
nand U13286 (N_13286,N_9675,N_11486);
nand U13287 (N_13287,N_9973,N_9203);
or U13288 (N_13288,N_9118,N_11608);
nand U13289 (N_13289,N_10019,N_8381);
or U13290 (N_13290,N_8193,N_10470);
or U13291 (N_13291,N_8583,N_8292);
nor U13292 (N_13292,N_10248,N_11822);
nand U13293 (N_13293,N_10054,N_8516);
or U13294 (N_13294,N_10124,N_10108);
and U13295 (N_13295,N_10654,N_9280);
or U13296 (N_13296,N_11690,N_10743);
nand U13297 (N_13297,N_10685,N_10361);
nand U13298 (N_13298,N_10882,N_9039);
nand U13299 (N_13299,N_11863,N_8584);
or U13300 (N_13300,N_11854,N_8043);
and U13301 (N_13301,N_10754,N_11198);
and U13302 (N_13302,N_9414,N_11253);
nand U13303 (N_13303,N_10349,N_8469);
and U13304 (N_13304,N_11865,N_11885);
and U13305 (N_13305,N_11648,N_9849);
nor U13306 (N_13306,N_9240,N_9852);
nand U13307 (N_13307,N_11076,N_11783);
nor U13308 (N_13308,N_9592,N_8754);
xor U13309 (N_13309,N_9757,N_10550);
nand U13310 (N_13310,N_10893,N_9766);
xor U13311 (N_13311,N_10437,N_8667);
xnor U13312 (N_13312,N_10384,N_11957);
nor U13313 (N_13313,N_9895,N_11726);
or U13314 (N_13314,N_9394,N_9956);
or U13315 (N_13315,N_8909,N_10747);
and U13316 (N_13316,N_10611,N_9644);
and U13317 (N_13317,N_9532,N_8901);
or U13318 (N_13318,N_11573,N_10768);
and U13319 (N_13319,N_8768,N_9444);
or U13320 (N_13320,N_10812,N_10566);
nor U13321 (N_13321,N_9116,N_8081);
nor U13322 (N_13322,N_8431,N_9094);
nand U13323 (N_13323,N_11421,N_10197);
and U13324 (N_13324,N_8034,N_8401);
nand U13325 (N_13325,N_9211,N_9563);
and U13326 (N_13326,N_9256,N_10044);
nand U13327 (N_13327,N_9271,N_11688);
and U13328 (N_13328,N_8932,N_11873);
or U13329 (N_13329,N_10439,N_9872);
and U13330 (N_13330,N_8925,N_10644);
or U13331 (N_13331,N_8156,N_11519);
nor U13332 (N_13332,N_9035,N_9914);
and U13333 (N_13333,N_8748,N_9238);
nor U13334 (N_13334,N_11866,N_11313);
nor U13335 (N_13335,N_9097,N_8899);
nand U13336 (N_13336,N_8848,N_8053);
and U13337 (N_13337,N_11808,N_11338);
or U13338 (N_13338,N_11674,N_9085);
nor U13339 (N_13339,N_10178,N_10777);
nor U13340 (N_13340,N_11721,N_8332);
or U13341 (N_13341,N_8885,N_11412);
nand U13342 (N_13342,N_9617,N_9919);
xor U13343 (N_13343,N_9722,N_9688);
or U13344 (N_13344,N_8705,N_9086);
or U13345 (N_13345,N_10835,N_10030);
nand U13346 (N_13346,N_9950,N_9833);
nor U13347 (N_13347,N_10409,N_8849);
or U13348 (N_13348,N_8738,N_10805);
or U13349 (N_13349,N_9262,N_11819);
xnor U13350 (N_13350,N_10520,N_10872);
or U13351 (N_13351,N_10016,N_11797);
or U13352 (N_13352,N_8550,N_11052);
nor U13353 (N_13353,N_11583,N_10070);
xor U13354 (N_13354,N_9264,N_11827);
nor U13355 (N_13355,N_9941,N_10590);
and U13356 (N_13356,N_9034,N_10843);
nor U13357 (N_13357,N_8628,N_9630);
and U13358 (N_13358,N_10091,N_9799);
and U13359 (N_13359,N_10099,N_9254);
nand U13360 (N_13360,N_9940,N_11535);
nor U13361 (N_13361,N_9643,N_10833);
nor U13362 (N_13362,N_8505,N_9893);
nand U13363 (N_13363,N_11407,N_10347);
or U13364 (N_13364,N_11946,N_11017);
nand U13365 (N_13365,N_9691,N_8683);
and U13366 (N_13366,N_9550,N_10261);
nand U13367 (N_13367,N_10509,N_11616);
nor U13368 (N_13368,N_11334,N_8347);
or U13369 (N_13369,N_11324,N_9736);
or U13370 (N_13370,N_9048,N_10949);
or U13371 (N_13371,N_8717,N_11890);
nor U13372 (N_13372,N_9587,N_9857);
or U13373 (N_13373,N_10818,N_11295);
or U13374 (N_13374,N_9121,N_8370);
nand U13375 (N_13375,N_11159,N_11225);
or U13376 (N_13376,N_8011,N_8556);
xnor U13377 (N_13377,N_10809,N_10139);
or U13378 (N_13378,N_10653,N_10615);
nor U13379 (N_13379,N_8099,N_9590);
nor U13380 (N_13380,N_8568,N_10026);
nor U13381 (N_13381,N_11332,N_9571);
nand U13382 (N_13382,N_10972,N_9927);
and U13383 (N_13383,N_9811,N_8176);
nand U13384 (N_13384,N_10485,N_10110);
nand U13385 (N_13385,N_11221,N_10703);
nand U13386 (N_13386,N_9937,N_10641);
and U13387 (N_13387,N_11182,N_8826);
or U13388 (N_13388,N_9252,N_10947);
or U13389 (N_13389,N_11515,N_8024);
nor U13390 (N_13390,N_9157,N_11394);
or U13391 (N_13391,N_10857,N_11214);
and U13392 (N_13392,N_9535,N_9074);
or U13393 (N_13393,N_9952,N_10948);
or U13394 (N_13394,N_8821,N_10959);
nor U13395 (N_13395,N_10063,N_8124);
xnor U13396 (N_13396,N_8893,N_9702);
or U13397 (N_13397,N_9968,N_8051);
or U13398 (N_13398,N_11250,N_9652);
or U13399 (N_13399,N_10406,N_9489);
or U13400 (N_13400,N_11943,N_11262);
xnor U13401 (N_13401,N_10962,N_11557);
and U13402 (N_13402,N_9417,N_8593);
and U13403 (N_13403,N_8766,N_11257);
nor U13404 (N_13404,N_8993,N_9006);
nand U13405 (N_13405,N_9689,N_8987);
and U13406 (N_13406,N_9181,N_10418);
nand U13407 (N_13407,N_10173,N_8722);
nand U13408 (N_13408,N_8953,N_10999);
nand U13409 (N_13409,N_11024,N_9794);
or U13410 (N_13410,N_10060,N_11368);
and U13411 (N_13411,N_9840,N_11493);
and U13412 (N_13412,N_11770,N_11450);
nor U13413 (N_13413,N_11994,N_10081);
nand U13414 (N_13414,N_8151,N_9797);
nor U13415 (N_13415,N_10806,N_10697);
and U13416 (N_13416,N_10337,N_9909);
nand U13417 (N_13417,N_10627,N_10477);
or U13418 (N_13418,N_9141,N_8730);
nand U13419 (N_13419,N_10629,N_9132);
or U13420 (N_13420,N_10491,N_10390);
nand U13421 (N_13421,N_10655,N_8484);
nor U13422 (N_13422,N_8355,N_9205);
nor U13423 (N_13423,N_8592,N_11189);
xnor U13424 (N_13424,N_8554,N_10880);
nor U13425 (N_13425,N_10921,N_10829);
nand U13426 (N_13426,N_8153,N_8745);
nor U13427 (N_13427,N_10010,N_10588);
and U13428 (N_13428,N_10822,N_11498);
nand U13429 (N_13429,N_8598,N_11032);
nor U13430 (N_13430,N_9421,N_10565);
nand U13431 (N_13431,N_10218,N_11879);
nand U13432 (N_13432,N_8540,N_9407);
and U13433 (N_13433,N_11033,N_11431);
xnor U13434 (N_13434,N_9647,N_10048);
xor U13435 (N_13435,N_10868,N_8389);
nand U13436 (N_13436,N_8892,N_11187);
xor U13437 (N_13437,N_11124,N_10631);
nand U13438 (N_13438,N_11956,N_11568);
xnor U13439 (N_13439,N_8066,N_8980);
nor U13440 (N_13440,N_11481,N_11989);
nor U13441 (N_13441,N_11846,N_11658);
nand U13442 (N_13442,N_10027,N_8876);
nand U13443 (N_13443,N_9555,N_10129);
nor U13444 (N_13444,N_10736,N_9488);
and U13445 (N_13445,N_10333,N_10622);
nor U13446 (N_13446,N_11403,N_10133);
or U13447 (N_13447,N_9522,N_9765);
nand U13448 (N_13448,N_10304,N_9834);
or U13449 (N_13449,N_10772,N_9007);
nor U13450 (N_13450,N_10486,N_10497);
and U13451 (N_13451,N_8262,N_9805);
and U13452 (N_13452,N_11702,N_10667);
and U13453 (N_13453,N_11506,N_11461);
and U13454 (N_13454,N_9478,N_10267);
nor U13455 (N_13455,N_11197,N_8915);
and U13456 (N_13456,N_11162,N_9897);
or U13457 (N_13457,N_9574,N_10103);
and U13458 (N_13458,N_10957,N_11195);
nand U13459 (N_13459,N_11675,N_8191);
nand U13460 (N_13460,N_11383,N_8860);
and U13461 (N_13461,N_10557,N_9810);
or U13462 (N_13462,N_11787,N_10977);
nand U13463 (N_13463,N_10901,N_9124);
or U13464 (N_13464,N_8740,N_10240);
and U13465 (N_13465,N_9838,N_11530);
nor U13466 (N_13466,N_8111,N_11862);
nor U13467 (N_13467,N_10719,N_8776);
or U13468 (N_13468,N_10558,N_10440);
or U13469 (N_13469,N_9494,N_10411);
and U13470 (N_13470,N_9296,N_9257);
nand U13471 (N_13471,N_9277,N_10774);
and U13472 (N_13472,N_8390,N_9525);
nor U13473 (N_13473,N_10944,N_9509);
xor U13474 (N_13474,N_9904,N_9720);
xnor U13475 (N_13475,N_10394,N_11222);
nand U13476 (N_13476,N_11701,N_10906);
and U13477 (N_13477,N_11718,N_9977);
and U13478 (N_13478,N_10392,N_8320);
or U13479 (N_13479,N_8727,N_9798);
or U13480 (N_13480,N_10179,N_11417);
or U13481 (N_13481,N_11907,N_9547);
nor U13482 (N_13482,N_9322,N_9348);
or U13483 (N_13483,N_9175,N_10369);
xor U13484 (N_13484,N_11130,N_8457);
xnor U13485 (N_13485,N_10953,N_10018);
and U13486 (N_13486,N_10795,N_10453);
nor U13487 (N_13487,N_9789,N_11668);
or U13488 (N_13488,N_9359,N_11739);
nand U13489 (N_13489,N_10076,N_8928);
and U13490 (N_13490,N_11930,N_11305);
xor U13491 (N_13491,N_9345,N_8453);
and U13492 (N_13492,N_9243,N_8843);
or U13493 (N_13493,N_11382,N_11676);
or U13494 (N_13494,N_9943,N_8448);
nor U13495 (N_13495,N_11309,N_9832);
or U13496 (N_13496,N_10981,N_9650);
or U13497 (N_13497,N_11213,N_10169);
nor U13498 (N_13498,N_11191,N_8400);
xor U13499 (N_13499,N_10814,N_8247);
and U13500 (N_13500,N_11545,N_11791);
and U13501 (N_13501,N_8914,N_8101);
or U13502 (N_13502,N_10605,N_8587);
and U13503 (N_13503,N_8039,N_11704);
and U13504 (N_13504,N_11501,N_9185);
nand U13505 (N_13505,N_10691,N_8661);
and U13506 (N_13506,N_9796,N_8582);
and U13507 (N_13507,N_11803,N_9112);
nor U13508 (N_13508,N_8663,N_11769);
and U13509 (N_13509,N_9373,N_10084);
and U13510 (N_13510,N_9520,N_8171);
xnor U13511 (N_13511,N_11695,N_11379);
nor U13512 (N_13512,N_8157,N_10350);
or U13513 (N_13513,N_11362,N_9431);
nor U13514 (N_13514,N_9877,N_9876);
and U13515 (N_13515,N_10219,N_11181);
nand U13516 (N_13516,N_8972,N_8468);
and U13517 (N_13517,N_10984,N_11260);
and U13518 (N_13518,N_11649,N_10260);
or U13519 (N_13519,N_10994,N_10396);
or U13520 (N_13520,N_10113,N_11388);
and U13521 (N_13521,N_10930,N_10597);
nand U13522 (N_13522,N_10189,N_8040);
and U13523 (N_13523,N_8348,N_8756);
or U13524 (N_13524,N_8104,N_9892);
nand U13525 (N_13525,N_9901,N_10784);
xor U13526 (N_13526,N_10681,N_8534);
or U13527 (N_13527,N_10824,N_10954);
and U13528 (N_13528,N_10996,N_8817);
and U13529 (N_13529,N_9795,N_9773);
nand U13530 (N_13530,N_8737,N_9651);
nand U13531 (N_13531,N_10208,N_9779);
and U13532 (N_13532,N_11543,N_8963);
or U13533 (N_13533,N_10728,N_10209);
nand U13534 (N_13534,N_9786,N_9615);
or U13535 (N_13535,N_10792,N_9780);
and U13536 (N_13536,N_8508,N_11308);
and U13537 (N_13537,N_8325,N_10188);
and U13538 (N_13538,N_11491,N_11730);
or U13539 (N_13539,N_8619,N_11143);
nor U13540 (N_13540,N_11467,N_8781);
or U13541 (N_13541,N_10495,N_11553);
and U13542 (N_13542,N_10638,N_10726);
or U13543 (N_13543,N_10738,N_10634);
and U13544 (N_13544,N_8708,N_8062);
nand U13545 (N_13545,N_9082,N_11210);
and U13546 (N_13546,N_8702,N_10779);
nor U13547 (N_13547,N_11365,N_11513);
or U13548 (N_13548,N_9200,N_9939);
nand U13549 (N_13549,N_9847,N_10819);
and U13550 (N_13550,N_11555,N_8423);
nor U13551 (N_13551,N_8811,N_10966);
or U13552 (N_13552,N_11132,N_8657);
xor U13553 (N_13553,N_10938,N_9481);
or U13554 (N_13554,N_9501,N_10800);
and U13555 (N_13555,N_8602,N_10690);
nor U13556 (N_13556,N_9450,N_10143);
xor U13557 (N_13557,N_8890,N_8642);
nand U13558 (N_13558,N_11270,N_10321);
nand U13559 (N_13559,N_11081,N_8601);
and U13560 (N_13560,N_11073,N_10983);
or U13561 (N_13561,N_8946,N_8533);
or U13562 (N_13562,N_10790,N_9863);
and U13563 (N_13563,N_9392,N_9503);
nor U13564 (N_13564,N_11069,N_11310);
and U13565 (N_13565,N_9046,N_10849);
nor U13566 (N_13566,N_10289,N_11537);
or U13567 (N_13567,N_9065,N_10589);
and U13568 (N_13568,N_10153,N_11889);
and U13569 (N_13569,N_10542,N_10057);
and U13570 (N_13570,N_9829,N_11973);
nand U13571 (N_13571,N_8596,N_10435);
nand U13572 (N_13572,N_8825,N_9479);
xnor U13573 (N_13573,N_9305,N_11780);
xnor U13574 (N_13574,N_9347,N_9059);
xnor U13575 (N_13575,N_10522,N_11320);
nor U13576 (N_13576,N_8309,N_10871);
nor U13577 (N_13577,N_10714,N_11013);
or U13578 (N_13578,N_10686,N_11782);
nor U13579 (N_13579,N_11845,N_9870);
nor U13580 (N_13580,N_11578,N_11325);
or U13581 (N_13581,N_8116,N_11398);
nand U13582 (N_13582,N_9098,N_8947);
or U13583 (N_13583,N_10923,N_11948);
and U13584 (N_13584,N_9173,N_9866);
or U13585 (N_13585,N_10791,N_11796);
nor U13586 (N_13586,N_9680,N_9869);
nand U13587 (N_13587,N_11965,N_11451);
nand U13588 (N_13588,N_10262,N_11836);
nand U13589 (N_13589,N_10033,N_8019);
nor U13590 (N_13590,N_9299,N_8887);
or U13591 (N_13591,N_11888,N_8974);
or U13592 (N_13592,N_8075,N_10723);
nand U13593 (N_13593,N_9202,N_11952);
nor U13594 (N_13594,N_10532,N_8036);
and U13595 (N_13595,N_11772,N_8403);
nor U13596 (N_13596,N_9304,N_10928);
or U13597 (N_13597,N_9130,N_10832);
and U13598 (N_13598,N_11048,N_11974);
xnor U13599 (N_13599,N_11204,N_10932);
or U13600 (N_13600,N_9117,N_10122);
xor U13601 (N_13601,N_9750,N_10493);
nand U13602 (N_13602,N_8989,N_10618);
nand U13603 (N_13603,N_10666,N_9423);
nor U13604 (N_13604,N_10410,N_8139);
or U13605 (N_13605,N_9206,N_8356);
or U13606 (N_13606,N_10053,N_10905);
and U13607 (N_13607,N_8302,N_10846);
nor U13608 (N_13608,N_8828,N_9380);
and U13609 (N_13609,N_9077,N_9183);
nor U13610 (N_13610,N_9954,N_11321);
and U13611 (N_13611,N_10309,N_10889);
nand U13612 (N_13612,N_9312,N_11326);
xor U13613 (N_13613,N_9516,N_10202);
or U13614 (N_13614,N_8223,N_8217);
or U13615 (N_13615,N_11987,N_11874);
or U13616 (N_13616,N_8954,N_9490);
and U13617 (N_13617,N_11153,N_11356);
and U13618 (N_13618,N_10551,N_10707);
or U13619 (N_13619,N_9033,N_11194);
nand U13620 (N_13620,N_10939,N_10389);
or U13621 (N_13621,N_11168,N_11717);
xor U13622 (N_13622,N_9045,N_11914);
or U13623 (N_13623,N_10925,N_8475);
or U13624 (N_13624,N_11918,N_10864);
or U13625 (N_13625,N_8788,N_9683);
or U13626 (N_13626,N_8490,N_10244);
and U13627 (N_13627,N_8650,N_8357);
nor U13628 (N_13628,N_11286,N_11805);
nor U13629 (N_13629,N_10062,N_9374);
nand U13630 (N_13630,N_9527,N_10138);
or U13631 (N_13631,N_8155,N_9760);
nor U13632 (N_13632,N_8634,N_10859);
or U13633 (N_13633,N_10436,N_9878);
and U13634 (N_13634,N_10803,N_10069);
and U13635 (N_13635,N_10191,N_11528);
or U13636 (N_13636,N_10319,N_10271);
nor U13637 (N_13637,N_8012,N_8573);
and U13638 (N_13638,N_11765,N_11910);
nor U13639 (N_13639,N_11152,N_10257);
or U13640 (N_13640,N_11605,N_8412);
or U13641 (N_13641,N_11025,N_9236);
nor U13642 (N_13642,N_10035,N_8365);
or U13643 (N_13643,N_9014,N_11653);
nand U13644 (N_13644,N_11115,N_11525);
and U13645 (N_13645,N_10722,N_11223);
nor U13646 (N_13646,N_9709,N_10273);
nand U13647 (N_13647,N_11816,N_10141);
nor U13648 (N_13648,N_10595,N_11410);
nor U13649 (N_13649,N_9697,N_10763);
nand U13650 (N_13650,N_10288,N_8284);
and U13651 (N_13651,N_9936,N_10345);
and U13652 (N_13652,N_8986,N_10005);
or U13653 (N_13653,N_11127,N_8548);
xor U13654 (N_13654,N_9545,N_8378);
or U13655 (N_13655,N_11297,N_9616);
and U13656 (N_13656,N_9978,N_9739);
or U13657 (N_13657,N_9498,N_11010);
nand U13658 (N_13658,N_8406,N_10412);
and U13659 (N_13659,N_10762,N_11738);
xnor U13660 (N_13660,N_10575,N_9108);
xor U13661 (N_13661,N_11691,N_10072);
or U13662 (N_13662,N_10498,N_11007);
nand U13663 (N_13663,N_8945,N_8149);
and U13664 (N_13664,N_9443,N_8030);
nand U13665 (N_13665,N_10936,N_8046);
nor U13666 (N_13666,N_11171,N_11856);
and U13667 (N_13667,N_9674,N_9357);
and U13668 (N_13668,N_11839,N_8281);
and U13669 (N_13669,N_8961,N_8366);
nand U13670 (N_13670,N_8820,N_8326);
xor U13671 (N_13671,N_9042,N_11057);
and U13672 (N_13672,N_11799,N_11719);
nor U13673 (N_13673,N_8090,N_9218);
nand U13674 (N_13674,N_8267,N_11849);
nor U13675 (N_13675,N_11452,N_8287);
and U13676 (N_13676,N_9196,N_11074);
or U13677 (N_13677,N_10821,N_11218);
nor U13678 (N_13678,N_11434,N_10372);
nand U13679 (N_13679,N_11361,N_10471);
and U13680 (N_13680,N_9462,N_11119);
or U13681 (N_13681,N_10383,N_9449);
xnor U13682 (N_13682,N_8314,N_11934);
nand U13683 (N_13683,N_9287,N_9603);
or U13684 (N_13684,N_11380,N_11328);
nand U13685 (N_13685,N_8699,N_11705);
and U13686 (N_13686,N_10741,N_10326);
xor U13687 (N_13687,N_10039,N_11241);
and U13688 (N_13688,N_8553,N_11692);
and U13689 (N_13689,N_11544,N_9024);
and U13690 (N_13690,N_8035,N_11020);
nor U13691 (N_13691,N_9237,N_9245);
nand U13692 (N_13692,N_9924,N_8246);
and U13693 (N_13693,N_9292,N_8810);
or U13694 (N_13694,N_9586,N_11289);
or U13695 (N_13695,N_11268,N_11287);
or U13696 (N_13696,N_11216,N_11697);
and U13697 (N_13697,N_9687,N_10603);
or U13698 (N_13698,N_9028,N_11318);
and U13699 (N_13699,N_10712,N_11179);
nor U13700 (N_13700,N_9229,N_10428);
nand U13701 (N_13701,N_9177,N_9542);
nand U13702 (N_13702,N_9519,N_8404);
and U13703 (N_13703,N_10067,N_10370);
and U13704 (N_13704,N_10106,N_11916);
and U13705 (N_13705,N_9341,N_9974);
nand U13706 (N_13706,N_9061,N_11405);
nand U13707 (N_13707,N_11459,N_10662);
nand U13708 (N_13708,N_10185,N_8387);
nand U13709 (N_13709,N_8793,N_10844);
or U13710 (N_13710,N_8279,N_11556);
nor U13711 (N_13711,N_11899,N_10904);
or U13712 (N_13712,N_10459,N_9764);
or U13713 (N_13713,N_8943,N_11606);
or U13714 (N_13714,N_9184,N_11971);
or U13715 (N_13715,N_9961,N_9638);
nor U13716 (N_13716,N_10127,N_9645);
or U13717 (N_13717,N_9931,N_8360);
nor U13718 (N_13718,N_9808,N_11546);
nand U13719 (N_13719,N_8496,N_10755);
nor U13720 (N_13720,N_9073,N_10187);
nor U13721 (N_13721,N_11004,N_10109);
or U13722 (N_13722,N_8798,N_10604);
nor U13723 (N_13723,N_8631,N_8033);
nand U13724 (N_13724,N_10167,N_9569);
nand U13725 (N_13725,N_11414,N_8927);
or U13726 (N_13726,N_8495,N_11455);
nor U13727 (N_13727,N_10675,N_11128);
and U13728 (N_13728,N_11588,N_9631);
nand U13729 (N_13729,N_10156,N_9686);
nand U13730 (N_13730,N_9989,N_10855);
nor U13731 (N_13731,N_11188,N_9746);
nand U13732 (N_13732,N_9099,N_9963);
xor U13733 (N_13733,N_8603,N_11436);
nand U13734 (N_13734,N_9844,N_11173);
nor U13735 (N_13735,N_9197,N_11864);
and U13736 (N_13736,N_11922,N_8778);
and U13737 (N_13737,N_10657,N_8352);
or U13738 (N_13738,N_11118,N_9485);
xnor U13739 (N_13739,N_11085,N_11524);
and U13740 (N_13740,N_9151,N_9096);
nand U13741 (N_13741,N_10320,N_11369);
or U13742 (N_13742,N_10585,N_8353);
or U13743 (N_13743,N_9837,N_8715);
nand U13744 (N_13744,N_10718,N_11733);
nand U13745 (N_13745,N_10243,N_9871);
or U13746 (N_13746,N_8413,N_9475);
nand U13747 (N_13747,N_8829,N_10277);
nand U13748 (N_13748,N_11773,N_8454);
and U13749 (N_13749,N_11597,N_11016);
or U13750 (N_13750,N_11244,N_9419);
xnor U13751 (N_13751,N_11790,N_11527);
nor U13752 (N_13752,N_11298,N_10159);
or U13753 (N_13753,N_11550,N_11667);
and U13754 (N_13754,N_8098,N_8021);
and U13755 (N_13755,N_10838,N_8809);
or U13756 (N_13756,N_11713,N_11729);
nor U13757 (N_13757,N_10694,N_8180);
nand U13758 (N_13758,N_9453,N_9965);
nor U13759 (N_13759,N_9148,N_10549);
and U13760 (N_13760,N_8379,N_8446);
nand U13761 (N_13761,N_10701,N_8115);
nor U13762 (N_13762,N_11154,N_8572);
xor U13763 (N_13763,N_9907,N_8800);
nand U13764 (N_13764,N_9678,N_10365);
xor U13765 (N_13765,N_8000,N_9530);
nor U13766 (N_13766,N_10121,N_9803);
nor U13767 (N_13767,N_9428,N_11002);
nor U13768 (N_13768,N_8935,N_8965);
and U13769 (N_13769,N_11180,N_9628);
and U13770 (N_13770,N_8574,N_8983);
or U13771 (N_13771,N_8520,N_10464);
xor U13772 (N_13772,N_9783,N_11438);
or U13773 (N_13773,N_9290,N_10236);
or U13774 (N_13774,N_9663,N_8823);
nand U13775 (N_13775,N_10913,N_8982);
or U13776 (N_13776,N_9339,N_11399);
nor U13777 (N_13777,N_10894,N_9057);
xnor U13778 (N_13778,N_11906,N_10166);
nor U13779 (N_13779,N_8949,N_8922);
nand U13780 (N_13780,N_11215,N_10991);
and U13781 (N_13781,N_10978,N_10748);
and U13782 (N_13782,N_8301,N_10732);
or U13783 (N_13783,N_9333,N_10340);
or U13784 (N_13784,N_11745,N_10668);
nor U13785 (N_13785,N_11446,N_10642);
nor U13786 (N_13786,N_10645,N_10303);
or U13787 (N_13787,N_8872,N_8970);
and U13788 (N_13788,N_11637,N_9772);
or U13789 (N_13789,N_11497,N_9513);
or U13790 (N_13790,N_10206,N_11861);
or U13791 (N_13791,N_9860,N_10131);
and U13792 (N_13792,N_10385,N_11283);
nand U13793 (N_13793,N_9861,N_11641);
and U13794 (N_13794,N_10285,N_8542);
nor U13795 (N_13795,N_10003,N_10756);
and U13796 (N_13796,N_9103,N_10620);
and U13797 (N_13797,N_8121,N_8884);
or U13798 (N_13798,N_11442,N_10573);
nand U13799 (N_13799,N_9957,N_9585);
nor U13800 (N_13800,N_9167,N_11883);
nand U13801 (N_13801,N_8186,N_9350);
nor U13802 (N_13802,N_8211,N_9217);
nor U13803 (N_13803,N_8321,N_8822);
nand U13804 (N_13804,N_11441,N_8135);
nand U13805 (N_13805,N_9707,N_8785);
nor U13806 (N_13806,N_9758,N_11129);
or U13807 (N_13807,N_10811,N_10503);
and U13808 (N_13808,N_11503,N_8263);
or U13809 (N_13809,N_8942,N_10170);
nor U13810 (N_13810,N_10658,N_10371);
or U13811 (N_13811,N_8169,N_10374);
or U13812 (N_13812,N_9626,N_10876);
nor U13813 (N_13813,N_9168,N_9070);
nor U13814 (N_13814,N_8489,N_9037);
xor U13815 (N_13815,N_11507,N_9988);
nand U13816 (N_13816,N_9429,N_10927);
or U13817 (N_13817,N_11687,N_10265);
and U13818 (N_13818,N_10086,N_10322);
or U13819 (N_13819,N_9465,N_11229);
and U13820 (N_13820,N_10529,N_10487);
or U13821 (N_13821,N_9476,N_11323);
and U13822 (N_13822,N_11249,N_9980);
nor U13823 (N_13823,N_11000,N_8559);
nor U13824 (N_13824,N_8257,N_9546);
or U13825 (N_13825,N_10788,N_9122);
or U13826 (N_13826,N_8830,N_11061);
nor U13827 (N_13827,N_8270,N_8862);
and U13828 (N_13828,N_8969,N_9286);
xor U13829 (N_13829,N_9285,N_11104);
nand U13830 (N_13830,N_11841,N_11831);
nand U13831 (N_13831,N_8513,N_8576);
or U13832 (N_13832,N_9640,N_8710);
xnor U13833 (N_13833,N_9036,N_10830);
and U13834 (N_13834,N_10576,N_8177);
or U13835 (N_13835,N_10778,N_9923);
nand U13836 (N_13836,N_9387,N_9681);
nor U13837 (N_13837,N_11912,N_11752);
nand U13838 (N_13838,N_10973,N_10580);
or U13839 (N_13839,N_9551,N_8994);
and U13840 (N_13840,N_8227,N_9754);
nor U13841 (N_13841,N_8886,N_10980);
or U13842 (N_13842,N_10101,N_9041);
nand U13843 (N_13843,N_8437,N_10461);
and U13844 (N_13844,N_11454,N_10914);
xor U13845 (N_13845,N_11012,N_8244);
or U13846 (N_13846,N_10651,N_10313);
nand U13847 (N_13847,N_9411,N_11416);
or U13848 (N_13848,N_9508,N_9223);
and U13849 (N_13849,N_9969,N_11817);
nor U13850 (N_13850,N_8258,N_11391);
or U13851 (N_13851,N_8443,N_11722);
or U13852 (N_13852,N_9749,N_9993);
and U13853 (N_13853,N_11015,N_9676);
or U13854 (N_13854,N_9180,N_10567);
nand U13855 (N_13855,N_11961,N_8122);
nor U13856 (N_13856,N_9268,N_10286);
nor U13857 (N_13857,N_8249,N_8273);
nand U13858 (N_13858,N_11638,N_9696);
nand U13859 (N_13859,N_8692,N_11895);
nor U13860 (N_13860,N_10987,N_9611);
or U13861 (N_13861,N_8853,N_11094);
and U13862 (N_13862,N_9745,N_11341);
or U13863 (N_13863,N_9568,N_11754);
nand U13864 (N_13864,N_10148,N_11255);
or U13865 (N_13865,N_8594,N_8324);
or U13866 (N_13866,N_11901,N_10960);
nand U13867 (N_13867,N_10896,N_8751);
and U13868 (N_13868,N_10280,N_9856);
or U13869 (N_13869,N_8316,N_11510);
nor U13870 (N_13870,N_11285,N_11100);
xor U13871 (N_13871,N_9917,N_9911);
nor U13872 (N_13872,N_8633,N_8445);
and U13873 (N_13873,N_8844,N_10664);
nand U13874 (N_13874,N_8686,N_11709);
and U13875 (N_13875,N_8907,N_9715);
nor U13876 (N_13876,N_10183,N_11474);
and U13877 (N_13877,N_10083,N_8205);
nand U13878 (N_13878,N_10400,N_11990);
nand U13879 (N_13879,N_10699,N_8575);
nand U13880 (N_13880,N_9864,N_10028);
and U13881 (N_13881,N_11601,N_11072);
and U13882 (N_13882,N_8861,N_11141);
xor U13883 (N_13883,N_10279,N_10596);
and U13884 (N_13884,N_10446,N_11366);
nand U13885 (N_13885,N_10004,N_10841);
nor U13886 (N_13886,N_10186,N_8623);
or U13887 (N_13887,N_9473,N_8865);
or U13888 (N_13888,N_9171,N_11208);
nand U13889 (N_13889,N_9016,N_10414);
and U13890 (N_13890,N_8760,N_11986);
and U13891 (N_13891,N_10210,N_9504);
xnor U13892 (N_13892,N_9382,N_8767);
nor U13893 (N_13893,N_10140,N_10112);
nand U13894 (N_13894,N_9900,N_11681);
xnor U13895 (N_13895,N_11470,N_8979);
nor U13896 (N_13896,N_9673,N_10460);
xnor U13897 (N_13897,N_9378,N_8581);
or U13898 (N_13898,N_10633,N_9087);
and U13899 (N_13899,N_10355,N_10164);
nor U13900 (N_13900,N_8998,N_8718);
nor U13901 (N_13901,N_10017,N_8092);
and U13902 (N_13902,N_9582,N_10327);
nand U13903 (N_13903,N_8192,N_9403);
nand U13904 (N_13904,N_8990,N_8202);
nand U13905 (N_13905,N_10080,N_9409);
nand U13906 (N_13906,N_9541,N_9990);
nor U13907 (N_13907,N_10781,N_10556);
or U13908 (N_13908,N_11619,N_11047);
xnor U13909 (N_13909,N_9370,N_8426);
or U13910 (N_13910,N_10933,N_10956);
or U13911 (N_13911,N_10292,N_8616);
nor U13912 (N_13912,N_11804,N_8673);
or U13913 (N_13913,N_8511,N_10066);
nor U13914 (N_13914,N_9439,N_9671);
or U13915 (N_13915,N_9867,N_11521);
and U13916 (N_13916,N_10794,N_9017);
nor U13917 (N_13917,N_10104,N_9748);
or U13918 (N_13918,N_8229,N_10182);
nor U13919 (N_13919,N_8741,N_11661);
or U13920 (N_13920,N_8563,N_11489);
nor U13921 (N_13921,N_9510,N_10344);
nand U13922 (N_13922,N_9328,N_10229);
nor U13923 (N_13923,N_11534,N_8930);
nand U13924 (N_13924,N_8440,N_9507);
and U13925 (N_13925,N_9410,N_10834);
xnor U13926 (N_13926,N_9533,N_9249);
or U13927 (N_13927,N_8866,N_10619);
or U13928 (N_13928,N_9868,N_9775);
xnor U13929 (N_13929,N_9885,N_11514);
or U13930 (N_13930,N_8163,N_10346);
nor U13931 (N_13931,N_10637,N_10047);
nand U13932 (N_13932,N_9078,N_10125);
or U13933 (N_13933,N_11996,N_11809);
nor U13934 (N_13934,N_11381,N_11411);
and U13935 (N_13935,N_9152,N_11625);
and U13936 (N_13936,N_8498,N_8870);
nand U13937 (N_13937,N_10941,N_9340);
nand U13938 (N_13938,N_10483,N_10474);
nand U13939 (N_13939,N_8805,N_9771);
and U13940 (N_13940,N_8212,N_11447);
nor U13941 (N_13941,N_8790,N_8242);
nand U13942 (N_13942,N_11540,N_10282);
and U13943 (N_13943,N_11938,N_11319);
xnor U13944 (N_13944,N_10943,N_9812);
nor U13945 (N_13945,N_8233,N_10425);
or U13946 (N_13946,N_10096,N_8769);
nand U13947 (N_13947,N_10672,N_9172);
nand U13948 (N_13948,N_11107,N_10881);
and U13949 (N_13949,N_9506,N_9306);
or U13950 (N_13950,N_11247,N_8750);
and U13951 (N_13951,N_10508,N_8855);
nor U13952 (N_13952,N_8154,N_9199);
and U13953 (N_13953,N_9412,N_10256);
nand U13954 (N_13954,N_9906,N_8351);
xnor U13955 (N_13955,N_10395,N_10810);
or U13956 (N_13956,N_9372,N_10910);
and U13957 (N_13957,N_9971,N_10569);
nand U13958 (N_13958,N_8646,N_9875);
nand U13959 (N_13959,N_8241,N_9999);
nor U13960 (N_13960,N_9260,N_10302);
and U13961 (N_13961,N_8999,N_8430);
nand U13962 (N_13962,N_11372,N_11192);
nor U13963 (N_13963,N_10480,N_10481);
or U13964 (N_13964,N_8757,N_9219);
nor U13965 (N_13965,N_11516,N_8436);
or U13966 (N_13966,N_10920,N_11842);
or U13967 (N_13967,N_8130,N_8607);
or U13968 (N_13968,N_10599,N_9538);
nand U13969 (N_13969,N_10144,N_8409);
or U13970 (N_13970,N_8160,N_9272);
and U13971 (N_13971,N_9352,N_9499);
nor U13972 (N_13972,N_9300,N_10869);
nor U13973 (N_13973,N_10336,N_8867);
xnor U13974 (N_13974,N_9553,N_11360);
nand U13975 (N_13975,N_9949,N_11672);
nor U13976 (N_13976,N_10284,N_11877);
nor U13977 (N_13977,N_8685,N_8260);
and U13978 (N_13978,N_9753,N_9910);
and U13979 (N_13979,N_9920,N_10393);
or U13980 (N_13980,N_10023,N_9930);
or U13981 (N_13981,N_10042,N_9579);
nor U13982 (N_13982,N_10274,N_11109);
or U13983 (N_13983,N_8546,N_9733);
or U13984 (N_13984,N_8020,N_10434);
and U13985 (N_13985,N_8138,N_11219);
nor U13986 (N_13986,N_9246,N_11378);
and U13987 (N_13987,N_11766,N_8076);
nand U13988 (N_13988,N_9466,N_10364);
and U13989 (N_13989,N_9463,N_11598);
and U13990 (N_13990,N_9657,N_9813);
xor U13991 (N_13991,N_11774,N_9889);
or U13992 (N_13992,N_8466,N_9090);
nor U13993 (N_13993,N_11640,N_9027);
nor U13994 (N_13994,N_9135,N_8146);
nand U13995 (N_13995,N_8773,N_10237);
nor U13996 (N_13996,N_8442,N_9188);
nand U13997 (N_13997,N_10692,N_9726);
and U13998 (N_13998,N_11066,N_10659);
nor U13999 (N_13999,N_9807,N_9377);
and U14000 (N_14000,N_9490,N_9752);
or U14001 (N_14001,N_11840,N_8937);
or U14002 (N_14002,N_11485,N_9930);
nand U14003 (N_14003,N_8493,N_9301);
and U14004 (N_14004,N_11678,N_10256);
nand U14005 (N_14005,N_10047,N_10134);
nand U14006 (N_14006,N_10325,N_11219);
nand U14007 (N_14007,N_10839,N_8147);
xor U14008 (N_14008,N_11363,N_9192);
nand U14009 (N_14009,N_11033,N_9045);
or U14010 (N_14010,N_10738,N_11509);
nand U14011 (N_14011,N_11811,N_9693);
or U14012 (N_14012,N_9502,N_10734);
xnor U14013 (N_14013,N_9056,N_8721);
nand U14014 (N_14014,N_8365,N_9090);
and U14015 (N_14015,N_11726,N_10969);
or U14016 (N_14016,N_11136,N_9656);
and U14017 (N_14017,N_10573,N_11538);
or U14018 (N_14018,N_10324,N_9513);
nor U14019 (N_14019,N_10360,N_8770);
xnor U14020 (N_14020,N_10906,N_9365);
or U14021 (N_14021,N_11680,N_10396);
nand U14022 (N_14022,N_11272,N_10730);
nand U14023 (N_14023,N_10062,N_8980);
nor U14024 (N_14024,N_10787,N_10273);
nor U14025 (N_14025,N_11668,N_10661);
or U14026 (N_14026,N_8324,N_8237);
or U14027 (N_14027,N_11162,N_8037);
nor U14028 (N_14028,N_11176,N_8376);
nor U14029 (N_14029,N_8075,N_9461);
or U14030 (N_14030,N_8723,N_8391);
or U14031 (N_14031,N_10522,N_9114);
nor U14032 (N_14032,N_11427,N_10989);
and U14033 (N_14033,N_11125,N_11848);
nand U14034 (N_14034,N_10258,N_10303);
xor U14035 (N_14035,N_9108,N_11604);
or U14036 (N_14036,N_9877,N_8260);
nand U14037 (N_14037,N_10516,N_10733);
or U14038 (N_14038,N_9576,N_9355);
and U14039 (N_14039,N_10657,N_11916);
nor U14040 (N_14040,N_10257,N_9573);
xor U14041 (N_14041,N_10987,N_10983);
nor U14042 (N_14042,N_8627,N_11827);
or U14043 (N_14043,N_9638,N_10368);
or U14044 (N_14044,N_8363,N_8274);
nor U14045 (N_14045,N_9073,N_10742);
and U14046 (N_14046,N_11297,N_10370);
or U14047 (N_14047,N_8393,N_10954);
and U14048 (N_14048,N_11741,N_9873);
nand U14049 (N_14049,N_8056,N_9510);
nand U14050 (N_14050,N_8786,N_10917);
or U14051 (N_14051,N_8157,N_9095);
nand U14052 (N_14052,N_9361,N_8772);
xnor U14053 (N_14053,N_8068,N_10480);
and U14054 (N_14054,N_11488,N_9552);
nor U14055 (N_14055,N_10942,N_11485);
nand U14056 (N_14056,N_11602,N_11813);
xnor U14057 (N_14057,N_8451,N_9156);
or U14058 (N_14058,N_9892,N_10574);
and U14059 (N_14059,N_10146,N_9918);
nor U14060 (N_14060,N_9881,N_10373);
nand U14061 (N_14061,N_8726,N_10524);
and U14062 (N_14062,N_11731,N_11251);
or U14063 (N_14063,N_9726,N_9074);
and U14064 (N_14064,N_9110,N_8769);
or U14065 (N_14065,N_9423,N_8378);
or U14066 (N_14066,N_11660,N_11767);
nor U14067 (N_14067,N_9222,N_8875);
and U14068 (N_14068,N_8572,N_11188);
nand U14069 (N_14069,N_11546,N_8203);
nor U14070 (N_14070,N_9640,N_10252);
nor U14071 (N_14071,N_8393,N_10357);
and U14072 (N_14072,N_9418,N_9028);
nor U14073 (N_14073,N_9372,N_10182);
nand U14074 (N_14074,N_8472,N_11707);
nor U14075 (N_14075,N_8869,N_10050);
nor U14076 (N_14076,N_8313,N_8930);
nor U14077 (N_14077,N_8828,N_9570);
and U14078 (N_14078,N_8504,N_9705);
nor U14079 (N_14079,N_11480,N_11160);
nor U14080 (N_14080,N_8621,N_10421);
nand U14081 (N_14081,N_10563,N_8993);
and U14082 (N_14082,N_8137,N_10256);
nor U14083 (N_14083,N_8791,N_10521);
and U14084 (N_14084,N_10072,N_9447);
nor U14085 (N_14085,N_8577,N_11257);
and U14086 (N_14086,N_9638,N_9860);
or U14087 (N_14087,N_11589,N_10703);
nand U14088 (N_14088,N_11150,N_9880);
or U14089 (N_14089,N_11764,N_9253);
and U14090 (N_14090,N_11688,N_11915);
or U14091 (N_14091,N_11867,N_8627);
and U14092 (N_14092,N_10108,N_9346);
nor U14093 (N_14093,N_11836,N_8362);
or U14094 (N_14094,N_8629,N_10645);
nand U14095 (N_14095,N_10979,N_11105);
nor U14096 (N_14096,N_10102,N_11691);
nor U14097 (N_14097,N_10697,N_10448);
nor U14098 (N_14098,N_11351,N_8975);
nand U14099 (N_14099,N_9507,N_9523);
xnor U14100 (N_14100,N_8782,N_9526);
or U14101 (N_14101,N_8957,N_9050);
nor U14102 (N_14102,N_8522,N_11980);
nand U14103 (N_14103,N_9250,N_9781);
nand U14104 (N_14104,N_9392,N_10075);
or U14105 (N_14105,N_9936,N_10918);
and U14106 (N_14106,N_10535,N_11045);
and U14107 (N_14107,N_11759,N_9957);
and U14108 (N_14108,N_11495,N_11255);
nor U14109 (N_14109,N_9249,N_9394);
or U14110 (N_14110,N_11918,N_10165);
or U14111 (N_14111,N_11878,N_11182);
nor U14112 (N_14112,N_10190,N_10908);
or U14113 (N_14113,N_9667,N_9262);
nand U14114 (N_14114,N_11192,N_10375);
xor U14115 (N_14115,N_11418,N_11426);
or U14116 (N_14116,N_9052,N_10490);
nand U14117 (N_14117,N_8023,N_8971);
and U14118 (N_14118,N_8037,N_11726);
and U14119 (N_14119,N_10322,N_8229);
and U14120 (N_14120,N_10724,N_11581);
or U14121 (N_14121,N_8073,N_8718);
nor U14122 (N_14122,N_10570,N_8408);
xor U14123 (N_14123,N_8154,N_8250);
or U14124 (N_14124,N_10476,N_9410);
or U14125 (N_14125,N_11090,N_10678);
and U14126 (N_14126,N_11654,N_8899);
and U14127 (N_14127,N_8715,N_9768);
nor U14128 (N_14128,N_8275,N_10536);
or U14129 (N_14129,N_11764,N_11979);
or U14130 (N_14130,N_9987,N_10708);
and U14131 (N_14131,N_9860,N_8661);
xnor U14132 (N_14132,N_11195,N_11710);
xnor U14133 (N_14133,N_8529,N_11231);
and U14134 (N_14134,N_11882,N_8968);
and U14135 (N_14135,N_8096,N_8666);
nor U14136 (N_14136,N_10817,N_10728);
and U14137 (N_14137,N_9822,N_10020);
or U14138 (N_14138,N_11303,N_8576);
nand U14139 (N_14139,N_11795,N_11829);
xnor U14140 (N_14140,N_10997,N_10311);
or U14141 (N_14141,N_9082,N_11752);
nand U14142 (N_14142,N_10362,N_10082);
nor U14143 (N_14143,N_9924,N_9380);
and U14144 (N_14144,N_8584,N_9742);
nor U14145 (N_14145,N_8938,N_8786);
and U14146 (N_14146,N_11356,N_10350);
nor U14147 (N_14147,N_10638,N_9235);
nor U14148 (N_14148,N_10182,N_10697);
or U14149 (N_14149,N_10699,N_11843);
and U14150 (N_14150,N_9610,N_11476);
or U14151 (N_14151,N_11690,N_8354);
nand U14152 (N_14152,N_11018,N_10358);
nand U14153 (N_14153,N_8384,N_11722);
and U14154 (N_14154,N_10484,N_8733);
and U14155 (N_14155,N_11855,N_10423);
or U14156 (N_14156,N_8120,N_10724);
and U14157 (N_14157,N_11930,N_10850);
nand U14158 (N_14158,N_8357,N_11508);
or U14159 (N_14159,N_10439,N_11214);
nor U14160 (N_14160,N_10287,N_8600);
nand U14161 (N_14161,N_8163,N_8217);
nand U14162 (N_14162,N_8617,N_8941);
and U14163 (N_14163,N_11176,N_11682);
or U14164 (N_14164,N_10741,N_8131);
and U14165 (N_14165,N_9606,N_8723);
nand U14166 (N_14166,N_10176,N_8167);
and U14167 (N_14167,N_11040,N_10545);
nor U14168 (N_14168,N_8932,N_10454);
nor U14169 (N_14169,N_11438,N_8898);
or U14170 (N_14170,N_8093,N_11243);
nor U14171 (N_14171,N_11526,N_11172);
nand U14172 (N_14172,N_11470,N_10059);
and U14173 (N_14173,N_11717,N_11031);
nor U14174 (N_14174,N_9029,N_9931);
nor U14175 (N_14175,N_8441,N_9416);
or U14176 (N_14176,N_8209,N_10733);
nand U14177 (N_14177,N_8810,N_10959);
or U14178 (N_14178,N_11903,N_10419);
or U14179 (N_14179,N_11883,N_8263);
and U14180 (N_14180,N_10902,N_8219);
or U14181 (N_14181,N_11891,N_11628);
nor U14182 (N_14182,N_10430,N_8714);
nand U14183 (N_14183,N_9544,N_10996);
nand U14184 (N_14184,N_11511,N_8528);
nor U14185 (N_14185,N_9321,N_8625);
and U14186 (N_14186,N_11937,N_9446);
nand U14187 (N_14187,N_9343,N_8797);
nand U14188 (N_14188,N_11071,N_8153);
nand U14189 (N_14189,N_8521,N_9531);
and U14190 (N_14190,N_9418,N_10435);
and U14191 (N_14191,N_11958,N_8807);
nand U14192 (N_14192,N_8344,N_9170);
and U14193 (N_14193,N_10802,N_10029);
nand U14194 (N_14194,N_8850,N_9008);
nor U14195 (N_14195,N_8017,N_9705);
nor U14196 (N_14196,N_8359,N_8450);
nand U14197 (N_14197,N_10285,N_11843);
nor U14198 (N_14198,N_10583,N_9539);
or U14199 (N_14199,N_10172,N_9942);
xnor U14200 (N_14200,N_10878,N_9527);
nor U14201 (N_14201,N_8518,N_8877);
xor U14202 (N_14202,N_9577,N_10483);
nand U14203 (N_14203,N_8829,N_8527);
or U14204 (N_14204,N_9191,N_10429);
nand U14205 (N_14205,N_9965,N_8557);
and U14206 (N_14206,N_10648,N_9236);
or U14207 (N_14207,N_9674,N_11150);
nor U14208 (N_14208,N_9966,N_10418);
and U14209 (N_14209,N_10017,N_11411);
nand U14210 (N_14210,N_9920,N_10318);
xor U14211 (N_14211,N_10938,N_10432);
or U14212 (N_14212,N_8912,N_8612);
or U14213 (N_14213,N_9887,N_8666);
nand U14214 (N_14214,N_8193,N_8543);
and U14215 (N_14215,N_8764,N_11348);
nand U14216 (N_14216,N_11970,N_8559);
nand U14217 (N_14217,N_9960,N_8005);
nor U14218 (N_14218,N_11309,N_9677);
nand U14219 (N_14219,N_9486,N_9515);
nand U14220 (N_14220,N_8560,N_9317);
or U14221 (N_14221,N_9709,N_8273);
and U14222 (N_14222,N_9111,N_10496);
and U14223 (N_14223,N_9874,N_10917);
and U14224 (N_14224,N_8578,N_8406);
nor U14225 (N_14225,N_8735,N_10142);
or U14226 (N_14226,N_8758,N_10632);
nand U14227 (N_14227,N_11563,N_11451);
nand U14228 (N_14228,N_9332,N_11685);
nor U14229 (N_14229,N_11980,N_9887);
nand U14230 (N_14230,N_10773,N_8830);
and U14231 (N_14231,N_11146,N_10454);
nor U14232 (N_14232,N_8232,N_10599);
and U14233 (N_14233,N_9965,N_11449);
nor U14234 (N_14234,N_10962,N_10862);
or U14235 (N_14235,N_11672,N_11611);
nand U14236 (N_14236,N_8164,N_8388);
nor U14237 (N_14237,N_10493,N_8991);
nand U14238 (N_14238,N_8892,N_9264);
nand U14239 (N_14239,N_11543,N_8449);
nor U14240 (N_14240,N_9815,N_10961);
or U14241 (N_14241,N_8976,N_8814);
or U14242 (N_14242,N_8297,N_8493);
or U14243 (N_14243,N_8414,N_8272);
nand U14244 (N_14244,N_8289,N_10706);
nor U14245 (N_14245,N_11464,N_9851);
or U14246 (N_14246,N_8221,N_10389);
or U14247 (N_14247,N_9737,N_8748);
and U14248 (N_14248,N_10077,N_8030);
or U14249 (N_14249,N_11714,N_10310);
and U14250 (N_14250,N_11117,N_9015);
nor U14251 (N_14251,N_8675,N_8969);
or U14252 (N_14252,N_10669,N_10722);
nand U14253 (N_14253,N_8331,N_9905);
and U14254 (N_14254,N_8223,N_8541);
and U14255 (N_14255,N_11561,N_9755);
nor U14256 (N_14256,N_8184,N_11995);
or U14257 (N_14257,N_9409,N_10702);
or U14258 (N_14258,N_8530,N_8662);
nor U14259 (N_14259,N_10577,N_8997);
or U14260 (N_14260,N_9477,N_11270);
or U14261 (N_14261,N_8195,N_11880);
or U14262 (N_14262,N_8713,N_8682);
nand U14263 (N_14263,N_10656,N_8443);
xnor U14264 (N_14264,N_10204,N_10160);
nand U14265 (N_14265,N_11383,N_9824);
nor U14266 (N_14266,N_9913,N_8394);
and U14267 (N_14267,N_8963,N_8016);
or U14268 (N_14268,N_9153,N_11461);
nor U14269 (N_14269,N_9624,N_8635);
or U14270 (N_14270,N_11613,N_11508);
and U14271 (N_14271,N_11790,N_9708);
or U14272 (N_14272,N_9937,N_9266);
xor U14273 (N_14273,N_9155,N_10371);
nand U14274 (N_14274,N_10993,N_9028);
and U14275 (N_14275,N_11287,N_10877);
or U14276 (N_14276,N_8890,N_11017);
nand U14277 (N_14277,N_9214,N_8821);
nand U14278 (N_14278,N_8803,N_11993);
or U14279 (N_14279,N_8391,N_9168);
nor U14280 (N_14280,N_8486,N_8840);
nand U14281 (N_14281,N_11112,N_8511);
nor U14282 (N_14282,N_11096,N_9307);
nor U14283 (N_14283,N_8693,N_8996);
nor U14284 (N_14284,N_11492,N_10399);
and U14285 (N_14285,N_10530,N_8862);
nor U14286 (N_14286,N_8433,N_8303);
and U14287 (N_14287,N_10747,N_8893);
nand U14288 (N_14288,N_8755,N_8183);
nor U14289 (N_14289,N_8729,N_11278);
or U14290 (N_14290,N_9298,N_10382);
nand U14291 (N_14291,N_10334,N_10396);
and U14292 (N_14292,N_10045,N_10975);
xor U14293 (N_14293,N_11895,N_11659);
nand U14294 (N_14294,N_8708,N_11077);
xnor U14295 (N_14295,N_10932,N_11497);
nand U14296 (N_14296,N_10705,N_8044);
nor U14297 (N_14297,N_11169,N_10702);
and U14298 (N_14298,N_11537,N_8531);
and U14299 (N_14299,N_10144,N_10959);
nand U14300 (N_14300,N_10251,N_9336);
nand U14301 (N_14301,N_9165,N_10727);
nor U14302 (N_14302,N_8951,N_8159);
nand U14303 (N_14303,N_9636,N_9224);
and U14304 (N_14304,N_9617,N_11921);
nand U14305 (N_14305,N_10395,N_8443);
nor U14306 (N_14306,N_11366,N_10762);
or U14307 (N_14307,N_10776,N_9873);
xor U14308 (N_14308,N_8336,N_8138);
nor U14309 (N_14309,N_8903,N_10839);
or U14310 (N_14310,N_9701,N_9607);
or U14311 (N_14311,N_10847,N_9257);
or U14312 (N_14312,N_10953,N_11588);
or U14313 (N_14313,N_11287,N_8990);
nor U14314 (N_14314,N_8459,N_10983);
nand U14315 (N_14315,N_11731,N_9857);
and U14316 (N_14316,N_8035,N_9687);
and U14317 (N_14317,N_9455,N_9325);
and U14318 (N_14318,N_9173,N_8206);
nand U14319 (N_14319,N_10650,N_8504);
or U14320 (N_14320,N_9190,N_11475);
nor U14321 (N_14321,N_9596,N_10451);
and U14322 (N_14322,N_10413,N_11992);
xnor U14323 (N_14323,N_10713,N_9566);
and U14324 (N_14324,N_8140,N_9727);
nand U14325 (N_14325,N_11933,N_10060);
xor U14326 (N_14326,N_9505,N_11126);
nand U14327 (N_14327,N_9793,N_8483);
and U14328 (N_14328,N_9810,N_10788);
xor U14329 (N_14329,N_11564,N_10542);
nor U14330 (N_14330,N_11238,N_8904);
and U14331 (N_14331,N_11698,N_10225);
xor U14332 (N_14332,N_11983,N_10472);
and U14333 (N_14333,N_11734,N_8734);
xor U14334 (N_14334,N_11655,N_9424);
xnor U14335 (N_14335,N_11630,N_9829);
nor U14336 (N_14336,N_8110,N_11445);
or U14337 (N_14337,N_11688,N_10896);
nor U14338 (N_14338,N_11592,N_11769);
nand U14339 (N_14339,N_8948,N_8557);
nor U14340 (N_14340,N_10921,N_10177);
and U14341 (N_14341,N_9872,N_8633);
nand U14342 (N_14342,N_10553,N_11290);
nand U14343 (N_14343,N_8975,N_8594);
xnor U14344 (N_14344,N_10457,N_8856);
xnor U14345 (N_14345,N_9490,N_11405);
and U14346 (N_14346,N_8275,N_11967);
nand U14347 (N_14347,N_9639,N_10827);
nor U14348 (N_14348,N_10823,N_8999);
and U14349 (N_14349,N_9143,N_8541);
and U14350 (N_14350,N_10609,N_10740);
or U14351 (N_14351,N_8028,N_11604);
and U14352 (N_14352,N_9754,N_8452);
and U14353 (N_14353,N_9200,N_8119);
and U14354 (N_14354,N_11452,N_9431);
nor U14355 (N_14355,N_8764,N_8242);
nand U14356 (N_14356,N_9876,N_8056);
and U14357 (N_14357,N_8648,N_8202);
nand U14358 (N_14358,N_9617,N_9532);
or U14359 (N_14359,N_11304,N_11806);
nor U14360 (N_14360,N_11405,N_8966);
and U14361 (N_14361,N_10218,N_11497);
or U14362 (N_14362,N_9065,N_8997);
nor U14363 (N_14363,N_8776,N_11699);
and U14364 (N_14364,N_11074,N_10849);
nor U14365 (N_14365,N_10841,N_10137);
nor U14366 (N_14366,N_11900,N_8695);
nor U14367 (N_14367,N_8611,N_9176);
nor U14368 (N_14368,N_9296,N_8248);
xor U14369 (N_14369,N_10763,N_10484);
nor U14370 (N_14370,N_9120,N_11832);
nand U14371 (N_14371,N_9528,N_11986);
nor U14372 (N_14372,N_11192,N_11204);
or U14373 (N_14373,N_10237,N_8041);
nand U14374 (N_14374,N_10934,N_11988);
nand U14375 (N_14375,N_9915,N_9423);
nor U14376 (N_14376,N_9988,N_9980);
nor U14377 (N_14377,N_11128,N_9155);
nor U14378 (N_14378,N_11030,N_10288);
xnor U14379 (N_14379,N_11276,N_10027);
nand U14380 (N_14380,N_9709,N_8405);
and U14381 (N_14381,N_8949,N_10370);
and U14382 (N_14382,N_9325,N_8322);
and U14383 (N_14383,N_9357,N_11621);
xor U14384 (N_14384,N_9180,N_10354);
nand U14385 (N_14385,N_8228,N_11907);
or U14386 (N_14386,N_10668,N_9239);
nand U14387 (N_14387,N_8502,N_9231);
and U14388 (N_14388,N_8446,N_8238);
nand U14389 (N_14389,N_11714,N_9443);
or U14390 (N_14390,N_10263,N_9857);
and U14391 (N_14391,N_8282,N_11932);
or U14392 (N_14392,N_8460,N_11840);
and U14393 (N_14393,N_11100,N_8896);
nand U14394 (N_14394,N_9006,N_11020);
or U14395 (N_14395,N_10715,N_8772);
nor U14396 (N_14396,N_9199,N_9165);
or U14397 (N_14397,N_11248,N_11109);
xnor U14398 (N_14398,N_9493,N_8216);
or U14399 (N_14399,N_10033,N_9831);
nand U14400 (N_14400,N_8782,N_9449);
nor U14401 (N_14401,N_9181,N_11921);
and U14402 (N_14402,N_8238,N_8833);
nor U14403 (N_14403,N_8063,N_10855);
nand U14404 (N_14404,N_10880,N_8395);
nor U14405 (N_14405,N_8024,N_10495);
nand U14406 (N_14406,N_10850,N_9844);
or U14407 (N_14407,N_10104,N_8531);
nor U14408 (N_14408,N_9025,N_10936);
nand U14409 (N_14409,N_9925,N_9398);
nor U14410 (N_14410,N_8756,N_11170);
nor U14411 (N_14411,N_11812,N_11888);
nor U14412 (N_14412,N_8402,N_8976);
or U14413 (N_14413,N_10996,N_8334);
or U14414 (N_14414,N_10829,N_9151);
nor U14415 (N_14415,N_10936,N_9189);
nand U14416 (N_14416,N_8017,N_9101);
or U14417 (N_14417,N_11507,N_11221);
and U14418 (N_14418,N_8261,N_11908);
nor U14419 (N_14419,N_11865,N_9719);
nor U14420 (N_14420,N_9245,N_11946);
or U14421 (N_14421,N_10270,N_8677);
or U14422 (N_14422,N_10592,N_8985);
nand U14423 (N_14423,N_9961,N_8043);
nand U14424 (N_14424,N_9914,N_11809);
nand U14425 (N_14425,N_9333,N_9526);
nor U14426 (N_14426,N_8727,N_8384);
or U14427 (N_14427,N_9458,N_10604);
and U14428 (N_14428,N_11775,N_10704);
nand U14429 (N_14429,N_8719,N_9592);
nor U14430 (N_14430,N_10840,N_8624);
or U14431 (N_14431,N_11860,N_11808);
and U14432 (N_14432,N_9484,N_11683);
and U14433 (N_14433,N_11627,N_8130);
or U14434 (N_14434,N_9127,N_10438);
and U14435 (N_14435,N_11748,N_8791);
and U14436 (N_14436,N_8823,N_10449);
and U14437 (N_14437,N_8182,N_11294);
nand U14438 (N_14438,N_8461,N_8268);
or U14439 (N_14439,N_9198,N_11131);
or U14440 (N_14440,N_9501,N_11024);
or U14441 (N_14441,N_8869,N_11917);
and U14442 (N_14442,N_11338,N_10881);
nand U14443 (N_14443,N_10497,N_9112);
xor U14444 (N_14444,N_8343,N_8996);
nor U14445 (N_14445,N_10953,N_10133);
xnor U14446 (N_14446,N_10723,N_11810);
nand U14447 (N_14447,N_9949,N_9854);
xnor U14448 (N_14448,N_10887,N_10356);
xnor U14449 (N_14449,N_9629,N_9223);
nand U14450 (N_14450,N_8686,N_11688);
nand U14451 (N_14451,N_9292,N_11055);
nor U14452 (N_14452,N_11886,N_10536);
nand U14453 (N_14453,N_9992,N_9777);
nand U14454 (N_14454,N_8736,N_11049);
or U14455 (N_14455,N_11695,N_8890);
nor U14456 (N_14456,N_9014,N_9981);
nand U14457 (N_14457,N_11197,N_10302);
and U14458 (N_14458,N_8587,N_11685);
and U14459 (N_14459,N_11712,N_9411);
nand U14460 (N_14460,N_8216,N_8682);
nand U14461 (N_14461,N_11609,N_10529);
or U14462 (N_14462,N_11421,N_8380);
nand U14463 (N_14463,N_10592,N_10014);
or U14464 (N_14464,N_8552,N_11046);
and U14465 (N_14465,N_8694,N_8066);
and U14466 (N_14466,N_8192,N_10880);
nand U14467 (N_14467,N_8889,N_11779);
or U14468 (N_14468,N_10117,N_11345);
and U14469 (N_14469,N_11945,N_8933);
nand U14470 (N_14470,N_10033,N_9802);
or U14471 (N_14471,N_8569,N_8533);
nand U14472 (N_14472,N_9213,N_10538);
or U14473 (N_14473,N_8897,N_11087);
and U14474 (N_14474,N_8566,N_11243);
nand U14475 (N_14475,N_11093,N_10299);
or U14476 (N_14476,N_10838,N_8639);
and U14477 (N_14477,N_9088,N_8781);
nor U14478 (N_14478,N_9742,N_10007);
nor U14479 (N_14479,N_9620,N_10060);
nor U14480 (N_14480,N_11367,N_11315);
xor U14481 (N_14481,N_9268,N_8337);
nand U14482 (N_14482,N_10556,N_9663);
nand U14483 (N_14483,N_11271,N_11970);
nor U14484 (N_14484,N_10568,N_11878);
nand U14485 (N_14485,N_10035,N_8459);
nor U14486 (N_14486,N_9444,N_10364);
nand U14487 (N_14487,N_10513,N_10224);
or U14488 (N_14488,N_11387,N_9648);
nor U14489 (N_14489,N_11405,N_9779);
or U14490 (N_14490,N_8072,N_11349);
and U14491 (N_14491,N_11240,N_11027);
and U14492 (N_14492,N_8514,N_8229);
nor U14493 (N_14493,N_10370,N_9109);
and U14494 (N_14494,N_11605,N_8467);
or U14495 (N_14495,N_9584,N_10276);
or U14496 (N_14496,N_11743,N_10266);
nand U14497 (N_14497,N_10688,N_10486);
and U14498 (N_14498,N_11811,N_9878);
or U14499 (N_14499,N_11646,N_11472);
or U14500 (N_14500,N_9492,N_8019);
xnor U14501 (N_14501,N_10611,N_10534);
xor U14502 (N_14502,N_11666,N_10726);
and U14503 (N_14503,N_11487,N_10546);
nor U14504 (N_14504,N_11319,N_10850);
and U14505 (N_14505,N_9242,N_10257);
xor U14506 (N_14506,N_8476,N_10997);
xnor U14507 (N_14507,N_8685,N_11615);
and U14508 (N_14508,N_11718,N_10239);
or U14509 (N_14509,N_9041,N_9064);
and U14510 (N_14510,N_11077,N_11359);
and U14511 (N_14511,N_10400,N_11349);
and U14512 (N_14512,N_9442,N_10595);
xnor U14513 (N_14513,N_11452,N_10792);
nand U14514 (N_14514,N_10404,N_9829);
and U14515 (N_14515,N_10857,N_11670);
nand U14516 (N_14516,N_10300,N_10482);
nor U14517 (N_14517,N_11018,N_9151);
nor U14518 (N_14518,N_9366,N_8316);
or U14519 (N_14519,N_11793,N_11646);
or U14520 (N_14520,N_8069,N_8473);
nand U14521 (N_14521,N_9950,N_8995);
or U14522 (N_14522,N_8098,N_9963);
nor U14523 (N_14523,N_11056,N_11987);
or U14524 (N_14524,N_11225,N_10997);
and U14525 (N_14525,N_8481,N_9462);
and U14526 (N_14526,N_11506,N_9824);
nor U14527 (N_14527,N_11350,N_11358);
or U14528 (N_14528,N_10863,N_11381);
nor U14529 (N_14529,N_11509,N_11818);
or U14530 (N_14530,N_8170,N_8503);
nand U14531 (N_14531,N_9313,N_8067);
xnor U14532 (N_14532,N_9187,N_10575);
nand U14533 (N_14533,N_11857,N_9843);
nand U14534 (N_14534,N_10082,N_10610);
and U14535 (N_14535,N_11324,N_8022);
nor U14536 (N_14536,N_8738,N_11803);
and U14537 (N_14537,N_8223,N_9899);
nand U14538 (N_14538,N_8497,N_10355);
nand U14539 (N_14539,N_9198,N_9797);
and U14540 (N_14540,N_11864,N_10687);
nor U14541 (N_14541,N_9809,N_9852);
nand U14542 (N_14542,N_11743,N_10554);
and U14543 (N_14543,N_8128,N_10308);
nand U14544 (N_14544,N_11808,N_8830);
nor U14545 (N_14545,N_9505,N_10645);
and U14546 (N_14546,N_8073,N_9799);
nor U14547 (N_14547,N_10629,N_9443);
xor U14548 (N_14548,N_8064,N_11185);
or U14549 (N_14549,N_9087,N_11304);
nor U14550 (N_14550,N_11934,N_9617);
or U14551 (N_14551,N_11015,N_9056);
and U14552 (N_14552,N_8805,N_8374);
and U14553 (N_14553,N_9336,N_8564);
nand U14554 (N_14554,N_9102,N_11759);
nor U14555 (N_14555,N_9634,N_10047);
or U14556 (N_14556,N_8155,N_11291);
and U14557 (N_14557,N_8597,N_11892);
nand U14558 (N_14558,N_9221,N_8595);
or U14559 (N_14559,N_11195,N_9713);
nand U14560 (N_14560,N_11336,N_11438);
or U14561 (N_14561,N_9721,N_11716);
and U14562 (N_14562,N_10912,N_10330);
or U14563 (N_14563,N_11987,N_9900);
nor U14564 (N_14564,N_11610,N_10360);
nand U14565 (N_14565,N_11957,N_8570);
nand U14566 (N_14566,N_9257,N_10860);
or U14567 (N_14567,N_9482,N_11651);
xnor U14568 (N_14568,N_8362,N_10271);
nor U14569 (N_14569,N_8253,N_10230);
nand U14570 (N_14570,N_9377,N_9013);
and U14571 (N_14571,N_8578,N_8757);
nor U14572 (N_14572,N_8815,N_11449);
nor U14573 (N_14573,N_10368,N_9953);
nor U14574 (N_14574,N_10453,N_10496);
nor U14575 (N_14575,N_10576,N_10064);
and U14576 (N_14576,N_10252,N_8687);
nor U14577 (N_14577,N_10682,N_10468);
and U14578 (N_14578,N_8624,N_9110);
or U14579 (N_14579,N_9369,N_9232);
nand U14580 (N_14580,N_8127,N_11269);
xnor U14581 (N_14581,N_9668,N_9100);
nor U14582 (N_14582,N_11179,N_8598);
nand U14583 (N_14583,N_10209,N_11603);
nand U14584 (N_14584,N_9683,N_11179);
and U14585 (N_14585,N_10138,N_8659);
and U14586 (N_14586,N_8311,N_9833);
nand U14587 (N_14587,N_11899,N_11322);
nor U14588 (N_14588,N_10428,N_9734);
nand U14589 (N_14589,N_8104,N_11019);
nor U14590 (N_14590,N_11923,N_8355);
nand U14591 (N_14591,N_11485,N_11221);
and U14592 (N_14592,N_8109,N_9914);
or U14593 (N_14593,N_8971,N_8950);
nand U14594 (N_14594,N_8687,N_8098);
xnor U14595 (N_14595,N_9458,N_11144);
nand U14596 (N_14596,N_10948,N_11966);
or U14597 (N_14597,N_10721,N_11939);
or U14598 (N_14598,N_11010,N_9065);
nor U14599 (N_14599,N_9210,N_11809);
nor U14600 (N_14600,N_10589,N_11381);
or U14601 (N_14601,N_8958,N_9539);
xor U14602 (N_14602,N_11617,N_10091);
nand U14603 (N_14603,N_9590,N_10222);
xnor U14604 (N_14604,N_8481,N_11584);
nand U14605 (N_14605,N_8146,N_9271);
or U14606 (N_14606,N_9955,N_11692);
and U14607 (N_14607,N_10831,N_9793);
nor U14608 (N_14608,N_8787,N_9901);
nand U14609 (N_14609,N_11282,N_9701);
nand U14610 (N_14610,N_9731,N_9390);
or U14611 (N_14611,N_9434,N_9686);
or U14612 (N_14612,N_11289,N_8860);
or U14613 (N_14613,N_11952,N_8775);
nor U14614 (N_14614,N_9928,N_8669);
xnor U14615 (N_14615,N_9772,N_10417);
nand U14616 (N_14616,N_10810,N_8871);
nor U14617 (N_14617,N_8219,N_9483);
or U14618 (N_14618,N_11658,N_11458);
or U14619 (N_14619,N_11059,N_9254);
and U14620 (N_14620,N_10634,N_8058);
nor U14621 (N_14621,N_11174,N_10052);
or U14622 (N_14622,N_10515,N_10926);
nor U14623 (N_14623,N_8653,N_9646);
xnor U14624 (N_14624,N_10534,N_10411);
xnor U14625 (N_14625,N_10353,N_10575);
or U14626 (N_14626,N_9231,N_10550);
nor U14627 (N_14627,N_11578,N_9006);
nor U14628 (N_14628,N_8258,N_9124);
and U14629 (N_14629,N_11953,N_8337);
nor U14630 (N_14630,N_10197,N_8377);
and U14631 (N_14631,N_11813,N_9589);
and U14632 (N_14632,N_11434,N_11684);
and U14633 (N_14633,N_10536,N_8726);
and U14634 (N_14634,N_8553,N_11268);
or U14635 (N_14635,N_9160,N_10723);
nand U14636 (N_14636,N_11580,N_11931);
nand U14637 (N_14637,N_10272,N_8827);
or U14638 (N_14638,N_8016,N_11754);
and U14639 (N_14639,N_8593,N_11108);
or U14640 (N_14640,N_11198,N_9204);
or U14641 (N_14641,N_8391,N_11797);
nor U14642 (N_14642,N_10535,N_8561);
xnor U14643 (N_14643,N_11867,N_9415);
nor U14644 (N_14644,N_9625,N_8020);
xnor U14645 (N_14645,N_11768,N_8412);
nand U14646 (N_14646,N_11100,N_10964);
and U14647 (N_14647,N_9179,N_9417);
nor U14648 (N_14648,N_8265,N_9445);
xor U14649 (N_14649,N_11403,N_11414);
or U14650 (N_14650,N_8248,N_9943);
and U14651 (N_14651,N_11451,N_9711);
nand U14652 (N_14652,N_8474,N_8273);
or U14653 (N_14653,N_9182,N_11930);
nor U14654 (N_14654,N_9237,N_11137);
nor U14655 (N_14655,N_9735,N_9739);
nand U14656 (N_14656,N_11617,N_10159);
and U14657 (N_14657,N_9004,N_11020);
nand U14658 (N_14658,N_10218,N_8754);
and U14659 (N_14659,N_8961,N_9171);
or U14660 (N_14660,N_8099,N_9765);
nor U14661 (N_14661,N_9737,N_9799);
nand U14662 (N_14662,N_9305,N_9335);
or U14663 (N_14663,N_11530,N_10854);
and U14664 (N_14664,N_9263,N_9221);
nand U14665 (N_14665,N_11851,N_8700);
and U14666 (N_14666,N_10777,N_9327);
nand U14667 (N_14667,N_9540,N_10049);
and U14668 (N_14668,N_10818,N_11723);
nand U14669 (N_14669,N_11803,N_9996);
nor U14670 (N_14670,N_8835,N_10995);
nor U14671 (N_14671,N_8969,N_11538);
xnor U14672 (N_14672,N_8006,N_8941);
nand U14673 (N_14673,N_8251,N_11310);
or U14674 (N_14674,N_8159,N_9541);
nor U14675 (N_14675,N_10475,N_10238);
nand U14676 (N_14676,N_10742,N_9177);
nand U14677 (N_14677,N_9647,N_10614);
nor U14678 (N_14678,N_11179,N_11002);
and U14679 (N_14679,N_10353,N_10274);
nand U14680 (N_14680,N_9335,N_10214);
nor U14681 (N_14681,N_10639,N_10479);
or U14682 (N_14682,N_11025,N_10386);
nand U14683 (N_14683,N_9293,N_8261);
nor U14684 (N_14684,N_11756,N_8397);
nand U14685 (N_14685,N_11176,N_9544);
or U14686 (N_14686,N_9161,N_11092);
nand U14687 (N_14687,N_9225,N_9667);
and U14688 (N_14688,N_10479,N_9185);
or U14689 (N_14689,N_10526,N_10037);
nor U14690 (N_14690,N_10411,N_10317);
nand U14691 (N_14691,N_9212,N_11966);
xor U14692 (N_14692,N_10447,N_11215);
xor U14693 (N_14693,N_8717,N_9232);
and U14694 (N_14694,N_8400,N_9214);
nor U14695 (N_14695,N_11205,N_10272);
nand U14696 (N_14696,N_9763,N_10581);
nand U14697 (N_14697,N_11072,N_8444);
and U14698 (N_14698,N_9348,N_8965);
and U14699 (N_14699,N_10499,N_9600);
nand U14700 (N_14700,N_10769,N_10693);
and U14701 (N_14701,N_8044,N_10867);
and U14702 (N_14702,N_9820,N_8704);
and U14703 (N_14703,N_9149,N_10043);
nand U14704 (N_14704,N_9079,N_9997);
nor U14705 (N_14705,N_11611,N_9806);
or U14706 (N_14706,N_9802,N_11762);
or U14707 (N_14707,N_11188,N_8053);
and U14708 (N_14708,N_10045,N_9445);
and U14709 (N_14709,N_8771,N_10175);
or U14710 (N_14710,N_11772,N_10931);
nand U14711 (N_14711,N_8948,N_9711);
nand U14712 (N_14712,N_11798,N_8722);
nor U14713 (N_14713,N_11345,N_11740);
or U14714 (N_14714,N_10820,N_10749);
nand U14715 (N_14715,N_10505,N_9053);
xnor U14716 (N_14716,N_10006,N_11999);
or U14717 (N_14717,N_10609,N_9588);
or U14718 (N_14718,N_8737,N_8311);
nor U14719 (N_14719,N_9253,N_8470);
and U14720 (N_14720,N_9834,N_10313);
or U14721 (N_14721,N_10453,N_8014);
and U14722 (N_14722,N_10793,N_8680);
or U14723 (N_14723,N_9281,N_10097);
or U14724 (N_14724,N_10179,N_8370);
nand U14725 (N_14725,N_8425,N_10085);
nand U14726 (N_14726,N_8449,N_11115);
and U14727 (N_14727,N_10234,N_9446);
or U14728 (N_14728,N_9506,N_11871);
nand U14729 (N_14729,N_11161,N_10332);
and U14730 (N_14730,N_11627,N_11413);
nor U14731 (N_14731,N_8696,N_9001);
or U14732 (N_14732,N_9608,N_8729);
or U14733 (N_14733,N_10646,N_8850);
or U14734 (N_14734,N_9136,N_9799);
and U14735 (N_14735,N_8997,N_11392);
nand U14736 (N_14736,N_9649,N_11311);
nand U14737 (N_14737,N_8083,N_11699);
and U14738 (N_14738,N_10041,N_8654);
nand U14739 (N_14739,N_9619,N_8146);
and U14740 (N_14740,N_10747,N_10471);
or U14741 (N_14741,N_9987,N_8205);
nor U14742 (N_14742,N_11765,N_9106);
and U14743 (N_14743,N_10396,N_8504);
xor U14744 (N_14744,N_9195,N_11402);
nand U14745 (N_14745,N_9148,N_8033);
and U14746 (N_14746,N_9170,N_9475);
and U14747 (N_14747,N_10933,N_10592);
nand U14748 (N_14748,N_9981,N_8198);
nand U14749 (N_14749,N_8729,N_8356);
or U14750 (N_14750,N_8066,N_9714);
xnor U14751 (N_14751,N_9668,N_9277);
xor U14752 (N_14752,N_11074,N_10083);
and U14753 (N_14753,N_9679,N_8063);
and U14754 (N_14754,N_10542,N_8581);
or U14755 (N_14755,N_10574,N_11673);
and U14756 (N_14756,N_11095,N_10360);
nor U14757 (N_14757,N_8103,N_9269);
nor U14758 (N_14758,N_11877,N_11081);
and U14759 (N_14759,N_9187,N_11620);
nand U14760 (N_14760,N_9464,N_10315);
and U14761 (N_14761,N_8257,N_11958);
nand U14762 (N_14762,N_10656,N_9029);
and U14763 (N_14763,N_11562,N_8648);
or U14764 (N_14764,N_9623,N_10689);
nor U14765 (N_14765,N_10564,N_8442);
nand U14766 (N_14766,N_9076,N_10502);
nand U14767 (N_14767,N_11213,N_10118);
and U14768 (N_14768,N_9233,N_9712);
nand U14769 (N_14769,N_8111,N_9845);
nand U14770 (N_14770,N_9064,N_10605);
or U14771 (N_14771,N_10497,N_8145);
and U14772 (N_14772,N_8616,N_9907);
and U14773 (N_14773,N_8998,N_11717);
nand U14774 (N_14774,N_9296,N_10445);
or U14775 (N_14775,N_9805,N_10150);
nand U14776 (N_14776,N_10938,N_9938);
or U14777 (N_14777,N_8249,N_9596);
and U14778 (N_14778,N_11097,N_8223);
or U14779 (N_14779,N_10436,N_10668);
nor U14780 (N_14780,N_9370,N_8931);
and U14781 (N_14781,N_8350,N_10034);
nand U14782 (N_14782,N_9240,N_9490);
nand U14783 (N_14783,N_11282,N_11585);
and U14784 (N_14784,N_8304,N_10850);
nand U14785 (N_14785,N_10379,N_9889);
xor U14786 (N_14786,N_10723,N_10094);
nand U14787 (N_14787,N_9687,N_9365);
nor U14788 (N_14788,N_11299,N_10481);
nor U14789 (N_14789,N_11623,N_9167);
and U14790 (N_14790,N_10914,N_8697);
or U14791 (N_14791,N_11140,N_8880);
nand U14792 (N_14792,N_8115,N_10137);
or U14793 (N_14793,N_8480,N_9056);
or U14794 (N_14794,N_8053,N_9842);
nor U14795 (N_14795,N_8163,N_10479);
nand U14796 (N_14796,N_8800,N_9220);
or U14797 (N_14797,N_10420,N_10588);
nor U14798 (N_14798,N_9064,N_11224);
or U14799 (N_14799,N_8950,N_8960);
and U14800 (N_14800,N_11474,N_10300);
nand U14801 (N_14801,N_9872,N_10956);
or U14802 (N_14802,N_10611,N_9010);
or U14803 (N_14803,N_8603,N_8644);
and U14804 (N_14804,N_11637,N_11708);
and U14805 (N_14805,N_10642,N_8198);
and U14806 (N_14806,N_10601,N_10899);
nor U14807 (N_14807,N_10390,N_8096);
nand U14808 (N_14808,N_9662,N_8834);
nor U14809 (N_14809,N_11595,N_11820);
nand U14810 (N_14810,N_11086,N_8855);
or U14811 (N_14811,N_10361,N_10896);
or U14812 (N_14812,N_8097,N_11892);
and U14813 (N_14813,N_11627,N_10018);
and U14814 (N_14814,N_9068,N_8824);
xnor U14815 (N_14815,N_9620,N_11846);
and U14816 (N_14816,N_11299,N_9772);
nand U14817 (N_14817,N_9299,N_8898);
nand U14818 (N_14818,N_9457,N_9147);
and U14819 (N_14819,N_9275,N_10586);
nand U14820 (N_14820,N_9588,N_8422);
and U14821 (N_14821,N_8283,N_10906);
or U14822 (N_14822,N_9688,N_11755);
and U14823 (N_14823,N_8072,N_9797);
and U14824 (N_14824,N_11007,N_10691);
or U14825 (N_14825,N_11198,N_11141);
nor U14826 (N_14826,N_10283,N_11598);
nor U14827 (N_14827,N_8774,N_10764);
and U14828 (N_14828,N_11177,N_9859);
and U14829 (N_14829,N_8761,N_9214);
nor U14830 (N_14830,N_9201,N_9687);
or U14831 (N_14831,N_11960,N_8643);
or U14832 (N_14832,N_8729,N_10532);
or U14833 (N_14833,N_9695,N_11357);
nand U14834 (N_14834,N_10494,N_9468);
or U14835 (N_14835,N_11890,N_10393);
or U14836 (N_14836,N_10515,N_9968);
and U14837 (N_14837,N_9298,N_9536);
nor U14838 (N_14838,N_8752,N_10256);
nor U14839 (N_14839,N_9104,N_10858);
or U14840 (N_14840,N_10162,N_9466);
and U14841 (N_14841,N_11254,N_10136);
nand U14842 (N_14842,N_10290,N_9169);
xnor U14843 (N_14843,N_10549,N_11916);
or U14844 (N_14844,N_8729,N_10970);
nand U14845 (N_14845,N_8247,N_11280);
and U14846 (N_14846,N_11776,N_8205);
nand U14847 (N_14847,N_10335,N_8209);
or U14848 (N_14848,N_8191,N_9974);
or U14849 (N_14849,N_8501,N_11993);
or U14850 (N_14850,N_8287,N_10056);
nand U14851 (N_14851,N_9577,N_11022);
nor U14852 (N_14852,N_10205,N_9809);
nand U14853 (N_14853,N_11373,N_8538);
and U14854 (N_14854,N_9399,N_8519);
or U14855 (N_14855,N_8122,N_8906);
and U14856 (N_14856,N_11691,N_8429);
or U14857 (N_14857,N_11192,N_11789);
or U14858 (N_14858,N_10307,N_10002);
and U14859 (N_14859,N_9523,N_11261);
nand U14860 (N_14860,N_10962,N_9092);
xnor U14861 (N_14861,N_9192,N_11925);
or U14862 (N_14862,N_9011,N_11799);
nand U14863 (N_14863,N_10962,N_9990);
nor U14864 (N_14864,N_9412,N_8049);
nor U14865 (N_14865,N_10235,N_11371);
nor U14866 (N_14866,N_10676,N_10366);
or U14867 (N_14867,N_11494,N_9895);
or U14868 (N_14868,N_9292,N_8033);
nand U14869 (N_14869,N_8241,N_11389);
and U14870 (N_14870,N_8815,N_8810);
or U14871 (N_14871,N_11813,N_8125);
or U14872 (N_14872,N_10635,N_8194);
nand U14873 (N_14873,N_9307,N_10253);
nand U14874 (N_14874,N_11592,N_9408);
and U14875 (N_14875,N_11101,N_11074);
or U14876 (N_14876,N_10743,N_11220);
nand U14877 (N_14877,N_10091,N_9936);
and U14878 (N_14878,N_11193,N_8365);
or U14879 (N_14879,N_10241,N_9340);
and U14880 (N_14880,N_8012,N_11544);
nor U14881 (N_14881,N_9321,N_9717);
xnor U14882 (N_14882,N_9893,N_10647);
and U14883 (N_14883,N_10750,N_9855);
xor U14884 (N_14884,N_10651,N_11214);
or U14885 (N_14885,N_9313,N_10232);
nand U14886 (N_14886,N_11600,N_8752);
nand U14887 (N_14887,N_10979,N_11922);
and U14888 (N_14888,N_8543,N_9049);
and U14889 (N_14889,N_11091,N_11260);
or U14890 (N_14890,N_8239,N_8289);
or U14891 (N_14891,N_10838,N_8452);
xor U14892 (N_14892,N_9468,N_11353);
nand U14893 (N_14893,N_8728,N_9418);
or U14894 (N_14894,N_10093,N_11918);
nor U14895 (N_14895,N_11245,N_10811);
xor U14896 (N_14896,N_9063,N_11958);
nor U14897 (N_14897,N_10555,N_11453);
nand U14898 (N_14898,N_11779,N_10531);
nand U14899 (N_14899,N_10294,N_9657);
and U14900 (N_14900,N_8832,N_9966);
and U14901 (N_14901,N_11148,N_11427);
nor U14902 (N_14902,N_8116,N_9795);
nor U14903 (N_14903,N_10322,N_9465);
nor U14904 (N_14904,N_8051,N_10282);
or U14905 (N_14905,N_11565,N_9693);
or U14906 (N_14906,N_9232,N_8975);
nand U14907 (N_14907,N_10924,N_8119);
and U14908 (N_14908,N_9067,N_8052);
or U14909 (N_14909,N_9228,N_9579);
nand U14910 (N_14910,N_8608,N_9498);
nor U14911 (N_14911,N_11344,N_8182);
and U14912 (N_14912,N_8745,N_11454);
nand U14913 (N_14913,N_11986,N_10316);
nand U14914 (N_14914,N_9317,N_9655);
or U14915 (N_14915,N_11033,N_9938);
or U14916 (N_14916,N_8422,N_11358);
nand U14917 (N_14917,N_10575,N_8719);
and U14918 (N_14918,N_11699,N_8003);
nand U14919 (N_14919,N_9006,N_8815);
or U14920 (N_14920,N_10206,N_10226);
nor U14921 (N_14921,N_10341,N_11798);
or U14922 (N_14922,N_11012,N_11490);
nor U14923 (N_14923,N_11237,N_11535);
or U14924 (N_14924,N_10698,N_10515);
or U14925 (N_14925,N_9048,N_10748);
or U14926 (N_14926,N_11000,N_8473);
nor U14927 (N_14927,N_11063,N_11742);
nor U14928 (N_14928,N_9761,N_9585);
nand U14929 (N_14929,N_10103,N_11137);
nor U14930 (N_14930,N_10249,N_10059);
or U14931 (N_14931,N_11491,N_9700);
and U14932 (N_14932,N_8959,N_9236);
or U14933 (N_14933,N_11287,N_9519);
nand U14934 (N_14934,N_8655,N_10933);
and U14935 (N_14935,N_9657,N_9622);
or U14936 (N_14936,N_10622,N_10697);
xnor U14937 (N_14937,N_11381,N_8725);
nand U14938 (N_14938,N_10000,N_11940);
nand U14939 (N_14939,N_9164,N_8813);
and U14940 (N_14940,N_9509,N_11469);
nand U14941 (N_14941,N_9844,N_8677);
xnor U14942 (N_14942,N_9711,N_8889);
nor U14943 (N_14943,N_8816,N_8052);
or U14944 (N_14944,N_11278,N_9265);
nand U14945 (N_14945,N_11519,N_8394);
nor U14946 (N_14946,N_8407,N_9818);
or U14947 (N_14947,N_9284,N_9524);
or U14948 (N_14948,N_10620,N_8842);
nor U14949 (N_14949,N_11420,N_11288);
or U14950 (N_14950,N_10981,N_8047);
xor U14951 (N_14951,N_10115,N_9041);
nor U14952 (N_14952,N_10133,N_10530);
and U14953 (N_14953,N_11404,N_11715);
and U14954 (N_14954,N_8072,N_11388);
or U14955 (N_14955,N_8214,N_9451);
and U14956 (N_14956,N_8119,N_9668);
and U14957 (N_14957,N_9602,N_9434);
and U14958 (N_14958,N_8427,N_9925);
xor U14959 (N_14959,N_8246,N_9457);
and U14960 (N_14960,N_9825,N_11812);
or U14961 (N_14961,N_8438,N_9443);
and U14962 (N_14962,N_11633,N_10625);
nand U14963 (N_14963,N_9426,N_10115);
nor U14964 (N_14964,N_8149,N_8300);
or U14965 (N_14965,N_8679,N_8647);
and U14966 (N_14966,N_9466,N_11160);
nor U14967 (N_14967,N_11766,N_10005);
nand U14968 (N_14968,N_9572,N_8473);
nand U14969 (N_14969,N_8020,N_8168);
and U14970 (N_14970,N_10237,N_9569);
nand U14971 (N_14971,N_8149,N_8594);
or U14972 (N_14972,N_10828,N_10751);
and U14973 (N_14973,N_10570,N_8619);
or U14974 (N_14974,N_10087,N_11012);
nor U14975 (N_14975,N_11116,N_10551);
and U14976 (N_14976,N_8011,N_11420);
nor U14977 (N_14977,N_8094,N_9427);
xnor U14978 (N_14978,N_8851,N_9003);
nor U14979 (N_14979,N_8590,N_11779);
nand U14980 (N_14980,N_11648,N_8871);
xor U14981 (N_14981,N_8697,N_8227);
xnor U14982 (N_14982,N_8757,N_8915);
nand U14983 (N_14983,N_9686,N_8973);
nand U14984 (N_14984,N_11356,N_8949);
and U14985 (N_14985,N_10961,N_8901);
nand U14986 (N_14986,N_11299,N_9461);
nor U14987 (N_14987,N_10844,N_10464);
or U14988 (N_14988,N_9611,N_11824);
nor U14989 (N_14989,N_11146,N_11829);
nand U14990 (N_14990,N_10531,N_11965);
xnor U14991 (N_14991,N_9014,N_10131);
nor U14992 (N_14992,N_8854,N_11215);
and U14993 (N_14993,N_10661,N_8925);
or U14994 (N_14994,N_9277,N_11898);
or U14995 (N_14995,N_10350,N_11141);
or U14996 (N_14996,N_11736,N_8584);
xnor U14997 (N_14997,N_10982,N_9093);
or U14998 (N_14998,N_8608,N_10846);
or U14999 (N_14999,N_9865,N_9620);
nand U15000 (N_15000,N_8221,N_11779);
nor U15001 (N_15001,N_10918,N_10891);
and U15002 (N_15002,N_10761,N_9794);
xnor U15003 (N_15003,N_11821,N_8882);
nand U15004 (N_15004,N_11444,N_8864);
and U15005 (N_15005,N_10285,N_11135);
or U15006 (N_15006,N_10038,N_11817);
or U15007 (N_15007,N_8090,N_9460);
or U15008 (N_15008,N_11895,N_9739);
or U15009 (N_15009,N_9112,N_11705);
nand U15010 (N_15010,N_9319,N_11071);
and U15011 (N_15011,N_8890,N_8672);
and U15012 (N_15012,N_10880,N_11889);
or U15013 (N_15013,N_11781,N_11405);
nor U15014 (N_15014,N_8350,N_11679);
nor U15015 (N_15015,N_9927,N_8236);
nand U15016 (N_15016,N_9883,N_10672);
and U15017 (N_15017,N_10564,N_11298);
and U15018 (N_15018,N_10773,N_11885);
and U15019 (N_15019,N_11168,N_10467);
or U15020 (N_15020,N_11104,N_8940);
nor U15021 (N_15021,N_10971,N_11092);
nor U15022 (N_15022,N_10452,N_8477);
nor U15023 (N_15023,N_10882,N_11498);
nand U15024 (N_15024,N_8731,N_9076);
nand U15025 (N_15025,N_9590,N_10490);
nand U15026 (N_15026,N_8036,N_10942);
xnor U15027 (N_15027,N_8882,N_9510);
nand U15028 (N_15028,N_10559,N_11660);
nor U15029 (N_15029,N_10597,N_10384);
nor U15030 (N_15030,N_10465,N_11122);
and U15031 (N_15031,N_8621,N_10999);
nand U15032 (N_15032,N_11005,N_9678);
nand U15033 (N_15033,N_11186,N_8542);
or U15034 (N_15034,N_11456,N_10660);
and U15035 (N_15035,N_11113,N_8597);
nand U15036 (N_15036,N_8705,N_10586);
nand U15037 (N_15037,N_10320,N_11784);
nor U15038 (N_15038,N_9643,N_10616);
nor U15039 (N_15039,N_8558,N_8760);
and U15040 (N_15040,N_8417,N_8638);
nand U15041 (N_15041,N_8135,N_10495);
nand U15042 (N_15042,N_10859,N_10932);
and U15043 (N_15043,N_11963,N_9615);
or U15044 (N_15044,N_9922,N_11986);
nand U15045 (N_15045,N_9926,N_11350);
or U15046 (N_15046,N_10196,N_9894);
and U15047 (N_15047,N_10644,N_9754);
nand U15048 (N_15048,N_11170,N_11525);
nor U15049 (N_15049,N_8561,N_10568);
nor U15050 (N_15050,N_9643,N_11307);
or U15051 (N_15051,N_9162,N_10402);
or U15052 (N_15052,N_9693,N_8098);
nand U15053 (N_15053,N_11685,N_8994);
nand U15054 (N_15054,N_9251,N_8097);
xnor U15055 (N_15055,N_9149,N_8372);
nor U15056 (N_15056,N_11465,N_11221);
and U15057 (N_15057,N_8663,N_9223);
and U15058 (N_15058,N_11014,N_8005);
xor U15059 (N_15059,N_10327,N_11577);
xor U15060 (N_15060,N_8609,N_10112);
or U15061 (N_15061,N_8730,N_8804);
and U15062 (N_15062,N_11975,N_10956);
or U15063 (N_15063,N_11784,N_10772);
nand U15064 (N_15064,N_8942,N_9198);
nand U15065 (N_15065,N_9939,N_11403);
and U15066 (N_15066,N_11846,N_11653);
nand U15067 (N_15067,N_11355,N_10533);
nand U15068 (N_15068,N_10575,N_11039);
nand U15069 (N_15069,N_8291,N_9872);
xor U15070 (N_15070,N_10839,N_9965);
and U15071 (N_15071,N_10702,N_8856);
or U15072 (N_15072,N_8619,N_10393);
nor U15073 (N_15073,N_10070,N_10867);
and U15074 (N_15074,N_9522,N_11884);
or U15075 (N_15075,N_8929,N_9530);
nand U15076 (N_15076,N_11508,N_9858);
and U15077 (N_15077,N_10029,N_9656);
and U15078 (N_15078,N_11998,N_10901);
nand U15079 (N_15079,N_10510,N_10670);
nand U15080 (N_15080,N_8733,N_10428);
nand U15081 (N_15081,N_10525,N_11615);
nor U15082 (N_15082,N_11022,N_10374);
and U15083 (N_15083,N_8851,N_11841);
nor U15084 (N_15084,N_8236,N_11918);
nor U15085 (N_15085,N_8187,N_8808);
and U15086 (N_15086,N_11941,N_8784);
nand U15087 (N_15087,N_11884,N_9566);
or U15088 (N_15088,N_8904,N_10317);
nor U15089 (N_15089,N_10089,N_9968);
and U15090 (N_15090,N_8670,N_10417);
and U15091 (N_15091,N_8107,N_10546);
or U15092 (N_15092,N_11188,N_11299);
or U15093 (N_15093,N_9550,N_10976);
nand U15094 (N_15094,N_10088,N_11163);
nand U15095 (N_15095,N_9734,N_10160);
or U15096 (N_15096,N_9169,N_9553);
and U15097 (N_15097,N_10433,N_11158);
nand U15098 (N_15098,N_8522,N_10460);
and U15099 (N_15099,N_9881,N_8533);
or U15100 (N_15100,N_9955,N_8925);
and U15101 (N_15101,N_10905,N_10369);
xnor U15102 (N_15102,N_10425,N_11441);
or U15103 (N_15103,N_10329,N_11651);
nand U15104 (N_15104,N_8290,N_10043);
and U15105 (N_15105,N_9962,N_8250);
nor U15106 (N_15106,N_11946,N_11239);
and U15107 (N_15107,N_11598,N_8045);
or U15108 (N_15108,N_8412,N_10283);
nand U15109 (N_15109,N_9283,N_10218);
nor U15110 (N_15110,N_11513,N_9123);
nand U15111 (N_15111,N_9206,N_11678);
nor U15112 (N_15112,N_11720,N_11221);
nor U15113 (N_15113,N_11001,N_11674);
nand U15114 (N_15114,N_9344,N_10882);
nand U15115 (N_15115,N_8255,N_8265);
nand U15116 (N_15116,N_11392,N_10745);
or U15117 (N_15117,N_11818,N_11812);
or U15118 (N_15118,N_9245,N_8444);
nor U15119 (N_15119,N_9686,N_9380);
nand U15120 (N_15120,N_8783,N_10460);
and U15121 (N_15121,N_9100,N_8921);
and U15122 (N_15122,N_9526,N_10372);
nand U15123 (N_15123,N_11595,N_10146);
or U15124 (N_15124,N_8741,N_9984);
or U15125 (N_15125,N_8607,N_9436);
nand U15126 (N_15126,N_10144,N_9679);
xor U15127 (N_15127,N_10328,N_8929);
nand U15128 (N_15128,N_9698,N_11986);
or U15129 (N_15129,N_10630,N_11921);
nor U15130 (N_15130,N_8473,N_8270);
xnor U15131 (N_15131,N_11069,N_10538);
nor U15132 (N_15132,N_9172,N_9743);
nor U15133 (N_15133,N_11840,N_8549);
and U15134 (N_15134,N_9001,N_8948);
nand U15135 (N_15135,N_10406,N_9239);
or U15136 (N_15136,N_10301,N_9012);
and U15137 (N_15137,N_10746,N_10343);
or U15138 (N_15138,N_8482,N_11475);
and U15139 (N_15139,N_10801,N_10508);
or U15140 (N_15140,N_8804,N_11420);
nor U15141 (N_15141,N_9843,N_11013);
nand U15142 (N_15142,N_9832,N_10860);
and U15143 (N_15143,N_9602,N_9808);
and U15144 (N_15144,N_10340,N_10221);
nand U15145 (N_15145,N_9882,N_8963);
nand U15146 (N_15146,N_10534,N_11484);
or U15147 (N_15147,N_8270,N_9149);
nand U15148 (N_15148,N_9743,N_9409);
nor U15149 (N_15149,N_8575,N_9204);
or U15150 (N_15150,N_10628,N_11605);
xor U15151 (N_15151,N_8550,N_9331);
nand U15152 (N_15152,N_8668,N_10267);
nand U15153 (N_15153,N_10601,N_10161);
nor U15154 (N_15154,N_10509,N_9966);
nor U15155 (N_15155,N_8330,N_8900);
nor U15156 (N_15156,N_11441,N_11667);
nor U15157 (N_15157,N_8124,N_8692);
nand U15158 (N_15158,N_8607,N_9042);
xnor U15159 (N_15159,N_8375,N_9642);
or U15160 (N_15160,N_10749,N_10045);
and U15161 (N_15161,N_8256,N_11986);
and U15162 (N_15162,N_11417,N_10979);
or U15163 (N_15163,N_9904,N_10482);
nor U15164 (N_15164,N_9195,N_10990);
and U15165 (N_15165,N_11137,N_9693);
and U15166 (N_15166,N_9501,N_8097);
nor U15167 (N_15167,N_10543,N_9859);
or U15168 (N_15168,N_9298,N_10705);
nor U15169 (N_15169,N_10476,N_11819);
xor U15170 (N_15170,N_9865,N_8011);
xor U15171 (N_15171,N_9600,N_8276);
or U15172 (N_15172,N_10733,N_9375);
nand U15173 (N_15173,N_9283,N_8829);
and U15174 (N_15174,N_10618,N_10885);
or U15175 (N_15175,N_8752,N_11898);
or U15176 (N_15176,N_10852,N_10014);
nor U15177 (N_15177,N_9109,N_11062);
nor U15178 (N_15178,N_8055,N_9869);
nor U15179 (N_15179,N_9540,N_8797);
nand U15180 (N_15180,N_9216,N_11079);
nor U15181 (N_15181,N_8923,N_10533);
nor U15182 (N_15182,N_8125,N_9930);
nor U15183 (N_15183,N_10992,N_8043);
nand U15184 (N_15184,N_11152,N_11025);
nor U15185 (N_15185,N_9786,N_9451);
nor U15186 (N_15186,N_8416,N_9927);
nand U15187 (N_15187,N_11832,N_8493);
nand U15188 (N_15188,N_11987,N_10316);
or U15189 (N_15189,N_11890,N_8082);
and U15190 (N_15190,N_8749,N_9868);
nor U15191 (N_15191,N_10277,N_11093);
or U15192 (N_15192,N_10042,N_8471);
nand U15193 (N_15193,N_8871,N_10459);
or U15194 (N_15194,N_10143,N_10325);
or U15195 (N_15195,N_8367,N_8375);
xor U15196 (N_15196,N_10516,N_11528);
and U15197 (N_15197,N_11833,N_9518);
or U15198 (N_15198,N_8991,N_10057);
nor U15199 (N_15199,N_8893,N_10072);
xnor U15200 (N_15200,N_11691,N_8586);
nor U15201 (N_15201,N_11230,N_9177);
nor U15202 (N_15202,N_9536,N_11268);
or U15203 (N_15203,N_10903,N_8602);
nor U15204 (N_15204,N_10732,N_11107);
xor U15205 (N_15205,N_9540,N_9639);
or U15206 (N_15206,N_9459,N_9841);
nand U15207 (N_15207,N_8904,N_11194);
nor U15208 (N_15208,N_9986,N_8177);
nand U15209 (N_15209,N_8081,N_8012);
nand U15210 (N_15210,N_10347,N_8676);
and U15211 (N_15211,N_9087,N_8640);
or U15212 (N_15212,N_10133,N_10989);
and U15213 (N_15213,N_10318,N_9616);
or U15214 (N_15214,N_10008,N_8209);
nor U15215 (N_15215,N_10317,N_11351);
nand U15216 (N_15216,N_10384,N_11456);
or U15217 (N_15217,N_10860,N_11372);
nand U15218 (N_15218,N_10703,N_10382);
nor U15219 (N_15219,N_10323,N_9675);
nor U15220 (N_15220,N_10846,N_11927);
nand U15221 (N_15221,N_9492,N_11169);
and U15222 (N_15222,N_8888,N_8727);
xnor U15223 (N_15223,N_10467,N_9736);
nand U15224 (N_15224,N_10060,N_8387);
nand U15225 (N_15225,N_11119,N_8096);
and U15226 (N_15226,N_9014,N_9057);
nand U15227 (N_15227,N_11899,N_10429);
xor U15228 (N_15228,N_11948,N_11830);
nor U15229 (N_15229,N_9075,N_8370);
xor U15230 (N_15230,N_11232,N_10805);
and U15231 (N_15231,N_8380,N_10355);
nor U15232 (N_15232,N_9586,N_11719);
xnor U15233 (N_15233,N_9987,N_9761);
and U15234 (N_15234,N_9260,N_9508);
and U15235 (N_15235,N_10893,N_10769);
nand U15236 (N_15236,N_11762,N_9328);
nor U15237 (N_15237,N_9303,N_10524);
and U15238 (N_15238,N_9244,N_11279);
or U15239 (N_15239,N_8854,N_8469);
xnor U15240 (N_15240,N_8223,N_9268);
nand U15241 (N_15241,N_8242,N_10545);
nor U15242 (N_15242,N_11628,N_11650);
or U15243 (N_15243,N_8068,N_9616);
nor U15244 (N_15244,N_9739,N_9291);
and U15245 (N_15245,N_11169,N_11229);
nor U15246 (N_15246,N_10098,N_8906);
and U15247 (N_15247,N_10472,N_9217);
nand U15248 (N_15248,N_9804,N_11740);
nor U15249 (N_15249,N_10544,N_8518);
or U15250 (N_15250,N_9934,N_11423);
and U15251 (N_15251,N_8542,N_9486);
xor U15252 (N_15252,N_11526,N_11755);
and U15253 (N_15253,N_10876,N_11499);
or U15254 (N_15254,N_9376,N_9049);
nand U15255 (N_15255,N_11381,N_10741);
nor U15256 (N_15256,N_11803,N_10427);
nor U15257 (N_15257,N_8864,N_11558);
nand U15258 (N_15258,N_11643,N_8113);
or U15259 (N_15259,N_8004,N_8208);
nor U15260 (N_15260,N_8420,N_9059);
nor U15261 (N_15261,N_8292,N_11645);
and U15262 (N_15262,N_9564,N_9377);
xor U15263 (N_15263,N_9563,N_10338);
nand U15264 (N_15264,N_9124,N_10816);
and U15265 (N_15265,N_10049,N_10019);
or U15266 (N_15266,N_8140,N_8228);
nand U15267 (N_15267,N_10273,N_11476);
nand U15268 (N_15268,N_11886,N_8857);
nor U15269 (N_15269,N_9481,N_11415);
or U15270 (N_15270,N_10187,N_10375);
or U15271 (N_15271,N_8673,N_11858);
or U15272 (N_15272,N_8983,N_9389);
and U15273 (N_15273,N_11231,N_8397);
and U15274 (N_15274,N_9224,N_10387);
nor U15275 (N_15275,N_8812,N_8745);
and U15276 (N_15276,N_11515,N_9980);
nand U15277 (N_15277,N_10299,N_10996);
nand U15278 (N_15278,N_8530,N_8868);
nand U15279 (N_15279,N_10013,N_10321);
nor U15280 (N_15280,N_9240,N_8332);
or U15281 (N_15281,N_8607,N_8037);
or U15282 (N_15282,N_11857,N_10499);
or U15283 (N_15283,N_9547,N_9905);
and U15284 (N_15284,N_10088,N_8475);
nand U15285 (N_15285,N_11457,N_9980);
and U15286 (N_15286,N_9906,N_10263);
or U15287 (N_15287,N_9493,N_9451);
nand U15288 (N_15288,N_8097,N_11570);
or U15289 (N_15289,N_11522,N_8992);
nor U15290 (N_15290,N_9507,N_9623);
and U15291 (N_15291,N_11787,N_10465);
nand U15292 (N_15292,N_9563,N_9356);
or U15293 (N_15293,N_8068,N_8589);
nor U15294 (N_15294,N_10508,N_10483);
nor U15295 (N_15295,N_8951,N_10074);
nand U15296 (N_15296,N_9338,N_11146);
nor U15297 (N_15297,N_9740,N_11443);
or U15298 (N_15298,N_9836,N_11132);
nor U15299 (N_15299,N_9484,N_11291);
nand U15300 (N_15300,N_9396,N_11102);
xnor U15301 (N_15301,N_8139,N_11957);
nand U15302 (N_15302,N_11333,N_10273);
and U15303 (N_15303,N_9727,N_11385);
nor U15304 (N_15304,N_10541,N_8737);
and U15305 (N_15305,N_8985,N_9646);
nor U15306 (N_15306,N_11545,N_11469);
and U15307 (N_15307,N_10309,N_9460);
nor U15308 (N_15308,N_11014,N_11425);
and U15309 (N_15309,N_8885,N_10801);
and U15310 (N_15310,N_8535,N_10037);
and U15311 (N_15311,N_11800,N_9128);
nand U15312 (N_15312,N_10676,N_11309);
and U15313 (N_15313,N_9561,N_8138);
or U15314 (N_15314,N_11323,N_10271);
and U15315 (N_15315,N_8744,N_8627);
nor U15316 (N_15316,N_10952,N_8854);
and U15317 (N_15317,N_9635,N_9064);
or U15318 (N_15318,N_9482,N_9129);
or U15319 (N_15319,N_11402,N_10371);
nor U15320 (N_15320,N_9995,N_11124);
nand U15321 (N_15321,N_10175,N_8189);
or U15322 (N_15322,N_10710,N_10551);
nor U15323 (N_15323,N_8133,N_10186);
xor U15324 (N_15324,N_10379,N_11051);
or U15325 (N_15325,N_11541,N_11317);
nand U15326 (N_15326,N_10838,N_8118);
and U15327 (N_15327,N_10656,N_8841);
nand U15328 (N_15328,N_11686,N_10624);
xor U15329 (N_15329,N_10684,N_9725);
and U15330 (N_15330,N_8292,N_9902);
xor U15331 (N_15331,N_10083,N_10170);
and U15332 (N_15332,N_11341,N_8593);
or U15333 (N_15333,N_8069,N_11779);
and U15334 (N_15334,N_8596,N_8184);
or U15335 (N_15335,N_10497,N_11835);
and U15336 (N_15336,N_9350,N_8123);
nor U15337 (N_15337,N_8484,N_8674);
and U15338 (N_15338,N_9754,N_8193);
or U15339 (N_15339,N_11410,N_10954);
nand U15340 (N_15340,N_9202,N_10672);
or U15341 (N_15341,N_8318,N_10596);
nor U15342 (N_15342,N_10708,N_8361);
or U15343 (N_15343,N_11527,N_8554);
or U15344 (N_15344,N_11755,N_11926);
and U15345 (N_15345,N_8435,N_9144);
nor U15346 (N_15346,N_8269,N_11770);
and U15347 (N_15347,N_9880,N_11550);
and U15348 (N_15348,N_11187,N_10404);
or U15349 (N_15349,N_9644,N_10778);
or U15350 (N_15350,N_10731,N_8835);
or U15351 (N_15351,N_8818,N_8261);
and U15352 (N_15352,N_10634,N_10504);
nor U15353 (N_15353,N_8908,N_8932);
nor U15354 (N_15354,N_9387,N_8601);
xnor U15355 (N_15355,N_8988,N_11509);
xor U15356 (N_15356,N_9656,N_9930);
or U15357 (N_15357,N_10148,N_10777);
nand U15358 (N_15358,N_10768,N_11593);
and U15359 (N_15359,N_10564,N_11905);
nand U15360 (N_15360,N_10646,N_10529);
nor U15361 (N_15361,N_11003,N_10340);
or U15362 (N_15362,N_11518,N_11044);
and U15363 (N_15363,N_8187,N_11710);
xnor U15364 (N_15364,N_11564,N_8452);
xor U15365 (N_15365,N_8439,N_8215);
or U15366 (N_15366,N_9182,N_8500);
nor U15367 (N_15367,N_11989,N_11892);
or U15368 (N_15368,N_11119,N_8078);
nand U15369 (N_15369,N_10534,N_11155);
nor U15370 (N_15370,N_8445,N_11071);
and U15371 (N_15371,N_8026,N_11803);
xnor U15372 (N_15372,N_9237,N_9953);
nor U15373 (N_15373,N_9624,N_9282);
nor U15374 (N_15374,N_8785,N_8940);
or U15375 (N_15375,N_11339,N_8842);
or U15376 (N_15376,N_9017,N_8232);
and U15377 (N_15377,N_8233,N_9143);
and U15378 (N_15378,N_9468,N_8890);
nand U15379 (N_15379,N_10532,N_8236);
xor U15380 (N_15380,N_11662,N_9749);
or U15381 (N_15381,N_11992,N_8131);
and U15382 (N_15382,N_10625,N_11596);
and U15383 (N_15383,N_8930,N_9495);
and U15384 (N_15384,N_11599,N_8639);
xor U15385 (N_15385,N_11476,N_8270);
or U15386 (N_15386,N_11675,N_8403);
nor U15387 (N_15387,N_9663,N_8392);
or U15388 (N_15388,N_9471,N_11625);
xor U15389 (N_15389,N_9436,N_11367);
or U15390 (N_15390,N_11737,N_10784);
nand U15391 (N_15391,N_8525,N_10229);
nand U15392 (N_15392,N_8329,N_11704);
nand U15393 (N_15393,N_9061,N_11726);
and U15394 (N_15394,N_8510,N_10720);
and U15395 (N_15395,N_11756,N_10165);
and U15396 (N_15396,N_8552,N_9887);
or U15397 (N_15397,N_9046,N_11742);
nor U15398 (N_15398,N_9006,N_10919);
nand U15399 (N_15399,N_8638,N_8029);
nor U15400 (N_15400,N_8980,N_11285);
or U15401 (N_15401,N_9574,N_8964);
or U15402 (N_15402,N_8766,N_10711);
and U15403 (N_15403,N_11301,N_10414);
nor U15404 (N_15404,N_11399,N_10817);
and U15405 (N_15405,N_11865,N_10187);
and U15406 (N_15406,N_9917,N_10246);
or U15407 (N_15407,N_9538,N_8183);
or U15408 (N_15408,N_8111,N_11089);
xnor U15409 (N_15409,N_9951,N_8798);
nand U15410 (N_15410,N_8348,N_9655);
nand U15411 (N_15411,N_10080,N_10150);
nand U15412 (N_15412,N_8288,N_11233);
and U15413 (N_15413,N_10432,N_8048);
and U15414 (N_15414,N_8640,N_9475);
nand U15415 (N_15415,N_8198,N_10064);
nand U15416 (N_15416,N_10600,N_9271);
nor U15417 (N_15417,N_9230,N_11503);
nor U15418 (N_15418,N_8448,N_10542);
nand U15419 (N_15419,N_11503,N_10298);
nor U15420 (N_15420,N_11598,N_9619);
and U15421 (N_15421,N_10626,N_8395);
xnor U15422 (N_15422,N_8153,N_8139);
and U15423 (N_15423,N_10797,N_9847);
nor U15424 (N_15424,N_11832,N_10230);
or U15425 (N_15425,N_11650,N_8635);
and U15426 (N_15426,N_9894,N_8439);
nand U15427 (N_15427,N_10397,N_11774);
nand U15428 (N_15428,N_10598,N_8177);
and U15429 (N_15429,N_8413,N_11540);
nand U15430 (N_15430,N_9978,N_10520);
nand U15431 (N_15431,N_8121,N_9510);
nor U15432 (N_15432,N_11180,N_8723);
nor U15433 (N_15433,N_11345,N_9350);
and U15434 (N_15434,N_8961,N_9846);
or U15435 (N_15435,N_9722,N_8563);
nor U15436 (N_15436,N_9778,N_10508);
xnor U15437 (N_15437,N_11683,N_11731);
xnor U15438 (N_15438,N_10338,N_8332);
or U15439 (N_15439,N_8363,N_11700);
nand U15440 (N_15440,N_11673,N_11488);
nand U15441 (N_15441,N_9949,N_11671);
nand U15442 (N_15442,N_11457,N_10113);
xor U15443 (N_15443,N_11053,N_11377);
nor U15444 (N_15444,N_9795,N_9142);
nand U15445 (N_15445,N_11997,N_8484);
nor U15446 (N_15446,N_10735,N_8867);
or U15447 (N_15447,N_10936,N_11899);
and U15448 (N_15448,N_8363,N_8120);
or U15449 (N_15449,N_8386,N_10706);
and U15450 (N_15450,N_10516,N_11606);
nor U15451 (N_15451,N_9473,N_9608);
and U15452 (N_15452,N_11761,N_8762);
nor U15453 (N_15453,N_11643,N_11984);
nand U15454 (N_15454,N_11846,N_11013);
nand U15455 (N_15455,N_9403,N_11836);
xor U15456 (N_15456,N_10694,N_11765);
nor U15457 (N_15457,N_8705,N_9716);
and U15458 (N_15458,N_8175,N_10068);
xnor U15459 (N_15459,N_9807,N_9679);
nand U15460 (N_15460,N_9697,N_11028);
and U15461 (N_15461,N_10069,N_8077);
nand U15462 (N_15462,N_10444,N_9434);
nand U15463 (N_15463,N_10769,N_9192);
nand U15464 (N_15464,N_10816,N_8366);
nand U15465 (N_15465,N_9350,N_11414);
nand U15466 (N_15466,N_8930,N_10959);
or U15467 (N_15467,N_10571,N_8676);
xor U15468 (N_15468,N_8957,N_11004);
and U15469 (N_15469,N_11995,N_9464);
or U15470 (N_15470,N_9733,N_11084);
or U15471 (N_15471,N_8540,N_11185);
xor U15472 (N_15472,N_8658,N_11388);
xnor U15473 (N_15473,N_9604,N_11743);
or U15474 (N_15474,N_8018,N_11706);
nor U15475 (N_15475,N_8098,N_9011);
nor U15476 (N_15476,N_11808,N_11525);
or U15477 (N_15477,N_10139,N_9703);
xor U15478 (N_15478,N_8619,N_9488);
nor U15479 (N_15479,N_8061,N_9071);
nor U15480 (N_15480,N_10587,N_8999);
nand U15481 (N_15481,N_9143,N_8269);
and U15482 (N_15482,N_9928,N_11612);
nand U15483 (N_15483,N_8989,N_11248);
nor U15484 (N_15484,N_8845,N_10735);
and U15485 (N_15485,N_9453,N_9549);
nand U15486 (N_15486,N_11693,N_10667);
nand U15487 (N_15487,N_11930,N_8475);
or U15488 (N_15488,N_11556,N_10791);
or U15489 (N_15489,N_9118,N_8267);
and U15490 (N_15490,N_9890,N_8994);
nor U15491 (N_15491,N_11357,N_9905);
xnor U15492 (N_15492,N_10324,N_9243);
xnor U15493 (N_15493,N_9289,N_9401);
xor U15494 (N_15494,N_10107,N_10294);
or U15495 (N_15495,N_9070,N_11263);
nand U15496 (N_15496,N_10059,N_8653);
or U15497 (N_15497,N_10176,N_9357);
nand U15498 (N_15498,N_8211,N_9713);
and U15499 (N_15499,N_9528,N_9614);
nand U15500 (N_15500,N_9506,N_10162);
and U15501 (N_15501,N_9674,N_10355);
nand U15502 (N_15502,N_8206,N_11374);
or U15503 (N_15503,N_10669,N_11147);
and U15504 (N_15504,N_10738,N_8319);
nor U15505 (N_15505,N_8634,N_10385);
or U15506 (N_15506,N_11951,N_9538);
nor U15507 (N_15507,N_10709,N_8353);
and U15508 (N_15508,N_8601,N_8243);
and U15509 (N_15509,N_8156,N_8041);
or U15510 (N_15510,N_11783,N_11151);
and U15511 (N_15511,N_10296,N_10487);
nor U15512 (N_15512,N_10524,N_9636);
nor U15513 (N_15513,N_8126,N_9780);
nor U15514 (N_15514,N_8293,N_11217);
or U15515 (N_15515,N_10142,N_11961);
nand U15516 (N_15516,N_10329,N_10817);
and U15517 (N_15517,N_11458,N_9191);
and U15518 (N_15518,N_11113,N_11186);
nor U15519 (N_15519,N_10601,N_10764);
nand U15520 (N_15520,N_9209,N_8350);
and U15521 (N_15521,N_11493,N_10444);
xnor U15522 (N_15522,N_8214,N_11353);
or U15523 (N_15523,N_10417,N_9462);
nand U15524 (N_15524,N_11424,N_11621);
or U15525 (N_15525,N_9570,N_9859);
nand U15526 (N_15526,N_9241,N_9435);
and U15527 (N_15527,N_10360,N_9283);
nor U15528 (N_15528,N_11128,N_10140);
nand U15529 (N_15529,N_8567,N_10898);
nor U15530 (N_15530,N_9173,N_9959);
and U15531 (N_15531,N_9632,N_10676);
nor U15532 (N_15532,N_10002,N_9637);
nand U15533 (N_15533,N_10815,N_9668);
and U15534 (N_15534,N_8010,N_9783);
nand U15535 (N_15535,N_9149,N_8652);
xor U15536 (N_15536,N_8203,N_8920);
nand U15537 (N_15537,N_11009,N_11547);
or U15538 (N_15538,N_10843,N_11319);
and U15539 (N_15539,N_9049,N_10627);
and U15540 (N_15540,N_9409,N_11652);
and U15541 (N_15541,N_9088,N_8893);
and U15542 (N_15542,N_10106,N_9208);
nor U15543 (N_15543,N_11720,N_9955);
nor U15544 (N_15544,N_8930,N_9804);
nor U15545 (N_15545,N_9224,N_8792);
nor U15546 (N_15546,N_10896,N_9356);
nand U15547 (N_15547,N_10039,N_11582);
nor U15548 (N_15548,N_8371,N_10738);
nor U15549 (N_15549,N_10070,N_10569);
xnor U15550 (N_15550,N_10355,N_10875);
and U15551 (N_15551,N_10860,N_11977);
or U15552 (N_15552,N_8319,N_8167);
and U15553 (N_15553,N_8639,N_8018);
nor U15554 (N_15554,N_8881,N_8752);
and U15555 (N_15555,N_8890,N_11008);
nor U15556 (N_15556,N_11395,N_11101);
and U15557 (N_15557,N_9637,N_10302);
and U15558 (N_15558,N_9245,N_8106);
and U15559 (N_15559,N_8833,N_9017);
or U15560 (N_15560,N_11158,N_8308);
nand U15561 (N_15561,N_9893,N_9534);
nand U15562 (N_15562,N_8237,N_10692);
and U15563 (N_15563,N_9275,N_11941);
or U15564 (N_15564,N_11988,N_9059);
nor U15565 (N_15565,N_10899,N_11819);
nand U15566 (N_15566,N_8073,N_10524);
or U15567 (N_15567,N_9793,N_11242);
nor U15568 (N_15568,N_10505,N_11795);
nor U15569 (N_15569,N_11183,N_11195);
or U15570 (N_15570,N_10234,N_11402);
or U15571 (N_15571,N_11435,N_11776);
nand U15572 (N_15572,N_11590,N_11192);
and U15573 (N_15573,N_11073,N_9144);
nand U15574 (N_15574,N_11728,N_10785);
xor U15575 (N_15575,N_9952,N_10403);
and U15576 (N_15576,N_9822,N_8408);
nand U15577 (N_15577,N_10911,N_11181);
nand U15578 (N_15578,N_9972,N_8695);
or U15579 (N_15579,N_9111,N_8671);
nor U15580 (N_15580,N_11642,N_9716);
nor U15581 (N_15581,N_9300,N_11988);
nor U15582 (N_15582,N_10904,N_11246);
nand U15583 (N_15583,N_8561,N_8753);
nand U15584 (N_15584,N_10535,N_10459);
or U15585 (N_15585,N_10900,N_11692);
nor U15586 (N_15586,N_9639,N_8306);
nand U15587 (N_15587,N_9766,N_9276);
nand U15588 (N_15588,N_10476,N_8791);
or U15589 (N_15589,N_8618,N_8757);
and U15590 (N_15590,N_10794,N_8214);
nand U15591 (N_15591,N_8499,N_11281);
or U15592 (N_15592,N_9885,N_9335);
nand U15593 (N_15593,N_9624,N_10745);
and U15594 (N_15594,N_9902,N_11819);
nor U15595 (N_15595,N_9683,N_9700);
xnor U15596 (N_15596,N_9755,N_8592);
nor U15597 (N_15597,N_8576,N_8235);
xnor U15598 (N_15598,N_9746,N_10743);
and U15599 (N_15599,N_8751,N_10142);
and U15600 (N_15600,N_11011,N_8242);
or U15601 (N_15601,N_11299,N_9207);
and U15602 (N_15602,N_8003,N_8206);
nand U15603 (N_15603,N_8181,N_9114);
nor U15604 (N_15604,N_8267,N_9315);
and U15605 (N_15605,N_11166,N_10448);
nor U15606 (N_15606,N_9730,N_8850);
or U15607 (N_15607,N_11176,N_11381);
or U15608 (N_15608,N_11822,N_11877);
xnor U15609 (N_15609,N_8861,N_9948);
nor U15610 (N_15610,N_8000,N_10398);
or U15611 (N_15611,N_11952,N_11559);
nand U15612 (N_15612,N_10172,N_9560);
nand U15613 (N_15613,N_11151,N_11519);
xor U15614 (N_15614,N_9355,N_8296);
nor U15615 (N_15615,N_8421,N_10476);
xnor U15616 (N_15616,N_10345,N_8100);
or U15617 (N_15617,N_10661,N_9578);
nor U15618 (N_15618,N_10560,N_8084);
nor U15619 (N_15619,N_11511,N_8167);
nor U15620 (N_15620,N_8939,N_10266);
nor U15621 (N_15621,N_8783,N_8046);
or U15622 (N_15622,N_10967,N_10381);
nor U15623 (N_15623,N_10975,N_10707);
nand U15624 (N_15624,N_9594,N_11063);
and U15625 (N_15625,N_10325,N_10952);
and U15626 (N_15626,N_11559,N_10089);
nor U15627 (N_15627,N_8831,N_11147);
or U15628 (N_15628,N_8208,N_10037);
or U15629 (N_15629,N_11302,N_9239);
nor U15630 (N_15630,N_9772,N_11400);
nand U15631 (N_15631,N_10828,N_11124);
or U15632 (N_15632,N_10459,N_8955);
nand U15633 (N_15633,N_11798,N_8696);
and U15634 (N_15634,N_8266,N_8068);
or U15635 (N_15635,N_11646,N_11807);
and U15636 (N_15636,N_9079,N_11050);
nand U15637 (N_15637,N_8779,N_10619);
or U15638 (N_15638,N_10076,N_8229);
nor U15639 (N_15639,N_10308,N_9117);
and U15640 (N_15640,N_9445,N_8352);
and U15641 (N_15641,N_8085,N_9721);
xor U15642 (N_15642,N_8838,N_11412);
nor U15643 (N_15643,N_11519,N_8172);
and U15644 (N_15644,N_10260,N_11074);
nor U15645 (N_15645,N_10466,N_10924);
or U15646 (N_15646,N_9774,N_8259);
nor U15647 (N_15647,N_8250,N_11448);
nand U15648 (N_15648,N_8948,N_9010);
nand U15649 (N_15649,N_8978,N_8179);
and U15650 (N_15650,N_9089,N_10467);
xnor U15651 (N_15651,N_9298,N_10555);
nand U15652 (N_15652,N_11711,N_11748);
or U15653 (N_15653,N_11958,N_10519);
nor U15654 (N_15654,N_11429,N_10915);
and U15655 (N_15655,N_8001,N_8153);
nor U15656 (N_15656,N_8639,N_8788);
nor U15657 (N_15657,N_8189,N_10375);
xor U15658 (N_15658,N_10336,N_11807);
nand U15659 (N_15659,N_9161,N_11961);
or U15660 (N_15660,N_9110,N_9383);
nor U15661 (N_15661,N_10034,N_8011);
nand U15662 (N_15662,N_11910,N_8341);
nor U15663 (N_15663,N_8500,N_10311);
nand U15664 (N_15664,N_11220,N_8670);
and U15665 (N_15665,N_9355,N_10345);
nand U15666 (N_15666,N_9591,N_9177);
nand U15667 (N_15667,N_10053,N_9870);
xnor U15668 (N_15668,N_9008,N_8168);
nor U15669 (N_15669,N_8608,N_10004);
nor U15670 (N_15670,N_10949,N_11182);
and U15671 (N_15671,N_11496,N_11584);
or U15672 (N_15672,N_11442,N_10281);
or U15673 (N_15673,N_10555,N_11667);
and U15674 (N_15674,N_8108,N_10510);
xnor U15675 (N_15675,N_11356,N_11033);
or U15676 (N_15676,N_10291,N_10803);
nand U15677 (N_15677,N_10098,N_11757);
or U15678 (N_15678,N_11331,N_8148);
nor U15679 (N_15679,N_9725,N_11230);
or U15680 (N_15680,N_10778,N_11833);
nor U15681 (N_15681,N_8051,N_11492);
or U15682 (N_15682,N_10480,N_11428);
or U15683 (N_15683,N_8987,N_9922);
or U15684 (N_15684,N_9229,N_10961);
and U15685 (N_15685,N_11417,N_11095);
and U15686 (N_15686,N_8885,N_9795);
nor U15687 (N_15687,N_9146,N_9287);
nand U15688 (N_15688,N_8147,N_10850);
nand U15689 (N_15689,N_11747,N_11017);
or U15690 (N_15690,N_9842,N_8359);
or U15691 (N_15691,N_10772,N_10925);
or U15692 (N_15692,N_11630,N_10037);
and U15693 (N_15693,N_11435,N_8327);
and U15694 (N_15694,N_10621,N_10430);
nand U15695 (N_15695,N_8115,N_10686);
xor U15696 (N_15696,N_10325,N_9402);
xor U15697 (N_15697,N_10437,N_11422);
or U15698 (N_15698,N_11486,N_9967);
and U15699 (N_15699,N_11344,N_10529);
nand U15700 (N_15700,N_8266,N_8674);
nor U15701 (N_15701,N_9767,N_10222);
or U15702 (N_15702,N_8190,N_10637);
or U15703 (N_15703,N_9538,N_10181);
xor U15704 (N_15704,N_10812,N_11965);
and U15705 (N_15705,N_10849,N_8111);
and U15706 (N_15706,N_11086,N_8785);
and U15707 (N_15707,N_9203,N_11211);
and U15708 (N_15708,N_9652,N_10952);
or U15709 (N_15709,N_8512,N_10408);
and U15710 (N_15710,N_10209,N_8837);
or U15711 (N_15711,N_10276,N_10468);
nand U15712 (N_15712,N_8060,N_8767);
nand U15713 (N_15713,N_10066,N_11551);
nor U15714 (N_15714,N_9307,N_9039);
nor U15715 (N_15715,N_11093,N_8624);
and U15716 (N_15716,N_8463,N_8783);
or U15717 (N_15717,N_11385,N_11859);
nor U15718 (N_15718,N_10706,N_11889);
or U15719 (N_15719,N_8298,N_8197);
and U15720 (N_15720,N_10291,N_11742);
nor U15721 (N_15721,N_8033,N_11072);
nor U15722 (N_15722,N_8762,N_8469);
xnor U15723 (N_15723,N_9262,N_11437);
xnor U15724 (N_15724,N_10161,N_9251);
nor U15725 (N_15725,N_10969,N_11979);
or U15726 (N_15726,N_11940,N_11491);
and U15727 (N_15727,N_10253,N_10143);
or U15728 (N_15728,N_11102,N_8206);
nand U15729 (N_15729,N_11502,N_11348);
or U15730 (N_15730,N_11504,N_8895);
nor U15731 (N_15731,N_10179,N_9259);
nor U15732 (N_15732,N_9845,N_11392);
or U15733 (N_15733,N_10567,N_9633);
nand U15734 (N_15734,N_9049,N_11699);
and U15735 (N_15735,N_8645,N_10800);
or U15736 (N_15736,N_10393,N_8389);
nor U15737 (N_15737,N_8423,N_9587);
and U15738 (N_15738,N_9324,N_8900);
xnor U15739 (N_15739,N_10198,N_9711);
or U15740 (N_15740,N_10973,N_8737);
or U15741 (N_15741,N_10433,N_10952);
or U15742 (N_15742,N_10854,N_10579);
nand U15743 (N_15743,N_8576,N_9242);
or U15744 (N_15744,N_10048,N_10663);
nand U15745 (N_15745,N_8377,N_10343);
and U15746 (N_15746,N_8062,N_10431);
nand U15747 (N_15747,N_10573,N_10718);
or U15748 (N_15748,N_9213,N_9453);
nand U15749 (N_15749,N_9079,N_10910);
nand U15750 (N_15750,N_10424,N_8473);
xor U15751 (N_15751,N_11749,N_11933);
and U15752 (N_15752,N_10892,N_10946);
or U15753 (N_15753,N_10737,N_9888);
or U15754 (N_15754,N_11385,N_11067);
nand U15755 (N_15755,N_9943,N_10056);
nor U15756 (N_15756,N_9732,N_11646);
nand U15757 (N_15757,N_11327,N_11359);
or U15758 (N_15758,N_11086,N_9850);
nand U15759 (N_15759,N_10357,N_11461);
nand U15760 (N_15760,N_9919,N_8219);
and U15761 (N_15761,N_9264,N_9318);
and U15762 (N_15762,N_11061,N_8618);
nor U15763 (N_15763,N_8222,N_11617);
and U15764 (N_15764,N_10365,N_8237);
nor U15765 (N_15765,N_8618,N_9447);
nor U15766 (N_15766,N_8059,N_10623);
nor U15767 (N_15767,N_11108,N_8451);
nor U15768 (N_15768,N_10263,N_11729);
nor U15769 (N_15769,N_11867,N_8343);
and U15770 (N_15770,N_10998,N_11432);
nor U15771 (N_15771,N_8241,N_10035);
or U15772 (N_15772,N_9260,N_8144);
nand U15773 (N_15773,N_8833,N_9174);
or U15774 (N_15774,N_10100,N_11996);
or U15775 (N_15775,N_10607,N_9722);
or U15776 (N_15776,N_11422,N_11242);
or U15777 (N_15777,N_11758,N_9695);
nand U15778 (N_15778,N_8915,N_11366);
nor U15779 (N_15779,N_8110,N_11813);
or U15780 (N_15780,N_9839,N_9493);
nand U15781 (N_15781,N_11877,N_11622);
nor U15782 (N_15782,N_9359,N_10192);
nor U15783 (N_15783,N_8275,N_9196);
or U15784 (N_15784,N_10960,N_8254);
xor U15785 (N_15785,N_9298,N_11784);
nor U15786 (N_15786,N_9903,N_11477);
xor U15787 (N_15787,N_9125,N_10634);
or U15788 (N_15788,N_10956,N_9016);
nand U15789 (N_15789,N_10001,N_8961);
and U15790 (N_15790,N_8811,N_10579);
xor U15791 (N_15791,N_10496,N_10744);
or U15792 (N_15792,N_9904,N_9809);
and U15793 (N_15793,N_10216,N_9119);
and U15794 (N_15794,N_10347,N_10853);
or U15795 (N_15795,N_10028,N_10629);
and U15796 (N_15796,N_11749,N_10645);
nor U15797 (N_15797,N_11016,N_9209);
nand U15798 (N_15798,N_10898,N_9589);
nor U15799 (N_15799,N_11714,N_8809);
nand U15800 (N_15800,N_9614,N_10517);
xnor U15801 (N_15801,N_11462,N_10715);
xor U15802 (N_15802,N_8458,N_10059);
nor U15803 (N_15803,N_11381,N_9485);
xor U15804 (N_15804,N_11284,N_10305);
or U15805 (N_15805,N_9218,N_8065);
or U15806 (N_15806,N_11743,N_8229);
or U15807 (N_15807,N_9302,N_11165);
or U15808 (N_15808,N_10755,N_10145);
xor U15809 (N_15809,N_11211,N_10200);
nand U15810 (N_15810,N_11712,N_11485);
nor U15811 (N_15811,N_8033,N_10730);
or U15812 (N_15812,N_9894,N_11921);
nor U15813 (N_15813,N_8930,N_9136);
and U15814 (N_15814,N_9329,N_8770);
or U15815 (N_15815,N_9820,N_9436);
nand U15816 (N_15816,N_10397,N_11244);
nand U15817 (N_15817,N_11841,N_10011);
nand U15818 (N_15818,N_11457,N_9016);
and U15819 (N_15819,N_8188,N_9988);
and U15820 (N_15820,N_9058,N_11832);
xor U15821 (N_15821,N_10310,N_11381);
nand U15822 (N_15822,N_8427,N_10507);
nand U15823 (N_15823,N_8220,N_8346);
or U15824 (N_15824,N_9700,N_11289);
and U15825 (N_15825,N_8965,N_8704);
nand U15826 (N_15826,N_11252,N_9792);
nand U15827 (N_15827,N_8772,N_9999);
nor U15828 (N_15828,N_9042,N_8641);
and U15829 (N_15829,N_9296,N_9675);
xnor U15830 (N_15830,N_10607,N_11080);
nor U15831 (N_15831,N_10257,N_10683);
and U15832 (N_15832,N_10754,N_9975);
or U15833 (N_15833,N_10845,N_8769);
or U15834 (N_15834,N_11228,N_9881);
or U15835 (N_15835,N_9061,N_10913);
and U15836 (N_15836,N_9635,N_9141);
and U15837 (N_15837,N_11885,N_8371);
nor U15838 (N_15838,N_11162,N_9593);
or U15839 (N_15839,N_11213,N_9056);
nand U15840 (N_15840,N_8600,N_11589);
nand U15841 (N_15841,N_9256,N_10767);
xnor U15842 (N_15842,N_11610,N_9158);
nand U15843 (N_15843,N_8776,N_9636);
nor U15844 (N_15844,N_8136,N_8885);
or U15845 (N_15845,N_9482,N_11367);
nor U15846 (N_15846,N_8755,N_8897);
nand U15847 (N_15847,N_11706,N_9369);
nor U15848 (N_15848,N_9744,N_8500);
and U15849 (N_15849,N_9515,N_11356);
and U15850 (N_15850,N_11833,N_10644);
and U15851 (N_15851,N_11882,N_9004);
or U15852 (N_15852,N_10206,N_10117);
nand U15853 (N_15853,N_8671,N_8755);
and U15854 (N_15854,N_8305,N_8748);
or U15855 (N_15855,N_8990,N_8843);
and U15856 (N_15856,N_8541,N_10179);
and U15857 (N_15857,N_8415,N_11415);
and U15858 (N_15858,N_9356,N_8664);
xnor U15859 (N_15859,N_8304,N_9537);
or U15860 (N_15860,N_11215,N_8040);
and U15861 (N_15861,N_8905,N_10317);
or U15862 (N_15862,N_10176,N_10985);
nor U15863 (N_15863,N_9923,N_10325);
or U15864 (N_15864,N_10884,N_8674);
or U15865 (N_15865,N_9916,N_10169);
nand U15866 (N_15866,N_9978,N_8975);
nand U15867 (N_15867,N_11136,N_11148);
or U15868 (N_15868,N_8253,N_10035);
nor U15869 (N_15869,N_10305,N_10815);
nand U15870 (N_15870,N_10417,N_9834);
and U15871 (N_15871,N_11852,N_9283);
nor U15872 (N_15872,N_8453,N_9605);
nand U15873 (N_15873,N_9470,N_10283);
nor U15874 (N_15874,N_11313,N_9418);
and U15875 (N_15875,N_10531,N_11208);
or U15876 (N_15876,N_10579,N_9749);
or U15877 (N_15877,N_11967,N_10647);
or U15878 (N_15878,N_8670,N_10948);
nor U15879 (N_15879,N_9798,N_8871);
and U15880 (N_15880,N_8503,N_11930);
and U15881 (N_15881,N_11292,N_11127);
nand U15882 (N_15882,N_11258,N_8789);
or U15883 (N_15883,N_8216,N_11343);
and U15884 (N_15884,N_11334,N_10311);
xnor U15885 (N_15885,N_9176,N_11511);
and U15886 (N_15886,N_10251,N_11978);
or U15887 (N_15887,N_9514,N_9745);
nor U15888 (N_15888,N_9228,N_11431);
nand U15889 (N_15889,N_10468,N_10606);
or U15890 (N_15890,N_8869,N_9918);
and U15891 (N_15891,N_11575,N_8985);
or U15892 (N_15892,N_10844,N_8518);
nand U15893 (N_15893,N_8095,N_8456);
and U15894 (N_15894,N_9279,N_8050);
nand U15895 (N_15895,N_9059,N_8722);
and U15896 (N_15896,N_8884,N_8408);
and U15897 (N_15897,N_10248,N_8105);
nor U15898 (N_15898,N_10230,N_9701);
or U15899 (N_15899,N_9102,N_10905);
or U15900 (N_15900,N_8421,N_11805);
xnor U15901 (N_15901,N_8720,N_10081);
nor U15902 (N_15902,N_8832,N_8640);
nand U15903 (N_15903,N_11017,N_11189);
nor U15904 (N_15904,N_10571,N_9768);
and U15905 (N_15905,N_10985,N_9639);
nand U15906 (N_15906,N_11980,N_9817);
and U15907 (N_15907,N_9556,N_10800);
nand U15908 (N_15908,N_11152,N_11499);
nand U15909 (N_15909,N_8755,N_8928);
and U15910 (N_15910,N_10773,N_9400);
and U15911 (N_15911,N_8931,N_11665);
nand U15912 (N_15912,N_9690,N_10104);
and U15913 (N_15913,N_11549,N_8884);
and U15914 (N_15914,N_10319,N_11000);
and U15915 (N_15915,N_9122,N_10939);
xor U15916 (N_15916,N_9615,N_11760);
nor U15917 (N_15917,N_11878,N_8407);
nand U15918 (N_15918,N_8710,N_11685);
and U15919 (N_15919,N_10576,N_10385);
nand U15920 (N_15920,N_8610,N_11330);
nor U15921 (N_15921,N_8631,N_10982);
nor U15922 (N_15922,N_10116,N_8472);
nor U15923 (N_15923,N_9557,N_8539);
nand U15924 (N_15924,N_8724,N_9456);
and U15925 (N_15925,N_8306,N_11567);
nand U15926 (N_15926,N_8663,N_9240);
nor U15927 (N_15927,N_9298,N_8831);
xnor U15928 (N_15928,N_10122,N_8270);
or U15929 (N_15929,N_8990,N_8425);
or U15930 (N_15930,N_10603,N_11376);
and U15931 (N_15931,N_11238,N_9095);
nand U15932 (N_15932,N_10400,N_9052);
nor U15933 (N_15933,N_8023,N_10280);
xnor U15934 (N_15934,N_9724,N_8667);
nand U15935 (N_15935,N_11114,N_8764);
or U15936 (N_15936,N_11077,N_11158);
and U15937 (N_15937,N_11938,N_9361);
nand U15938 (N_15938,N_9468,N_11062);
or U15939 (N_15939,N_11480,N_8534);
and U15940 (N_15940,N_8253,N_8938);
nand U15941 (N_15941,N_11648,N_10940);
nand U15942 (N_15942,N_11048,N_10363);
or U15943 (N_15943,N_8091,N_10803);
xor U15944 (N_15944,N_10012,N_9161);
xnor U15945 (N_15945,N_9521,N_8400);
or U15946 (N_15946,N_9221,N_8954);
nor U15947 (N_15947,N_10235,N_8553);
nor U15948 (N_15948,N_8336,N_9057);
or U15949 (N_15949,N_9455,N_11123);
or U15950 (N_15950,N_9424,N_10143);
nand U15951 (N_15951,N_11477,N_8792);
or U15952 (N_15952,N_8356,N_9697);
nand U15953 (N_15953,N_10024,N_11374);
and U15954 (N_15954,N_11171,N_9096);
nand U15955 (N_15955,N_11528,N_8593);
nand U15956 (N_15956,N_9110,N_9048);
and U15957 (N_15957,N_8977,N_9414);
or U15958 (N_15958,N_8431,N_9579);
nor U15959 (N_15959,N_9058,N_9828);
or U15960 (N_15960,N_10020,N_10401);
nor U15961 (N_15961,N_9419,N_8739);
nor U15962 (N_15962,N_8964,N_9295);
or U15963 (N_15963,N_8114,N_9131);
nor U15964 (N_15964,N_8217,N_8965);
xor U15965 (N_15965,N_9757,N_8010);
nor U15966 (N_15966,N_9111,N_10419);
nor U15967 (N_15967,N_9696,N_8762);
and U15968 (N_15968,N_8317,N_9836);
nand U15969 (N_15969,N_8069,N_9910);
nor U15970 (N_15970,N_10349,N_10075);
nand U15971 (N_15971,N_9856,N_9919);
or U15972 (N_15972,N_8053,N_10400);
xnor U15973 (N_15973,N_9873,N_10964);
or U15974 (N_15974,N_9565,N_9825);
and U15975 (N_15975,N_11567,N_11884);
and U15976 (N_15976,N_11124,N_8756);
nand U15977 (N_15977,N_11465,N_10963);
or U15978 (N_15978,N_11543,N_8953);
nor U15979 (N_15979,N_8223,N_11391);
and U15980 (N_15980,N_11381,N_11806);
xor U15981 (N_15981,N_10930,N_11272);
nand U15982 (N_15982,N_8526,N_11879);
nor U15983 (N_15983,N_8745,N_8099);
nor U15984 (N_15984,N_8182,N_10160);
or U15985 (N_15985,N_9466,N_8945);
or U15986 (N_15986,N_9812,N_10628);
or U15987 (N_15987,N_9564,N_9534);
nand U15988 (N_15988,N_10849,N_9241);
nand U15989 (N_15989,N_10926,N_8459);
or U15990 (N_15990,N_9600,N_9639);
or U15991 (N_15991,N_10050,N_10494);
nor U15992 (N_15992,N_9058,N_11376);
xnor U15993 (N_15993,N_8500,N_8426);
nor U15994 (N_15994,N_11391,N_8976);
or U15995 (N_15995,N_11334,N_8937);
and U15996 (N_15996,N_8185,N_9099);
or U15997 (N_15997,N_10350,N_10325);
nand U15998 (N_15998,N_8294,N_8154);
or U15999 (N_15999,N_11400,N_9949);
and U16000 (N_16000,N_13042,N_14912);
and U16001 (N_16001,N_15165,N_14178);
nor U16002 (N_16002,N_15519,N_14360);
and U16003 (N_16003,N_14816,N_14530);
xor U16004 (N_16004,N_12541,N_15436);
and U16005 (N_16005,N_15791,N_12552);
nand U16006 (N_16006,N_12377,N_12427);
or U16007 (N_16007,N_12472,N_15920);
or U16008 (N_16008,N_13079,N_15777);
nor U16009 (N_16009,N_13271,N_14999);
and U16010 (N_16010,N_15578,N_14885);
nor U16011 (N_16011,N_13788,N_15250);
nand U16012 (N_16012,N_13145,N_15941);
nor U16013 (N_16013,N_15674,N_15807);
nand U16014 (N_16014,N_13744,N_12771);
nand U16015 (N_16015,N_12682,N_14297);
xor U16016 (N_16016,N_14015,N_13436);
nor U16017 (N_16017,N_14818,N_12575);
nor U16018 (N_16018,N_14992,N_15369);
and U16019 (N_16019,N_13600,N_12261);
xor U16020 (N_16020,N_15365,N_15762);
xor U16021 (N_16021,N_13994,N_13093);
and U16022 (N_16022,N_14058,N_14959);
or U16023 (N_16023,N_15890,N_12819);
or U16024 (N_16024,N_14591,N_12964);
xnor U16025 (N_16025,N_15735,N_15356);
or U16026 (N_16026,N_14018,N_14861);
nand U16027 (N_16027,N_14216,N_14917);
and U16028 (N_16028,N_13048,N_14499);
nor U16029 (N_16029,N_14248,N_14078);
xnor U16030 (N_16030,N_12580,N_14919);
and U16031 (N_16031,N_13414,N_12642);
and U16032 (N_16032,N_15399,N_15146);
or U16033 (N_16033,N_13303,N_15912);
or U16034 (N_16034,N_15390,N_13666);
and U16035 (N_16035,N_14199,N_12816);
and U16036 (N_16036,N_12500,N_14269);
nand U16037 (N_16037,N_14024,N_13964);
nand U16038 (N_16038,N_13512,N_12911);
xor U16039 (N_16039,N_15852,N_13819);
or U16040 (N_16040,N_15232,N_13888);
nor U16041 (N_16041,N_13517,N_12561);
nand U16042 (N_16042,N_15543,N_13368);
or U16043 (N_16043,N_12968,N_13711);
or U16044 (N_16044,N_15593,N_15228);
and U16045 (N_16045,N_14138,N_15123);
and U16046 (N_16046,N_13805,N_14004);
nor U16047 (N_16047,N_14082,N_13510);
xnor U16048 (N_16048,N_13919,N_13406);
or U16049 (N_16049,N_13698,N_12509);
nand U16050 (N_16050,N_13962,N_15427);
or U16051 (N_16051,N_13828,N_15893);
nor U16052 (N_16052,N_15013,N_12923);
and U16053 (N_16053,N_12846,N_15090);
nor U16054 (N_16054,N_15173,N_13551);
xnor U16055 (N_16055,N_12494,N_15631);
or U16056 (N_16056,N_14697,N_14643);
and U16057 (N_16057,N_14104,N_15114);
xnor U16058 (N_16058,N_12461,N_14839);
nor U16059 (N_16059,N_14169,N_12961);
and U16060 (N_16060,N_14034,N_14096);
nor U16061 (N_16061,N_13712,N_12656);
or U16062 (N_16062,N_15469,N_14937);
and U16063 (N_16063,N_15715,N_13416);
nor U16064 (N_16064,N_13185,N_14606);
nand U16065 (N_16065,N_12717,N_13362);
and U16066 (N_16066,N_15281,N_12939);
or U16067 (N_16067,N_12808,N_12707);
and U16068 (N_16068,N_12774,N_14484);
xor U16069 (N_16069,N_13315,N_13407);
and U16070 (N_16070,N_15122,N_15442);
nor U16071 (N_16071,N_14263,N_12845);
nand U16072 (N_16072,N_12936,N_13216);
or U16073 (N_16073,N_13080,N_12640);
nor U16074 (N_16074,N_12438,N_13864);
nor U16075 (N_16075,N_15499,N_15358);
or U16076 (N_16076,N_12834,N_13261);
xor U16077 (N_16077,N_12206,N_12768);
nand U16078 (N_16078,N_13404,N_12751);
nor U16079 (N_16079,N_14645,N_12013);
and U16080 (N_16080,N_12087,N_13892);
nor U16081 (N_16081,N_15311,N_15523);
and U16082 (N_16082,N_14671,N_13931);
nor U16083 (N_16083,N_15875,N_14105);
and U16084 (N_16084,N_13942,N_14116);
or U16085 (N_16085,N_15615,N_12841);
nand U16086 (N_16086,N_12007,N_15301);
nand U16087 (N_16087,N_15116,N_12047);
nor U16088 (N_16088,N_15803,N_15914);
xnor U16089 (N_16089,N_12130,N_13502);
nor U16090 (N_16090,N_12770,N_14927);
nand U16091 (N_16091,N_14422,N_12594);
or U16092 (N_16092,N_14056,N_13693);
nand U16093 (N_16093,N_13907,N_14930);
xnor U16094 (N_16094,N_12672,N_12673);
nand U16095 (N_16095,N_13287,N_15848);
nand U16096 (N_16096,N_14938,N_14909);
xor U16097 (N_16097,N_15098,N_14650);
nor U16098 (N_16098,N_12071,N_12873);
nand U16099 (N_16099,N_12003,N_12469);
nand U16100 (N_16100,N_14412,N_15838);
nand U16101 (N_16101,N_15647,N_14546);
or U16102 (N_16102,N_14906,N_14226);
or U16103 (N_16103,N_14145,N_15652);
nand U16104 (N_16104,N_12838,N_14177);
nand U16105 (N_16105,N_15425,N_12467);
or U16106 (N_16106,N_15298,N_15183);
nand U16107 (N_16107,N_12277,N_15610);
or U16108 (N_16108,N_15211,N_14803);
nand U16109 (N_16109,N_14130,N_14785);
and U16110 (N_16110,N_14842,N_14021);
or U16111 (N_16111,N_13408,N_12378);
and U16112 (N_16112,N_15397,N_13754);
nand U16113 (N_16113,N_15200,N_12022);
xor U16114 (N_16114,N_14743,N_14010);
nand U16115 (N_16115,N_14005,N_13121);
nand U16116 (N_16116,N_15789,N_14037);
xnor U16117 (N_16117,N_15625,N_13196);
and U16118 (N_16118,N_15790,N_14926);
nand U16119 (N_16119,N_14060,N_15672);
nor U16120 (N_16120,N_14717,N_14899);
and U16121 (N_16121,N_15573,N_15779);
and U16122 (N_16122,N_14398,N_13629);
or U16123 (N_16123,N_12918,N_14332);
nand U16124 (N_16124,N_13901,N_15457);
and U16125 (N_16125,N_13974,N_12014);
nand U16126 (N_16126,N_15704,N_14473);
nor U16127 (N_16127,N_12476,N_13178);
xor U16128 (N_16128,N_12522,N_12898);
nor U16129 (N_16129,N_14335,N_15225);
xnor U16130 (N_16130,N_14465,N_14866);
and U16131 (N_16131,N_12681,N_15468);
and U16132 (N_16132,N_12966,N_12443);
or U16133 (N_16133,N_12279,N_12927);
and U16134 (N_16134,N_15651,N_12394);
or U16135 (N_16135,N_13365,N_15565);
nor U16136 (N_16136,N_12492,N_13897);
or U16137 (N_16137,N_14515,N_14444);
and U16138 (N_16138,N_12689,N_13138);
or U16139 (N_16139,N_13797,N_12280);
xor U16140 (N_16140,N_12629,N_15881);
and U16141 (N_16141,N_13949,N_13215);
nand U16142 (N_16142,N_12767,N_13734);
or U16143 (N_16143,N_13356,N_12214);
nor U16144 (N_16144,N_15895,N_15248);
and U16145 (N_16145,N_15039,N_13043);
or U16146 (N_16146,N_12411,N_12638);
nand U16147 (N_16147,N_12262,N_15155);
nand U16148 (N_16148,N_12082,N_13473);
nand U16149 (N_16149,N_12074,N_15398);
or U16150 (N_16150,N_15581,N_13589);
nand U16151 (N_16151,N_12035,N_15574);
nor U16152 (N_16152,N_15361,N_13274);
or U16153 (N_16153,N_13978,N_14517);
nor U16154 (N_16154,N_14521,N_13300);
nor U16155 (N_16155,N_13321,N_14958);
xnor U16156 (N_16156,N_15821,N_13339);
xor U16157 (N_16157,N_13157,N_14485);
or U16158 (N_16158,N_12941,N_15420);
and U16159 (N_16159,N_15302,N_14993);
or U16160 (N_16160,N_12112,N_13598);
or U16161 (N_16161,N_15156,N_14298);
and U16162 (N_16162,N_13490,N_12077);
nand U16163 (N_16163,N_12899,N_12361);
nand U16164 (N_16164,N_14972,N_12789);
and U16165 (N_16165,N_15926,N_14222);
and U16166 (N_16166,N_14935,N_14132);
or U16167 (N_16167,N_12205,N_15108);
and U16168 (N_16168,N_12307,N_14529);
nor U16169 (N_16169,N_12231,N_13470);
nor U16170 (N_16170,N_15406,N_15632);
and U16171 (N_16171,N_13397,N_13072);
nor U16172 (N_16172,N_14090,N_13681);
xnor U16173 (N_16173,N_15150,N_15772);
nor U16174 (N_16174,N_15115,N_13085);
nor U16175 (N_16175,N_14008,N_14244);
or U16176 (N_16176,N_13433,N_13278);
nor U16177 (N_16177,N_13735,N_12316);
nor U16178 (N_16178,N_13767,N_15382);
or U16179 (N_16179,N_12148,N_13521);
nand U16180 (N_16180,N_12983,N_13582);
nor U16181 (N_16181,N_15255,N_13903);
xnor U16182 (N_16182,N_15564,N_12286);
or U16183 (N_16183,N_14735,N_14555);
xnor U16184 (N_16184,N_12713,N_13979);
or U16185 (N_16185,N_12348,N_14512);
nor U16186 (N_16186,N_14769,N_12422);
xnor U16187 (N_16187,N_13289,N_15247);
nand U16188 (N_16188,N_13984,N_12926);
nor U16189 (N_16189,N_13799,N_15238);
or U16190 (N_16190,N_13933,N_15755);
nand U16191 (N_16191,N_15990,N_14347);
and U16192 (N_16192,N_12581,N_12624);
nand U16193 (N_16193,N_13493,N_14794);
nor U16194 (N_16194,N_12753,N_15995);
nand U16195 (N_16195,N_13911,N_12473);
nand U16196 (N_16196,N_13899,N_12989);
nand U16197 (N_16197,N_14337,N_13239);
and U16198 (N_16198,N_13360,N_13509);
nand U16199 (N_16199,N_12048,N_12298);
xnor U16200 (N_16200,N_12912,N_13625);
nand U16201 (N_16201,N_14148,N_12134);
or U16202 (N_16202,N_12549,N_14914);
or U16203 (N_16203,N_12437,N_13202);
or U16204 (N_16204,N_12894,N_13181);
nand U16205 (N_16205,N_12612,N_15078);
xnor U16206 (N_16206,N_13120,N_12216);
nand U16207 (N_16207,N_15191,N_12371);
or U16208 (N_16208,N_12879,N_12024);
nor U16209 (N_16209,N_14857,N_15186);
xor U16210 (N_16210,N_15166,N_14257);
and U16211 (N_16211,N_12357,N_15510);
nand U16212 (N_16212,N_12779,N_15158);
xor U16213 (N_16213,N_14789,N_13817);
nand U16214 (N_16214,N_15592,N_15252);
or U16215 (N_16215,N_15375,N_14406);
nand U16216 (N_16216,N_13420,N_14224);
nor U16217 (N_16217,N_14136,N_13373);
nand U16218 (N_16218,N_13870,N_12744);
nand U16219 (N_16219,N_12142,N_14664);
nand U16220 (N_16220,N_12023,N_14641);
or U16221 (N_16221,N_12881,N_14193);
nand U16222 (N_16222,N_13444,N_14330);
nand U16223 (N_16223,N_15962,N_12046);
nand U16224 (N_16224,N_13078,N_12765);
nor U16225 (N_16225,N_13268,N_14210);
nand U16226 (N_16226,N_13855,N_13111);
or U16227 (N_16227,N_14623,N_15571);
and U16228 (N_16228,N_15068,N_15045);
or U16229 (N_16229,N_12972,N_13527);
and U16230 (N_16230,N_12554,N_12855);
nand U16231 (N_16231,N_12419,N_13272);
nor U16232 (N_16232,N_12706,N_12167);
or U16233 (N_16233,N_14071,N_14172);
and U16234 (N_16234,N_14504,N_15575);
nor U16235 (N_16235,N_13658,N_14679);
nor U16236 (N_16236,N_13168,N_14251);
and U16237 (N_16237,N_14538,N_15272);
nand U16238 (N_16238,N_14859,N_14036);
nand U16239 (N_16239,N_13124,N_13208);
or U16240 (N_16240,N_15580,N_14590);
nor U16241 (N_16241,N_13973,N_12274);
nand U16242 (N_16242,N_14062,N_14092);
nor U16243 (N_16243,N_15378,N_13662);
xnor U16244 (N_16244,N_14585,N_14513);
and U16245 (N_16245,N_12909,N_15371);
nor U16246 (N_16246,N_13661,N_13818);
nand U16247 (N_16247,N_13602,N_13467);
and U16248 (N_16248,N_12959,N_13566);
xnor U16249 (N_16249,N_12539,N_13027);
or U16250 (N_16250,N_14615,N_15389);
nor U16251 (N_16251,N_15088,N_13677);
and U16252 (N_16252,N_13084,N_14001);
nand U16253 (N_16253,N_13190,N_12527);
nand U16254 (N_16254,N_13013,N_15874);
nor U16255 (N_16255,N_15682,N_13789);
nor U16256 (N_16256,N_13354,N_15133);
and U16257 (N_16257,N_12452,N_14273);
nand U16258 (N_16258,N_15143,N_12096);
nand U16259 (N_16259,N_13366,N_14173);
or U16260 (N_16260,N_12997,N_14271);
xnor U16261 (N_16261,N_12017,N_13073);
or U16262 (N_16262,N_12868,N_13871);
nor U16263 (N_16263,N_15236,N_12871);
xor U16264 (N_16264,N_12127,N_15760);
or U16265 (N_16265,N_12658,N_12268);
or U16266 (N_16266,N_14441,N_12585);
and U16267 (N_16267,N_13466,N_12178);
or U16268 (N_16268,N_12693,N_14532);
xor U16269 (N_16269,N_12141,N_12556);
nand U16270 (N_16270,N_12407,N_12697);
or U16271 (N_16271,N_12632,N_14265);
nor U16272 (N_16272,N_15027,N_13655);
nand U16273 (N_16273,N_15545,N_12347);
nand U16274 (N_16274,N_15898,N_13905);
or U16275 (N_16275,N_12525,N_15500);
or U16276 (N_16276,N_13573,N_15986);
or U16277 (N_16277,N_13972,N_14170);
nand U16278 (N_16278,N_14491,N_13916);
and U16279 (N_16279,N_13721,N_13331);
nor U16280 (N_16280,N_15982,N_13358);
nand U16281 (N_16281,N_15983,N_15911);
or U16282 (N_16282,N_13612,N_14647);
or U16283 (N_16283,N_15638,N_13488);
and U16284 (N_16284,N_15071,N_13890);
and U16285 (N_16285,N_15826,N_12172);
or U16286 (N_16286,N_15612,N_15641);
and U16287 (N_16287,N_15555,N_14738);
nor U16288 (N_16288,N_15622,N_13813);
nor U16289 (N_16289,N_12932,N_14890);
and U16290 (N_16290,N_14159,N_13590);
nor U16291 (N_16291,N_15100,N_12054);
nand U16292 (N_16292,N_14617,N_14425);
nor U16293 (N_16293,N_13485,N_14845);
nor U16294 (N_16294,N_15325,N_13513);
or U16295 (N_16295,N_14597,N_13082);
nor U16296 (N_16296,N_15263,N_14605);
and U16297 (N_16297,N_15416,N_14728);
nor U16298 (N_16298,N_14581,N_14374);
or U16299 (N_16299,N_13447,N_12062);
and U16300 (N_16300,N_12576,N_15554);
or U16301 (N_16301,N_13494,N_12613);
nand U16302 (N_16302,N_12780,N_13529);
nor U16303 (N_16303,N_12115,N_15728);
nor U16304 (N_16304,N_15331,N_15832);
and U16305 (N_16305,N_14762,N_12812);
and U16306 (N_16306,N_15797,N_13346);
nand U16307 (N_16307,N_13793,N_14046);
nor U16308 (N_16308,N_13379,N_15835);
nor U16309 (N_16309,N_12109,N_14867);
nor U16310 (N_16310,N_12244,N_15258);
or U16311 (N_16311,N_12353,N_13839);
nor U16312 (N_16312,N_14653,N_12967);
nor U16313 (N_16313,N_12907,N_15805);
nor U16314 (N_16314,N_13282,N_13332);
or U16315 (N_16315,N_15703,N_12844);
xor U16316 (N_16316,N_13647,N_14793);
and U16317 (N_16317,N_15992,N_15597);
nand U16318 (N_16318,N_13955,N_13099);
and U16319 (N_16319,N_14835,N_15276);
xnor U16320 (N_16320,N_12573,N_14883);
or U16321 (N_16321,N_15501,N_12444);
or U16322 (N_16322,N_12884,N_15530);
nor U16323 (N_16323,N_13290,N_15182);
and U16324 (N_16324,N_14249,N_12579);
and U16325 (N_16325,N_14250,N_15814);
and U16326 (N_16326,N_14746,N_12466);
nand U16327 (N_16327,N_14611,N_15199);
or U16328 (N_16328,N_14573,N_12042);
and U16329 (N_16329,N_14516,N_12962);
or U16330 (N_16330,N_12691,N_12839);
nor U16331 (N_16331,N_15877,N_14955);
xnor U16332 (N_16332,N_12451,N_15600);
or U16333 (N_16333,N_14439,N_13900);
and U16334 (N_16334,N_14457,N_13659);
nor U16335 (N_16335,N_12182,N_13320);
or U16336 (N_16336,N_12542,N_15752);
or U16337 (N_16337,N_14527,N_14236);
and U16338 (N_16338,N_14840,N_14979);
nand U16339 (N_16339,N_13259,N_12160);
or U16340 (N_16340,N_14002,N_14272);
or U16341 (N_16341,N_14213,N_14276);
and U16342 (N_16342,N_15010,N_15937);
nor U16343 (N_16343,N_12275,N_13001);
nand U16344 (N_16344,N_15538,N_15148);
or U16345 (N_16345,N_15285,N_12595);
or U16346 (N_16346,N_15967,N_12343);
nand U16347 (N_16347,N_12002,N_14299);
nor U16348 (N_16348,N_13774,N_14450);
or U16349 (N_16349,N_15536,N_14990);
or U16350 (N_16350,N_12931,N_15957);
nand U16351 (N_16351,N_14328,N_15900);
and U16352 (N_16352,N_15411,N_12184);
nor U16353 (N_16353,N_12583,N_13096);
xor U16354 (N_16354,N_13090,N_14395);
nand U16355 (N_16355,N_13419,N_13562);
and U16356 (N_16356,N_12795,N_15294);
nor U16357 (N_16357,N_13227,N_15401);
nor U16358 (N_16358,N_12135,N_13577);
and U16359 (N_16359,N_12462,N_12450);
or U16360 (N_16360,N_15707,N_12196);
nand U16361 (N_16361,N_14414,N_14825);
or U16362 (N_16362,N_13400,N_13234);
or U16363 (N_16363,N_15443,N_15453);
and U16364 (N_16364,N_14634,N_14290);
nor U16365 (N_16365,N_15084,N_13807);
and U16366 (N_16366,N_12031,N_14327);
xor U16367 (N_16367,N_13306,N_14201);
or U16368 (N_16368,N_12725,N_15408);
and U16369 (N_16369,N_12916,N_14542);
nor U16370 (N_16370,N_14855,N_12193);
nand U16371 (N_16371,N_15241,N_12772);
nand U16372 (N_16372,N_13389,N_13830);
nor U16373 (N_16373,N_15717,N_12039);
nor U16374 (N_16374,N_14241,N_15346);
nor U16375 (N_16375,N_13349,N_12705);
xnor U16376 (N_16376,N_12677,N_14106);
and U16377 (N_16377,N_13175,N_12714);
or U16378 (N_16378,N_12053,N_13731);
nor U16379 (N_16379,N_15393,N_13755);
or U16380 (N_16380,N_13434,N_13141);
nor U16381 (N_16381,N_12766,N_14903);
nand U16382 (N_16382,N_14551,N_13352);
xor U16383 (N_16383,N_14892,N_15763);
and U16384 (N_16384,N_14753,N_15337);
and U16385 (N_16385,N_12416,N_13055);
or U16386 (N_16386,N_14121,N_15491);
or U16387 (N_16387,N_13547,N_12732);
and U16388 (N_16388,N_12258,N_15840);
or U16389 (N_16389,N_15660,N_12091);
nand U16390 (N_16390,N_14278,N_13125);
nand U16391 (N_16391,N_15976,N_15938);
or U16392 (N_16392,N_14716,N_13772);
nor U16393 (N_16393,N_12558,N_15861);
or U16394 (N_16394,N_15781,N_13425);
nor U16395 (N_16395,N_15105,N_13429);
nand U16396 (N_16396,N_15945,N_13587);
xnor U16397 (N_16397,N_12238,N_12584);
nor U16398 (N_16398,N_15765,N_13336);
and U16399 (N_16399,N_14316,N_14287);
nor U16400 (N_16400,N_12257,N_12914);
nand U16401 (N_16401,N_12938,N_15894);
nand U16402 (N_16402,N_14695,N_12530);
nor U16403 (N_16403,N_12028,N_14811);
or U16404 (N_16404,N_12337,N_13476);
nand U16405 (N_16405,N_14809,N_13743);
nor U16406 (N_16406,N_13110,N_13136);
and U16407 (N_16407,N_12987,N_12078);
nand U16408 (N_16408,N_13249,N_13391);
nor U16409 (N_16409,N_13275,N_14792);
and U16410 (N_16410,N_15198,N_15452);
and U16411 (N_16411,N_15506,N_12308);
or U16412 (N_16412,N_12719,N_14045);
nand U16413 (N_16413,N_13804,N_15277);
and U16414 (N_16414,N_14974,N_12519);
nor U16415 (N_16415,N_12072,N_15730);
and U16416 (N_16416,N_12954,N_15630);
xnor U16417 (N_16417,N_15423,N_13236);
nor U16418 (N_16418,N_14949,N_14787);
xor U16419 (N_16419,N_14127,N_14771);
nand U16420 (N_16420,N_13155,N_12301);
or U16421 (N_16421,N_14920,N_15267);
nor U16422 (N_16422,N_14757,N_14505);
nand U16423 (N_16423,N_14514,N_14942);
xnor U16424 (N_16424,N_15395,N_12920);
nor U16425 (N_16425,N_15541,N_13678);
or U16426 (N_16426,N_14583,N_15194);
nor U16427 (N_16427,N_15761,N_14548);
and U16428 (N_16428,N_14747,N_12230);
nor U16429 (N_16429,N_13708,N_13238);
or U16430 (N_16430,N_13832,N_13671);
nand U16431 (N_16431,N_15409,N_14943);
and U16432 (N_16432,N_13646,N_15209);
nand U16433 (N_16433,N_12708,N_13390);
nand U16434 (N_16434,N_13019,N_13684);
or U16435 (N_16435,N_14913,N_15724);
nor U16436 (N_16436,N_15322,N_12496);
nand U16437 (N_16437,N_13049,N_14295);
nand U16438 (N_16438,N_13947,N_15218);
or U16439 (N_16439,N_15496,N_13021);
or U16440 (N_16440,N_15847,N_14904);
and U16441 (N_16441,N_14537,N_13538);
or U16442 (N_16442,N_13318,N_14989);
and U16443 (N_16443,N_12081,N_14593);
nor U16444 (N_16444,N_12250,N_15801);
or U16445 (N_16445,N_13226,N_14503);
nor U16446 (N_16446,N_14508,N_13615);
nor U16447 (N_16447,N_15429,N_13847);
nand U16448 (N_16448,N_13197,N_15745);
and U16449 (N_16449,N_14150,N_14688);
or U16450 (N_16450,N_14519,N_13139);
and U16451 (N_16451,N_12226,N_12123);
nor U16452 (N_16452,N_15953,N_12646);
or U16453 (N_16453,N_14985,N_12327);
nand U16454 (N_16454,N_14874,N_14385);
nand U16455 (N_16455,N_15678,N_15015);
or U16456 (N_16456,N_13965,N_13245);
nor U16457 (N_16457,N_14091,N_15863);
and U16458 (N_16458,N_12557,N_15141);
or U16459 (N_16459,N_13187,N_15658);
or U16460 (N_16460,N_13980,N_15869);
or U16461 (N_16461,N_13343,N_15112);
nand U16462 (N_16462,N_15074,N_15918);
and U16463 (N_16463,N_13308,N_15954);
nand U16464 (N_16464,N_14739,N_12571);
and U16465 (N_16465,N_14834,N_15036);
or U16466 (N_16466,N_14939,N_12246);
nor U16467 (N_16467,N_14559,N_12477);
nor U16468 (N_16468,N_13291,N_15721);
or U16469 (N_16469,N_13607,N_13829);
and U16470 (N_16470,N_13987,N_12104);
nor U16471 (N_16471,N_14107,N_12090);
nor U16472 (N_16472,N_12299,N_15726);
nand U16473 (N_16473,N_13191,N_14007);
nor U16474 (N_16474,N_15579,N_13727);
nand U16475 (N_16475,N_14858,N_14714);
nor U16476 (N_16476,N_13811,N_13667);
xor U16477 (N_16477,N_13388,N_14836);
and U16478 (N_16478,N_13382,N_13802);
and U16479 (N_16479,N_13653,N_15201);
xnor U16480 (N_16480,N_13702,N_15283);
or U16481 (N_16481,N_15534,N_13976);
and U16482 (N_16482,N_14802,N_12928);
and U16483 (N_16483,N_15739,N_13951);
nor U16484 (N_16484,N_14326,N_12190);
nand U16485 (N_16485,N_13293,N_14701);
or U16486 (N_16486,N_15160,N_14042);
and U16487 (N_16487,N_13355,N_13394);
or U16488 (N_16488,N_15539,N_13594);
xor U16489 (N_16489,N_12041,N_12146);
nor U16490 (N_16490,N_13679,N_13182);
xnor U16491 (N_16491,N_14409,N_13621);
nor U16492 (N_16492,N_14351,N_12864);
or U16493 (N_16493,N_13747,N_15226);
nand U16494 (N_16494,N_12102,N_14191);
nand U16495 (N_16495,N_15362,N_13761);
nand U16496 (N_16496,N_13775,N_12953);
nor U16497 (N_16497,N_13025,N_12153);
xor U16498 (N_16498,N_13007,N_14399);
or U16499 (N_16499,N_15537,N_13252);
nor U16500 (N_16500,N_14604,N_14182);
nand U16501 (N_16501,N_12040,N_13061);
nand U16502 (N_16502,N_14808,N_15246);
nand U16503 (N_16503,N_15109,N_13690);
and U16504 (N_16504,N_12164,N_12326);
or U16505 (N_16505,N_12797,N_12752);
nor U16506 (N_16506,N_12156,N_12428);
nor U16507 (N_16507,N_12034,N_12475);
nand U16508 (N_16508,N_15603,N_14511);
nor U16509 (N_16509,N_12630,N_13917);
nand U16510 (N_16510,N_15775,N_15125);
and U16511 (N_16511,N_15670,N_12796);
nor U16512 (N_16512,N_13045,N_14479);
nand U16513 (N_16513,N_13203,N_15430);
nand U16514 (N_16514,N_15619,N_12222);
and U16515 (N_16515,N_12290,N_14578);
or U16516 (N_16516,N_14383,N_13053);
nor U16517 (N_16517,N_13022,N_15551);
and U16518 (N_16518,N_15507,N_15136);
xor U16519 (N_16519,N_12215,N_12080);
and U16520 (N_16520,N_13288,N_13651);
nor U16521 (N_16521,N_12322,N_14194);
nor U16522 (N_16522,N_13132,N_12933);
nor U16523 (N_16523,N_13652,N_14049);
nand U16524 (N_16524,N_14097,N_14324);
nor U16525 (N_16525,N_13363,N_12482);
or U16526 (N_16526,N_13656,N_15007);
nor U16527 (N_16527,N_15489,N_12066);
xnor U16528 (N_16528,N_12934,N_13704);
and U16529 (N_16529,N_15134,N_13446);
or U16530 (N_16530,N_15870,N_15662);
and U16531 (N_16531,N_13322,N_13119);
nor U16532 (N_16532,N_13956,N_12903);
and U16533 (N_16533,N_12536,N_13581);
nor U16534 (N_16534,N_13044,N_15367);
and U16535 (N_16535,N_13569,N_14750);
nor U16536 (N_16536,N_13777,N_14626);
nor U16537 (N_16537,N_12850,N_15041);
xor U16538 (N_16538,N_12060,N_12978);
and U16539 (N_16539,N_14011,N_15035);
nand U16540 (N_16540,N_14970,N_13280);
or U16541 (N_16541,N_15683,N_12221);
xnor U16542 (N_16542,N_13489,N_15655);
nor U16543 (N_16543,N_14921,N_12151);
nand U16544 (N_16544,N_13012,N_13552);
xnor U16545 (N_16545,N_12203,N_15694);
nor U16546 (N_16546,N_14402,N_12370);
xnor U16547 (N_16547,N_15278,N_13867);
or U16548 (N_16548,N_14987,N_15341);
nand U16549 (N_16549,N_12075,N_14164);
nand U16550 (N_16550,N_15720,N_14065);
and U16551 (N_16551,N_12448,N_13134);
nand U16552 (N_16552,N_15697,N_15386);
or U16553 (N_16553,N_14427,N_13995);
or U16554 (N_16554,N_15618,N_15000);
nor U16555 (N_16555,N_14322,N_13159);
or U16556 (N_16556,N_15913,N_15486);
and U16557 (N_16557,N_14448,N_12463);
nand U16558 (N_16558,N_14415,N_12490);
nor U16559 (N_16559,N_12809,N_12293);
nor U16560 (N_16560,N_14779,N_14202);
nor U16561 (N_16561,N_14431,N_12947);
nand U16562 (N_16562,N_14539,N_12061);
or U16563 (N_16563,N_12833,N_14038);
nand U16564 (N_16564,N_13330,N_13403);
xnor U16565 (N_16565,N_14554,N_13849);
nand U16566 (N_16566,N_13455,N_13872);
and U16567 (N_16567,N_15271,N_14751);
nand U16568 (N_16568,N_12303,N_15607);
and U16569 (N_16569,N_13633,N_12567);
and U16570 (N_16570,N_15985,N_15930);
nand U16571 (N_16571,N_14397,N_12587);
and U16572 (N_16572,N_14873,N_12069);
nor U16573 (N_16573,N_14531,N_15048);
or U16574 (N_16574,N_15206,N_13458);
nor U16575 (N_16575,N_15640,N_14214);
and U16576 (N_16576,N_12424,N_15927);
xnor U16577 (N_16577,N_15628,N_14575);
nand U16578 (N_16578,N_14584,N_13885);
nor U16579 (N_16579,N_15586,N_14629);
and U16580 (N_16580,N_13398,N_14497);
nand U16581 (N_16581,N_14352,N_12999);
and U16582 (N_16582,N_15352,N_14693);
nor U16583 (N_16583,N_15946,N_13622);
nand U16584 (N_16584,N_14242,N_13840);
and U16585 (N_16585,N_14536,N_12212);
nor U16586 (N_16586,N_12234,N_15296);
nor U16587 (N_16587,N_15971,N_13639);
xnor U16588 (N_16588,N_14783,N_14986);
nor U16589 (N_16589,N_12996,N_13927);
and U16590 (N_16590,N_14944,N_13877);
nand U16591 (N_16591,N_12908,N_14733);
nand U16592 (N_16592,N_15403,N_12985);
nor U16593 (N_16593,N_14969,N_12175);
and U16594 (N_16594,N_14622,N_13768);
and U16595 (N_16595,N_14325,N_14123);
or U16596 (N_16596,N_14156,N_12895);
or U16597 (N_16597,N_13058,N_13592);
xnor U16598 (N_16598,N_15091,N_14962);
and U16599 (N_16599,N_14331,N_14195);
and U16600 (N_16600,N_14960,N_13483);
nand U16601 (N_16601,N_15069,N_13486);
or U16602 (N_16602,N_13235,N_15381);
or U16603 (N_16603,N_12217,N_12545);
nor U16604 (N_16604,N_15439,N_14988);
xor U16605 (N_16605,N_14219,N_15606);
xor U16606 (N_16606,N_13014,N_12946);
or U16607 (N_16607,N_13062,N_14160);
or U16608 (N_16608,N_13889,N_14703);
xor U16609 (N_16609,N_14149,N_13500);
nand U16610 (N_16610,N_14764,N_15157);
and U16611 (N_16611,N_14953,N_13195);
and U16612 (N_16612,N_15216,N_15103);
nand U16613 (N_16613,N_14947,N_12271);
xnor U16614 (N_16614,N_15679,N_13172);
and U16615 (N_16615,N_12239,N_12345);
nor U16616 (N_16616,N_13200,N_15659);
nand U16617 (N_16617,N_13454,N_12384);
or U16618 (N_16618,N_14680,N_14722);
or U16619 (N_16619,N_12826,N_14526);
nand U16620 (N_16620,N_13457,N_14685);
nor U16621 (N_16621,N_12517,N_12641);
or U16622 (N_16622,N_13162,N_12950);
xor U16623 (N_16623,N_12344,N_15195);
and U16624 (N_16624,N_14570,N_13514);
nand U16625 (N_16625,N_14209,N_14997);
or U16626 (N_16626,N_12396,N_12548);
and U16627 (N_16627,N_14469,N_12032);
nor U16628 (N_16628,N_14378,N_12568);
xor U16629 (N_16629,N_14040,N_12764);
nor U16630 (N_16630,N_14110,N_15653);
and U16631 (N_16631,N_14778,N_15623);
nor U16632 (N_16632,N_15964,N_13123);
nand U16633 (N_16633,N_12349,N_15701);
and U16634 (N_16634,N_13683,N_14403);
or U16635 (N_16635,N_13593,N_15584);
or U16636 (N_16636,N_15588,N_15117);
nor U16637 (N_16637,N_15667,N_15328);
or U16638 (N_16638,N_12199,N_14013);
nand U16639 (N_16639,N_14541,N_12661);
and U16640 (N_16640,N_12982,N_14487);
nor U16641 (N_16641,N_14852,N_14948);
and U16642 (N_16642,N_15958,N_15259);
and U16643 (N_16643,N_14261,N_12281);
and U16644 (N_16644,N_12897,N_12990);
and U16645 (N_16645,N_12524,N_14141);
nand U16646 (N_16646,N_14462,N_12674);
xnor U16647 (N_16647,N_12784,N_14870);
nand U16648 (N_16648,N_12169,N_13105);
nor U16649 (N_16649,N_13285,N_15513);
nor U16650 (N_16650,N_13542,N_12101);
and U16651 (N_16651,N_15079,N_12792);
and U16652 (N_16652,N_15925,N_12866);
or U16653 (N_16653,N_12389,N_13431);
nor U16654 (N_16654,N_14931,N_15208);
and U16655 (N_16655,N_14819,N_13660);
and U16656 (N_16656,N_13932,N_13359);
nor U16657 (N_16657,N_13101,N_13334);
or U16658 (N_16658,N_15274,N_15989);
nor U16659 (N_16659,N_15664,N_14983);
nand U16660 (N_16660,N_12533,N_15239);
nor U16661 (N_16661,N_15152,N_12940);
and U16662 (N_16662,N_13760,N_14708);
or U16663 (N_16663,N_15360,N_13904);
xnor U16664 (N_16664,N_15340,N_14118);
or U16665 (N_16665,N_15055,N_15014);
and U16666 (N_16666,N_13179,N_14343);
xnor U16667 (N_16667,N_14627,N_15016);
and U16668 (N_16668,N_14245,N_14369);
nand U16669 (N_16669,N_15891,N_15065);
nor U16670 (N_16670,N_12393,N_13461);
nand U16671 (N_16671,N_15922,N_14270);
nand U16672 (N_16672,N_15804,N_14044);
nor U16673 (N_16673,N_15076,N_15107);
xnor U16674 (N_16674,N_14731,N_12009);
or U16675 (N_16675,N_12659,N_13387);
and U16676 (N_16676,N_13224,N_12433);
or U16677 (N_16677,N_14994,N_13576);
nor U16678 (N_16678,N_14237,N_13674);
or U16679 (N_16679,N_12975,N_14940);
xnor U16680 (N_16680,N_14658,N_15189);
nor U16681 (N_16681,N_14232,N_13481);
nand U16682 (N_16682,N_14371,N_12597);
nor U16683 (N_16683,N_15560,N_12511);
nor U16684 (N_16684,N_13626,N_13383);
nor U16685 (N_16685,N_13596,N_15106);
nand U16686 (N_16686,N_15461,N_15407);
and U16687 (N_16687,N_14599,N_13170);
nor U16688 (N_16688,N_15478,N_15810);
nand U16689 (N_16689,N_15994,N_12731);
nand U16690 (N_16690,N_13153,N_12773);
xor U16691 (N_16691,N_15865,N_12255);
and U16692 (N_16692,N_12008,N_12056);
nand U16693 (N_16693,N_12037,N_12488);
nand U16694 (N_16694,N_15509,N_14644);
nor U16695 (N_16695,N_15960,N_14752);
nor U16696 (N_16696,N_14543,N_12586);
nor U16697 (N_16697,N_13729,N_14361);
and U16698 (N_16698,N_14660,N_15264);
xnor U16699 (N_16699,N_12405,N_15947);
nor U16700 (N_16700,N_13737,N_15860);
or U16701 (N_16701,N_12313,N_14375);
or U16702 (N_16702,N_13853,N_12949);
nor U16703 (N_16703,N_15326,N_13498);
and U16704 (N_16704,N_12386,N_13010);
and U16705 (N_16705,N_15737,N_12198);
xnor U16706 (N_16706,N_13097,N_14296);
nor U16707 (N_16707,N_15601,N_15943);
nand U16708 (N_16708,N_13201,N_14190);
and U16709 (N_16709,N_14081,N_12620);
nand U16710 (N_16710,N_15680,N_13199);
and U16711 (N_16711,N_12880,N_12232);
or U16712 (N_16712,N_14126,N_14509);
nand U16713 (N_16713,N_15729,N_14152);
nor U16714 (N_16714,N_13881,N_15394);
nor U16715 (N_16715,N_12098,N_15043);
or U16716 (N_16716,N_14657,N_14568);
and U16717 (N_16717,N_14689,N_12696);
nor U16718 (N_16718,N_15502,N_13395);
nand U16719 (N_16719,N_15567,N_13753);
nor U16720 (N_16720,N_13472,N_14321);
nand U16721 (N_16721,N_15719,N_14311);
nand U16722 (N_16722,N_14128,N_14984);
and U16723 (N_16723,N_15230,N_15793);
nor U16724 (N_16724,N_14767,N_15753);
or U16725 (N_16725,N_15351,N_13827);
or U16726 (N_16726,N_15636,N_15942);
or U16727 (N_16727,N_15313,N_15526);
xnor U16728 (N_16728,N_15059,N_12055);
or U16729 (N_16729,N_12700,N_14907);
xnor U16730 (N_16730,N_14877,N_15663);
nor U16731 (N_16731,N_15177,N_12197);
or U16732 (N_16732,N_15323,N_15227);
or U16733 (N_16733,N_15268,N_12011);
or U16734 (N_16734,N_12088,N_15621);
and U16735 (N_16735,N_13415,N_14745);
and U16736 (N_16736,N_14613,N_14453);
nor U16737 (N_16737,N_14871,N_12363);
xor U16738 (N_16738,N_14064,N_13757);
and U16739 (N_16739,N_13535,N_13148);
nor U16740 (N_16740,N_14329,N_13628);
or U16741 (N_16741,N_13005,N_13723);
and U16742 (N_16742,N_15193,N_12382);
and U16743 (N_16743,N_14493,N_12431);
or U16744 (N_16744,N_12029,N_14279);
or U16745 (N_16745,N_14829,N_14387);
and U16746 (N_16746,N_12319,N_13939);
or U16747 (N_16747,N_14699,N_15347);
or U16748 (N_16748,N_13294,N_15689);
xnor U16749 (N_16749,N_13545,N_15768);
and U16750 (N_16750,N_12885,N_14725);
nor U16751 (N_16751,N_12667,N_12671);
and U16752 (N_16752,N_13675,N_13051);
nor U16753 (N_16753,N_15288,N_15487);
nor U16754 (N_16754,N_14507,N_12742);
nor U16755 (N_16755,N_14633,N_15306);
xor U16756 (N_16756,N_14359,N_14346);
nor U16757 (N_16757,N_13109,N_15237);
nor U16758 (N_16758,N_15092,N_12489);
nor U16759 (N_16759,N_15656,N_12265);
nand U16760 (N_16760,N_15727,N_13077);
and U16761 (N_16761,N_14309,N_12577);
nor U16762 (N_16762,N_14975,N_13525);
and U16763 (N_16763,N_13207,N_13841);
and U16764 (N_16764,N_12177,N_13015);
xor U16765 (N_16765,N_13838,N_13026);
and U16766 (N_16766,N_13624,N_14791);
nor U16767 (N_16767,N_12550,N_14355);
nand U16768 (N_16768,N_13113,N_12603);
or U16769 (N_16769,N_15939,N_13060);
xor U16770 (N_16770,N_13225,N_14492);
or U16771 (N_16771,N_14596,N_13011);
and U16772 (N_16772,N_14313,N_12016);
nand U16773 (N_16773,N_15072,N_14965);
nand U16774 (N_16774,N_12922,N_14486);
xnor U16775 (N_16775,N_12817,N_15096);
nor U16776 (N_16776,N_12976,N_13848);
or U16777 (N_16777,N_12683,N_14678);
nor U16778 (N_16778,N_14929,N_12304);
nor U16779 (N_16779,N_13851,N_14820);
nor U16780 (N_16780,N_12644,N_12183);
nor U16781 (N_16781,N_13971,N_14882);
and U16782 (N_16782,N_15970,N_12333);
nand U16783 (N_16783,N_13020,N_14934);
or U16784 (N_16784,N_13808,N_14610);
and U16785 (N_16785,N_15540,N_14982);
or U16786 (N_16786,N_15005,N_13710);
and U16787 (N_16787,N_15149,N_15451);
and U16788 (N_16788,N_14677,N_13967);
nor U16789 (N_16789,N_12079,N_14200);
and U16790 (N_16790,N_15254,N_14307);
or U16791 (N_16791,N_14482,N_13518);
nor U16792 (N_16792,N_14977,N_12684);
and U16793 (N_16793,N_15514,N_15853);
xor U16794 (N_16794,N_14589,N_13924);
nand U16795 (N_16795,N_13887,N_13393);
or U16796 (N_16796,N_14922,N_14300);
or U16797 (N_16797,N_12486,N_12403);
nor U16798 (N_16798,N_12388,N_12295);
and U16799 (N_16799,N_12690,N_14267);
nand U16800 (N_16800,N_14282,N_14340);
or U16801 (N_16801,N_15661,N_13244);
nand U16802 (N_16802,N_12830,N_14086);
nand U16803 (N_16803,N_12836,N_13815);
or U16804 (N_16804,N_12692,N_15978);
nor U16805 (N_16805,N_12560,N_15466);
or U16806 (N_16806,N_12617,N_12588);
xnor U16807 (N_16807,N_13559,N_12325);
nand U16808 (N_16808,N_14162,N_13118);
and U16809 (N_16809,N_14954,N_14085);
or U16810 (N_16810,N_15746,N_15144);
nor U16811 (N_16811,N_15479,N_15290);
nor U16812 (N_16812,N_14243,N_12678);
xnor U16813 (N_16813,N_13686,N_12651);
or U16814 (N_16814,N_13948,N_12351);
nand U16815 (N_16815,N_15883,N_13990);
nand U16816 (N_16816,N_13114,N_13836);
nand U16817 (N_16817,N_13324,N_12179);
nor U16818 (N_16818,N_13350,N_14916);
or U16819 (N_16819,N_12759,N_14449);
nand U16820 (N_16820,N_12804,N_14831);
nand U16821 (N_16821,N_14456,N_15187);
or U16822 (N_16822,N_12191,N_15711);
or U16823 (N_16823,N_13893,N_14619);
or U16824 (N_16824,N_13209,N_13742);
nor U16825 (N_16825,N_12979,N_15759);
nand U16826 (N_16826,N_12703,N_12366);
nor U16827 (N_16827,N_15676,N_15110);
and U16828 (N_16828,N_12018,N_12149);
nand U16829 (N_16829,N_13206,N_12487);
xnor U16830 (N_16830,N_13663,N_12170);
nand U16831 (N_16831,N_13773,N_15033);
and U16832 (N_16832,N_14252,N_12064);
nand U16833 (N_16833,N_14967,N_15410);
and U16834 (N_16834,N_15882,N_13254);
nand U16835 (N_16835,N_13374,N_15441);
and U16836 (N_16836,N_12137,N_15857);
or U16837 (N_16837,N_13564,N_12263);
or U16838 (N_16838,N_15314,N_15511);
and U16839 (N_16839,N_14665,N_13692);
and U16840 (N_16840,N_13765,N_12249);
nor U16841 (N_16841,N_12902,N_13325);
and U16842 (N_16842,N_13642,N_14628);
nor U16843 (N_16843,N_14824,N_15731);
nand U16844 (N_16844,N_15696,N_13649);
or U16845 (N_16845,N_13353,N_13076);
nand U16846 (N_16846,N_12485,N_14095);
xnor U16847 (N_16847,N_12831,N_12952);
and U16848 (N_16848,N_14277,N_15687);
nand U16849 (N_16849,N_12663,N_12910);
nand U16850 (N_16850,N_14404,N_12970);
nor U16851 (N_16851,N_12716,N_13304);
and U16852 (N_16852,N_12284,N_12019);
or U16853 (N_16853,N_15368,N_14288);
xnor U16854 (N_16854,N_12501,N_15244);
and U16855 (N_16855,N_12745,N_15903);
nor U16856 (N_16856,N_12633,N_12317);
or U16857 (N_16857,N_14238,N_15716);
or U16858 (N_16858,N_12173,N_14998);
and U16859 (N_16859,N_12757,N_15851);
nand U16860 (N_16860,N_13796,N_14721);
nand U16861 (N_16861,N_14853,N_14968);
nor U16862 (N_16862,N_12698,N_12832);
and U16863 (N_16863,N_15018,N_13557);
nor U16864 (N_16864,N_13122,N_12562);
or U16865 (N_16865,N_14365,N_15334);
xnor U16866 (N_16866,N_12685,N_14886);
nand U16867 (N_16867,N_14142,N_15415);
and U16868 (N_16868,N_14391,N_14592);
nand U16869 (N_16869,N_15137,N_13295);
and U16870 (N_16870,N_15372,N_12657);
nor U16871 (N_16871,N_12676,N_15384);
or U16872 (N_16872,N_13714,N_13426);
nor U16873 (N_16873,N_14759,N_13140);
nor U16874 (N_16874,N_15700,N_15448);
and U16875 (N_16875,N_12128,N_13724);
and U16876 (N_16876,N_14995,N_12125);
xnor U16877 (N_16877,N_13198,N_14120);
nor U16878 (N_16878,N_15587,N_15585);
and U16879 (N_16879,N_15093,N_15508);
nor U16880 (N_16880,N_12951,N_12610);
or U16881 (N_16881,N_12516,N_12094);
and U16882 (N_16882,N_15188,N_12122);
and U16883 (N_16883,N_15126,N_14734);
nand U16884 (N_16884,N_15907,N_14715);
nand U16885 (N_16885,N_15822,N_13459);
nand U16886 (N_16886,N_13083,N_15404);
nand U16887 (N_16887,N_14319,N_13780);
nor U16888 (N_16888,N_15080,N_14698);
nand U16889 (N_16889,N_13707,N_14996);
and U16890 (N_16890,N_12171,N_15047);
nor U16891 (N_16891,N_12900,N_15030);
nor U16892 (N_16892,N_13722,N_14174);
nand U16893 (N_16893,N_14668,N_14227);
or U16894 (N_16894,N_13725,N_12455);
nand U16895 (N_16895,N_14155,N_14893);
nor U16896 (N_16896,N_15725,N_12207);
or U16897 (N_16897,N_15529,N_12848);
and U16898 (N_16898,N_13469,N_12645);
xnor U16899 (N_16899,N_14868,N_14171);
and U16900 (N_16900,N_15289,N_14719);
xor U16901 (N_16901,N_13066,N_15796);
nor U16902 (N_16902,N_15533,N_15355);
and U16903 (N_16903,N_13879,N_12110);
nand U16904 (N_16904,N_12373,N_14786);
and U16905 (N_16905,N_15798,N_14911);
and U16906 (N_16906,N_14524,N_15952);
and U16907 (N_16907,N_12810,N_12253);
nand U16908 (N_16908,N_12593,N_12468);
and U16909 (N_16909,N_12418,N_12572);
nand U16910 (N_16910,N_15896,N_15935);
and U16911 (N_16911,N_14452,N_13608);
nand U16912 (N_16912,N_14609,N_13484);
and U16913 (N_16913,N_14639,N_12605);
or U16914 (N_16914,N_13220,N_15923);
nor U16915 (N_16915,N_15494,N_12491);
nor U16916 (N_16916,N_13137,N_15396);
and U16917 (N_16917,N_15295,N_12737);
nor U16918 (N_16918,N_15624,N_13165);
nor U16919 (N_16919,N_15598,N_15897);
or U16920 (N_16920,N_14872,N_12241);
and U16921 (N_16921,N_13654,N_13378);
or U16922 (N_16922,N_13597,N_15431);
nor U16923 (N_16923,N_12718,N_12166);
or U16924 (N_16924,N_13739,N_15138);
and U16925 (N_16925,N_12086,N_13409);
xnor U16926 (N_16926,N_12869,N_13070);
nand U16927 (N_16927,N_14534,N_14389);
nand U16928 (N_16928,N_13413,N_15032);
and U16929 (N_16929,N_15419,N_13543);
xor U16930 (N_16930,N_15799,N_12276);
xor U16931 (N_16931,N_14255,N_13998);
or U16932 (N_16932,N_12459,N_12777);
nand U16933 (N_16933,N_13344,N_12420);
nor U16934 (N_16934,N_13309,N_13064);
and U16935 (N_16935,N_12600,N_14754);
nand U16936 (N_16936,N_15974,N_14125);
nor U16937 (N_16937,N_15180,N_15335);
nand U16938 (N_16938,N_12408,N_12748);
or U16939 (N_16939,N_12248,N_14557);
or U16940 (N_16940,N_13863,N_14135);
nor U16941 (N_16941,N_15308,N_14663);
nor U16942 (N_16942,N_15026,N_15374);
xnor U16943 (N_16943,N_14562,N_15495);
and U16944 (N_16944,N_12944,N_12800);
nand U16945 (N_16945,N_15712,N_14362);
and U16946 (N_16946,N_12650,N_13834);
or U16947 (N_16947,N_13632,N_13161);
nand U16948 (N_16948,N_13763,N_15317);
nor U16949 (N_16949,N_12302,N_12935);
or U16950 (N_16950,N_12120,N_13301);
or U16951 (N_16951,N_12105,N_14586);
nor U16952 (N_16952,N_13380,N_12240);
or U16953 (N_16953,N_15673,N_13981);
nand U16954 (N_16954,N_12315,N_12038);
nand U16955 (N_16955,N_14518,N_14447);
or U16956 (N_16956,N_13563,N_15159);
nor U16957 (N_16957,N_12824,N_15740);
nor U16958 (N_16958,N_14229,N_13218);
and U16959 (N_16959,N_12224,N_15280);
and U16960 (N_16960,N_13539,N_13730);
or U16961 (N_16961,N_15644,N_15969);
and U16962 (N_16962,N_13277,N_14614);
and U16963 (N_16963,N_14020,N_14849);
nor U16964 (N_16964,N_12412,N_13950);
or U16965 (N_16965,N_15140,N_12729);
and U16966 (N_16966,N_15884,N_14780);
nand U16967 (N_16967,N_15792,N_15286);
nand U16968 (N_16968,N_12311,N_12878);
nand U16969 (N_16969,N_12460,N_13925);
or U16970 (N_16970,N_15997,N_12504);
xnor U16971 (N_16971,N_13800,N_12449);
or U16972 (N_16972,N_13610,N_13283);
and U16973 (N_16973,N_14259,N_15129);
and U16974 (N_16974,N_13479,N_15359);
nand U16975 (N_16975,N_15906,N_14776);
nand U16976 (N_16976,N_13116,N_13549);
or U16977 (N_16977,N_12870,N_12945);
nand U16978 (N_16978,N_14342,N_15433);
nand U16979 (N_16979,N_12905,N_12859);
or U16980 (N_16980,N_13865,N_15470);
or U16981 (N_16981,N_13627,N_15836);
nor U16982 (N_16982,N_12758,N_13748);
nor U16983 (N_16983,N_13574,N_12103);
nor U16984 (N_16984,N_13826,N_15979);
nor U16985 (N_16985,N_12709,N_12746);
and U16986 (N_16986,N_14083,N_15748);
nand U16987 (N_16987,N_14736,N_13620);
nand U16988 (N_16988,N_12030,N_14436);
xnor U16989 (N_16989,N_12876,N_12336);
nand U16990 (N_16990,N_13749,N_15073);
or U16991 (N_16991,N_15788,N_12743);
nand U16992 (N_16992,N_12842,N_14050);
nor U16993 (N_16993,N_12998,N_12306);
or U16994 (N_16994,N_13131,N_14687);
nor U16995 (N_16995,N_15544,N_15101);
or U16996 (N_16996,N_12986,N_12528);
and U16997 (N_16997,N_12592,N_14292);
nand U16998 (N_16998,N_12722,N_14467);
and U16999 (N_16999,N_13936,N_14880);
and U17000 (N_17000,N_15060,N_14476);
xnor U17001 (N_17001,N_15097,N_13882);
or U17002 (N_17002,N_13107,N_14401);
xor U17003 (N_17003,N_13558,N_12465);
and U17004 (N_17004,N_14055,N_13613);
and U17005 (N_17005,N_12085,N_14964);
and U17006 (N_17006,N_14827,N_15710);
xor U17007 (N_17007,N_14129,N_12379);
and U17008 (N_17008,N_12606,N_13709);
nand U17009 (N_17009,N_12497,N_12470);
or U17010 (N_17010,N_13791,N_15202);
or U17011 (N_17011,N_15284,N_14800);
or U17012 (N_17012,N_12761,N_14830);
and U17013 (N_17013,N_12329,N_13074);
nand U17014 (N_17014,N_12512,N_15858);
nor U17015 (N_17015,N_15245,N_14247);
and U17016 (N_17016,N_15981,N_14410);
nand U17017 (N_17017,N_12180,N_15344);
or U17018 (N_17018,N_13063,N_12825);
and U17019 (N_17019,N_12006,N_12863);
xnor U17020 (N_17020,N_14556,N_13126);
nand U17021 (N_17021,N_13617,N_14897);
xnor U17022 (N_17022,N_14221,N_13237);
nor U17023 (N_17023,N_14720,N_12464);
xnor U17024 (N_17024,N_14284,N_12442);
or U17025 (N_17025,N_13641,N_13522);
or U17026 (N_17026,N_14167,N_15319);
nor U17027 (N_17027,N_14694,N_12223);
or U17028 (N_17028,N_14094,N_15795);
or U17029 (N_17029,N_12152,N_12155);
and U17030 (N_17030,N_12202,N_14344);
xnor U17031 (N_17031,N_13528,N_12694);
nand U17032 (N_17032,N_15559,N_14052);
or U17033 (N_17033,N_14723,N_15872);
and U17034 (N_17034,N_15757,N_15657);
nor U17035 (N_17035,N_14063,N_15521);
xnor U17036 (N_17036,N_15732,N_12887);
nand U17037 (N_17037,N_12332,N_15028);
or U17038 (N_17038,N_15966,N_14165);
nor U17039 (N_17039,N_12654,N_15400);
nand U17040 (N_17040,N_15275,N_15984);
or U17041 (N_17041,N_14881,N_13251);
nor U17042 (N_17042,N_12805,N_15082);
nor U17043 (N_17043,N_12245,N_14451);
and U17044 (N_17044,N_12358,N_14370);
nor U17045 (N_17045,N_14446,N_13689);
nand U17046 (N_17046,N_13694,N_14702);
and U17047 (N_17047,N_14027,N_15392);
nor U17048 (N_17048,N_15050,N_13006);
nor U17049 (N_17049,N_13375,N_14782);
nor U17050 (N_17050,N_13319,N_13385);
and U17051 (N_17051,N_12799,N_15418);
and U17052 (N_17052,N_12387,N_15493);
or U17053 (N_17053,N_15975,N_14233);
nand U17054 (N_17054,N_13717,N_14246);
and U17055 (N_17055,N_13194,N_13957);
nor U17056 (N_17056,N_14798,N_15916);
nand U17057 (N_17057,N_13174,N_12334);
and U17058 (N_17058,N_14367,N_14574);
nand U17059 (N_17059,N_13367,N_13524);
and U17060 (N_17060,N_12647,N_13586);
xor U17061 (N_17061,N_13384,N_13214);
or U17062 (N_17062,N_15197,N_14718);
and U17063 (N_17063,N_14183,N_12793);
nor U17064 (N_17064,N_15681,N_14433);
nor U17065 (N_17065,N_13842,N_15176);
and U17066 (N_17066,N_13668,N_13738);
nand U17067 (N_17067,N_14266,N_13664);
or U17068 (N_17068,N_12523,N_15965);
or U17069 (N_17069,N_15940,N_14775);
and U17070 (N_17070,N_12117,N_15061);
and U17071 (N_17071,N_13229,N_12305);
and U17072 (N_17072,N_15162,N_15888);
or U17073 (N_17073,N_15262,N_12631);
and U17074 (N_17074,N_12818,N_13432);
and U17075 (N_17075,N_14602,N_12392);
or U17076 (N_17076,N_13696,N_14197);
nor U17077 (N_17077,N_15558,N_14131);
and U17078 (N_17078,N_14280,N_15695);
nor U17079 (N_17079,N_13776,N_14624);
and U17080 (N_17080,N_14192,N_15932);
nand U17081 (N_17081,N_13790,N_13523);
nand U17082 (N_17082,N_12665,N_12445);
nand U17083 (N_17083,N_13002,N_15482);
xor U17084 (N_17084,N_15377,N_15528);
and U17085 (N_17085,N_13691,N_12318);
or U17086 (N_17086,N_12108,N_14844);
nor U17087 (N_17087,N_13801,N_15570);
nor U17088 (N_17088,N_12121,N_13039);
and U17089 (N_17089,N_13634,N_13150);
nand U17090 (N_17090,N_12192,N_13423);
nor U17091 (N_17091,N_15261,N_15312);
or U17092 (N_17092,N_14674,N_12484);
nand U17093 (N_17093,N_14396,N_15214);
nor U17094 (N_17094,N_12237,N_12296);
nand U17095 (N_17095,N_13144,N_15062);
and U17096 (N_17096,N_15111,N_15871);
nand U17097 (N_17097,N_12331,N_14860);
or U17098 (N_17098,N_15233,N_12020);
xnor U17099 (N_17099,N_14041,N_13327);
nor U17100 (N_17100,N_12131,N_12874);
nor U17101 (N_17101,N_13531,N_13741);
and U17102 (N_17102,N_15462,N_13944);
nand U17103 (N_17103,N_15025,N_15635);
or U17104 (N_17104,N_14686,N_15594);
nor U17105 (N_17105,N_15809,N_13784);
or U17106 (N_17106,N_15446,N_13695);
and U17107 (N_17107,N_15190,N_15566);
nand U17108 (N_17108,N_12021,N_12749);
and U17109 (N_17109,N_15044,N_14423);
or U17110 (N_17110,N_12555,N_13405);
nand U17111 (N_17111,N_12837,N_13418);
and U17112 (N_17112,N_14498,N_14748);
and U17113 (N_17113,N_12994,N_13183);
or U17114 (N_17114,N_14978,N_12350);
nand U17115 (N_17115,N_14019,N_13969);
nor U17116 (N_17116,N_12247,N_13030);
nand U17117 (N_17117,N_15669,N_14413);
xor U17118 (N_17118,N_15161,N_13785);
nor U17119 (N_17119,N_14435,N_14260);
or U17120 (N_17120,N_15944,N_15310);
and U17121 (N_17121,N_15063,N_14638);
and U17122 (N_17122,N_13928,N_13312);
nor U17123 (N_17123,N_12188,N_12145);
xnor U17124 (N_17124,N_15023,N_13792);
nand U17125 (N_17125,N_14442,N_14478);
or U17126 (N_17126,N_14823,N_12520);
and U17127 (N_17127,N_14832,N_14601);
and U17128 (N_17128,N_12404,N_14826);
nand U17129 (N_17129,N_13507,N_14134);
or U17130 (N_17130,N_14817,N_15650);
xor U17131 (N_17131,N_15388,N_14729);
nand U17132 (N_17132,N_13716,N_15643);
nor U17133 (N_17133,N_15666,N_12636);
nand U17134 (N_17134,N_13396,N_12385);
or U17135 (N_17135,N_12113,N_12243);
and U17136 (N_17136,N_13158,N_14048);
or U17137 (N_17137,N_13604,N_15304);
nor U17138 (N_17138,N_14198,N_12901);
nand U17139 (N_17139,N_15154,N_15366);
or U17140 (N_17140,N_13102,N_13823);
nor U17141 (N_17141,N_13794,N_14124);
nor U17142 (N_17142,N_13719,N_15145);
or U17143 (N_17143,N_12794,N_15709);
nand U17144 (N_17144,N_12679,N_13875);
and U17145 (N_17145,N_12354,N_15736);
nand U17146 (N_17146,N_12049,N_13004);
and U17147 (N_17147,N_12957,N_15391);
and U17148 (N_17148,N_15629,N_12168);
and U17149 (N_17149,N_12776,N_14308);
nor U17150 (N_17150,N_14496,N_14281);
nor U17151 (N_17151,N_12702,N_12189);
xnor U17152 (N_17152,N_13682,N_15488);
xor U17153 (N_17153,N_13029,N_13670);
or U17154 (N_17154,N_15831,N_12415);
and U17155 (N_17155,N_15605,N_12724);
or U17156 (N_17156,N_14579,N_12829);
nand U17157 (N_17157,N_14683,N_14026);
or U17158 (N_17158,N_15864,N_14087);
or U17159 (N_17159,N_12896,N_12390);
nand U17160 (N_17160,N_15842,N_13862);
or U17161 (N_17161,N_13970,N_15303);
nand U17162 (N_17162,N_13333,N_14067);
nor U17163 (N_17163,N_14077,N_13439);
and U17164 (N_17164,N_14407,N_15034);
or U17165 (N_17165,N_15800,N_15645);
or U17166 (N_17166,N_12447,N_12930);
or U17167 (N_17167,N_13036,N_13635);
and U17168 (N_17168,N_13345,N_15616);
and U17169 (N_17169,N_14612,N_15617);
or U17170 (N_17170,N_12204,N_12383);
and U17171 (N_17171,N_14656,N_15477);
and U17172 (N_17172,N_13920,N_13856);
xnor U17173 (N_17173,N_13898,N_12626);
nand U17174 (N_17174,N_12278,N_13128);
nor U17175 (N_17175,N_15020,N_14813);
and U17176 (N_17176,N_12111,N_15196);
nor U17177 (N_17177,N_14179,N_12015);
or U17178 (N_17178,N_15602,N_12067);
nor U17179 (N_17179,N_13501,N_12309);
and U17180 (N_17180,N_13601,N_13231);
nand U17181 (N_17181,N_13341,N_13764);
or U17182 (N_17182,N_14025,N_15021);
nand U17183 (N_17183,N_14108,N_14477);
and U17184 (N_17184,N_12680,N_13733);
and U17185 (N_17185,N_13565,N_14189);
nor U17186 (N_17186,N_14418,N_14682);
and U17187 (N_17187,N_14293,N_15332);
xnor U17188 (N_17188,N_15119,N_15758);
nand U17189 (N_17189,N_14372,N_13266);
and U17190 (N_17190,N_15234,N_13445);
nor U17191 (N_17191,N_14704,N_12143);
xnor U17192 (N_17192,N_13438,N_15009);
xor U17193 (N_17193,N_13024,N_14713);
and U17194 (N_17194,N_12948,N_12251);
nor U17195 (N_17195,N_12675,N_13089);
nor U17196 (N_17196,N_13258,N_14523);
nor U17197 (N_17197,N_12782,N_14569);
xnor U17198 (N_17198,N_12712,N_15802);
xnor U17199 (N_17199,N_13894,N_12139);
nor U17200 (N_17200,N_14766,N_12297);
nand U17201 (N_17201,N_15012,N_15668);
or U17202 (N_17202,N_12045,N_14147);
and U17203 (N_17203,N_14380,N_12161);
nor U17204 (N_17204,N_15124,N_14706);
and U17205 (N_17205,N_15385,N_14463);
nor U17206 (N_17206,N_14305,N_14426);
and U17207 (N_17207,N_15693,N_13427);
nor U17208 (N_17208,N_12283,N_15928);
or U17209 (N_17209,N_13770,N_13448);
nor U17210 (N_17210,N_12057,N_13779);
nand U17211 (N_17211,N_15557,N_14133);
and U17212 (N_17212,N_14039,N_12854);
nor U17213 (N_17213,N_13534,N_15620);
nand U17214 (N_17214,N_12735,N_13392);
nor U17215 (N_17215,N_15449,N_15878);
nor U17216 (N_17216,N_14936,N_14690);
or U17217 (N_17217,N_15130,N_13213);
and U17218 (N_17218,N_15873,N_12441);
xor U17219 (N_17219,N_15424,N_12346);
nor U17220 (N_17220,N_13934,N_13985);
and U17221 (N_17221,N_14341,N_15774);
nand U17222 (N_17222,N_13503,N_14846);
nand U17223 (N_17223,N_13003,N_12655);
or U17224 (N_17224,N_15993,N_13837);
and U17225 (N_17225,N_14339,N_12956);
and U17226 (N_17226,N_12359,N_14744);
xor U17227 (N_17227,N_14742,N_15767);
nand U17228 (N_17228,N_13171,N_14066);
nor U17229 (N_17229,N_13991,N_15204);
and U17230 (N_17230,N_15257,N_13583);
nand U17231 (N_17231,N_13992,N_14726);
and U17232 (N_17232,N_15933,N_15771);
and U17233 (N_17233,N_14394,N_13940);
and U17234 (N_17234,N_13579,N_12840);
nand U17235 (N_17235,N_12668,N_13474);
nand U17236 (N_17236,N_12619,N_14971);
nor U17237 (N_17237,N_13286,N_15463);
or U17238 (N_17238,N_13328,N_12000);
nor U17239 (N_17239,N_13313,N_14286);
nor U17240 (N_17240,N_14796,N_12502);
nor U17241 (N_17241,N_12582,N_13381);
and U17242 (N_17242,N_15577,N_12856);
xor U17243 (N_17243,N_15474,N_14891);
nor U17244 (N_17244,N_14901,N_14168);
and U17245 (N_17245,N_14563,N_14923);
nor U17246 (N_17246,N_14217,N_15817);
or U17247 (N_17247,N_15634,N_12095);
or U17248 (N_17248,N_12364,N_15207);
or U17249 (N_17249,N_14595,N_15812);
nor U17250 (N_17250,N_12723,N_13606);
xnor U17251 (N_17251,N_12052,N_15698);
nor U17252 (N_17252,N_13876,N_14408);
and U17253 (N_17253,N_13591,N_13499);
nand U17254 (N_17254,N_12704,N_15699);
or U17255 (N_17255,N_14068,N_14203);
or U17256 (N_17256,N_13585,N_13611);
nand U17257 (N_17257,N_12314,N_13988);
nor U17258 (N_17258,N_12294,N_12507);
xor U17259 (N_17259,N_14981,N_13810);
and U17260 (N_17260,N_15549,N_15490);
and U17261 (N_17261,N_14033,N_14419);
and U17262 (N_17262,N_13108,N_13253);
or U17263 (N_17263,N_14100,N_15339);
and U17264 (N_17264,N_15151,N_14032);
and U17265 (N_17265,N_13152,N_15741);
nand U17266 (N_17266,N_14661,N_13560);
nor U17267 (N_17267,N_13993,N_14878);
nor U17268 (N_17268,N_14231,N_14289);
nand U17269 (N_17269,N_13908,N_14520);
xnor U17270 (N_17270,N_15754,N_13745);
nand U17271 (N_17271,N_12044,N_15973);
xnor U17272 (N_17272,N_15417,N_15131);
nor U17273 (N_17273,N_15713,N_12259);
and U17274 (N_17274,N_13609,N_13603);
nor U17275 (N_17275,N_15049,N_14662);
or U17276 (N_17276,N_14057,N_13262);
and U17277 (N_17277,N_12929,N_13449);
nand U17278 (N_17278,N_15329,N_12495);
xnor U17279 (N_17279,N_15604,N_15440);
or U17280 (N_17280,N_14963,N_12919);
or U17281 (N_17281,N_13081,N_14673);
and U17282 (N_17282,N_12330,N_15094);
nand U17283 (N_17283,N_12589,N_15040);
and U17284 (N_17284,N_15846,N_12960);
xor U17285 (N_17285,N_13705,N_12570);
nand U17286 (N_17286,N_13149,N_12843);
and U17287 (N_17287,N_14763,N_12036);
or U17288 (N_17288,N_15349,N_15008);
xnor U17289 (N_17289,N_15671,N_12977);
or U17290 (N_17290,N_12740,N_15504);
or U17291 (N_17291,N_14336,N_14945);
nor U17292 (N_17292,N_13550,N_14807);
nand U17293 (N_17293,N_13100,N_12406);
nand U17294 (N_17294,N_12106,N_13437);
and U17295 (N_17295,N_12176,N_13167);
xor U17296 (N_17296,N_13644,N_12513);
nand U17297 (N_17297,N_12747,N_14070);
xnor U17298 (N_17298,N_13732,N_15987);
nor U17299 (N_17299,N_13492,N_13242);
nand U17300 (N_17300,N_15808,N_14470);
or U17301 (N_17301,N_13540,N_13769);
nor U17302 (N_17302,N_14047,N_15242);
nand U17303 (N_17303,N_13648,N_14828);
and U17304 (N_17304,N_12369,N_12807);
nor U17305 (N_17305,N_14691,N_12505);
nor U17306 (N_17306,N_13424,N_15179);
nor U17307 (N_17307,N_13766,N_14240);
xnor U17308 (N_17308,N_13930,N_14884);
nor U17309 (N_17309,N_15829,N_12292);
and U17310 (N_17310,N_12531,N_14205);
xor U17311 (N_17311,N_12417,N_13977);
or U17312 (N_17312,N_13243,N_14950);
nor U17313 (N_17313,N_14157,N_12738);
and U17314 (N_17314,N_13302,N_15834);
nand U17315 (N_17315,N_13023,N_15435);
xnor U17316 (N_17316,N_12288,N_14302);
nand U17317 (N_17317,N_14781,N_14895);
or U17318 (N_17318,N_12360,N_13417);
xor U17319 (N_17319,N_12425,N_12852);
or U17320 (N_17320,N_13180,N_14544);
nor U17321 (N_17321,N_14561,N_12604);
nand U17322 (N_17322,N_12801,N_12446);
and U17323 (N_17323,N_15075,N_12526);
nand U17324 (N_17324,N_14669,N_14758);
nand U17325 (N_17325,N_12988,N_13861);
nor U17326 (N_17326,N_15708,N_12849);
and U17327 (N_17327,N_15213,N_12958);
nand U17328 (N_17328,N_14566,N_15902);
nand U17329 (N_17329,N_15054,N_13462);
and U17330 (N_17330,N_14710,N_14770);
nor U17331 (N_17331,N_13056,N_15095);
nand U17332 (N_17332,N_13204,N_13316);
xor U17333 (N_17333,N_12551,N_14636);
nor U17334 (N_17334,N_12602,N_13273);
nand U17335 (N_17335,N_14139,N_15910);
and U17336 (N_17336,N_12219,N_13151);
nand U17337 (N_17337,N_14973,N_12666);
nor U17338 (N_17338,N_14188,N_15056);
xnor U17339 (N_17339,N_14220,N_12942);
nor U17340 (N_17340,N_12565,N_12711);
nand U17341 (N_17341,N_15181,N_13075);
nor U17342 (N_17342,N_13361,N_14620);
or U17343 (N_17343,N_12775,N_12499);
and U17344 (N_17344,N_12566,N_15472);
nor U17345 (N_17345,N_14006,N_12649);
nand U17346 (N_17346,N_14483,N_15516);
nand U17347 (N_17347,N_13572,N_14430);
or U17348 (N_17348,N_15782,N_13335);
and U17349 (N_17349,N_14187,N_15465);
and U17350 (N_17350,N_14889,N_14547);
nand U17351 (N_17351,N_13511,N_15066);
and U17352 (N_17352,N_15185,N_15691);
nor U17353 (N_17353,N_12235,N_13912);
nand U17354 (N_17354,N_15843,N_14400);
nand U17355 (N_17355,N_15077,N_15841);
nand U17356 (N_17356,N_13034,N_13480);
xor U17357 (N_17357,N_14014,N_15649);
nand U17358 (N_17358,N_15563,N_13803);
and U17359 (N_17359,N_13891,N_12734);
and U17360 (N_17360,N_13401,N_13781);
and U17361 (N_17361,N_12355,N_12157);
nor U17362 (N_17362,N_14291,N_14490);
nand U17363 (N_17363,N_15243,N_15338);
or U17364 (N_17364,N_13952,N_13211);
and U17365 (N_17365,N_15749,N_15854);
or U17366 (N_17366,N_15287,N_13584);
nor U17367 (N_17367,N_14667,N_15524);
nand U17368 (N_17368,N_12506,N_13442);
or U17369 (N_17369,N_15968,N_12687);
and U17370 (N_17370,N_12653,N_13812);
or U17371 (N_17371,N_13866,N_12043);
xor U17372 (N_17372,N_14466,N_13989);
nand U17373 (N_17373,N_12553,N_15291);
nand U17374 (N_17374,N_13217,N_12187);
and U17375 (N_17375,N_12851,N_14549);
nor U17376 (N_17376,N_12229,N_13205);
and U17377 (N_17377,N_14961,N_14349);
nand U17378 (N_17378,N_15794,N_12627);
or U17379 (N_17379,N_12564,N_14393);
nand U17380 (N_17380,N_15885,N_15471);
nor U17381 (N_17381,N_12534,N_14111);
and U17382 (N_17382,N_14760,N_13376);
or U17383 (N_17383,N_12059,N_12891);
nor U17384 (N_17384,N_12917,N_12256);
and U17385 (N_17385,N_15889,N_12599);
and U17386 (N_17386,N_12686,N_13868);
nor U17387 (N_17387,N_12107,N_14822);
nand U17388 (N_17388,N_13267,N_14864);
or U17389 (N_17389,N_14956,N_12615);
and U17390 (N_17390,N_13506,N_13843);
nor U17391 (N_17391,N_12399,N_14675);
and U17392 (N_17392,N_12213,N_12340);
nand U17393 (N_17393,N_13047,N_13103);
and U17394 (N_17394,N_13926,N_13129);
or U17395 (N_17395,N_15004,N_15249);
or U17396 (N_17396,N_13623,N_12875);
or U17397 (N_17397,N_13298,N_14186);
nand U17398 (N_17398,N_15168,N_14709);
xor U17399 (N_17399,N_13537,N_12338);
nand U17400 (N_17400,N_12185,N_13578);
nor U17401 (N_17401,N_15876,N_15299);
or U17402 (N_17402,N_15590,N_12372);
xnor U17403 (N_17403,N_15948,N_15692);
and U17404 (N_17404,N_14114,N_12853);
or U17405 (N_17405,N_14806,N_14137);
nand U17406 (N_17406,N_12715,N_15336);
nand U17407 (N_17407,N_13311,N_14898);
or U17408 (N_17408,N_12264,N_14761);
and U17409 (N_17409,N_14966,N_12969);
nand U17410 (N_17410,N_15784,N_15221);
nor U17411 (N_17411,N_14681,N_15128);
nor U17412 (N_17412,N_12435,N_13910);
and U17413 (N_17413,N_14016,N_14093);
or U17414 (N_17414,N_14991,N_14345);
nand U17415 (N_17415,N_13687,N_15053);
or U17416 (N_17416,N_13771,N_13657);
or U17417 (N_17417,N_14119,N_13338);
and U17418 (N_17418,N_15081,N_12820);
nor U17419 (N_17419,N_15046,N_12068);
nor U17420 (N_17420,N_14454,N_13351);
or U17421 (N_17421,N_14376,N_15414);
nand U17422 (N_17422,N_13975,N_12559);
xor U17423 (N_17423,N_13147,N_12521);
nand U17424 (N_17424,N_15099,N_12342);
or U17425 (N_17425,N_15576,N_12339);
nor U17426 (N_17426,N_12413,N_15688);
and U17427 (N_17427,N_14420,N_12786);
xnor U17428 (N_17428,N_14815,N_14712);
nor U17429 (N_17429,N_13676,N_15350);
nand U17430 (N_17430,N_14749,N_13713);
or U17431 (N_17431,N_12886,N_13347);
or U17432 (N_17432,N_14637,N_15648);
nand U17433 (N_17433,N_12165,N_14876);
and U17434 (N_17434,N_13412,N_15387);
nand U17435 (N_17435,N_12287,N_12025);
nor U17436 (N_17436,N_13605,N_15153);
nor U17437 (N_17437,N_15102,N_15120);
nand U17438 (N_17438,N_12242,N_14887);
nor U17439 (N_17439,N_13706,N_14804);
or U17440 (N_17440,N_14528,N_14558);
and U17441 (N_17441,N_12033,N_15833);
and U17442 (N_17442,N_14799,N_13637);
or U17443 (N_17443,N_12479,N_14655);
and U17444 (N_17444,N_13314,N_15300);
or U17445 (N_17445,N_13241,N_15222);
and U17446 (N_17446,N_14900,N_12374);
nand U17447 (N_17447,N_14109,N_15915);
nand U17448 (N_17448,N_15282,N_15256);
and U17449 (N_17449,N_14144,N_14363);
nand U17450 (N_17450,N_15909,N_13669);
and U17451 (N_17451,N_15742,N_15364);
or U17452 (N_17452,N_14810,N_15498);
nor U17453 (N_17453,N_13497,N_14741);
xnor U17454 (N_17454,N_12436,N_15999);
nor U17455 (N_17455,N_14651,N_14384);
and U17456 (N_17456,N_15476,N_13184);
nor U17457 (N_17457,N_12781,N_15455);
or U17458 (N_17458,N_12904,N_15518);
nand U17459 (N_17459,N_14812,N_15456);
nand U17460 (N_17460,N_13265,N_12906);
and U17461 (N_17461,N_13809,N_14618);
nor U17462 (N_17462,N_14358,N_15562);
nand U17463 (N_17463,N_13094,N_15899);
nand U17464 (N_17464,N_13163,N_13740);
or U17465 (N_17465,N_15991,N_15505);
nor U17466 (N_17466,N_13160,N_15626);
or U17467 (N_17467,N_14875,N_12400);
xor U17468 (N_17468,N_12026,N_12010);
or U17469 (N_17469,N_14206,N_15582);
and U17470 (N_17470,N_13130,N_14616);
xor U17471 (N_17471,N_15067,N_12529);
or U17472 (N_17472,N_14724,N_15599);
or U17473 (N_17473,N_15318,N_12596);
nor U17474 (N_17474,N_15951,N_14941);
or U17475 (N_17475,N_13451,N_14223);
and U17476 (N_17476,N_14185,N_13508);
or U17477 (N_17477,N_15085,N_12609);
xor U17478 (N_17478,N_12783,N_15665);
nor U17479 (N_17479,N_15217,N_15769);
or U17480 (N_17480,N_14317,N_12623);
nor U17481 (N_17481,N_14176,N_14184);
xnor U17482 (N_17482,N_15723,N_15330);
nor U17483 (N_17483,N_15357,N_12458);
or U17484 (N_17484,N_14869,N_13782);
xor U17485 (N_17485,N_13850,N_15333);
nor U17486 (N_17486,N_13348,N_13938);
nor U17487 (N_17487,N_12474,N_14784);
nor U17488 (N_17488,N_14275,N_12591);
or U17489 (N_17489,N_12273,N_15633);
nand U17490 (N_17490,N_12785,N_14797);
or U17491 (N_17491,N_13223,N_13256);
nand U17492 (N_17492,N_15042,N_15305);
xor U17493 (N_17493,N_14468,N_15827);
or U17494 (N_17494,N_12368,N_14234);
nand U17495 (N_17495,N_14350,N_13115);
nor U17496 (N_17496,N_15844,N_13546);
or U17497 (N_17497,N_15959,N_12787);
or U17498 (N_17498,N_14207,N_13869);
nand U17499 (N_17499,N_15738,N_14035);
nor U17500 (N_17500,N_14642,N_13752);
or U17501 (N_17501,N_15744,N_12430);
nand U17502 (N_17502,N_14850,N_12083);
nor U17503 (N_17503,N_15824,N_13673);
or U17504 (N_17504,N_12211,N_15320);
nand U17505 (N_17505,N_13086,N_13264);
or U17506 (N_17506,N_14603,N_14676);
or U17507 (N_17507,N_13909,N_12209);
nor U17508 (N_17508,N_12925,N_14952);
xnor U17509 (N_17509,N_15766,N_14059);
or U17510 (N_17510,N_14790,N_12195);
or U17511 (N_17511,N_14553,N_14838);
xor U17512 (N_17512,N_14428,N_14888);
xnor U17513 (N_17513,N_12440,N_12621);
and U17514 (N_17514,N_14354,N_14847);
xnor U17515 (N_17515,N_13092,N_14023);
nor U17516 (N_17516,N_12254,N_12861);
and U17517 (N_17517,N_14630,N_12828);
nand U17518 (N_17518,N_13450,N_13762);
or U17519 (N_17519,N_15816,N_13599);
or U17520 (N_17520,N_15309,N_13645);
nor U17521 (N_17521,N_15839,N_13491);
and U17522 (N_17522,N_13323,N_15223);
and U17523 (N_17523,N_13281,N_12733);
and U17524 (N_17524,N_15837,N_14862);
and U17525 (N_17525,N_13038,N_13186);
and U17526 (N_17526,N_15038,N_14461);
or U17527 (N_17527,N_15373,N_12984);
or U17528 (N_17528,N_15642,N_12158);
xor U17529 (N_17529,N_13616,N_13880);
nand U17530 (N_17530,N_14801,N_15654);
and U17531 (N_17531,N_13270,N_15327);
nor U17532 (N_17532,N_13041,N_14088);
and U17533 (N_17533,N_14510,N_15266);
or U17534 (N_17534,N_12391,N_13533);
nand U17535 (N_17535,N_12320,N_15481);
or U17536 (N_17536,N_14294,N_14043);
nand U17537 (N_17537,N_14580,N_12233);
nand U17538 (N_17538,N_15532,N_15380);
xor U17539 (N_17539,N_15934,N_14009);
and U17540 (N_17540,N_14500,N_13816);
xor U17541 (N_17541,N_14382,N_13672);
nor U17542 (N_17542,N_12739,N_14103);
or U17543 (N_17543,N_14074,N_15070);
or U17544 (N_17544,N_12806,N_15253);
nor U17545 (N_17545,N_14905,N_15422);
nor U17546 (N_17546,N_14474,N_13953);
nand U17547 (N_17547,N_14550,N_15690);
and U17548 (N_17548,N_12544,N_13806);
nor U17549 (N_17549,N_15169,N_13247);
xnor U17550 (N_17550,N_15170,N_15850);
and U17551 (N_17551,N_15164,N_12778);
nor U17552 (N_17552,N_15820,N_13475);
or U17553 (N_17553,N_14843,N_14915);
or U17554 (N_17554,N_14196,N_15706);
and U17555 (N_17555,N_14334,N_14000);
and U17556 (N_17556,N_13884,N_12124);
and U17557 (N_17557,N_13982,N_15121);
and U17558 (N_17558,N_15480,N_15866);
xnor U17559 (N_17559,N_14310,N_13902);
and U17560 (N_17560,N_15497,N_13937);
and U17561 (N_17561,N_12637,N_15379);
or U17562 (N_17562,N_13688,N_12398);
nand U17563 (N_17563,N_14368,N_12432);
and U17564 (N_17564,N_13619,N_13164);
and U17565 (N_17565,N_12815,N_14700);
and U17566 (N_17566,N_12726,N_14577);
nand U17567 (N_17567,N_12367,N_14417);
or U17568 (N_17568,N_13906,N_13189);
nand U17569 (N_17569,N_15037,N_12788);
or U17570 (N_17570,N_14458,N_15972);
xnor U17571 (N_17571,N_15931,N_14851);
nor U17572 (N_17572,N_15017,N_13778);
nand U17573 (N_17573,N_15684,N_14705);
xnor U17574 (N_17574,N_15949,N_15147);
nor U17575 (N_17575,N_12291,N_13575);
or U17576 (N_17576,N_12607,N_14069);
nor U17577 (N_17577,N_14161,N_12973);
and U17578 (N_17578,N_12380,N_15292);
xor U17579 (N_17579,N_13854,N_12546);
and U17580 (N_17580,N_13873,N_14080);
or U17581 (N_17581,N_15880,N_14031);
and U17582 (N_17582,N_14494,N_13169);
nand U17583 (N_17583,N_14598,N_13758);
or U17584 (N_17584,N_15483,N_13154);
and U17585 (N_17585,N_12857,N_12401);
or U17586 (N_17586,N_14353,N_15342);
nor U17587 (N_17587,N_12439,N_14488);
nand U17588 (N_17588,N_14181,N_13037);
nor U17589 (N_17589,N_12648,N_12811);
and U17590 (N_17590,N_12643,N_14649);
xor U17591 (N_17591,N_14910,N_15210);
nand U17592 (N_17592,N_13720,N_13699);
nor U17593 (N_17593,N_13292,N_15353);
or U17594 (N_17594,N_13471,N_14460);
and U17595 (N_17595,N_13568,N_12867);
and U17596 (N_17596,N_14215,N_12943);
or U17597 (N_17597,N_15064,N_12547);
and U17598 (N_17598,N_12821,N_12119);
nor U17599 (N_17599,N_13305,N_15862);
nor U17600 (N_17600,N_14411,N_15002);
xnor U17601 (N_17601,N_14254,N_13087);
or U17602 (N_17602,N_14390,N_14274);
or U17603 (N_17603,N_15307,N_12688);
or U17604 (N_17604,N_13703,N_14648);
nand U17605 (N_17605,N_13456,N_15637);
nor U17606 (N_17606,N_14684,N_14756);
or U17607 (N_17607,N_14707,N_14022);
and U17608 (N_17608,N_14755,N_15996);
xor U17609 (N_17609,N_13958,N_14180);
or U17610 (N_17610,N_14424,N_12721);
nor U17611 (N_17611,N_13858,N_12965);
nor U17612 (N_17612,N_13824,N_14166);
or U17613 (N_17613,N_13878,N_13059);
or U17614 (N_17614,N_14030,N_13786);
nor U17615 (N_17615,N_15609,N_14204);
nor U17616 (N_17616,N_13650,N_13554);
and U17617 (N_17617,N_13248,N_15830);
xnor U17618 (N_17618,N_15905,N_12186);
nor U17619 (N_17619,N_12051,N_13913);
and U17620 (N_17620,N_12118,N_14560);
xor U17621 (N_17621,N_13541,N_14051);
and U17622 (N_17622,N_13443,N_12129);
and U17623 (N_17623,N_12076,N_12543);
nor U17624 (N_17624,N_15428,N_15955);
nand U17625 (N_17625,N_15828,N_12756);
nor U17626 (N_17626,N_14732,N_14833);
or U17627 (N_17627,N_13759,N_13246);
and U17628 (N_17628,N_12664,N_13018);
and U17629 (N_17629,N_14377,N_15269);
nand U17630 (N_17630,N_14416,N_12376);
nor U17631 (N_17631,N_14421,N_14576);
nand U17632 (N_17632,N_15686,N_13463);
nor U17633 (N_17633,N_13307,N_15178);
nand U17634 (N_17634,N_15608,N_15542);
or U17635 (N_17635,N_15460,N_13067);
or U17636 (N_17636,N_15751,N_12710);
nand U17637 (N_17637,N_13588,N_15434);
xor U17638 (N_17638,N_12414,N_15458);
and U17639 (N_17639,N_12097,N_15432);
xor U17640 (N_17640,N_15192,N_14256);
or U17641 (N_17641,N_15977,N_15363);
nor U17642 (N_17642,N_13221,N_15776);
and U17643 (N_17643,N_12410,N_13040);
nor U17644 (N_17644,N_14471,N_14472);
nand U17645 (N_17645,N_15345,N_13337);
or U17646 (N_17646,N_15438,N_13728);
nand U17647 (N_17647,N_13555,N_15412);
or U17648 (N_17648,N_14545,N_12628);
xor U17649 (N_17649,N_15783,N_12662);
and U17650 (N_17650,N_14283,N_15904);
or U17651 (N_17651,N_15142,N_14879);
nand U17652 (N_17652,N_13477,N_13515);
nor U17653 (N_17653,N_14475,N_15980);
or U17654 (N_17654,N_15734,N_14440);
nand U17655 (N_17655,N_12140,N_13570);
or U17656 (N_17656,N_15685,N_12892);
or U17657 (N_17657,N_15343,N_13460);
nand U17658 (N_17658,N_15722,N_12356);
and U17659 (N_17659,N_15917,N_15089);
or U17660 (N_17660,N_12150,N_12285);
and U17661 (N_17661,N_13357,N_13883);
nand U17662 (N_17662,N_13859,N_14003);
and U17663 (N_17663,N_14053,N_13033);
nand U17664 (N_17664,N_14285,N_14632);
nand U17665 (N_17665,N_13269,N_13421);
nor U17666 (N_17666,N_13580,N_12089);
and U17667 (N_17667,N_12574,N_15421);
nor U17668 (N_17668,N_13279,N_15535);
and U17669 (N_17669,N_15919,N_12695);
and U17670 (N_17670,N_14506,N_15589);
nor U17671 (N_17671,N_14438,N_14153);
and U17672 (N_17672,N_12310,N_13233);
nor U17673 (N_17673,N_12493,N_13297);
nor U17674 (N_17674,N_12616,N_14572);
nor U17675 (N_17675,N_12508,N_14902);
nand U17676 (N_17676,N_14333,N_14101);
or U17677 (N_17677,N_12269,N_14652);
nand U17678 (N_17678,N_13795,N_15057);
or U17679 (N_17679,N_12012,N_14455);
and U17680 (N_17680,N_14098,N_12421);
nor U17681 (N_17681,N_14076,N_13618);
nor U17682 (N_17682,N_12429,N_14445);
nand U17683 (N_17683,N_14054,N_15215);
xnor U17684 (N_17684,N_15859,N_15316);
and U17685 (N_17685,N_12236,N_12608);
nand U17686 (N_17686,N_13364,N_12803);
and U17687 (N_17687,N_12065,N_13963);
or U17688 (N_17688,N_13342,N_15324);
nor U17689 (N_17689,N_14117,N_12754);
and U17690 (N_17690,N_14928,N_14437);
nand U17691 (N_17691,N_15595,N_14146);
and U17692 (N_17692,N_15868,N_12397);
and U17693 (N_17693,N_13028,N_12639);
nor U17694 (N_17694,N_13530,N_12569);
or U17695 (N_17695,N_15231,N_15845);
nor U17696 (N_17696,N_12937,N_15550);
and U17697 (N_17697,N_15273,N_15251);
or U17698 (N_17698,N_12312,N_12995);
and U17699 (N_17699,N_15520,N_14061);
and U17700 (N_17700,N_13176,N_14102);
or U17701 (N_17701,N_13787,N_15376);
and U17702 (N_17702,N_15770,N_12154);
and U17703 (N_17703,N_15003,N_12027);
and U17704 (N_17704,N_12614,N_12116);
and U17705 (N_17705,N_14253,N_15447);
or U17706 (N_17706,N_13017,N_14304);
nor U17707 (N_17707,N_12260,N_14154);
and U17708 (N_17708,N_12769,N_13465);
nand U17709 (N_17709,N_15464,N_15811);
nand U17710 (N_17710,N_14301,N_14837);
nand U17711 (N_17711,N_13561,N_12266);
nand U17712 (N_17712,N_15818,N_13402);
or U17713 (N_17713,N_12073,N_12611);
nand U17714 (N_17714,N_14112,N_13519);
and U17715 (N_17715,N_14163,N_13526);
xor U17716 (N_17716,N_14533,N_15819);
nand U17717 (N_17717,N_13943,N_13852);
nand U17718 (N_17718,N_14646,N_15029);
and U17719 (N_17719,N_15785,N_12478);
nand U17720 (N_17720,N_15270,N_15413);
nor U17721 (N_17721,N_13000,N_13482);
and U17722 (N_17722,N_13016,N_12883);
nand U17723 (N_17723,N_12272,N_12578);
or U17724 (N_17724,N_12835,N_12877);
and U17725 (N_17725,N_12481,N_13756);
nand U17726 (N_17726,N_13945,N_12453);
nand U17727 (N_17727,N_15747,N_13088);
nor U17728 (N_17728,N_15901,N_14175);
nor U17729 (N_17729,N_13310,N_13914);
and U17730 (N_17730,N_15988,N_15552);
and U17731 (N_17731,N_12225,N_15611);
or U17732 (N_17732,N_15743,N_15293);
nand U17733 (N_17733,N_15172,N_15548);
nand U17734 (N_17734,N_15426,N_15135);
and U17735 (N_17735,N_13614,N_13193);
nand U17736 (N_17736,N_15405,N_15475);
or U17737 (N_17737,N_12728,N_14388);
and U17738 (N_17738,N_12814,N_12618);
nand U17739 (N_17739,N_12872,N_14946);
or U17740 (N_17740,N_14588,N_14151);
and U17741 (N_17741,N_12323,N_14432);
nand U17742 (N_17742,N_12598,N_12375);
nor U17743 (N_17743,N_14670,N_12652);
nor U17744 (N_17744,N_12423,N_12456);
nor U17745 (N_17745,N_14788,N_15924);
and U17746 (N_17746,N_14143,N_14318);
nor U17747 (N_17747,N_12514,N_15646);
and U17748 (N_17748,N_15517,N_14306);
nand U17749 (N_17749,N_15348,N_13106);
xnor U17750 (N_17750,N_12532,N_13453);
nand U17751 (N_17751,N_14765,N_12457);
nand U17752 (N_17752,N_13009,N_13822);
xor U17753 (N_17753,N_14084,N_14268);
or U17754 (N_17754,N_13929,N_15572);
and U17755 (N_17755,N_13896,N_13329);
and U17756 (N_17756,N_14312,N_12063);
or U17757 (N_17757,N_15773,N_12730);
nor U17758 (N_17758,N_12300,N_15437);
xnor U17759 (N_17759,N_13464,N_14079);
xnor U17760 (N_17760,N_13399,N_12093);
xor U17761 (N_17761,N_14772,N_14841);
or U17762 (N_17762,N_13966,N_12395);
and U17763 (N_17763,N_15892,N_13232);
and U17764 (N_17764,N_12590,N_14017);
nor U17765 (N_17765,N_13146,N_15950);
or U17766 (N_17766,N_13946,N_13750);
and U17767 (N_17767,N_13643,N_13636);
nand U17768 (N_17768,N_14980,N_15556);
or U17769 (N_17769,N_12136,N_12890);
nor U17770 (N_17770,N_13959,N_13276);
and U17771 (N_17771,N_14379,N_12050);
nand U17772 (N_17772,N_14525,N_14540);
nand U17773 (N_17773,N_15086,N_13986);
nand U17774 (N_17774,N_13340,N_13680);
nor U17775 (N_17775,N_12755,N_14692);
nor U17776 (N_17776,N_14208,N_13571);
and U17777 (N_17777,N_13640,N_14495);
xnor U17778 (N_17778,N_12324,N_12822);
nand U17779 (N_17779,N_13212,N_14814);
or U17780 (N_17780,N_13104,N_14075);
nand U17781 (N_17781,N_12210,N_14356);
nand U17782 (N_17782,N_12471,N_13032);
or U17783 (N_17783,N_13496,N_14587);
nor U17784 (N_17784,N_14582,N_12181);
nand U17785 (N_17785,N_14211,N_13386);
and U17786 (N_17786,N_12510,N_12201);
or U17787 (N_17787,N_13008,N_12321);
nand U17788 (N_17788,N_13260,N_13372);
xnor U17789 (N_17789,N_12208,N_12882);
nor U17790 (N_17790,N_15132,N_14821);
nor U17791 (N_17791,N_12503,N_15052);
nor U17792 (N_17792,N_12084,N_12267);
or U17793 (N_17793,N_15454,N_14552);
nor U17794 (N_17794,N_12409,N_13895);
or U17795 (N_17795,N_14099,N_14727);
or U17796 (N_17796,N_12763,N_13411);
or U17797 (N_17797,N_13630,N_15596);
nor U17798 (N_17798,N_12227,N_13095);
nand U17799 (N_17799,N_13410,N_14115);
nand U17800 (N_17800,N_12741,N_15205);
or U17801 (N_17801,N_14625,N_12535);
nor U17802 (N_17802,N_12865,N_14522);
nor U17803 (N_17803,N_12974,N_12971);
and U17804 (N_17804,N_15886,N_13821);
and U17805 (N_17805,N_13052,N_13567);
xnor U17806 (N_17806,N_12980,N_15786);
nor U17807 (N_17807,N_12750,N_12924);
nor U17808 (N_17808,N_13857,N_15175);
nor U17809 (N_17809,N_15806,N_13046);
or U17810 (N_17810,N_13117,N_13505);
or U17811 (N_17811,N_14951,N_14711);
xor U17812 (N_17812,N_15639,N_13422);
nand U17813 (N_17813,N_12992,N_13263);
nand U17814 (N_17814,N_12991,N_14730);
and U17815 (N_17815,N_12893,N_12194);
or U17816 (N_17816,N_14357,N_13874);
or U17817 (N_17817,N_14856,N_15445);
nand U17818 (N_17818,N_14608,N_14366);
and U17819 (N_17819,N_12701,N_15127);
and U17820 (N_17820,N_15998,N_13941);
and U17821 (N_17821,N_14863,N_12092);
nor U17822 (N_17822,N_13143,N_15184);
xnor U17823 (N_17823,N_14235,N_15956);
nor U17824 (N_17824,N_12862,N_12498);
nor U17825 (N_17825,N_13071,N_12004);
or U17826 (N_17826,N_13548,N_13228);
nor U17827 (N_17827,N_15714,N_13142);
nand U17828 (N_17828,N_12802,N_14924);
nand U17829 (N_17829,N_15515,N_13886);
nor U17830 (N_17830,N_13441,N_12133);
or U17831 (N_17831,N_14429,N_13736);
nor U17832 (N_17832,N_13718,N_13685);
nor U17833 (N_17833,N_15825,N_12402);
or U17834 (N_17834,N_15459,N_12058);
or U17835 (N_17835,N_12790,N_15813);
xnor U17836 (N_17836,N_15503,N_15613);
or U17837 (N_17837,N_12070,N_13825);
nand U17838 (N_17838,N_15019,N_12352);
and U17839 (N_17839,N_14696,N_14303);
nor U17840 (N_17840,N_15220,N_15702);
nand U17841 (N_17841,N_14957,N_12827);
or U17842 (N_17842,N_13440,N_13188);
or U17843 (N_17843,N_15051,N_13697);
nor U17844 (N_17844,N_12736,N_14607);
or U17845 (N_17845,N_13127,N_13173);
nor U17846 (N_17846,N_14230,N_14089);
nor U17847 (N_17847,N_15279,N_14654);
nand U17848 (N_17848,N_13961,N_12913);
and U17849 (N_17849,N_15224,N_13999);
xnor U17850 (N_17850,N_14434,N_12200);
nor U17851 (N_17851,N_12798,N_14073);
or U17852 (N_17852,N_13751,N_13299);
nand U17853 (N_17853,N_15677,N_15879);
or U17854 (N_17854,N_12921,N_15022);
or U17855 (N_17855,N_13833,N_13370);
nand U17856 (N_17856,N_12981,N_15614);
and U17857 (N_17857,N_14140,N_13452);
and U17858 (N_17858,N_14225,N_13701);
and U17859 (N_17859,N_12381,N_15787);
and U17860 (N_17860,N_13846,N_12635);
and U17861 (N_17861,N_15113,N_13371);
and U17862 (N_17862,N_13069,N_14122);
or U17863 (N_17863,N_12335,N_12220);
or U17864 (N_17864,N_13783,N_13516);
nand U17865 (N_17865,N_15001,N_13430);
nand U17866 (N_17866,N_12159,N_13935);
and U17867 (N_17867,N_12005,N_12762);
or U17868 (N_17868,N_15174,N_15627);
nand U17869 (N_17869,N_12660,N_13050);
xor U17870 (N_17870,N_13504,N_13495);
nand U17871 (N_17871,N_13726,N_13135);
nand U17872 (N_17872,N_15929,N_14464);
and U17873 (N_17873,N_13296,N_12813);
or U17874 (N_17874,N_12426,N_12126);
and U17875 (N_17875,N_14672,N_14459);
and U17876 (N_17876,N_13544,N_15219);
nand U17877 (N_17877,N_14854,N_12138);
nor U17878 (N_17878,N_12365,N_14564);
nor U17879 (N_17879,N_14072,N_14364);
nand U17880 (N_17880,N_13996,N_12144);
nor U17881 (N_17881,N_14443,N_12362);
nor U17882 (N_17882,N_15370,N_14737);
nor U17883 (N_17883,N_15354,N_13166);
nor U17884 (N_17884,N_14635,N_13997);
nand U17885 (N_17885,N_13532,N_12699);
nor U17886 (N_17886,N_13091,N_14218);
and U17887 (N_17887,N_12289,N_15492);
nor U17888 (N_17888,N_13631,N_14740);
nand U17889 (N_17889,N_12563,N_13845);
nor U17890 (N_17890,N_14012,N_13192);
or U17891 (N_17891,N_15167,N_14774);
nor U17892 (N_17892,N_13222,N_14631);
or U17893 (N_17893,N_14768,N_14028);
nand U17894 (N_17894,N_12622,N_15260);
and U17895 (N_17895,N_15321,N_13133);
and U17896 (N_17896,N_15467,N_13230);
nand U17897 (N_17897,N_12162,N_15921);
nor U17898 (N_17898,N_12480,N_13820);
or U17899 (N_17899,N_15315,N_14386);
nand U17900 (N_17900,N_14314,N_12100);
nand U17901 (N_17901,N_12228,N_12669);
or U17902 (N_17902,N_12860,N_15855);
and U17903 (N_17903,N_15553,N_15778);
and U17904 (N_17904,N_13638,N_13257);
and U17905 (N_17905,N_12915,N_14925);
xor U17906 (N_17906,N_14323,N_13715);
or U17907 (N_17907,N_15104,N_15823);
nor U17908 (N_17908,N_15867,N_12001);
nand U17909 (N_17909,N_13844,N_12537);
and U17910 (N_17910,N_13255,N_13054);
xor U17911 (N_17911,N_13210,N_13068);
and U17912 (N_17912,N_13057,N_14502);
nor U17913 (N_17913,N_15087,N_13665);
or U17914 (N_17914,N_14405,N_12888);
xor U17915 (N_17915,N_15849,N_12454);
and U17916 (N_17916,N_13031,N_14489);
nor U17917 (N_17917,N_15887,N_12483);
xor U17918 (N_17918,N_12791,N_15815);
nand U17919 (N_17919,N_14894,N_13468);
nand U17920 (N_17920,N_13746,N_14848);
nor U17921 (N_17921,N_14381,N_14795);
nor U17922 (N_17922,N_14348,N_12760);
or U17923 (N_17923,N_14565,N_15512);
and U17924 (N_17924,N_15568,N_14029);
or U17925 (N_17925,N_14481,N_15212);
and U17926 (N_17926,N_15058,N_12538);
and U17927 (N_17927,N_14258,N_12823);
or U17928 (N_17928,N_14228,N_12858);
and U17929 (N_17929,N_13317,N_13860);
and U17930 (N_17930,N_12540,N_15235);
and U17931 (N_17931,N_13478,N_15171);
nand U17932 (N_17932,N_13284,N_14666);
nor U17933 (N_17933,N_14933,N_12601);
nand U17934 (N_17934,N_14773,N_15139);
and U17935 (N_17935,N_15203,N_14640);
nand U17936 (N_17936,N_14594,N_14501);
nand U17937 (N_17937,N_15163,N_14392);
and U17938 (N_17938,N_14918,N_12727);
or U17939 (N_17939,N_15522,N_15546);
nand U17940 (N_17940,N_14338,N_14805);
or U17941 (N_17941,N_15936,N_14896);
nor U17942 (N_17942,N_14373,N_13369);
and U17943 (N_17943,N_15705,N_15265);
and U17944 (N_17944,N_15525,N_15485);
xor U17945 (N_17945,N_13177,N_13968);
and U17946 (N_17946,N_12270,N_14659);
or U17947 (N_17947,N_15006,N_15531);
and U17948 (N_17948,N_15750,N_13520);
or U17949 (N_17949,N_13065,N_12218);
or U17950 (N_17950,N_13922,N_13250);
or U17951 (N_17951,N_13035,N_14262);
and U17952 (N_17952,N_13983,N_12434);
and U17953 (N_17953,N_14600,N_15547);
or U17954 (N_17954,N_13915,N_13798);
or U17955 (N_17955,N_14212,N_14239);
and U17956 (N_17956,N_14480,N_13219);
nand U17957 (N_17957,N_15011,N_14571);
nand U17958 (N_17958,N_13923,N_13960);
nand U17959 (N_17959,N_13112,N_15561);
xnor U17960 (N_17960,N_12132,N_12174);
and U17961 (N_17961,N_12282,N_13536);
nor U17962 (N_17962,N_13831,N_13814);
and U17963 (N_17963,N_15780,N_13556);
and U17964 (N_17964,N_13156,N_15297);
and U17965 (N_17965,N_14320,N_13553);
nand U17966 (N_17966,N_15450,N_13921);
nand U17967 (N_17967,N_15569,N_12847);
or U17968 (N_17968,N_15402,N_12720);
xnor U17969 (N_17969,N_14865,N_12955);
nor U17970 (N_17970,N_13918,N_14908);
nor U17971 (N_17971,N_12099,N_13428);
nor U17972 (N_17972,N_12328,N_15229);
nor U17973 (N_17973,N_14264,N_14567);
and U17974 (N_17974,N_14158,N_15733);
xnor U17975 (N_17975,N_15118,N_15756);
nor U17976 (N_17976,N_12147,N_13240);
and U17977 (N_17977,N_12518,N_13595);
nand U17978 (N_17978,N_12634,N_13326);
nand U17979 (N_17979,N_13954,N_14976);
nor U17980 (N_17980,N_12341,N_12515);
and U17981 (N_17981,N_15591,N_12889);
nor U17982 (N_17982,N_15583,N_15484);
nand U17983 (N_17983,N_15083,N_13377);
or U17984 (N_17984,N_15718,N_15240);
nor U17985 (N_17985,N_13835,N_15383);
nand U17986 (N_17986,N_14621,N_15856);
nand U17987 (N_17987,N_13435,N_12670);
nand U17988 (N_17988,N_15675,N_15024);
or U17989 (N_17989,N_15908,N_15473);
xnor U17990 (N_17990,N_15031,N_15963);
nand U17991 (N_17991,N_14777,N_14535);
nor U17992 (N_17992,N_12252,N_12625);
nor U17993 (N_17993,N_12163,N_15527);
nor U17994 (N_17994,N_15764,N_14315);
nor U17995 (N_17995,N_12963,N_13487);
nand U17996 (N_17996,N_12114,N_15444);
nand U17997 (N_17997,N_14113,N_12993);
xnor U17998 (N_17998,N_14932,N_15961);
nor U17999 (N_17999,N_13700,N_13098);
nand U18000 (N_18000,N_12329,N_14022);
and U18001 (N_18001,N_12911,N_12528);
nand U18002 (N_18002,N_14217,N_15300);
or U18003 (N_18003,N_15040,N_12283);
and U18004 (N_18004,N_13806,N_13001);
nand U18005 (N_18005,N_13155,N_13270);
and U18006 (N_18006,N_15025,N_13257);
xnor U18007 (N_18007,N_13419,N_12320);
and U18008 (N_18008,N_14911,N_12668);
and U18009 (N_18009,N_15321,N_15564);
or U18010 (N_18010,N_13831,N_12221);
or U18011 (N_18011,N_12094,N_13880);
nor U18012 (N_18012,N_15698,N_14619);
nand U18013 (N_18013,N_15117,N_15734);
nor U18014 (N_18014,N_12496,N_12728);
and U18015 (N_18015,N_12806,N_12395);
nor U18016 (N_18016,N_15587,N_14086);
and U18017 (N_18017,N_15928,N_14931);
or U18018 (N_18018,N_14643,N_14080);
nand U18019 (N_18019,N_13611,N_12652);
nor U18020 (N_18020,N_13083,N_15737);
and U18021 (N_18021,N_14866,N_13665);
and U18022 (N_18022,N_12841,N_15295);
and U18023 (N_18023,N_12275,N_12834);
xnor U18024 (N_18024,N_14456,N_12764);
and U18025 (N_18025,N_15220,N_14017);
and U18026 (N_18026,N_14860,N_13604);
xnor U18027 (N_18027,N_15802,N_12728);
nand U18028 (N_18028,N_14767,N_15429);
nand U18029 (N_18029,N_12400,N_15187);
or U18030 (N_18030,N_12642,N_12269);
nor U18031 (N_18031,N_13423,N_14144);
nand U18032 (N_18032,N_12471,N_14009);
nor U18033 (N_18033,N_14197,N_14995);
and U18034 (N_18034,N_12827,N_15078);
nand U18035 (N_18035,N_14211,N_14677);
or U18036 (N_18036,N_15005,N_12660);
or U18037 (N_18037,N_12100,N_13629);
nor U18038 (N_18038,N_12258,N_13857);
xor U18039 (N_18039,N_14681,N_15527);
nand U18040 (N_18040,N_13395,N_14768);
nor U18041 (N_18041,N_12074,N_13300);
and U18042 (N_18042,N_13163,N_12603);
nor U18043 (N_18043,N_14887,N_15874);
nor U18044 (N_18044,N_13876,N_15715);
nand U18045 (N_18045,N_14087,N_15104);
and U18046 (N_18046,N_12190,N_15705);
nor U18047 (N_18047,N_14064,N_14097);
or U18048 (N_18048,N_12972,N_15491);
nand U18049 (N_18049,N_14373,N_12140);
nand U18050 (N_18050,N_15911,N_12186);
and U18051 (N_18051,N_13847,N_14090);
and U18052 (N_18052,N_14570,N_12281);
or U18053 (N_18053,N_14030,N_13469);
or U18054 (N_18054,N_15782,N_12069);
nand U18055 (N_18055,N_13384,N_13453);
or U18056 (N_18056,N_15089,N_12566);
nand U18057 (N_18057,N_12082,N_15771);
or U18058 (N_18058,N_15659,N_13789);
nand U18059 (N_18059,N_15794,N_15947);
nand U18060 (N_18060,N_15560,N_15455);
nor U18061 (N_18061,N_12567,N_14227);
and U18062 (N_18062,N_12864,N_14803);
nand U18063 (N_18063,N_14278,N_13296);
nor U18064 (N_18064,N_13286,N_12438);
nor U18065 (N_18065,N_12123,N_15887);
nand U18066 (N_18066,N_13422,N_15421);
nand U18067 (N_18067,N_12045,N_14250);
and U18068 (N_18068,N_12418,N_14320);
or U18069 (N_18069,N_13060,N_13586);
nand U18070 (N_18070,N_15692,N_15214);
and U18071 (N_18071,N_14034,N_15023);
and U18072 (N_18072,N_15309,N_12108);
and U18073 (N_18073,N_14545,N_13525);
nand U18074 (N_18074,N_15267,N_14962);
and U18075 (N_18075,N_14056,N_14920);
nor U18076 (N_18076,N_13702,N_14941);
nand U18077 (N_18077,N_13363,N_14574);
nor U18078 (N_18078,N_12851,N_14050);
nand U18079 (N_18079,N_13621,N_13204);
nand U18080 (N_18080,N_12925,N_14380);
and U18081 (N_18081,N_15695,N_14161);
nand U18082 (N_18082,N_13019,N_14162);
nand U18083 (N_18083,N_13960,N_15333);
nand U18084 (N_18084,N_13455,N_15398);
and U18085 (N_18085,N_15558,N_12975);
or U18086 (N_18086,N_13822,N_14119);
or U18087 (N_18087,N_12199,N_15278);
or U18088 (N_18088,N_13453,N_13718);
or U18089 (N_18089,N_14859,N_15549);
xor U18090 (N_18090,N_12404,N_13072);
nor U18091 (N_18091,N_12673,N_13160);
or U18092 (N_18092,N_13683,N_12886);
nor U18093 (N_18093,N_12103,N_14033);
or U18094 (N_18094,N_13757,N_14141);
xnor U18095 (N_18095,N_13604,N_14490);
nand U18096 (N_18096,N_15620,N_15562);
nor U18097 (N_18097,N_15988,N_13491);
nor U18098 (N_18098,N_12596,N_12427);
or U18099 (N_18099,N_15215,N_15525);
and U18100 (N_18100,N_15970,N_15160);
and U18101 (N_18101,N_13588,N_12981);
or U18102 (N_18102,N_12135,N_12031);
nand U18103 (N_18103,N_14166,N_13729);
xnor U18104 (N_18104,N_15711,N_13628);
nor U18105 (N_18105,N_15743,N_14249);
xor U18106 (N_18106,N_15342,N_15431);
and U18107 (N_18107,N_15870,N_13517);
nor U18108 (N_18108,N_13412,N_13265);
nand U18109 (N_18109,N_14462,N_12585);
nand U18110 (N_18110,N_14628,N_15125);
or U18111 (N_18111,N_15623,N_12962);
or U18112 (N_18112,N_15187,N_15933);
nand U18113 (N_18113,N_15169,N_12293);
or U18114 (N_18114,N_14817,N_13696);
and U18115 (N_18115,N_14811,N_14095);
or U18116 (N_18116,N_13532,N_13936);
and U18117 (N_18117,N_12669,N_12899);
and U18118 (N_18118,N_13894,N_14151);
xnor U18119 (N_18119,N_12943,N_14147);
xnor U18120 (N_18120,N_13873,N_12840);
nand U18121 (N_18121,N_15101,N_13713);
nor U18122 (N_18122,N_12099,N_13773);
nand U18123 (N_18123,N_13473,N_12692);
nand U18124 (N_18124,N_12785,N_12436);
nand U18125 (N_18125,N_14619,N_14197);
nand U18126 (N_18126,N_12160,N_15596);
nand U18127 (N_18127,N_13508,N_12878);
and U18128 (N_18128,N_15525,N_15908);
nand U18129 (N_18129,N_15715,N_15149);
xnor U18130 (N_18130,N_12505,N_12049);
nand U18131 (N_18131,N_15721,N_14094);
or U18132 (N_18132,N_14435,N_13666);
nor U18133 (N_18133,N_13032,N_14455);
nor U18134 (N_18134,N_13669,N_13688);
or U18135 (N_18135,N_14799,N_14676);
and U18136 (N_18136,N_15105,N_13706);
nor U18137 (N_18137,N_13651,N_14655);
and U18138 (N_18138,N_15705,N_15177);
and U18139 (N_18139,N_12209,N_13755);
nand U18140 (N_18140,N_15776,N_15315);
nand U18141 (N_18141,N_14583,N_12051);
nand U18142 (N_18142,N_14236,N_13490);
nand U18143 (N_18143,N_12547,N_15107);
nand U18144 (N_18144,N_14304,N_15878);
nand U18145 (N_18145,N_13364,N_13998);
and U18146 (N_18146,N_13216,N_12385);
nand U18147 (N_18147,N_13219,N_15740);
nand U18148 (N_18148,N_13322,N_15251);
nor U18149 (N_18149,N_13126,N_14149);
xor U18150 (N_18150,N_13131,N_14580);
or U18151 (N_18151,N_15264,N_14858);
and U18152 (N_18152,N_12492,N_13521);
and U18153 (N_18153,N_15173,N_15201);
nor U18154 (N_18154,N_14751,N_14142);
and U18155 (N_18155,N_15457,N_13250);
xnor U18156 (N_18156,N_14821,N_12388);
xnor U18157 (N_18157,N_12617,N_13653);
or U18158 (N_18158,N_13388,N_13096);
and U18159 (N_18159,N_12935,N_12278);
xnor U18160 (N_18160,N_14812,N_13170);
xnor U18161 (N_18161,N_14206,N_12566);
or U18162 (N_18162,N_13530,N_12125);
xor U18163 (N_18163,N_12171,N_12923);
nor U18164 (N_18164,N_15984,N_12588);
nand U18165 (N_18165,N_13195,N_13308);
nor U18166 (N_18166,N_12493,N_13381);
or U18167 (N_18167,N_15659,N_13634);
xnor U18168 (N_18168,N_13112,N_15583);
xnor U18169 (N_18169,N_14385,N_12396);
or U18170 (N_18170,N_12200,N_13215);
nor U18171 (N_18171,N_13991,N_13067);
xnor U18172 (N_18172,N_14683,N_12055);
and U18173 (N_18173,N_15310,N_14522);
nand U18174 (N_18174,N_13895,N_14692);
and U18175 (N_18175,N_12387,N_12435);
or U18176 (N_18176,N_13756,N_14091);
or U18177 (N_18177,N_15536,N_15262);
and U18178 (N_18178,N_12721,N_15520);
nand U18179 (N_18179,N_15197,N_15380);
or U18180 (N_18180,N_15458,N_14966);
and U18181 (N_18181,N_13293,N_13736);
nor U18182 (N_18182,N_13928,N_15873);
or U18183 (N_18183,N_13477,N_15833);
or U18184 (N_18184,N_12375,N_15610);
nand U18185 (N_18185,N_15709,N_14776);
nand U18186 (N_18186,N_12793,N_15714);
and U18187 (N_18187,N_12979,N_14364);
nor U18188 (N_18188,N_12963,N_12564);
and U18189 (N_18189,N_13589,N_15579);
nand U18190 (N_18190,N_13272,N_15431);
and U18191 (N_18191,N_12938,N_12430);
or U18192 (N_18192,N_14133,N_12195);
and U18193 (N_18193,N_13545,N_12646);
nor U18194 (N_18194,N_12918,N_15177);
nor U18195 (N_18195,N_15469,N_14795);
nand U18196 (N_18196,N_15673,N_15624);
nand U18197 (N_18197,N_12123,N_14478);
nand U18198 (N_18198,N_15490,N_15660);
or U18199 (N_18199,N_15580,N_13638);
and U18200 (N_18200,N_12135,N_12713);
or U18201 (N_18201,N_13528,N_15089);
and U18202 (N_18202,N_14014,N_12727);
nand U18203 (N_18203,N_13994,N_15819);
nand U18204 (N_18204,N_15302,N_12067);
or U18205 (N_18205,N_14115,N_12448);
or U18206 (N_18206,N_13519,N_13878);
xnor U18207 (N_18207,N_14135,N_14299);
nand U18208 (N_18208,N_14602,N_15717);
nand U18209 (N_18209,N_13162,N_15700);
and U18210 (N_18210,N_12206,N_15882);
nand U18211 (N_18211,N_15660,N_13799);
nor U18212 (N_18212,N_15500,N_14188);
or U18213 (N_18213,N_13851,N_13089);
or U18214 (N_18214,N_14447,N_13955);
xnor U18215 (N_18215,N_13660,N_15376);
nand U18216 (N_18216,N_13262,N_12406);
and U18217 (N_18217,N_14506,N_13421);
and U18218 (N_18218,N_13791,N_12610);
nand U18219 (N_18219,N_12014,N_13254);
nand U18220 (N_18220,N_14798,N_12631);
nor U18221 (N_18221,N_13360,N_14329);
nand U18222 (N_18222,N_15181,N_14937);
nor U18223 (N_18223,N_15080,N_14343);
or U18224 (N_18224,N_13085,N_12367);
or U18225 (N_18225,N_12117,N_15677);
nor U18226 (N_18226,N_13280,N_12543);
and U18227 (N_18227,N_13941,N_14225);
or U18228 (N_18228,N_13097,N_15964);
or U18229 (N_18229,N_15407,N_15318);
or U18230 (N_18230,N_15122,N_14245);
and U18231 (N_18231,N_15433,N_12232);
nand U18232 (N_18232,N_12522,N_15898);
nand U18233 (N_18233,N_15097,N_13435);
and U18234 (N_18234,N_15134,N_12250);
xnor U18235 (N_18235,N_13603,N_13714);
nand U18236 (N_18236,N_15308,N_12435);
nand U18237 (N_18237,N_12526,N_15042);
nor U18238 (N_18238,N_12142,N_12073);
or U18239 (N_18239,N_15040,N_15939);
nor U18240 (N_18240,N_12543,N_12151);
and U18241 (N_18241,N_13699,N_15318);
and U18242 (N_18242,N_13937,N_14348);
or U18243 (N_18243,N_14607,N_14928);
nor U18244 (N_18244,N_14357,N_12800);
or U18245 (N_18245,N_12788,N_14005);
nor U18246 (N_18246,N_14812,N_13089);
nand U18247 (N_18247,N_15207,N_14216);
nand U18248 (N_18248,N_12149,N_13441);
and U18249 (N_18249,N_12359,N_12652);
nand U18250 (N_18250,N_14020,N_13265);
or U18251 (N_18251,N_15922,N_12504);
or U18252 (N_18252,N_14013,N_14436);
nor U18253 (N_18253,N_13651,N_14881);
and U18254 (N_18254,N_13426,N_12755);
nor U18255 (N_18255,N_14551,N_15485);
nand U18256 (N_18256,N_13818,N_13598);
nor U18257 (N_18257,N_12150,N_13910);
nand U18258 (N_18258,N_12829,N_12911);
or U18259 (N_18259,N_14479,N_13849);
nand U18260 (N_18260,N_14166,N_13550);
nor U18261 (N_18261,N_14162,N_15538);
nor U18262 (N_18262,N_14197,N_13147);
nand U18263 (N_18263,N_15060,N_13391);
nor U18264 (N_18264,N_15680,N_13783);
nor U18265 (N_18265,N_12651,N_15187);
nand U18266 (N_18266,N_15491,N_15370);
and U18267 (N_18267,N_13440,N_13544);
or U18268 (N_18268,N_13649,N_14428);
xor U18269 (N_18269,N_14839,N_12032);
nor U18270 (N_18270,N_13332,N_15648);
or U18271 (N_18271,N_13098,N_12305);
nand U18272 (N_18272,N_13535,N_14543);
or U18273 (N_18273,N_13151,N_13661);
and U18274 (N_18274,N_13825,N_14592);
and U18275 (N_18275,N_12078,N_15396);
nand U18276 (N_18276,N_12087,N_14881);
nand U18277 (N_18277,N_14724,N_15788);
nor U18278 (N_18278,N_13944,N_14455);
nor U18279 (N_18279,N_14070,N_12660);
or U18280 (N_18280,N_13982,N_15671);
and U18281 (N_18281,N_12706,N_13067);
or U18282 (N_18282,N_15908,N_13510);
and U18283 (N_18283,N_14285,N_14967);
nor U18284 (N_18284,N_13776,N_13653);
and U18285 (N_18285,N_13197,N_12976);
or U18286 (N_18286,N_13903,N_13066);
nand U18287 (N_18287,N_13678,N_14884);
nor U18288 (N_18288,N_12728,N_15771);
xnor U18289 (N_18289,N_14127,N_13092);
and U18290 (N_18290,N_15440,N_13009);
and U18291 (N_18291,N_12228,N_12337);
nor U18292 (N_18292,N_12572,N_13030);
nand U18293 (N_18293,N_14255,N_13957);
and U18294 (N_18294,N_13718,N_12281);
or U18295 (N_18295,N_14823,N_14398);
nor U18296 (N_18296,N_12429,N_14869);
and U18297 (N_18297,N_13158,N_15216);
xnor U18298 (N_18298,N_15763,N_12834);
nand U18299 (N_18299,N_13566,N_14072);
nor U18300 (N_18300,N_15941,N_13370);
xnor U18301 (N_18301,N_13697,N_12239);
or U18302 (N_18302,N_14093,N_13075);
and U18303 (N_18303,N_14431,N_14913);
nor U18304 (N_18304,N_14547,N_14089);
nor U18305 (N_18305,N_15012,N_14829);
nor U18306 (N_18306,N_15470,N_14260);
xor U18307 (N_18307,N_12871,N_15301);
and U18308 (N_18308,N_12661,N_15897);
and U18309 (N_18309,N_13103,N_13288);
and U18310 (N_18310,N_12922,N_14739);
and U18311 (N_18311,N_15403,N_14448);
nor U18312 (N_18312,N_14561,N_12211);
nor U18313 (N_18313,N_12888,N_14765);
and U18314 (N_18314,N_13616,N_12451);
and U18315 (N_18315,N_13631,N_12205);
nor U18316 (N_18316,N_13255,N_12273);
nand U18317 (N_18317,N_14619,N_15554);
nand U18318 (N_18318,N_15886,N_13882);
or U18319 (N_18319,N_14900,N_13456);
nor U18320 (N_18320,N_13938,N_14202);
and U18321 (N_18321,N_14924,N_15838);
nor U18322 (N_18322,N_15137,N_15862);
nor U18323 (N_18323,N_15408,N_13024);
and U18324 (N_18324,N_12217,N_14643);
or U18325 (N_18325,N_14849,N_14112);
or U18326 (N_18326,N_14338,N_12723);
nor U18327 (N_18327,N_13452,N_15592);
nand U18328 (N_18328,N_14713,N_12780);
nand U18329 (N_18329,N_15763,N_13431);
and U18330 (N_18330,N_13046,N_12639);
nand U18331 (N_18331,N_13945,N_14167);
or U18332 (N_18332,N_12145,N_12350);
nor U18333 (N_18333,N_12410,N_14829);
nand U18334 (N_18334,N_13343,N_12203);
and U18335 (N_18335,N_14540,N_12903);
nor U18336 (N_18336,N_13806,N_15795);
xor U18337 (N_18337,N_14110,N_12945);
xor U18338 (N_18338,N_12931,N_12471);
and U18339 (N_18339,N_14707,N_13708);
nor U18340 (N_18340,N_15430,N_15753);
or U18341 (N_18341,N_15998,N_14799);
nor U18342 (N_18342,N_13430,N_14435);
nand U18343 (N_18343,N_12713,N_15607);
nand U18344 (N_18344,N_12141,N_14819);
nand U18345 (N_18345,N_12117,N_13635);
xnor U18346 (N_18346,N_14146,N_12498);
or U18347 (N_18347,N_12173,N_13449);
or U18348 (N_18348,N_14563,N_12211);
and U18349 (N_18349,N_15494,N_14380);
and U18350 (N_18350,N_14675,N_12962);
nand U18351 (N_18351,N_12041,N_13580);
or U18352 (N_18352,N_15774,N_15532);
xnor U18353 (N_18353,N_14299,N_12147);
xnor U18354 (N_18354,N_14639,N_14633);
and U18355 (N_18355,N_14141,N_14145);
and U18356 (N_18356,N_12519,N_13350);
nor U18357 (N_18357,N_15593,N_13471);
xnor U18358 (N_18358,N_15945,N_14375);
and U18359 (N_18359,N_15364,N_14978);
or U18360 (N_18360,N_13142,N_13977);
nand U18361 (N_18361,N_13910,N_13540);
xor U18362 (N_18362,N_13810,N_14372);
nand U18363 (N_18363,N_13989,N_12475);
or U18364 (N_18364,N_15331,N_14722);
nand U18365 (N_18365,N_12893,N_14369);
or U18366 (N_18366,N_13529,N_15305);
or U18367 (N_18367,N_12010,N_12265);
or U18368 (N_18368,N_15305,N_14228);
or U18369 (N_18369,N_13808,N_15680);
nor U18370 (N_18370,N_15294,N_14794);
or U18371 (N_18371,N_15251,N_12960);
xor U18372 (N_18372,N_15227,N_13683);
and U18373 (N_18373,N_14281,N_12035);
xor U18374 (N_18374,N_13497,N_13282);
nand U18375 (N_18375,N_13337,N_15872);
and U18376 (N_18376,N_15295,N_15252);
nand U18377 (N_18377,N_15123,N_13879);
and U18378 (N_18378,N_12638,N_14032);
xnor U18379 (N_18379,N_12996,N_12127);
or U18380 (N_18380,N_15610,N_12853);
or U18381 (N_18381,N_12772,N_15637);
and U18382 (N_18382,N_15444,N_14825);
nand U18383 (N_18383,N_13938,N_14717);
nor U18384 (N_18384,N_13857,N_12483);
nand U18385 (N_18385,N_15310,N_15115);
or U18386 (N_18386,N_12124,N_14745);
and U18387 (N_18387,N_15983,N_14570);
and U18388 (N_18388,N_15079,N_14206);
and U18389 (N_18389,N_12582,N_15086);
or U18390 (N_18390,N_14151,N_13645);
xor U18391 (N_18391,N_12393,N_12244);
or U18392 (N_18392,N_15544,N_13375);
or U18393 (N_18393,N_12917,N_12236);
and U18394 (N_18394,N_13933,N_13304);
nor U18395 (N_18395,N_14452,N_15651);
or U18396 (N_18396,N_12481,N_12232);
or U18397 (N_18397,N_14250,N_12933);
or U18398 (N_18398,N_13326,N_12109);
or U18399 (N_18399,N_13451,N_14772);
or U18400 (N_18400,N_15098,N_13684);
and U18401 (N_18401,N_12810,N_14031);
or U18402 (N_18402,N_14903,N_13317);
or U18403 (N_18403,N_13739,N_15035);
or U18404 (N_18404,N_13157,N_14752);
or U18405 (N_18405,N_13071,N_15449);
and U18406 (N_18406,N_12656,N_13569);
or U18407 (N_18407,N_15052,N_14912);
and U18408 (N_18408,N_15743,N_13648);
nand U18409 (N_18409,N_12775,N_12242);
or U18410 (N_18410,N_12117,N_15164);
nand U18411 (N_18411,N_15961,N_13847);
nor U18412 (N_18412,N_13250,N_14393);
xor U18413 (N_18413,N_14070,N_14727);
nor U18414 (N_18414,N_13485,N_15449);
xnor U18415 (N_18415,N_13227,N_13933);
nor U18416 (N_18416,N_12007,N_13199);
nand U18417 (N_18417,N_14364,N_12878);
or U18418 (N_18418,N_13558,N_12065);
nand U18419 (N_18419,N_15640,N_13697);
or U18420 (N_18420,N_13847,N_14578);
nor U18421 (N_18421,N_14972,N_15168);
or U18422 (N_18422,N_12062,N_15764);
xor U18423 (N_18423,N_13370,N_15878);
nor U18424 (N_18424,N_13900,N_15890);
or U18425 (N_18425,N_13317,N_12123);
or U18426 (N_18426,N_13586,N_12689);
or U18427 (N_18427,N_14317,N_12995);
nor U18428 (N_18428,N_13281,N_12226);
and U18429 (N_18429,N_13711,N_13907);
nand U18430 (N_18430,N_12613,N_13792);
and U18431 (N_18431,N_12534,N_13451);
and U18432 (N_18432,N_14189,N_13798);
xnor U18433 (N_18433,N_12282,N_13275);
or U18434 (N_18434,N_15897,N_14233);
or U18435 (N_18435,N_13703,N_14327);
nor U18436 (N_18436,N_15733,N_13142);
xnor U18437 (N_18437,N_15947,N_15730);
and U18438 (N_18438,N_14299,N_13921);
nand U18439 (N_18439,N_12033,N_14342);
or U18440 (N_18440,N_12174,N_13839);
or U18441 (N_18441,N_13875,N_15798);
and U18442 (N_18442,N_14925,N_12684);
nor U18443 (N_18443,N_13118,N_14234);
nor U18444 (N_18444,N_14240,N_14690);
nor U18445 (N_18445,N_12287,N_15698);
or U18446 (N_18446,N_12485,N_12571);
nor U18447 (N_18447,N_14000,N_14156);
nand U18448 (N_18448,N_13166,N_14411);
or U18449 (N_18449,N_12482,N_13571);
nand U18450 (N_18450,N_12268,N_13878);
nand U18451 (N_18451,N_12445,N_15334);
xor U18452 (N_18452,N_14661,N_13258);
and U18453 (N_18453,N_15298,N_13516);
nand U18454 (N_18454,N_14573,N_14330);
nand U18455 (N_18455,N_15503,N_13870);
nand U18456 (N_18456,N_15569,N_14754);
nand U18457 (N_18457,N_13672,N_13886);
and U18458 (N_18458,N_12307,N_13546);
or U18459 (N_18459,N_12834,N_12672);
nor U18460 (N_18460,N_14656,N_14749);
or U18461 (N_18461,N_14546,N_15718);
nor U18462 (N_18462,N_14892,N_14346);
nor U18463 (N_18463,N_12057,N_13057);
nor U18464 (N_18464,N_12165,N_14088);
and U18465 (N_18465,N_15463,N_15944);
and U18466 (N_18466,N_14092,N_12446);
nand U18467 (N_18467,N_15961,N_12880);
nand U18468 (N_18468,N_13416,N_15038);
nor U18469 (N_18469,N_14872,N_14877);
and U18470 (N_18470,N_15648,N_15479);
and U18471 (N_18471,N_14312,N_14969);
or U18472 (N_18472,N_13427,N_13641);
and U18473 (N_18473,N_12471,N_14896);
or U18474 (N_18474,N_14759,N_13044);
nor U18475 (N_18475,N_13878,N_14040);
nand U18476 (N_18476,N_13268,N_13236);
nand U18477 (N_18477,N_15169,N_14728);
nor U18478 (N_18478,N_12820,N_15952);
or U18479 (N_18479,N_13332,N_13952);
xor U18480 (N_18480,N_14916,N_12880);
nor U18481 (N_18481,N_13686,N_12608);
nor U18482 (N_18482,N_14197,N_15233);
and U18483 (N_18483,N_12563,N_13320);
nand U18484 (N_18484,N_15597,N_15027);
nand U18485 (N_18485,N_12572,N_15571);
and U18486 (N_18486,N_13707,N_15546);
and U18487 (N_18487,N_13641,N_14078);
xnor U18488 (N_18488,N_14709,N_14754);
or U18489 (N_18489,N_12670,N_12368);
nor U18490 (N_18490,N_14454,N_15390);
nor U18491 (N_18491,N_12508,N_14269);
nor U18492 (N_18492,N_15725,N_14647);
or U18493 (N_18493,N_12516,N_14935);
nor U18494 (N_18494,N_12005,N_13049);
or U18495 (N_18495,N_13772,N_14032);
and U18496 (N_18496,N_12219,N_14700);
and U18497 (N_18497,N_13290,N_13825);
nand U18498 (N_18498,N_12357,N_13672);
nand U18499 (N_18499,N_14357,N_15969);
nor U18500 (N_18500,N_12876,N_13986);
and U18501 (N_18501,N_13959,N_15974);
nor U18502 (N_18502,N_12511,N_14399);
or U18503 (N_18503,N_14544,N_15985);
xor U18504 (N_18504,N_13947,N_14853);
or U18505 (N_18505,N_12882,N_15830);
and U18506 (N_18506,N_13699,N_15058);
nand U18507 (N_18507,N_13948,N_14008);
xor U18508 (N_18508,N_13753,N_14539);
nand U18509 (N_18509,N_14656,N_15267);
nand U18510 (N_18510,N_15169,N_14648);
nand U18511 (N_18511,N_12898,N_12049);
and U18512 (N_18512,N_14150,N_15681);
or U18513 (N_18513,N_13264,N_14896);
nand U18514 (N_18514,N_15763,N_14320);
nand U18515 (N_18515,N_14299,N_14191);
nand U18516 (N_18516,N_13370,N_13043);
and U18517 (N_18517,N_13870,N_12018);
nand U18518 (N_18518,N_13245,N_14379);
nor U18519 (N_18519,N_12529,N_13734);
and U18520 (N_18520,N_13301,N_13311);
nand U18521 (N_18521,N_12449,N_14731);
and U18522 (N_18522,N_12983,N_15430);
nor U18523 (N_18523,N_14071,N_14821);
or U18524 (N_18524,N_15138,N_14837);
or U18525 (N_18525,N_13924,N_15868);
and U18526 (N_18526,N_15666,N_12630);
nand U18527 (N_18527,N_15638,N_15102);
nor U18528 (N_18528,N_15134,N_12345);
and U18529 (N_18529,N_14842,N_15661);
and U18530 (N_18530,N_13861,N_13730);
and U18531 (N_18531,N_14542,N_13454);
or U18532 (N_18532,N_15299,N_12149);
nand U18533 (N_18533,N_15152,N_12858);
nor U18534 (N_18534,N_15483,N_14056);
nand U18535 (N_18535,N_13404,N_13469);
nand U18536 (N_18536,N_13865,N_12541);
and U18537 (N_18537,N_14148,N_12131);
nor U18538 (N_18538,N_15063,N_15632);
and U18539 (N_18539,N_12245,N_15858);
and U18540 (N_18540,N_15049,N_13285);
or U18541 (N_18541,N_12632,N_15668);
and U18542 (N_18542,N_12758,N_12746);
or U18543 (N_18543,N_14622,N_15371);
xor U18544 (N_18544,N_12456,N_15428);
and U18545 (N_18545,N_13118,N_15960);
xor U18546 (N_18546,N_15102,N_12279);
nand U18547 (N_18547,N_15245,N_14451);
nand U18548 (N_18548,N_13628,N_14321);
and U18549 (N_18549,N_15274,N_15582);
xnor U18550 (N_18550,N_15678,N_13446);
nor U18551 (N_18551,N_13787,N_13972);
or U18552 (N_18552,N_13848,N_13092);
and U18553 (N_18553,N_14290,N_15813);
and U18554 (N_18554,N_15548,N_12204);
and U18555 (N_18555,N_15505,N_15176);
nand U18556 (N_18556,N_13241,N_14585);
nand U18557 (N_18557,N_15634,N_14435);
and U18558 (N_18558,N_14734,N_15700);
nor U18559 (N_18559,N_14287,N_12919);
nand U18560 (N_18560,N_14804,N_12508);
and U18561 (N_18561,N_12514,N_15857);
nor U18562 (N_18562,N_14383,N_14358);
nand U18563 (N_18563,N_14744,N_15211);
nor U18564 (N_18564,N_13409,N_13509);
or U18565 (N_18565,N_15115,N_13739);
or U18566 (N_18566,N_13242,N_14400);
and U18567 (N_18567,N_14088,N_14057);
nand U18568 (N_18568,N_14300,N_14233);
nor U18569 (N_18569,N_13023,N_15302);
nor U18570 (N_18570,N_14662,N_13565);
nand U18571 (N_18571,N_14667,N_12968);
and U18572 (N_18572,N_13064,N_13796);
and U18573 (N_18573,N_14767,N_13983);
nand U18574 (N_18574,N_15850,N_14695);
nand U18575 (N_18575,N_14691,N_15468);
and U18576 (N_18576,N_13004,N_14470);
nand U18577 (N_18577,N_13210,N_12353);
nand U18578 (N_18578,N_13287,N_14461);
or U18579 (N_18579,N_15236,N_12971);
xnor U18580 (N_18580,N_14265,N_13533);
nor U18581 (N_18581,N_12819,N_14034);
or U18582 (N_18582,N_13330,N_13574);
nand U18583 (N_18583,N_13260,N_14899);
nand U18584 (N_18584,N_12941,N_15170);
nand U18585 (N_18585,N_13820,N_14800);
nor U18586 (N_18586,N_12003,N_12788);
nand U18587 (N_18587,N_13381,N_14695);
and U18588 (N_18588,N_14382,N_13452);
nor U18589 (N_18589,N_12876,N_13328);
nand U18590 (N_18590,N_15040,N_14318);
or U18591 (N_18591,N_15623,N_12794);
nand U18592 (N_18592,N_14656,N_13744);
nor U18593 (N_18593,N_13762,N_13496);
nor U18594 (N_18594,N_13224,N_15880);
nand U18595 (N_18595,N_13491,N_15486);
nand U18596 (N_18596,N_15214,N_14155);
or U18597 (N_18597,N_13684,N_13094);
or U18598 (N_18598,N_13691,N_13387);
nand U18599 (N_18599,N_13623,N_15542);
and U18600 (N_18600,N_13774,N_13706);
nand U18601 (N_18601,N_12882,N_12387);
nand U18602 (N_18602,N_14949,N_15499);
xnor U18603 (N_18603,N_13444,N_15224);
xnor U18604 (N_18604,N_14644,N_15163);
and U18605 (N_18605,N_15544,N_12343);
and U18606 (N_18606,N_14294,N_14868);
or U18607 (N_18607,N_15992,N_15659);
or U18608 (N_18608,N_13607,N_15972);
nand U18609 (N_18609,N_15177,N_13660);
nand U18610 (N_18610,N_14806,N_14183);
and U18611 (N_18611,N_15138,N_12927);
nor U18612 (N_18612,N_14351,N_14756);
nor U18613 (N_18613,N_13016,N_13604);
nand U18614 (N_18614,N_14891,N_13436);
and U18615 (N_18615,N_12169,N_12779);
nor U18616 (N_18616,N_13997,N_14395);
and U18617 (N_18617,N_12135,N_14119);
nor U18618 (N_18618,N_14632,N_12213);
nand U18619 (N_18619,N_14815,N_12774);
or U18620 (N_18620,N_14931,N_13658);
nor U18621 (N_18621,N_13199,N_14111);
nand U18622 (N_18622,N_15317,N_12324);
nand U18623 (N_18623,N_15649,N_15854);
nor U18624 (N_18624,N_15753,N_13912);
and U18625 (N_18625,N_13072,N_12599);
or U18626 (N_18626,N_14223,N_15986);
nor U18627 (N_18627,N_12926,N_13295);
and U18628 (N_18628,N_14808,N_14388);
nand U18629 (N_18629,N_12122,N_14582);
and U18630 (N_18630,N_14680,N_13776);
nor U18631 (N_18631,N_12981,N_15362);
nor U18632 (N_18632,N_12981,N_15549);
xnor U18633 (N_18633,N_15059,N_12346);
nor U18634 (N_18634,N_15360,N_12698);
nor U18635 (N_18635,N_13781,N_14723);
nand U18636 (N_18636,N_13052,N_13953);
nor U18637 (N_18637,N_13053,N_14454);
nor U18638 (N_18638,N_13116,N_14089);
nand U18639 (N_18639,N_15802,N_13267);
nand U18640 (N_18640,N_15447,N_15749);
xor U18641 (N_18641,N_14630,N_14574);
and U18642 (N_18642,N_12888,N_14920);
or U18643 (N_18643,N_12016,N_15743);
xnor U18644 (N_18644,N_15288,N_14893);
nor U18645 (N_18645,N_13286,N_14098);
nor U18646 (N_18646,N_14033,N_14172);
and U18647 (N_18647,N_12204,N_13955);
nand U18648 (N_18648,N_13836,N_15356);
or U18649 (N_18649,N_14301,N_15296);
nor U18650 (N_18650,N_14036,N_14918);
nor U18651 (N_18651,N_13846,N_13529);
or U18652 (N_18652,N_15877,N_13093);
nor U18653 (N_18653,N_12967,N_14772);
and U18654 (N_18654,N_15203,N_14931);
or U18655 (N_18655,N_12757,N_12092);
nand U18656 (N_18656,N_12049,N_14665);
xnor U18657 (N_18657,N_14775,N_13346);
and U18658 (N_18658,N_15707,N_15541);
nand U18659 (N_18659,N_13200,N_14874);
or U18660 (N_18660,N_12560,N_13819);
and U18661 (N_18661,N_14008,N_15135);
and U18662 (N_18662,N_14315,N_15733);
nand U18663 (N_18663,N_13613,N_15701);
nand U18664 (N_18664,N_12972,N_14637);
or U18665 (N_18665,N_12938,N_12605);
nor U18666 (N_18666,N_14750,N_14123);
nor U18667 (N_18667,N_13810,N_13817);
and U18668 (N_18668,N_13981,N_12428);
or U18669 (N_18669,N_14829,N_12139);
and U18670 (N_18670,N_13351,N_12021);
and U18671 (N_18671,N_12260,N_13292);
or U18672 (N_18672,N_15165,N_12245);
and U18673 (N_18673,N_14983,N_14138);
and U18674 (N_18674,N_13579,N_13522);
and U18675 (N_18675,N_12632,N_15660);
xor U18676 (N_18676,N_12043,N_14309);
nand U18677 (N_18677,N_14260,N_13389);
nand U18678 (N_18678,N_15180,N_12219);
nor U18679 (N_18679,N_13127,N_15603);
or U18680 (N_18680,N_12069,N_15704);
or U18681 (N_18681,N_15597,N_12692);
and U18682 (N_18682,N_13170,N_14100);
nor U18683 (N_18683,N_13546,N_12275);
xnor U18684 (N_18684,N_12884,N_13481);
xnor U18685 (N_18685,N_14704,N_14855);
and U18686 (N_18686,N_13623,N_12217);
and U18687 (N_18687,N_12858,N_12325);
nor U18688 (N_18688,N_14063,N_13195);
nor U18689 (N_18689,N_13019,N_14005);
nor U18690 (N_18690,N_12967,N_12460);
and U18691 (N_18691,N_13417,N_12412);
xnor U18692 (N_18692,N_14745,N_14435);
or U18693 (N_18693,N_13079,N_13530);
nand U18694 (N_18694,N_12642,N_14696);
xor U18695 (N_18695,N_14458,N_14129);
nand U18696 (N_18696,N_13014,N_15391);
xor U18697 (N_18697,N_15914,N_14407);
nand U18698 (N_18698,N_13699,N_13817);
and U18699 (N_18699,N_15041,N_12162);
or U18700 (N_18700,N_12114,N_15041);
nor U18701 (N_18701,N_15572,N_12402);
and U18702 (N_18702,N_15557,N_15077);
or U18703 (N_18703,N_12764,N_13532);
nor U18704 (N_18704,N_15932,N_14978);
or U18705 (N_18705,N_15520,N_14246);
nor U18706 (N_18706,N_13098,N_13418);
xnor U18707 (N_18707,N_14430,N_13320);
and U18708 (N_18708,N_14695,N_12527);
or U18709 (N_18709,N_12689,N_14075);
nand U18710 (N_18710,N_13533,N_14041);
nor U18711 (N_18711,N_15107,N_12403);
nand U18712 (N_18712,N_13034,N_15908);
nor U18713 (N_18713,N_15000,N_15900);
and U18714 (N_18714,N_14950,N_13129);
and U18715 (N_18715,N_14495,N_15385);
or U18716 (N_18716,N_14554,N_15070);
nor U18717 (N_18717,N_14590,N_13377);
nor U18718 (N_18718,N_12628,N_15800);
or U18719 (N_18719,N_13555,N_12687);
and U18720 (N_18720,N_12733,N_13336);
or U18721 (N_18721,N_15268,N_12301);
xor U18722 (N_18722,N_15434,N_15549);
and U18723 (N_18723,N_13496,N_13181);
or U18724 (N_18724,N_13749,N_14790);
nand U18725 (N_18725,N_13140,N_14033);
and U18726 (N_18726,N_13379,N_13076);
nand U18727 (N_18727,N_14748,N_15982);
nor U18728 (N_18728,N_13804,N_14975);
xor U18729 (N_18729,N_13340,N_12025);
or U18730 (N_18730,N_12560,N_12541);
nand U18731 (N_18731,N_12463,N_13641);
nor U18732 (N_18732,N_13091,N_14777);
nor U18733 (N_18733,N_15272,N_13450);
nor U18734 (N_18734,N_15247,N_12915);
and U18735 (N_18735,N_12790,N_12975);
nand U18736 (N_18736,N_12457,N_13728);
or U18737 (N_18737,N_12316,N_13112);
nand U18738 (N_18738,N_12737,N_14590);
nor U18739 (N_18739,N_13901,N_12871);
nor U18740 (N_18740,N_13391,N_15900);
or U18741 (N_18741,N_12276,N_14289);
or U18742 (N_18742,N_14921,N_12221);
or U18743 (N_18743,N_12668,N_14765);
and U18744 (N_18744,N_12362,N_15116);
and U18745 (N_18745,N_12233,N_13361);
and U18746 (N_18746,N_13683,N_12461);
or U18747 (N_18747,N_12389,N_15450);
nor U18748 (N_18748,N_15491,N_13886);
or U18749 (N_18749,N_12779,N_15298);
nor U18750 (N_18750,N_15520,N_12165);
nor U18751 (N_18751,N_14502,N_13926);
xor U18752 (N_18752,N_12911,N_12930);
or U18753 (N_18753,N_13979,N_13620);
nand U18754 (N_18754,N_12428,N_13922);
and U18755 (N_18755,N_13041,N_14614);
xnor U18756 (N_18756,N_12572,N_13037);
xnor U18757 (N_18757,N_12293,N_14465);
nand U18758 (N_18758,N_15371,N_15579);
nand U18759 (N_18759,N_15874,N_12126);
and U18760 (N_18760,N_12992,N_13088);
nand U18761 (N_18761,N_12510,N_13218);
xnor U18762 (N_18762,N_13889,N_14506);
or U18763 (N_18763,N_15585,N_12794);
and U18764 (N_18764,N_14042,N_12568);
or U18765 (N_18765,N_15060,N_14100);
nor U18766 (N_18766,N_14078,N_14807);
nand U18767 (N_18767,N_15331,N_14504);
or U18768 (N_18768,N_12230,N_15553);
xor U18769 (N_18769,N_12406,N_14352);
nand U18770 (N_18770,N_13423,N_13955);
and U18771 (N_18771,N_13310,N_14052);
and U18772 (N_18772,N_12984,N_15839);
or U18773 (N_18773,N_15789,N_12432);
nor U18774 (N_18774,N_13166,N_14566);
and U18775 (N_18775,N_13052,N_15360);
xnor U18776 (N_18776,N_14830,N_12515);
and U18777 (N_18777,N_14969,N_15401);
xnor U18778 (N_18778,N_12940,N_14895);
or U18779 (N_18779,N_12479,N_13407);
or U18780 (N_18780,N_14952,N_14298);
or U18781 (N_18781,N_14142,N_14176);
xor U18782 (N_18782,N_12124,N_13556);
xnor U18783 (N_18783,N_12442,N_15349);
nand U18784 (N_18784,N_14324,N_14995);
xor U18785 (N_18785,N_15561,N_14872);
and U18786 (N_18786,N_13359,N_15708);
or U18787 (N_18787,N_12717,N_12927);
nand U18788 (N_18788,N_13152,N_12849);
nor U18789 (N_18789,N_13214,N_15397);
or U18790 (N_18790,N_15557,N_13061);
xnor U18791 (N_18791,N_15734,N_14853);
and U18792 (N_18792,N_12554,N_15790);
nand U18793 (N_18793,N_12710,N_12567);
or U18794 (N_18794,N_13334,N_14254);
nand U18795 (N_18795,N_13579,N_15805);
xor U18796 (N_18796,N_12573,N_13047);
nand U18797 (N_18797,N_12322,N_15331);
nand U18798 (N_18798,N_14025,N_13622);
and U18799 (N_18799,N_15738,N_13213);
xor U18800 (N_18800,N_15059,N_15620);
nand U18801 (N_18801,N_14325,N_12849);
or U18802 (N_18802,N_12122,N_14033);
nor U18803 (N_18803,N_15447,N_14741);
xor U18804 (N_18804,N_13730,N_13297);
nand U18805 (N_18805,N_12202,N_14946);
xor U18806 (N_18806,N_14886,N_15937);
xor U18807 (N_18807,N_14445,N_12598);
and U18808 (N_18808,N_15464,N_15643);
xor U18809 (N_18809,N_12541,N_14191);
nand U18810 (N_18810,N_15459,N_14919);
or U18811 (N_18811,N_13883,N_15179);
or U18812 (N_18812,N_12853,N_12765);
nor U18813 (N_18813,N_13342,N_13940);
and U18814 (N_18814,N_12434,N_13861);
or U18815 (N_18815,N_13964,N_14381);
nand U18816 (N_18816,N_12279,N_13924);
nor U18817 (N_18817,N_12000,N_15254);
or U18818 (N_18818,N_12364,N_12019);
and U18819 (N_18819,N_14770,N_15959);
and U18820 (N_18820,N_13491,N_14417);
and U18821 (N_18821,N_14019,N_13178);
or U18822 (N_18822,N_12945,N_13024);
nor U18823 (N_18823,N_14221,N_13942);
xnor U18824 (N_18824,N_13323,N_13460);
or U18825 (N_18825,N_13095,N_13698);
and U18826 (N_18826,N_13991,N_12464);
or U18827 (N_18827,N_12436,N_15764);
nand U18828 (N_18828,N_14711,N_13396);
or U18829 (N_18829,N_15953,N_14519);
nor U18830 (N_18830,N_14805,N_15505);
nand U18831 (N_18831,N_12369,N_15594);
nand U18832 (N_18832,N_14885,N_14092);
nor U18833 (N_18833,N_12567,N_12161);
and U18834 (N_18834,N_13258,N_13353);
or U18835 (N_18835,N_15517,N_12570);
nor U18836 (N_18836,N_12128,N_13143);
nand U18837 (N_18837,N_13748,N_13594);
nand U18838 (N_18838,N_14382,N_14788);
nand U18839 (N_18839,N_13177,N_15941);
nand U18840 (N_18840,N_15867,N_13917);
nand U18841 (N_18841,N_12813,N_12716);
nor U18842 (N_18842,N_12311,N_13826);
and U18843 (N_18843,N_14678,N_14908);
nor U18844 (N_18844,N_14465,N_15408);
nor U18845 (N_18845,N_12925,N_15067);
or U18846 (N_18846,N_13603,N_12246);
or U18847 (N_18847,N_12437,N_12025);
and U18848 (N_18848,N_15829,N_13043);
xnor U18849 (N_18849,N_14969,N_15753);
and U18850 (N_18850,N_13514,N_14839);
or U18851 (N_18851,N_13734,N_13778);
or U18852 (N_18852,N_13965,N_14013);
nor U18853 (N_18853,N_14317,N_13801);
nor U18854 (N_18854,N_12827,N_12058);
and U18855 (N_18855,N_15208,N_15706);
and U18856 (N_18856,N_14075,N_15699);
or U18857 (N_18857,N_12974,N_15851);
and U18858 (N_18858,N_14453,N_14270);
nand U18859 (N_18859,N_15749,N_15490);
nor U18860 (N_18860,N_14953,N_13931);
nor U18861 (N_18861,N_14265,N_15400);
xnor U18862 (N_18862,N_15873,N_13135);
nor U18863 (N_18863,N_12531,N_12713);
nand U18864 (N_18864,N_15222,N_14537);
and U18865 (N_18865,N_15621,N_12414);
or U18866 (N_18866,N_12844,N_14704);
nor U18867 (N_18867,N_12156,N_15794);
and U18868 (N_18868,N_14386,N_15616);
and U18869 (N_18869,N_15164,N_12325);
nor U18870 (N_18870,N_13190,N_12623);
nor U18871 (N_18871,N_14778,N_12543);
or U18872 (N_18872,N_15981,N_15754);
or U18873 (N_18873,N_12104,N_14561);
nand U18874 (N_18874,N_13072,N_12253);
nor U18875 (N_18875,N_13434,N_13084);
nand U18876 (N_18876,N_12335,N_14051);
or U18877 (N_18877,N_14936,N_15815);
nand U18878 (N_18878,N_13436,N_12421);
or U18879 (N_18879,N_15440,N_14159);
or U18880 (N_18880,N_12330,N_13748);
nor U18881 (N_18881,N_15712,N_15074);
nand U18882 (N_18882,N_15379,N_12962);
nand U18883 (N_18883,N_14762,N_13422);
nand U18884 (N_18884,N_13237,N_14245);
nand U18885 (N_18885,N_15282,N_14313);
and U18886 (N_18886,N_14727,N_14510);
nor U18887 (N_18887,N_15643,N_13319);
xnor U18888 (N_18888,N_15321,N_15612);
or U18889 (N_18889,N_15907,N_14190);
nor U18890 (N_18890,N_12713,N_12997);
nand U18891 (N_18891,N_14020,N_15581);
xor U18892 (N_18892,N_12100,N_15842);
or U18893 (N_18893,N_15423,N_14541);
and U18894 (N_18894,N_13615,N_12485);
and U18895 (N_18895,N_13726,N_12222);
nor U18896 (N_18896,N_14429,N_14948);
nand U18897 (N_18897,N_14398,N_12958);
xnor U18898 (N_18898,N_12986,N_13309);
and U18899 (N_18899,N_13543,N_15596);
nor U18900 (N_18900,N_13621,N_12770);
nand U18901 (N_18901,N_14731,N_12724);
nor U18902 (N_18902,N_14502,N_12760);
or U18903 (N_18903,N_15331,N_12255);
and U18904 (N_18904,N_15226,N_12459);
or U18905 (N_18905,N_13289,N_13347);
or U18906 (N_18906,N_15935,N_15500);
nand U18907 (N_18907,N_13893,N_14518);
nor U18908 (N_18908,N_14184,N_13526);
and U18909 (N_18909,N_14645,N_14013);
nand U18910 (N_18910,N_15718,N_13377);
or U18911 (N_18911,N_14392,N_15092);
nand U18912 (N_18912,N_13822,N_14184);
nand U18913 (N_18913,N_12304,N_14017);
nor U18914 (N_18914,N_12056,N_15755);
and U18915 (N_18915,N_15205,N_14017);
or U18916 (N_18916,N_13842,N_12390);
xnor U18917 (N_18917,N_15318,N_12097);
nor U18918 (N_18918,N_13450,N_12933);
and U18919 (N_18919,N_14294,N_15118);
nor U18920 (N_18920,N_13147,N_13759);
and U18921 (N_18921,N_12751,N_13424);
nor U18922 (N_18922,N_12088,N_14547);
nand U18923 (N_18923,N_13863,N_15858);
nand U18924 (N_18924,N_12325,N_13035);
xnor U18925 (N_18925,N_14310,N_15821);
nand U18926 (N_18926,N_15505,N_14342);
nor U18927 (N_18927,N_15290,N_12461);
or U18928 (N_18928,N_12681,N_14799);
and U18929 (N_18929,N_14404,N_14246);
xor U18930 (N_18930,N_13215,N_13730);
nor U18931 (N_18931,N_13326,N_13160);
and U18932 (N_18932,N_13853,N_15086);
and U18933 (N_18933,N_12168,N_14797);
or U18934 (N_18934,N_15448,N_12028);
and U18935 (N_18935,N_13613,N_15506);
nor U18936 (N_18936,N_15333,N_14790);
and U18937 (N_18937,N_15042,N_13159);
and U18938 (N_18938,N_12225,N_13351);
nor U18939 (N_18939,N_13511,N_14005);
or U18940 (N_18940,N_15897,N_12833);
or U18941 (N_18941,N_12831,N_13860);
nand U18942 (N_18942,N_15933,N_14820);
nor U18943 (N_18943,N_13820,N_12205);
nand U18944 (N_18944,N_15184,N_15697);
xor U18945 (N_18945,N_13523,N_12120);
nor U18946 (N_18946,N_12280,N_15057);
or U18947 (N_18947,N_15239,N_15533);
xnor U18948 (N_18948,N_14477,N_15524);
nor U18949 (N_18949,N_12825,N_13589);
or U18950 (N_18950,N_13637,N_13531);
nor U18951 (N_18951,N_12863,N_12834);
and U18952 (N_18952,N_12241,N_13181);
and U18953 (N_18953,N_13967,N_12736);
nor U18954 (N_18954,N_12040,N_13155);
or U18955 (N_18955,N_15390,N_13678);
and U18956 (N_18956,N_14895,N_13914);
nor U18957 (N_18957,N_15605,N_13281);
or U18958 (N_18958,N_13514,N_13835);
and U18959 (N_18959,N_14039,N_15834);
or U18960 (N_18960,N_12331,N_12241);
nand U18961 (N_18961,N_12888,N_13892);
nand U18962 (N_18962,N_13851,N_14667);
nor U18963 (N_18963,N_12227,N_14149);
and U18964 (N_18964,N_12726,N_14528);
or U18965 (N_18965,N_12877,N_15229);
or U18966 (N_18966,N_14559,N_12487);
or U18967 (N_18967,N_15341,N_12233);
xnor U18968 (N_18968,N_15593,N_15251);
nand U18969 (N_18969,N_13346,N_15188);
nand U18970 (N_18970,N_14006,N_12858);
or U18971 (N_18971,N_13212,N_13902);
nand U18972 (N_18972,N_15184,N_12886);
and U18973 (N_18973,N_15501,N_12872);
nand U18974 (N_18974,N_12252,N_14570);
nor U18975 (N_18975,N_14326,N_13628);
or U18976 (N_18976,N_12566,N_15071);
nor U18977 (N_18977,N_12667,N_14695);
and U18978 (N_18978,N_13525,N_13629);
and U18979 (N_18979,N_13041,N_13969);
or U18980 (N_18980,N_13807,N_13945);
xnor U18981 (N_18981,N_15513,N_14798);
and U18982 (N_18982,N_12303,N_12552);
nand U18983 (N_18983,N_15387,N_15050);
nand U18984 (N_18984,N_15047,N_15748);
or U18985 (N_18985,N_15010,N_14053);
nor U18986 (N_18986,N_15897,N_12634);
nand U18987 (N_18987,N_12108,N_15057);
or U18988 (N_18988,N_12465,N_12452);
and U18989 (N_18989,N_14407,N_12693);
nand U18990 (N_18990,N_12223,N_12827);
xor U18991 (N_18991,N_15476,N_13009);
nor U18992 (N_18992,N_15680,N_13323);
xor U18993 (N_18993,N_14654,N_12907);
nor U18994 (N_18994,N_13246,N_13700);
or U18995 (N_18995,N_15826,N_13863);
xnor U18996 (N_18996,N_14361,N_12398);
or U18997 (N_18997,N_15352,N_13893);
nor U18998 (N_18998,N_12529,N_13068);
nor U18999 (N_18999,N_12962,N_12279);
and U19000 (N_19000,N_14173,N_13428);
and U19001 (N_19001,N_15329,N_12707);
or U19002 (N_19002,N_15267,N_12145);
or U19003 (N_19003,N_13708,N_15171);
nor U19004 (N_19004,N_15814,N_12886);
nand U19005 (N_19005,N_15590,N_15218);
or U19006 (N_19006,N_12941,N_12190);
nor U19007 (N_19007,N_12775,N_12037);
nand U19008 (N_19008,N_15766,N_13401);
nand U19009 (N_19009,N_15586,N_13816);
and U19010 (N_19010,N_12128,N_13085);
or U19011 (N_19011,N_15613,N_13298);
xor U19012 (N_19012,N_14169,N_13919);
or U19013 (N_19013,N_13669,N_13430);
nor U19014 (N_19014,N_13043,N_15422);
or U19015 (N_19015,N_13039,N_14658);
or U19016 (N_19016,N_14460,N_12765);
and U19017 (N_19017,N_13172,N_15700);
nor U19018 (N_19018,N_13934,N_14199);
nor U19019 (N_19019,N_13058,N_15798);
nor U19020 (N_19020,N_12401,N_15779);
nand U19021 (N_19021,N_12075,N_14124);
xnor U19022 (N_19022,N_13921,N_13699);
nand U19023 (N_19023,N_12205,N_13520);
nor U19024 (N_19024,N_12888,N_13045);
or U19025 (N_19025,N_14408,N_13331);
nand U19026 (N_19026,N_14100,N_13613);
or U19027 (N_19027,N_15400,N_14195);
or U19028 (N_19028,N_13804,N_13995);
or U19029 (N_19029,N_14489,N_13471);
or U19030 (N_19030,N_14718,N_12624);
or U19031 (N_19031,N_13958,N_15453);
nand U19032 (N_19032,N_14943,N_13777);
and U19033 (N_19033,N_15465,N_13182);
nor U19034 (N_19034,N_15517,N_15453);
or U19035 (N_19035,N_12758,N_12788);
nor U19036 (N_19036,N_15432,N_12777);
nor U19037 (N_19037,N_13769,N_12324);
nor U19038 (N_19038,N_13929,N_15531);
nand U19039 (N_19039,N_14271,N_14929);
and U19040 (N_19040,N_12201,N_13786);
nor U19041 (N_19041,N_13490,N_13317);
nand U19042 (N_19042,N_15879,N_15288);
and U19043 (N_19043,N_15648,N_14757);
and U19044 (N_19044,N_12669,N_12535);
xor U19045 (N_19045,N_15992,N_13329);
nand U19046 (N_19046,N_12645,N_14938);
or U19047 (N_19047,N_12579,N_13927);
nor U19048 (N_19048,N_14362,N_13468);
xor U19049 (N_19049,N_12492,N_12572);
or U19050 (N_19050,N_13068,N_15225);
nand U19051 (N_19051,N_14413,N_12953);
and U19052 (N_19052,N_12231,N_14582);
nand U19053 (N_19053,N_15713,N_12339);
nor U19054 (N_19054,N_14875,N_15576);
and U19055 (N_19055,N_13887,N_12925);
or U19056 (N_19056,N_15021,N_14236);
xor U19057 (N_19057,N_15967,N_15459);
nor U19058 (N_19058,N_15392,N_13865);
and U19059 (N_19059,N_12668,N_14511);
nor U19060 (N_19060,N_15924,N_13870);
nand U19061 (N_19061,N_14777,N_12508);
nor U19062 (N_19062,N_15050,N_15078);
or U19063 (N_19063,N_13131,N_15060);
and U19064 (N_19064,N_14579,N_14518);
or U19065 (N_19065,N_12459,N_12350);
and U19066 (N_19066,N_15901,N_12011);
xor U19067 (N_19067,N_15611,N_13206);
or U19068 (N_19068,N_13449,N_15583);
and U19069 (N_19069,N_13683,N_12557);
nand U19070 (N_19070,N_13888,N_13002);
or U19071 (N_19071,N_13076,N_15117);
or U19072 (N_19072,N_13884,N_15566);
nor U19073 (N_19073,N_13296,N_15454);
or U19074 (N_19074,N_12467,N_14632);
or U19075 (N_19075,N_15200,N_15484);
nand U19076 (N_19076,N_13862,N_14277);
nand U19077 (N_19077,N_14108,N_15113);
xnor U19078 (N_19078,N_13827,N_13006);
nand U19079 (N_19079,N_15777,N_15614);
and U19080 (N_19080,N_12282,N_15997);
nor U19081 (N_19081,N_12724,N_14908);
and U19082 (N_19082,N_14840,N_14726);
nand U19083 (N_19083,N_12041,N_13941);
and U19084 (N_19084,N_14887,N_14941);
nand U19085 (N_19085,N_15262,N_14091);
or U19086 (N_19086,N_15959,N_14691);
or U19087 (N_19087,N_15807,N_13048);
nand U19088 (N_19088,N_13407,N_13955);
nor U19089 (N_19089,N_12660,N_15735);
or U19090 (N_19090,N_12189,N_13699);
and U19091 (N_19091,N_12825,N_15746);
nand U19092 (N_19092,N_12461,N_12843);
and U19093 (N_19093,N_15667,N_12015);
nor U19094 (N_19094,N_15199,N_12511);
nand U19095 (N_19095,N_15934,N_14377);
or U19096 (N_19096,N_14584,N_15948);
and U19097 (N_19097,N_13545,N_14133);
nor U19098 (N_19098,N_12466,N_14941);
nand U19099 (N_19099,N_15398,N_15271);
and U19100 (N_19100,N_14883,N_15260);
or U19101 (N_19101,N_15637,N_13911);
nor U19102 (N_19102,N_14838,N_13711);
or U19103 (N_19103,N_15393,N_14952);
and U19104 (N_19104,N_15478,N_12689);
nand U19105 (N_19105,N_13568,N_15742);
nor U19106 (N_19106,N_13658,N_12997);
nand U19107 (N_19107,N_14400,N_15254);
or U19108 (N_19108,N_14274,N_12632);
nand U19109 (N_19109,N_13898,N_14373);
or U19110 (N_19110,N_14567,N_12156);
and U19111 (N_19111,N_14703,N_15637);
nand U19112 (N_19112,N_13819,N_14123);
and U19113 (N_19113,N_14484,N_12299);
and U19114 (N_19114,N_13558,N_12835);
nand U19115 (N_19115,N_13791,N_13957);
and U19116 (N_19116,N_15335,N_13927);
nor U19117 (N_19117,N_12290,N_14318);
and U19118 (N_19118,N_13842,N_12584);
nand U19119 (N_19119,N_14519,N_13379);
or U19120 (N_19120,N_14678,N_14537);
or U19121 (N_19121,N_14956,N_12871);
xnor U19122 (N_19122,N_12448,N_12248);
and U19123 (N_19123,N_15100,N_13658);
nor U19124 (N_19124,N_13184,N_13010);
and U19125 (N_19125,N_14993,N_13165);
or U19126 (N_19126,N_15410,N_13763);
and U19127 (N_19127,N_15294,N_13016);
nand U19128 (N_19128,N_14212,N_12439);
nor U19129 (N_19129,N_15047,N_12856);
nor U19130 (N_19130,N_15786,N_13389);
nand U19131 (N_19131,N_12635,N_15267);
nand U19132 (N_19132,N_12661,N_13306);
nand U19133 (N_19133,N_15160,N_13795);
or U19134 (N_19134,N_13483,N_12551);
and U19135 (N_19135,N_13017,N_12177);
xor U19136 (N_19136,N_13524,N_14053);
nor U19137 (N_19137,N_14534,N_14171);
nor U19138 (N_19138,N_13281,N_15845);
nor U19139 (N_19139,N_12283,N_13817);
and U19140 (N_19140,N_15149,N_12196);
nor U19141 (N_19141,N_15765,N_15434);
nor U19142 (N_19142,N_12560,N_12344);
nand U19143 (N_19143,N_12952,N_14626);
nand U19144 (N_19144,N_12490,N_12272);
nor U19145 (N_19145,N_14600,N_13145);
or U19146 (N_19146,N_13234,N_15327);
and U19147 (N_19147,N_14533,N_13878);
xnor U19148 (N_19148,N_15629,N_13097);
nor U19149 (N_19149,N_14070,N_15386);
and U19150 (N_19150,N_13589,N_15010);
and U19151 (N_19151,N_13906,N_12744);
nand U19152 (N_19152,N_14065,N_14655);
nor U19153 (N_19153,N_13608,N_12467);
nor U19154 (N_19154,N_14049,N_12991);
or U19155 (N_19155,N_13539,N_12637);
and U19156 (N_19156,N_12095,N_12300);
nor U19157 (N_19157,N_13048,N_12133);
xnor U19158 (N_19158,N_15788,N_15998);
and U19159 (N_19159,N_12079,N_14951);
nor U19160 (N_19160,N_15904,N_14033);
or U19161 (N_19161,N_15817,N_15828);
nor U19162 (N_19162,N_12571,N_14273);
nor U19163 (N_19163,N_15255,N_13740);
or U19164 (N_19164,N_15011,N_14115);
or U19165 (N_19165,N_14913,N_14025);
and U19166 (N_19166,N_13884,N_15016);
or U19167 (N_19167,N_13837,N_14565);
nor U19168 (N_19168,N_12977,N_15618);
or U19169 (N_19169,N_13152,N_15092);
nand U19170 (N_19170,N_13139,N_15278);
or U19171 (N_19171,N_14389,N_12786);
nand U19172 (N_19172,N_13394,N_13379);
and U19173 (N_19173,N_14088,N_15657);
nor U19174 (N_19174,N_15315,N_13903);
nand U19175 (N_19175,N_15778,N_12862);
nand U19176 (N_19176,N_15271,N_15284);
and U19177 (N_19177,N_14445,N_13962);
or U19178 (N_19178,N_15687,N_13191);
nand U19179 (N_19179,N_14005,N_15464);
xor U19180 (N_19180,N_12604,N_15402);
nand U19181 (N_19181,N_15616,N_13238);
and U19182 (N_19182,N_12155,N_13721);
nand U19183 (N_19183,N_15491,N_15908);
xor U19184 (N_19184,N_14527,N_14932);
nand U19185 (N_19185,N_14996,N_13659);
nor U19186 (N_19186,N_15055,N_14719);
and U19187 (N_19187,N_13614,N_12938);
nand U19188 (N_19188,N_14881,N_13738);
and U19189 (N_19189,N_13384,N_15347);
or U19190 (N_19190,N_13043,N_13846);
and U19191 (N_19191,N_12442,N_14432);
and U19192 (N_19192,N_12970,N_13127);
nor U19193 (N_19193,N_14367,N_12346);
or U19194 (N_19194,N_13329,N_15387);
and U19195 (N_19195,N_12169,N_14878);
nand U19196 (N_19196,N_14853,N_14163);
nand U19197 (N_19197,N_15612,N_12488);
or U19198 (N_19198,N_15302,N_12465);
or U19199 (N_19199,N_14647,N_15630);
and U19200 (N_19200,N_15904,N_12621);
and U19201 (N_19201,N_15741,N_12162);
xor U19202 (N_19202,N_12752,N_15710);
nor U19203 (N_19203,N_12676,N_12228);
nor U19204 (N_19204,N_15068,N_15014);
or U19205 (N_19205,N_13155,N_14159);
nor U19206 (N_19206,N_15760,N_12003);
nand U19207 (N_19207,N_12247,N_12837);
and U19208 (N_19208,N_12231,N_12525);
and U19209 (N_19209,N_15258,N_12815);
or U19210 (N_19210,N_13682,N_14097);
nor U19211 (N_19211,N_13289,N_13969);
nand U19212 (N_19212,N_12735,N_13762);
nand U19213 (N_19213,N_15433,N_12458);
and U19214 (N_19214,N_14596,N_12902);
nor U19215 (N_19215,N_12846,N_13057);
or U19216 (N_19216,N_14667,N_12697);
nand U19217 (N_19217,N_14886,N_13501);
nor U19218 (N_19218,N_14023,N_15567);
and U19219 (N_19219,N_14686,N_13639);
nand U19220 (N_19220,N_13088,N_12096);
and U19221 (N_19221,N_14043,N_14458);
nor U19222 (N_19222,N_14659,N_15974);
and U19223 (N_19223,N_15161,N_15961);
nor U19224 (N_19224,N_15006,N_14317);
and U19225 (N_19225,N_15312,N_14157);
nor U19226 (N_19226,N_14802,N_13440);
nor U19227 (N_19227,N_14258,N_12516);
or U19228 (N_19228,N_12958,N_12837);
xor U19229 (N_19229,N_14067,N_15335);
nor U19230 (N_19230,N_15874,N_12149);
nor U19231 (N_19231,N_14682,N_15950);
nand U19232 (N_19232,N_12571,N_15457);
xnor U19233 (N_19233,N_14733,N_14857);
nand U19234 (N_19234,N_14971,N_13079);
or U19235 (N_19235,N_14896,N_12933);
nand U19236 (N_19236,N_14617,N_13288);
and U19237 (N_19237,N_13669,N_13987);
xnor U19238 (N_19238,N_15359,N_14881);
and U19239 (N_19239,N_12361,N_15406);
and U19240 (N_19240,N_15878,N_12052);
or U19241 (N_19241,N_14468,N_13967);
nor U19242 (N_19242,N_15737,N_15440);
and U19243 (N_19243,N_15497,N_12424);
nand U19244 (N_19244,N_12435,N_15975);
and U19245 (N_19245,N_15960,N_15151);
nor U19246 (N_19246,N_15395,N_13958);
nor U19247 (N_19247,N_12064,N_14561);
xor U19248 (N_19248,N_15067,N_13628);
nand U19249 (N_19249,N_13817,N_13793);
or U19250 (N_19250,N_12182,N_12267);
or U19251 (N_19251,N_14489,N_13959);
nor U19252 (N_19252,N_15799,N_12312);
xor U19253 (N_19253,N_13153,N_15615);
nor U19254 (N_19254,N_15338,N_15207);
nor U19255 (N_19255,N_15767,N_12684);
or U19256 (N_19256,N_15878,N_12674);
or U19257 (N_19257,N_15676,N_12636);
nor U19258 (N_19258,N_13818,N_12813);
or U19259 (N_19259,N_14209,N_12364);
nor U19260 (N_19260,N_12278,N_13969);
nand U19261 (N_19261,N_12792,N_15160);
and U19262 (N_19262,N_12184,N_12253);
nor U19263 (N_19263,N_15976,N_12193);
or U19264 (N_19264,N_15262,N_13874);
and U19265 (N_19265,N_13119,N_12552);
nand U19266 (N_19266,N_13103,N_13517);
and U19267 (N_19267,N_12406,N_13938);
and U19268 (N_19268,N_14675,N_12679);
and U19269 (N_19269,N_13159,N_14874);
nand U19270 (N_19270,N_12568,N_15459);
xor U19271 (N_19271,N_14184,N_14148);
or U19272 (N_19272,N_15214,N_13246);
or U19273 (N_19273,N_12705,N_13552);
nand U19274 (N_19274,N_14111,N_14429);
or U19275 (N_19275,N_15873,N_14942);
nand U19276 (N_19276,N_14426,N_13471);
or U19277 (N_19277,N_14320,N_12167);
nor U19278 (N_19278,N_12714,N_12548);
or U19279 (N_19279,N_14693,N_12925);
nor U19280 (N_19280,N_13052,N_15881);
or U19281 (N_19281,N_12298,N_12071);
or U19282 (N_19282,N_14103,N_15219);
nand U19283 (N_19283,N_12315,N_15514);
and U19284 (N_19284,N_12230,N_13517);
nor U19285 (N_19285,N_13905,N_13065);
nand U19286 (N_19286,N_15796,N_13764);
xnor U19287 (N_19287,N_15941,N_14123);
and U19288 (N_19288,N_15000,N_13785);
and U19289 (N_19289,N_15059,N_12166);
and U19290 (N_19290,N_13851,N_12287);
and U19291 (N_19291,N_15913,N_13105);
nor U19292 (N_19292,N_13519,N_12477);
nand U19293 (N_19293,N_14232,N_15499);
and U19294 (N_19294,N_12275,N_13727);
and U19295 (N_19295,N_13273,N_14620);
nand U19296 (N_19296,N_14507,N_14330);
or U19297 (N_19297,N_12575,N_14794);
or U19298 (N_19298,N_12469,N_13660);
or U19299 (N_19299,N_14320,N_15230);
nor U19300 (N_19300,N_15882,N_13398);
or U19301 (N_19301,N_14084,N_15232);
and U19302 (N_19302,N_15825,N_15149);
and U19303 (N_19303,N_15544,N_13067);
and U19304 (N_19304,N_13070,N_14409);
nand U19305 (N_19305,N_14692,N_12327);
and U19306 (N_19306,N_12336,N_12570);
and U19307 (N_19307,N_12096,N_15242);
and U19308 (N_19308,N_15829,N_14662);
xnor U19309 (N_19309,N_13216,N_12422);
nand U19310 (N_19310,N_15598,N_15687);
or U19311 (N_19311,N_14447,N_13275);
nand U19312 (N_19312,N_15023,N_12758);
and U19313 (N_19313,N_15084,N_15388);
nand U19314 (N_19314,N_13030,N_13416);
or U19315 (N_19315,N_14900,N_15744);
nand U19316 (N_19316,N_15847,N_14350);
or U19317 (N_19317,N_15662,N_15699);
or U19318 (N_19318,N_14378,N_15570);
or U19319 (N_19319,N_12201,N_13486);
or U19320 (N_19320,N_13978,N_12640);
or U19321 (N_19321,N_15224,N_15965);
and U19322 (N_19322,N_13341,N_13180);
and U19323 (N_19323,N_15964,N_13744);
xor U19324 (N_19324,N_15525,N_15791);
nand U19325 (N_19325,N_15562,N_15688);
and U19326 (N_19326,N_12253,N_13422);
nor U19327 (N_19327,N_12885,N_13413);
nand U19328 (N_19328,N_15071,N_12752);
nand U19329 (N_19329,N_12132,N_13336);
xor U19330 (N_19330,N_14708,N_12815);
or U19331 (N_19331,N_12803,N_13578);
or U19332 (N_19332,N_15059,N_12680);
and U19333 (N_19333,N_14705,N_13116);
or U19334 (N_19334,N_15034,N_15294);
nand U19335 (N_19335,N_14960,N_12615);
nor U19336 (N_19336,N_13255,N_12009);
and U19337 (N_19337,N_15854,N_12286);
nor U19338 (N_19338,N_15052,N_15909);
xnor U19339 (N_19339,N_15937,N_15317);
xnor U19340 (N_19340,N_15580,N_13758);
and U19341 (N_19341,N_14867,N_13506);
or U19342 (N_19342,N_15190,N_14039);
nand U19343 (N_19343,N_14911,N_12761);
and U19344 (N_19344,N_13966,N_15439);
and U19345 (N_19345,N_13834,N_13138);
and U19346 (N_19346,N_15424,N_12018);
nor U19347 (N_19347,N_14915,N_14190);
and U19348 (N_19348,N_14599,N_15446);
and U19349 (N_19349,N_15453,N_12966);
and U19350 (N_19350,N_14151,N_15193);
and U19351 (N_19351,N_14294,N_15480);
or U19352 (N_19352,N_12331,N_13492);
and U19353 (N_19353,N_13104,N_12546);
nand U19354 (N_19354,N_13310,N_12484);
nor U19355 (N_19355,N_12116,N_14629);
nor U19356 (N_19356,N_13232,N_12441);
nand U19357 (N_19357,N_12123,N_14832);
nand U19358 (N_19358,N_13668,N_12860);
or U19359 (N_19359,N_15978,N_14959);
and U19360 (N_19360,N_13025,N_15989);
nand U19361 (N_19361,N_14025,N_15609);
nand U19362 (N_19362,N_15583,N_12896);
nor U19363 (N_19363,N_13030,N_14777);
and U19364 (N_19364,N_15343,N_15158);
nor U19365 (N_19365,N_13136,N_15794);
and U19366 (N_19366,N_12052,N_15642);
and U19367 (N_19367,N_12525,N_15422);
xnor U19368 (N_19368,N_15957,N_13538);
and U19369 (N_19369,N_15747,N_14149);
and U19370 (N_19370,N_13037,N_15098);
or U19371 (N_19371,N_13024,N_15505);
or U19372 (N_19372,N_15586,N_13019);
xnor U19373 (N_19373,N_13076,N_14937);
xnor U19374 (N_19374,N_14966,N_14727);
nand U19375 (N_19375,N_15686,N_13223);
nor U19376 (N_19376,N_13831,N_14936);
xnor U19377 (N_19377,N_15147,N_13304);
or U19378 (N_19378,N_15312,N_14306);
and U19379 (N_19379,N_13812,N_14664);
nand U19380 (N_19380,N_15960,N_12706);
or U19381 (N_19381,N_15903,N_13823);
nor U19382 (N_19382,N_13946,N_12722);
and U19383 (N_19383,N_13779,N_15068);
or U19384 (N_19384,N_12412,N_14408);
and U19385 (N_19385,N_12629,N_12785);
nor U19386 (N_19386,N_12877,N_14823);
or U19387 (N_19387,N_14420,N_13596);
and U19388 (N_19388,N_13995,N_14874);
and U19389 (N_19389,N_15919,N_12064);
or U19390 (N_19390,N_14398,N_13826);
nor U19391 (N_19391,N_12056,N_15383);
nor U19392 (N_19392,N_12128,N_13299);
or U19393 (N_19393,N_12546,N_13042);
xor U19394 (N_19394,N_12210,N_15382);
and U19395 (N_19395,N_13024,N_12589);
and U19396 (N_19396,N_14454,N_12623);
nor U19397 (N_19397,N_13406,N_12532);
nand U19398 (N_19398,N_15088,N_14580);
nor U19399 (N_19399,N_14570,N_13348);
nor U19400 (N_19400,N_15290,N_15924);
and U19401 (N_19401,N_12372,N_14225);
nor U19402 (N_19402,N_14696,N_12429);
nor U19403 (N_19403,N_14176,N_13297);
nand U19404 (N_19404,N_14277,N_14481);
nand U19405 (N_19405,N_14429,N_15402);
and U19406 (N_19406,N_13193,N_15046);
and U19407 (N_19407,N_12313,N_14931);
and U19408 (N_19408,N_15836,N_15441);
nor U19409 (N_19409,N_15859,N_12803);
or U19410 (N_19410,N_14258,N_12582);
and U19411 (N_19411,N_12075,N_12082);
or U19412 (N_19412,N_13484,N_14424);
and U19413 (N_19413,N_15402,N_13462);
nand U19414 (N_19414,N_15120,N_13436);
nand U19415 (N_19415,N_13287,N_13481);
nor U19416 (N_19416,N_15054,N_15948);
nand U19417 (N_19417,N_13824,N_13532);
xnor U19418 (N_19418,N_12749,N_12150);
nand U19419 (N_19419,N_15630,N_14887);
xor U19420 (N_19420,N_14468,N_12397);
nand U19421 (N_19421,N_12876,N_12252);
xnor U19422 (N_19422,N_15438,N_14566);
and U19423 (N_19423,N_15480,N_13387);
or U19424 (N_19424,N_13810,N_13198);
or U19425 (N_19425,N_12208,N_15375);
or U19426 (N_19426,N_14394,N_12885);
and U19427 (N_19427,N_14730,N_13384);
nor U19428 (N_19428,N_12808,N_12794);
xor U19429 (N_19429,N_13901,N_12127);
and U19430 (N_19430,N_15935,N_15488);
and U19431 (N_19431,N_13300,N_13678);
nand U19432 (N_19432,N_12044,N_12969);
and U19433 (N_19433,N_15677,N_14032);
xnor U19434 (N_19434,N_12971,N_14910);
nor U19435 (N_19435,N_15979,N_14132);
nor U19436 (N_19436,N_12667,N_15022);
xnor U19437 (N_19437,N_13144,N_15845);
nand U19438 (N_19438,N_13946,N_14244);
xor U19439 (N_19439,N_14634,N_13501);
or U19440 (N_19440,N_12008,N_13299);
nor U19441 (N_19441,N_14686,N_12511);
and U19442 (N_19442,N_13702,N_12912);
nand U19443 (N_19443,N_12911,N_12145);
or U19444 (N_19444,N_12375,N_14901);
nor U19445 (N_19445,N_13874,N_14267);
nand U19446 (N_19446,N_13200,N_15419);
and U19447 (N_19447,N_14441,N_15915);
and U19448 (N_19448,N_12393,N_13567);
xor U19449 (N_19449,N_14536,N_14936);
nor U19450 (N_19450,N_15324,N_14774);
or U19451 (N_19451,N_13822,N_13164);
nand U19452 (N_19452,N_14208,N_15946);
or U19453 (N_19453,N_15592,N_12583);
and U19454 (N_19454,N_15182,N_12321);
nor U19455 (N_19455,N_14195,N_13600);
nor U19456 (N_19456,N_14958,N_12020);
nor U19457 (N_19457,N_15313,N_15725);
nor U19458 (N_19458,N_14751,N_12552);
nand U19459 (N_19459,N_12750,N_13287);
nand U19460 (N_19460,N_12214,N_13230);
nor U19461 (N_19461,N_14210,N_14807);
nor U19462 (N_19462,N_15381,N_12058);
nor U19463 (N_19463,N_14348,N_13461);
nand U19464 (N_19464,N_14863,N_13019);
and U19465 (N_19465,N_15788,N_12045);
or U19466 (N_19466,N_12080,N_13982);
xnor U19467 (N_19467,N_14101,N_12666);
nor U19468 (N_19468,N_15648,N_15364);
nor U19469 (N_19469,N_12471,N_15828);
or U19470 (N_19470,N_15300,N_15308);
xnor U19471 (N_19471,N_15575,N_13357);
and U19472 (N_19472,N_13479,N_15688);
xnor U19473 (N_19473,N_14257,N_12178);
or U19474 (N_19474,N_13817,N_15482);
nor U19475 (N_19475,N_14012,N_14324);
and U19476 (N_19476,N_13368,N_13945);
or U19477 (N_19477,N_15167,N_12178);
nand U19478 (N_19478,N_13208,N_15412);
and U19479 (N_19479,N_15462,N_14474);
nand U19480 (N_19480,N_15195,N_14878);
and U19481 (N_19481,N_13721,N_13879);
or U19482 (N_19482,N_14375,N_15883);
or U19483 (N_19483,N_13587,N_15547);
nand U19484 (N_19484,N_12447,N_15234);
nand U19485 (N_19485,N_13911,N_14876);
nor U19486 (N_19486,N_12700,N_13422);
or U19487 (N_19487,N_14079,N_12466);
and U19488 (N_19488,N_13931,N_15475);
nor U19489 (N_19489,N_15499,N_13670);
and U19490 (N_19490,N_12206,N_14214);
and U19491 (N_19491,N_14268,N_15177);
and U19492 (N_19492,N_13499,N_15250);
xnor U19493 (N_19493,N_12558,N_15344);
nand U19494 (N_19494,N_13108,N_13454);
or U19495 (N_19495,N_14622,N_14160);
nand U19496 (N_19496,N_14811,N_13784);
nand U19497 (N_19497,N_13313,N_13003);
or U19498 (N_19498,N_13252,N_12600);
or U19499 (N_19499,N_13848,N_13369);
nand U19500 (N_19500,N_14213,N_15021);
and U19501 (N_19501,N_15380,N_15992);
or U19502 (N_19502,N_15038,N_15718);
or U19503 (N_19503,N_12584,N_14453);
nand U19504 (N_19504,N_14090,N_12047);
xor U19505 (N_19505,N_13984,N_15265);
and U19506 (N_19506,N_13830,N_12399);
or U19507 (N_19507,N_13227,N_14902);
xnor U19508 (N_19508,N_15555,N_12662);
nor U19509 (N_19509,N_14418,N_15379);
nand U19510 (N_19510,N_13855,N_12745);
and U19511 (N_19511,N_12890,N_13632);
and U19512 (N_19512,N_15924,N_13225);
nor U19513 (N_19513,N_13012,N_14712);
or U19514 (N_19514,N_12673,N_13254);
or U19515 (N_19515,N_13442,N_13679);
or U19516 (N_19516,N_12037,N_13204);
nand U19517 (N_19517,N_14159,N_15813);
nand U19518 (N_19518,N_13291,N_12569);
nor U19519 (N_19519,N_13038,N_14783);
nor U19520 (N_19520,N_14579,N_15829);
or U19521 (N_19521,N_12758,N_14976);
xnor U19522 (N_19522,N_15694,N_12795);
nand U19523 (N_19523,N_13772,N_14105);
nor U19524 (N_19524,N_13230,N_13492);
and U19525 (N_19525,N_15070,N_15054);
xor U19526 (N_19526,N_13533,N_14954);
and U19527 (N_19527,N_14547,N_14063);
nor U19528 (N_19528,N_13875,N_13546);
or U19529 (N_19529,N_15019,N_13373);
and U19530 (N_19530,N_13217,N_13928);
or U19531 (N_19531,N_12037,N_15330);
xor U19532 (N_19532,N_14839,N_12102);
and U19533 (N_19533,N_14058,N_12087);
nor U19534 (N_19534,N_12927,N_12219);
and U19535 (N_19535,N_14131,N_14203);
and U19536 (N_19536,N_13368,N_15119);
xor U19537 (N_19537,N_15499,N_12658);
nand U19538 (N_19538,N_14741,N_12590);
nor U19539 (N_19539,N_13458,N_12726);
nand U19540 (N_19540,N_14026,N_12713);
or U19541 (N_19541,N_14801,N_14749);
or U19542 (N_19542,N_14395,N_15620);
and U19543 (N_19543,N_14462,N_14496);
nand U19544 (N_19544,N_15260,N_12992);
or U19545 (N_19545,N_13281,N_12817);
and U19546 (N_19546,N_15870,N_12425);
or U19547 (N_19547,N_15716,N_14334);
or U19548 (N_19548,N_13171,N_13302);
or U19549 (N_19549,N_14071,N_13749);
nor U19550 (N_19550,N_15469,N_14169);
and U19551 (N_19551,N_12191,N_12286);
nor U19552 (N_19552,N_12482,N_15543);
nor U19553 (N_19553,N_12417,N_12579);
and U19554 (N_19554,N_12173,N_14119);
nor U19555 (N_19555,N_13675,N_12635);
xor U19556 (N_19556,N_14031,N_14666);
or U19557 (N_19557,N_15964,N_12676);
or U19558 (N_19558,N_15162,N_15973);
nor U19559 (N_19559,N_14601,N_13384);
nor U19560 (N_19560,N_12231,N_12400);
nand U19561 (N_19561,N_13227,N_15046);
and U19562 (N_19562,N_12791,N_15269);
nor U19563 (N_19563,N_15361,N_15796);
and U19564 (N_19564,N_12241,N_13314);
nand U19565 (N_19565,N_15057,N_14004);
nand U19566 (N_19566,N_14030,N_15452);
or U19567 (N_19567,N_15889,N_13078);
nand U19568 (N_19568,N_12734,N_12779);
and U19569 (N_19569,N_13229,N_12046);
and U19570 (N_19570,N_13586,N_15599);
xnor U19571 (N_19571,N_14122,N_15065);
nor U19572 (N_19572,N_13925,N_12786);
nand U19573 (N_19573,N_12159,N_13186);
and U19574 (N_19574,N_15372,N_14057);
or U19575 (N_19575,N_15429,N_14418);
nor U19576 (N_19576,N_13893,N_14606);
nand U19577 (N_19577,N_15803,N_12121);
nand U19578 (N_19578,N_15159,N_15408);
and U19579 (N_19579,N_13494,N_13868);
xnor U19580 (N_19580,N_13938,N_14668);
nor U19581 (N_19581,N_14531,N_15273);
nand U19582 (N_19582,N_13498,N_13504);
and U19583 (N_19583,N_12584,N_14644);
nor U19584 (N_19584,N_14060,N_15436);
nand U19585 (N_19585,N_14519,N_12595);
nand U19586 (N_19586,N_12333,N_13336);
nor U19587 (N_19587,N_14332,N_15491);
nor U19588 (N_19588,N_14785,N_13642);
nand U19589 (N_19589,N_14847,N_12950);
nand U19590 (N_19590,N_15757,N_14062);
or U19591 (N_19591,N_13525,N_12086);
nand U19592 (N_19592,N_14795,N_13985);
nor U19593 (N_19593,N_12248,N_14221);
nand U19594 (N_19594,N_13530,N_14558);
nand U19595 (N_19595,N_12623,N_15578);
and U19596 (N_19596,N_13003,N_13879);
nand U19597 (N_19597,N_12527,N_13903);
or U19598 (N_19598,N_12414,N_15188);
and U19599 (N_19599,N_14389,N_12962);
nor U19600 (N_19600,N_12527,N_15495);
and U19601 (N_19601,N_14373,N_15886);
and U19602 (N_19602,N_13403,N_12666);
nor U19603 (N_19603,N_14530,N_12272);
nand U19604 (N_19604,N_13166,N_12635);
nor U19605 (N_19605,N_13582,N_15031);
and U19606 (N_19606,N_15008,N_15426);
xor U19607 (N_19607,N_13042,N_13720);
and U19608 (N_19608,N_13151,N_15904);
and U19609 (N_19609,N_13747,N_13652);
and U19610 (N_19610,N_15441,N_13129);
xnor U19611 (N_19611,N_12524,N_14618);
nor U19612 (N_19612,N_13758,N_15032);
xnor U19613 (N_19613,N_13400,N_13752);
or U19614 (N_19614,N_15265,N_14192);
nand U19615 (N_19615,N_14942,N_12210);
nor U19616 (N_19616,N_15553,N_13463);
nor U19617 (N_19617,N_15234,N_13514);
nand U19618 (N_19618,N_15901,N_13845);
and U19619 (N_19619,N_15169,N_13548);
nor U19620 (N_19620,N_12096,N_15772);
nand U19621 (N_19621,N_12139,N_14847);
or U19622 (N_19622,N_13894,N_13009);
xor U19623 (N_19623,N_12738,N_12991);
or U19624 (N_19624,N_15067,N_13613);
nand U19625 (N_19625,N_14287,N_15201);
or U19626 (N_19626,N_12998,N_12046);
and U19627 (N_19627,N_14676,N_15173);
nand U19628 (N_19628,N_12049,N_15702);
and U19629 (N_19629,N_13765,N_13617);
nand U19630 (N_19630,N_12709,N_12400);
nand U19631 (N_19631,N_13093,N_15577);
nand U19632 (N_19632,N_15716,N_14063);
and U19633 (N_19633,N_15951,N_12563);
nor U19634 (N_19634,N_14733,N_12198);
and U19635 (N_19635,N_13659,N_15656);
and U19636 (N_19636,N_12251,N_13618);
nand U19637 (N_19637,N_13098,N_15660);
nor U19638 (N_19638,N_12394,N_12686);
nor U19639 (N_19639,N_14160,N_13483);
nand U19640 (N_19640,N_12387,N_13391);
or U19641 (N_19641,N_14669,N_14330);
nor U19642 (N_19642,N_13901,N_15056);
and U19643 (N_19643,N_12428,N_14482);
or U19644 (N_19644,N_13023,N_12536);
nand U19645 (N_19645,N_12115,N_14941);
nand U19646 (N_19646,N_13041,N_12376);
or U19647 (N_19647,N_14051,N_15861);
xor U19648 (N_19648,N_13879,N_13183);
nor U19649 (N_19649,N_15510,N_15802);
xnor U19650 (N_19650,N_14379,N_15925);
or U19651 (N_19651,N_15678,N_15150);
nand U19652 (N_19652,N_12166,N_13684);
nor U19653 (N_19653,N_13589,N_14957);
and U19654 (N_19654,N_14564,N_12802);
and U19655 (N_19655,N_14217,N_12167);
nand U19656 (N_19656,N_14125,N_15840);
or U19657 (N_19657,N_12302,N_12993);
or U19658 (N_19658,N_13221,N_13156);
nand U19659 (N_19659,N_12123,N_15369);
xnor U19660 (N_19660,N_12135,N_14077);
nor U19661 (N_19661,N_15693,N_14058);
and U19662 (N_19662,N_15578,N_12842);
nor U19663 (N_19663,N_14846,N_15341);
nor U19664 (N_19664,N_14724,N_13441);
nor U19665 (N_19665,N_15218,N_15362);
nor U19666 (N_19666,N_14851,N_14536);
xnor U19667 (N_19667,N_13243,N_12775);
nor U19668 (N_19668,N_13915,N_13413);
or U19669 (N_19669,N_13372,N_13562);
or U19670 (N_19670,N_14739,N_12463);
xor U19671 (N_19671,N_12175,N_15056);
xnor U19672 (N_19672,N_14582,N_12029);
or U19673 (N_19673,N_13355,N_14878);
and U19674 (N_19674,N_15945,N_14329);
and U19675 (N_19675,N_14576,N_14480);
or U19676 (N_19676,N_14521,N_12500);
and U19677 (N_19677,N_12606,N_12566);
and U19678 (N_19678,N_14434,N_13150);
nor U19679 (N_19679,N_13859,N_13006);
and U19680 (N_19680,N_12526,N_14573);
and U19681 (N_19681,N_14981,N_14185);
or U19682 (N_19682,N_12668,N_13197);
nor U19683 (N_19683,N_12041,N_15021);
and U19684 (N_19684,N_12124,N_15751);
and U19685 (N_19685,N_12262,N_13904);
and U19686 (N_19686,N_13256,N_14366);
nand U19687 (N_19687,N_15382,N_14163);
nor U19688 (N_19688,N_15915,N_15334);
or U19689 (N_19689,N_12641,N_15353);
nor U19690 (N_19690,N_15373,N_13262);
and U19691 (N_19691,N_12957,N_13389);
nor U19692 (N_19692,N_13527,N_12962);
xor U19693 (N_19693,N_15035,N_15705);
or U19694 (N_19694,N_13861,N_12671);
and U19695 (N_19695,N_14968,N_14375);
nand U19696 (N_19696,N_15927,N_15263);
xor U19697 (N_19697,N_13598,N_13291);
nand U19698 (N_19698,N_14414,N_14141);
nor U19699 (N_19699,N_14799,N_12329);
nor U19700 (N_19700,N_13405,N_14346);
nand U19701 (N_19701,N_14454,N_12206);
or U19702 (N_19702,N_13768,N_12405);
or U19703 (N_19703,N_12675,N_12251);
nand U19704 (N_19704,N_14810,N_13653);
and U19705 (N_19705,N_14493,N_12659);
and U19706 (N_19706,N_15082,N_14009);
nor U19707 (N_19707,N_12803,N_14766);
nor U19708 (N_19708,N_14198,N_12762);
or U19709 (N_19709,N_15574,N_15270);
nand U19710 (N_19710,N_14341,N_15971);
xnor U19711 (N_19711,N_15249,N_15664);
nor U19712 (N_19712,N_15383,N_13658);
xor U19713 (N_19713,N_15991,N_12103);
or U19714 (N_19714,N_15794,N_15039);
or U19715 (N_19715,N_15413,N_13089);
nor U19716 (N_19716,N_15738,N_12614);
nor U19717 (N_19717,N_14057,N_15774);
nand U19718 (N_19718,N_13148,N_15175);
or U19719 (N_19719,N_14267,N_15128);
nand U19720 (N_19720,N_14739,N_13167);
or U19721 (N_19721,N_13124,N_14260);
and U19722 (N_19722,N_15489,N_13617);
nor U19723 (N_19723,N_15725,N_12407);
nor U19724 (N_19724,N_12835,N_15661);
or U19725 (N_19725,N_12992,N_12694);
nand U19726 (N_19726,N_13719,N_14334);
nor U19727 (N_19727,N_14314,N_13676);
nor U19728 (N_19728,N_13576,N_12354);
and U19729 (N_19729,N_13141,N_12909);
xor U19730 (N_19730,N_13538,N_13673);
xnor U19731 (N_19731,N_14147,N_12076);
and U19732 (N_19732,N_12697,N_14806);
nand U19733 (N_19733,N_15896,N_15537);
or U19734 (N_19734,N_12150,N_14420);
or U19735 (N_19735,N_14067,N_14408);
nand U19736 (N_19736,N_12372,N_13087);
nand U19737 (N_19737,N_14065,N_14473);
nor U19738 (N_19738,N_14412,N_12527);
nand U19739 (N_19739,N_13379,N_12400);
or U19740 (N_19740,N_14252,N_14571);
and U19741 (N_19741,N_15386,N_15764);
nand U19742 (N_19742,N_14553,N_14161);
nor U19743 (N_19743,N_13639,N_15455);
and U19744 (N_19744,N_15003,N_14982);
and U19745 (N_19745,N_15195,N_14438);
nand U19746 (N_19746,N_12595,N_14460);
nor U19747 (N_19747,N_13420,N_15403);
and U19748 (N_19748,N_14109,N_14015);
and U19749 (N_19749,N_15289,N_12592);
nand U19750 (N_19750,N_14673,N_12838);
and U19751 (N_19751,N_14210,N_14742);
nor U19752 (N_19752,N_15100,N_12102);
nor U19753 (N_19753,N_14160,N_13022);
or U19754 (N_19754,N_15496,N_14967);
nor U19755 (N_19755,N_12413,N_12231);
nor U19756 (N_19756,N_14573,N_13230);
or U19757 (N_19757,N_12263,N_14010);
nor U19758 (N_19758,N_12329,N_15834);
or U19759 (N_19759,N_15961,N_12986);
nand U19760 (N_19760,N_14734,N_15211);
nor U19761 (N_19761,N_15168,N_12221);
and U19762 (N_19762,N_13608,N_12827);
and U19763 (N_19763,N_14874,N_15248);
xnor U19764 (N_19764,N_15535,N_12704);
or U19765 (N_19765,N_15574,N_15036);
nand U19766 (N_19766,N_14754,N_15645);
xor U19767 (N_19767,N_14435,N_15941);
or U19768 (N_19768,N_12961,N_12697);
or U19769 (N_19769,N_15992,N_15278);
or U19770 (N_19770,N_15603,N_15677);
xnor U19771 (N_19771,N_13477,N_15162);
nand U19772 (N_19772,N_12044,N_14849);
and U19773 (N_19773,N_14259,N_14214);
nor U19774 (N_19774,N_13375,N_12780);
and U19775 (N_19775,N_14467,N_15067);
xor U19776 (N_19776,N_15769,N_12810);
or U19777 (N_19777,N_13908,N_12118);
nor U19778 (N_19778,N_12663,N_12156);
xnor U19779 (N_19779,N_12236,N_13209);
and U19780 (N_19780,N_14493,N_15258);
or U19781 (N_19781,N_15670,N_13847);
and U19782 (N_19782,N_14915,N_15235);
xor U19783 (N_19783,N_15490,N_13651);
nor U19784 (N_19784,N_15407,N_15433);
nand U19785 (N_19785,N_12556,N_13274);
nand U19786 (N_19786,N_13954,N_15172);
and U19787 (N_19787,N_15517,N_13668);
or U19788 (N_19788,N_15178,N_12181);
nor U19789 (N_19789,N_13493,N_14278);
nor U19790 (N_19790,N_15613,N_13358);
and U19791 (N_19791,N_15067,N_12069);
nor U19792 (N_19792,N_15722,N_14998);
and U19793 (N_19793,N_15593,N_12773);
xnor U19794 (N_19794,N_12226,N_13607);
and U19795 (N_19795,N_14335,N_12360);
nor U19796 (N_19796,N_14412,N_15856);
nand U19797 (N_19797,N_14641,N_12048);
or U19798 (N_19798,N_12839,N_12756);
xnor U19799 (N_19799,N_13030,N_14889);
nor U19800 (N_19800,N_13587,N_13200);
or U19801 (N_19801,N_15963,N_12582);
or U19802 (N_19802,N_14970,N_15637);
nand U19803 (N_19803,N_15673,N_13961);
or U19804 (N_19804,N_15151,N_12797);
nand U19805 (N_19805,N_12538,N_15130);
or U19806 (N_19806,N_13082,N_12310);
nor U19807 (N_19807,N_15019,N_14835);
xnor U19808 (N_19808,N_12915,N_12252);
nor U19809 (N_19809,N_12766,N_13747);
nor U19810 (N_19810,N_13263,N_13397);
nor U19811 (N_19811,N_14574,N_14225);
or U19812 (N_19812,N_12883,N_12334);
nand U19813 (N_19813,N_14551,N_13426);
or U19814 (N_19814,N_15588,N_14682);
and U19815 (N_19815,N_12956,N_14538);
nand U19816 (N_19816,N_15504,N_13360);
and U19817 (N_19817,N_13891,N_15528);
and U19818 (N_19818,N_14344,N_12942);
or U19819 (N_19819,N_14577,N_15449);
or U19820 (N_19820,N_13930,N_14090);
nand U19821 (N_19821,N_13886,N_13383);
or U19822 (N_19822,N_15990,N_15403);
nand U19823 (N_19823,N_13659,N_14421);
and U19824 (N_19824,N_14102,N_15865);
or U19825 (N_19825,N_13291,N_12065);
nor U19826 (N_19826,N_12339,N_14983);
or U19827 (N_19827,N_14066,N_15688);
nand U19828 (N_19828,N_13200,N_14531);
nand U19829 (N_19829,N_14287,N_12719);
nor U19830 (N_19830,N_14165,N_15591);
nand U19831 (N_19831,N_15275,N_12985);
and U19832 (N_19832,N_12948,N_12344);
or U19833 (N_19833,N_15140,N_13546);
nor U19834 (N_19834,N_13431,N_15222);
or U19835 (N_19835,N_13681,N_15453);
nor U19836 (N_19836,N_13080,N_14198);
xor U19837 (N_19837,N_15419,N_14169);
and U19838 (N_19838,N_13198,N_14613);
nor U19839 (N_19839,N_13855,N_14434);
nor U19840 (N_19840,N_15593,N_12930);
or U19841 (N_19841,N_14036,N_14620);
or U19842 (N_19842,N_15316,N_12229);
and U19843 (N_19843,N_13823,N_12115);
nor U19844 (N_19844,N_14058,N_12596);
or U19845 (N_19845,N_12074,N_14008);
and U19846 (N_19846,N_12694,N_14197);
and U19847 (N_19847,N_14480,N_15740);
or U19848 (N_19848,N_15980,N_12650);
nand U19849 (N_19849,N_15876,N_15308);
nand U19850 (N_19850,N_12216,N_15764);
or U19851 (N_19851,N_13053,N_13339);
nand U19852 (N_19852,N_13561,N_12039);
nand U19853 (N_19853,N_12983,N_13380);
nor U19854 (N_19854,N_12133,N_13412);
nand U19855 (N_19855,N_14730,N_15696);
nor U19856 (N_19856,N_13304,N_12127);
nor U19857 (N_19857,N_14322,N_14221);
and U19858 (N_19858,N_15882,N_14321);
nand U19859 (N_19859,N_12577,N_12554);
or U19860 (N_19860,N_13704,N_12071);
nand U19861 (N_19861,N_12390,N_15405);
nand U19862 (N_19862,N_12466,N_13371);
nor U19863 (N_19863,N_13373,N_14583);
and U19864 (N_19864,N_13791,N_15948);
and U19865 (N_19865,N_13623,N_14727);
and U19866 (N_19866,N_12551,N_14621);
nor U19867 (N_19867,N_14325,N_13154);
nor U19868 (N_19868,N_14148,N_12914);
xnor U19869 (N_19869,N_12767,N_13014);
nand U19870 (N_19870,N_13003,N_13037);
and U19871 (N_19871,N_13643,N_14823);
nor U19872 (N_19872,N_13342,N_15639);
xnor U19873 (N_19873,N_12648,N_15678);
nand U19874 (N_19874,N_14024,N_12914);
and U19875 (N_19875,N_15235,N_12799);
xnor U19876 (N_19876,N_12148,N_13686);
or U19877 (N_19877,N_14755,N_13919);
and U19878 (N_19878,N_12557,N_13686);
nand U19879 (N_19879,N_13205,N_13826);
and U19880 (N_19880,N_14116,N_12212);
nor U19881 (N_19881,N_13019,N_12612);
xor U19882 (N_19882,N_14239,N_12305);
nor U19883 (N_19883,N_13527,N_15102);
nor U19884 (N_19884,N_14168,N_12376);
and U19885 (N_19885,N_13351,N_12619);
xnor U19886 (N_19886,N_14283,N_12680);
nand U19887 (N_19887,N_14179,N_15818);
and U19888 (N_19888,N_12516,N_15843);
and U19889 (N_19889,N_13790,N_15132);
or U19890 (N_19890,N_15624,N_12416);
nor U19891 (N_19891,N_12190,N_14613);
or U19892 (N_19892,N_13182,N_13162);
nand U19893 (N_19893,N_14884,N_12893);
nor U19894 (N_19894,N_12286,N_15590);
nand U19895 (N_19895,N_14241,N_12366);
xnor U19896 (N_19896,N_15903,N_15876);
nand U19897 (N_19897,N_12207,N_14213);
nand U19898 (N_19898,N_15634,N_14562);
and U19899 (N_19899,N_13742,N_13164);
and U19900 (N_19900,N_13557,N_14364);
and U19901 (N_19901,N_12938,N_13131);
nor U19902 (N_19902,N_15943,N_14347);
nor U19903 (N_19903,N_12568,N_14598);
nor U19904 (N_19904,N_12790,N_14411);
or U19905 (N_19905,N_15501,N_14269);
nor U19906 (N_19906,N_14763,N_15938);
or U19907 (N_19907,N_12275,N_13257);
and U19908 (N_19908,N_13547,N_15059);
xnor U19909 (N_19909,N_13433,N_15478);
and U19910 (N_19910,N_12187,N_13842);
nand U19911 (N_19911,N_13486,N_15215);
or U19912 (N_19912,N_14691,N_13713);
nor U19913 (N_19913,N_13817,N_15771);
xnor U19914 (N_19914,N_14069,N_13716);
nand U19915 (N_19915,N_12153,N_13318);
or U19916 (N_19916,N_12706,N_12232);
nand U19917 (N_19917,N_13885,N_12144);
or U19918 (N_19918,N_15554,N_15408);
nor U19919 (N_19919,N_15772,N_15569);
xnor U19920 (N_19920,N_13724,N_15417);
nor U19921 (N_19921,N_15917,N_15942);
nor U19922 (N_19922,N_15382,N_12956);
nor U19923 (N_19923,N_15144,N_13391);
nand U19924 (N_19924,N_13506,N_14452);
nand U19925 (N_19925,N_14531,N_15711);
or U19926 (N_19926,N_13607,N_13203);
nor U19927 (N_19927,N_12311,N_15093);
and U19928 (N_19928,N_15208,N_12252);
or U19929 (N_19929,N_15327,N_13470);
or U19930 (N_19930,N_15310,N_14300);
and U19931 (N_19931,N_14259,N_13181);
nand U19932 (N_19932,N_12757,N_13050);
nand U19933 (N_19933,N_15884,N_14513);
or U19934 (N_19934,N_12197,N_13734);
or U19935 (N_19935,N_15171,N_12546);
nor U19936 (N_19936,N_15616,N_13468);
nor U19937 (N_19937,N_12129,N_12993);
nand U19938 (N_19938,N_12805,N_14874);
nand U19939 (N_19939,N_12938,N_14937);
nand U19940 (N_19940,N_13328,N_13125);
xor U19941 (N_19941,N_13419,N_13201);
and U19942 (N_19942,N_15714,N_14592);
nor U19943 (N_19943,N_12842,N_13240);
nand U19944 (N_19944,N_12900,N_14503);
and U19945 (N_19945,N_14058,N_12187);
or U19946 (N_19946,N_12921,N_14812);
xnor U19947 (N_19947,N_12417,N_13611);
nor U19948 (N_19948,N_13859,N_15973);
nor U19949 (N_19949,N_12334,N_15128);
and U19950 (N_19950,N_12689,N_14350);
or U19951 (N_19951,N_15454,N_12968);
nand U19952 (N_19952,N_12135,N_13098);
or U19953 (N_19953,N_12121,N_15615);
nand U19954 (N_19954,N_15641,N_13647);
or U19955 (N_19955,N_14438,N_12147);
and U19956 (N_19956,N_13231,N_12048);
nand U19957 (N_19957,N_13222,N_15972);
nor U19958 (N_19958,N_12808,N_12876);
and U19959 (N_19959,N_12842,N_13006);
or U19960 (N_19960,N_12947,N_12125);
nor U19961 (N_19961,N_12082,N_13536);
nand U19962 (N_19962,N_13729,N_14668);
nor U19963 (N_19963,N_13409,N_15728);
nand U19964 (N_19964,N_13050,N_12905);
or U19965 (N_19965,N_13201,N_15771);
or U19966 (N_19966,N_12721,N_15406);
and U19967 (N_19967,N_14369,N_13236);
and U19968 (N_19968,N_14995,N_14209);
or U19969 (N_19969,N_15158,N_12758);
and U19970 (N_19970,N_14773,N_14938);
nand U19971 (N_19971,N_12603,N_15295);
or U19972 (N_19972,N_13128,N_13415);
and U19973 (N_19973,N_15894,N_12813);
nand U19974 (N_19974,N_12341,N_13765);
and U19975 (N_19975,N_15635,N_14313);
or U19976 (N_19976,N_12002,N_13594);
nand U19977 (N_19977,N_12944,N_14548);
and U19978 (N_19978,N_13229,N_15795);
xnor U19979 (N_19979,N_14421,N_15725);
nand U19980 (N_19980,N_13813,N_13181);
nand U19981 (N_19981,N_13915,N_13021);
and U19982 (N_19982,N_15627,N_12516);
nand U19983 (N_19983,N_13854,N_15910);
nor U19984 (N_19984,N_13454,N_13621);
nand U19985 (N_19985,N_12508,N_13775);
and U19986 (N_19986,N_14948,N_14812);
or U19987 (N_19987,N_13054,N_13328);
or U19988 (N_19988,N_12646,N_15604);
nand U19989 (N_19989,N_13373,N_15852);
or U19990 (N_19990,N_15858,N_15282);
or U19991 (N_19991,N_13710,N_13469);
nor U19992 (N_19992,N_12549,N_14472);
nand U19993 (N_19993,N_12531,N_13705);
xnor U19994 (N_19994,N_15433,N_12605);
and U19995 (N_19995,N_14312,N_12840);
and U19996 (N_19996,N_14648,N_15097);
or U19997 (N_19997,N_15762,N_12127);
nor U19998 (N_19998,N_14648,N_14321);
nand U19999 (N_19999,N_12940,N_15045);
nor UO_0 (O_0,N_19158,N_16249);
xnor UO_1 (O_1,N_18864,N_19285);
and UO_2 (O_2,N_16560,N_19701);
or UO_3 (O_3,N_18507,N_16865);
nand UO_4 (O_4,N_16625,N_18474);
nand UO_5 (O_5,N_18367,N_17789);
nand UO_6 (O_6,N_16119,N_17103);
nand UO_7 (O_7,N_19626,N_19633);
nor UO_8 (O_8,N_17626,N_18301);
xor UO_9 (O_9,N_16878,N_16569);
and UO_10 (O_10,N_17247,N_16002);
nand UO_11 (O_11,N_16347,N_16449);
nand UO_12 (O_12,N_17479,N_17071);
or UO_13 (O_13,N_18799,N_16128);
and UO_14 (O_14,N_18838,N_16144);
nand UO_15 (O_15,N_19832,N_17457);
nor UO_16 (O_16,N_19241,N_18324);
nand UO_17 (O_17,N_17302,N_19900);
nor UO_18 (O_18,N_19096,N_18419);
nor UO_19 (O_19,N_19118,N_19151);
nand UO_20 (O_20,N_17577,N_18496);
nor UO_21 (O_21,N_17097,N_17051);
and UO_22 (O_22,N_17769,N_19177);
nor UO_23 (O_23,N_18498,N_18800);
nor UO_24 (O_24,N_17263,N_17284);
nand UO_25 (O_25,N_18738,N_17452);
nor UO_26 (O_26,N_16289,N_17370);
or UO_27 (O_27,N_19209,N_16621);
or UO_28 (O_28,N_16542,N_17440);
or UO_29 (O_29,N_17742,N_18717);
or UO_30 (O_30,N_16985,N_17035);
and UO_31 (O_31,N_19572,N_18068);
nand UO_32 (O_32,N_16054,N_17253);
or UO_33 (O_33,N_17733,N_16605);
nand UO_34 (O_34,N_18848,N_19875);
nand UO_35 (O_35,N_18416,N_17838);
and UO_36 (O_36,N_19051,N_18778);
xnor UO_37 (O_37,N_17488,N_18797);
nor UO_38 (O_38,N_18781,N_19665);
or UO_39 (O_39,N_17926,N_16643);
and UO_40 (O_40,N_19018,N_18779);
xnor UO_41 (O_41,N_16452,N_17456);
or UO_42 (O_42,N_19208,N_18308);
nor UO_43 (O_43,N_19358,N_16710);
xor UO_44 (O_44,N_19661,N_18270);
nor UO_45 (O_45,N_17857,N_19362);
or UO_46 (O_46,N_19270,N_18707);
and UO_47 (O_47,N_19152,N_18047);
xnor UO_48 (O_48,N_17165,N_17984);
xor UO_49 (O_49,N_19444,N_17996);
or UO_50 (O_50,N_18501,N_18348);
xor UO_51 (O_51,N_16165,N_16889);
and UO_52 (O_52,N_18294,N_17311);
and UO_53 (O_53,N_17227,N_18318);
nor UO_54 (O_54,N_18244,N_18150);
nor UO_55 (O_55,N_19433,N_16359);
nor UO_56 (O_56,N_19120,N_18414);
nor UO_57 (O_57,N_17008,N_18229);
and UO_58 (O_58,N_18786,N_16918);
nor UO_59 (O_59,N_19602,N_19275);
and UO_60 (O_60,N_17204,N_16770);
or UO_61 (O_61,N_19332,N_18311);
nor UO_62 (O_62,N_16399,N_18876);
and UO_63 (O_63,N_16582,N_18508);
xor UO_64 (O_64,N_17972,N_19599);
and UO_65 (O_65,N_17959,N_19729);
nor UO_66 (O_66,N_18827,N_16803);
or UO_67 (O_67,N_18636,N_19485);
nand UO_68 (O_68,N_19329,N_18731);
nand UO_69 (O_69,N_18382,N_19594);
and UO_70 (O_70,N_16283,N_16725);
and UO_71 (O_71,N_17631,N_19727);
or UO_72 (O_72,N_16444,N_18943);
nand UO_73 (O_73,N_19569,N_18551);
xnor UO_74 (O_74,N_17320,N_16245);
nand UO_75 (O_75,N_18836,N_17380);
or UO_76 (O_76,N_18834,N_16323);
and UO_77 (O_77,N_18368,N_17872);
nor UO_78 (O_78,N_18028,N_18587);
xor UO_79 (O_79,N_17550,N_17669);
nor UO_80 (O_80,N_19743,N_19678);
and UO_81 (O_81,N_19793,N_19331);
and UO_82 (O_82,N_17219,N_18926);
or UO_83 (O_83,N_17995,N_18693);
nor UO_84 (O_84,N_18662,N_18049);
nand UO_85 (O_85,N_16425,N_18100);
nor UO_86 (O_86,N_16113,N_17105);
nor UO_87 (O_87,N_17389,N_16860);
nor UO_88 (O_88,N_17060,N_18486);
and UO_89 (O_89,N_19767,N_17407);
nor UO_90 (O_90,N_16873,N_18166);
xnor UO_91 (O_91,N_18725,N_18819);
and UO_92 (O_92,N_17798,N_19979);
and UO_93 (O_93,N_19595,N_16185);
nor UO_94 (O_94,N_16816,N_18437);
nor UO_95 (O_95,N_16975,N_19176);
or UO_96 (O_96,N_18614,N_17442);
or UO_97 (O_97,N_16440,N_19983);
xnor UO_98 (O_98,N_18652,N_18116);
nand UO_99 (O_99,N_17428,N_17334);
nor UO_100 (O_100,N_17907,N_17718);
or UO_101 (O_101,N_16965,N_16272);
or UO_102 (O_102,N_18616,N_19293);
and UO_103 (O_103,N_17726,N_17684);
or UO_104 (O_104,N_18787,N_19029);
xor UO_105 (O_105,N_17374,N_16535);
or UO_106 (O_106,N_16180,N_19932);
and UO_107 (O_107,N_18405,N_17941);
or UO_108 (O_108,N_17388,N_18897);
nand UO_109 (O_109,N_16726,N_16084);
or UO_110 (O_110,N_17013,N_16663);
nor UO_111 (O_111,N_18687,N_18042);
and UO_112 (O_112,N_18647,N_17496);
xor UO_113 (O_113,N_17490,N_16291);
nand UO_114 (O_114,N_16281,N_18243);
or UO_115 (O_115,N_17588,N_16368);
nor UO_116 (O_116,N_19415,N_16817);
nor UO_117 (O_117,N_16278,N_17056);
and UO_118 (O_118,N_18059,N_19135);
and UO_119 (O_119,N_18095,N_17888);
or UO_120 (O_120,N_17729,N_16942);
nor UO_121 (O_121,N_17537,N_19340);
nor UO_122 (O_122,N_19884,N_18670);
or UO_123 (O_123,N_19373,N_19348);
or UO_124 (O_124,N_18928,N_19837);
nor UO_125 (O_125,N_18205,N_18742);
nand UO_126 (O_126,N_17472,N_18122);
nor UO_127 (O_127,N_16624,N_18334);
or UO_128 (O_128,N_16495,N_17672);
nand UO_129 (O_129,N_17702,N_16932);
nand UO_130 (O_130,N_19654,N_16698);
and UO_131 (O_131,N_18126,N_18760);
nand UO_132 (O_132,N_19377,N_17079);
and UO_133 (O_133,N_19730,N_18162);
or UO_134 (O_134,N_17159,N_17854);
and UO_135 (O_135,N_19213,N_19774);
nor UO_136 (O_136,N_19137,N_18165);
or UO_137 (O_137,N_17983,N_17605);
nor UO_138 (O_138,N_19423,N_19820);
and UO_139 (O_139,N_18478,N_16530);
nor UO_140 (O_140,N_19612,N_19789);
or UO_141 (O_141,N_19577,N_18950);
nand UO_142 (O_142,N_16564,N_16718);
and UO_143 (O_143,N_18350,N_19080);
nand UO_144 (O_144,N_18255,N_16253);
nand UO_145 (O_145,N_18690,N_17503);
or UO_146 (O_146,N_18306,N_16265);
or UO_147 (O_147,N_16315,N_17691);
nand UO_148 (O_148,N_17713,N_19801);
or UO_149 (O_149,N_19148,N_19345);
or UO_150 (O_150,N_17083,N_16929);
xnor UO_151 (O_151,N_17226,N_17610);
nor UO_152 (O_152,N_16472,N_19311);
nor UO_153 (O_153,N_16102,N_19129);
nand UO_154 (O_154,N_17009,N_19788);
nand UO_155 (O_155,N_17814,N_18328);
and UO_156 (O_156,N_16051,N_19061);
or UO_157 (O_157,N_16752,N_16615);
and UO_158 (O_158,N_16438,N_16243);
nand UO_159 (O_159,N_19307,N_16334);
and UO_160 (O_160,N_16343,N_19698);
and UO_161 (O_161,N_16383,N_17775);
nor UO_162 (O_162,N_17340,N_16740);
nor UO_163 (O_163,N_19397,N_19508);
nand UO_164 (O_164,N_16971,N_17939);
xor UO_165 (O_165,N_16130,N_16749);
xor UO_166 (O_166,N_17618,N_18624);
xnor UO_167 (O_167,N_19295,N_18724);
nand UO_168 (O_168,N_17381,N_19927);
nand UO_169 (O_169,N_18104,N_17205);
nand UO_170 (O_170,N_19658,N_18139);
nand UO_171 (O_171,N_16757,N_19778);
and UO_172 (O_172,N_18345,N_16040);
and UO_173 (O_173,N_19326,N_19179);
nand UO_174 (O_174,N_17192,N_16261);
or UO_175 (O_175,N_16514,N_17583);
nor UO_176 (O_176,N_17045,N_16636);
and UO_177 (O_177,N_17700,N_16125);
and UO_178 (O_178,N_18626,N_17243);
nor UO_179 (O_179,N_19552,N_17870);
xnor UO_180 (O_180,N_19609,N_17938);
and UO_181 (O_181,N_19145,N_16973);
nand UO_182 (O_182,N_17770,N_18110);
nor UO_183 (O_183,N_16462,N_18279);
nand UO_184 (O_184,N_16471,N_17688);
nor UO_185 (O_185,N_18176,N_17287);
and UO_186 (O_186,N_16677,N_19799);
or UO_187 (O_187,N_16519,N_18247);
nand UO_188 (O_188,N_18506,N_16198);
or UO_189 (O_189,N_18022,N_18712);
nor UO_190 (O_190,N_19053,N_17874);
nand UO_191 (O_191,N_17494,N_16487);
nor UO_192 (O_192,N_18347,N_17540);
or UO_193 (O_193,N_16976,N_19556);
nand UO_194 (O_194,N_19903,N_19703);
nand UO_195 (O_195,N_19598,N_19160);
or UO_196 (O_196,N_18954,N_19705);
or UO_197 (O_197,N_16910,N_19227);
and UO_198 (O_198,N_19829,N_16745);
xor UO_199 (O_199,N_17753,N_16786);
or UO_200 (O_200,N_17741,N_18806);
or UO_201 (O_201,N_17375,N_17639);
nand UO_202 (O_202,N_19310,N_17063);
and UO_203 (O_203,N_18004,N_19839);
and UO_204 (O_204,N_16262,N_19041);
or UO_205 (O_205,N_17924,N_19000);
and UO_206 (O_206,N_18676,N_18874);
nand UO_207 (O_207,N_18917,N_18429);
and UO_208 (O_208,N_19605,N_17262);
nor UO_209 (O_209,N_19369,N_17911);
nand UO_210 (O_210,N_19621,N_17273);
nand UO_211 (O_211,N_18451,N_17749);
and UO_212 (O_212,N_17853,N_17687);
or UO_213 (O_213,N_18445,N_17366);
or UO_214 (O_214,N_17716,N_16466);
and UO_215 (O_215,N_17176,N_17963);
nand UO_216 (O_216,N_17365,N_16345);
nand UO_217 (O_217,N_17068,N_17889);
xor UO_218 (O_218,N_19221,N_19885);
nand UO_219 (O_219,N_17135,N_19722);
nor UO_220 (O_220,N_16016,N_19883);
and UO_221 (O_221,N_19054,N_19800);
and UO_222 (O_222,N_16023,N_18591);
nor UO_223 (O_223,N_16746,N_16826);
nor UO_224 (O_224,N_16191,N_19680);
and UO_225 (O_225,N_18715,N_19472);
nor UO_226 (O_226,N_17506,N_18525);
xor UO_227 (O_227,N_18239,N_19264);
nand UO_228 (O_228,N_17113,N_16576);
nor UO_229 (O_229,N_18517,N_17714);
nand UO_230 (O_230,N_16839,N_16407);
nand UO_231 (O_231,N_17585,N_16657);
nor UO_232 (O_232,N_17112,N_17128);
and UO_233 (O_233,N_19744,N_19697);
nand UO_234 (O_234,N_16126,N_17676);
and UO_235 (O_235,N_19850,N_17796);
nor UO_236 (O_236,N_18857,N_17852);
or UO_237 (O_237,N_16597,N_18567);
and UO_238 (O_238,N_18331,N_18955);
nand UO_239 (O_239,N_18759,N_19024);
nor UO_240 (O_240,N_16818,N_19125);
nor UO_241 (O_241,N_18089,N_19814);
or UO_242 (O_242,N_18035,N_18489);
nand UO_243 (O_243,N_19775,N_17947);
nand UO_244 (O_244,N_16465,N_19781);
or UO_245 (O_245,N_17044,N_19030);
nor UO_246 (O_246,N_17988,N_18342);
nor UO_247 (O_247,N_17104,N_19312);
and UO_248 (O_248,N_16606,N_16142);
xor UO_249 (O_249,N_16993,N_16790);
and UO_250 (O_250,N_18862,N_16488);
xor UO_251 (O_251,N_17777,N_16441);
and UO_252 (O_252,N_17125,N_19381);
xnor UO_253 (O_253,N_19649,N_19498);
nor UO_254 (O_254,N_16046,N_18684);
nor UO_255 (O_255,N_17269,N_18262);
nor UO_256 (O_256,N_16800,N_19905);
nand UO_257 (O_257,N_18958,N_19175);
nand UO_258 (O_258,N_16493,N_18488);
and UO_259 (O_259,N_16073,N_17280);
or UO_260 (O_260,N_16139,N_18106);
nand UO_261 (O_261,N_17146,N_18384);
or UO_262 (O_262,N_17359,N_16335);
nand UO_263 (O_263,N_16913,N_16526);
xor UO_264 (O_264,N_17221,N_19407);
and UO_265 (O_265,N_17845,N_16206);
nor UO_266 (O_266,N_19763,N_19032);
nand UO_267 (O_267,N_17134,N_16732);
or UO_268 (O_268,N_16111,N_18067);
nand UO_269 (O_269,N_17039,N_16647);
or UO_270 (O_270,N_18091,N_18401);
xor UO_271 (O_271,N_16987,N_16109);
nor UO_272 (O_272,N_18070,N_19197);
and UO_273 (O_273,N_17641,N_19773);
or UO_274 (O_274,N_16885,N_18949);
nor UO_275 (O_275,N_18322,N_19116);
xor UO_276 (O_276,N_19561,N_19233);
or UO_277 (O_277,N_16492,N_17519);
and UO_278 (O_278,N_17945,N_18282);
nor UO_279 (O_279,N_17520,N_19013);
and UO_280 (O_280,N_18169,N_18397);
or UO_281 (O_281,N_18372,N_16485);
and UO_282 (O_282,N_16851,N_17073);
and UO_283 (O_283,N_16618,N_18538);
nand UO_284 (O_284,N_19857,N_18642);
xor UO_285 (O_285,N_18018,N_17834);
or UO_286 (O_286,N_19622,N_18271);
nand UO_287 (O_287,N_16326,N_19823);
nor UO_288 (O_288,N_16446,N_19828);
or UO_289 (O_289,N_16812,N_19974);
and UO_290 (O_290,N_18983,N_17444);
or UO_291 (O_291,N_18516,N_16617);
nor UO_292 (O_292,N_17871,N_17075);
and UO_293 (O_293,N_18889,N_17617);
or UO_294 (O_294,N_17774,N_19404);
and UO_295 (O_295,N_17484,N_18537);
or UO_296 (O_296,N_16434,N_18867);
xnor UO_297 (O_297,N_18761,N_17378);
nand UO_298 (O_298,N_18096,N_16908);
nor UO_299 (O_299,N_18298,N_19019);
and UO_300 (O_300,N_17771,N_17634);
and UO_301 (O_301,N_17461,N_19826);
nand UO_302 (O_302,N_18952,N_18562);
and UO_303 (O_303,N_16925,N_19586);
nor UO_304 (O_304,N_17455,N_19431);
xor UO_305 (O_305,N_19287,N_18393);
nand UO_306 (O_306,N_18034,N_16711);
xnor UO_307 (O_307,N_18805,N_17504);
or UO_308 (O_308,N_18029,N_19593);
or UO_309 (O_309,N_16979,N_18792);
or UO_310 (O_310,N_18154,N_16859);
nor UO_311 (O_311,N_16413,N_16880);
nor UO_312 (O_312,N_19534,N_17492);
and UO_313 (O_313,N_16149,N_17913);
nor UO_314 (O_314,N_17252,N_18597);
nand UO_315 (O_315,N_17141,N_18979);
xnor UO_316 (O_316,N_19025,N_19476);
and UO_317 (O_317,N_19717,N_16687);
and UO_318 (O_318,N_16264,N_17629);
and UO_319 (O_319,N_17211,N_19716);
or UO_320 (O_320,N_19110,N_19704);
or UO_321 (O_321,N_16696,N_17998);
and UO_322 (O_322,N_19503,N_18924);
nor UO_323 (O_323,N_18132,N_17756);
and UO_324 (O_324,N_18568,N_17795);
nor UO_325 (O_325,N_19993,N_18638);
nand UO_326 (O_326,N_18973,N_17481);
nand UO_327 (O_327,N_16948,N_19478);
nand UO_328 (O_328,N_16280,N_19222);
nand UO_329 (O_329,N_16823,N_16090);
nand UO_330 (O_330,N_18346,N_16238);
nand UO_331 (O_331,N_17685,N_18961);
nand UO_332 (O_332,N_17002,N_19999);
or UO_333 (O_333,N_16954,N_19591);
and UO_334 (O_334,N_16435,N_19853);
nor UO_335 (O_335,N_19634,N_17489);
nand UO_336 (O_336,N_18084,N_16121);
nand UO_337 (O_337,N_19147,N_16117);
nor UO_338 (O_338,N_18518,N_16221);
and UO_339 (O_339,N_17076,N_18899);
nor UO_340 (O_340,N_17040,N_17215);
and UO_341 (O_341,N_16502,N_16694);
nor UO_342 (O_342,N_19298,N_17092);
nand UO_343 (O_343,N_19164,N_19418);
nand UO_344 (O_344,N_18152,N_18793);
or UO_345 (O_345,N_19925,N_19426);
xnor UO_346 (O_346,N_18815,N_19059);
and UO_347 (O_347,N_16209,N_18410);
or UO_348 (O_348,N_18672,N_19901);
and UO_349 (O_349,N_16496,N_17430);
nor UO_350 (O_350,N_18181,N_17164);
or UO_351 (O_351,N_17940,N_18151);
xor UO_352 (O_352,N_19261,N_16251);
or UO_353 (O_353,N_19170,N_16388);
xnor UO_354 (O_354,N_16066,N_19475);
nand UO_355 (O_355,N_17750,N_16020);
nor UO_356 (O_356,N_18957,N_17014);
or UO_357 (O_357,N_16374,N_16683);
nor UO_358 (O_358,N_16742,N_19746);
or UO_359 (O_359,N_18714,N_18594);
nor UO_360 (O_360,N_16436,N_18558);
or UO_361 (O_361,N_16995,N_18530);
nand UO_362 (O_362,N_19628,N_19607);
and UO_363 (O_363,N_17169,N_17338);
and UO_364 (O_364,N_16268,N_16713);
or UO_365 (O_365,N_18751,N_19088);
nand UO_366 (O_366,N_16120,N_17579);
xnor UO_367 (O_367,N_17446,N_17783);
and UO_368 (O_368,N_17415,N_18058);
and UO_369 (O_369,N_17978,N_16288);
and UO_370 (O_370,N_18077,N_16849);
and UO_371 (O_371,N_17544,N_18448);
xnor UO_372 (O_372,N_18967,N_19245);
and UO_373 (O_373,N_17353,N_17842);
and UO_374 (O_374,N_18275,N_17233);
nor UO_375 (O_375,N_17239,N_18012);
nor UO_376 (O_376,N_19317,N_18025);
or UO_377 (O_377,N_18556,N_17763);
and UO_378 (O_378,N_19127,N_17348);
and UO_379 (O_379,N_17564,N_18400);
and UO_380 (O_380,N_17342,N_17188);
and UO_381 (O_381,N_17127,N_16899);
xor UO_382 (O_382,N_18098,N_18916);
or UO_383 (O_383,N_16834,N_17326);
xnor UO_384 (O_384,N_16775,N_16587);
or UO_385 (O_385,N_16646,N_18884);
or UO_386 (O_386,N_17546,N_17249);
xor UO_387 (O_387,N_19747,N_17208);
or UO_388 (O_388,N_16609,N_16372);
nor UO_389 (O_389,N_17566,N_16701);
nand UO_390 (O_390,N_17130,N_19690);
and UO_391 (O_391,N_19985,N_19263);
or UO_392 (O_392,N_17080,N_19846);
nand UO_393 (O_393,N_18998,N_18253);
nand UO_394 (O_394,N_17106,N_17882);
nor UO_395 (O_395,N_16961,N_18774);
or UO_396 (O_396,N_17553,N_18103);
nor UO_397 (O_397,N_19872,N_18728);
or UO_398 (O_398,N_17024,N_17514);
nand UO_399 (O_399,N_19074,N_19702);
and UO_400 (O_400,N_17194,N_18390);
and UO_401 (O_401,N_18119,N_16919);
nor UO_402 (O_402,N_17663,N_18529);
or UO_403 (O_403,N_17897,N_18056);
nor UO_404 (O_404,N_19419,N_18906);
xor UO_405 (O_405,N_17666,N_18560);
nor UO_406 (O_406,N_19689,N_17581);
nand UO_407 (O_407,N_17516,N_17743);
and UO_408 (O_408,N_18911,N_18804);
or UO_409 (O_409,N_18063,N_19174);
nor UO_410 (O_410,N_18534,N_17168);
or UO_411 (O_411,N_18005,N_19083);
xor UO_412 (O_412,N_16468,N_16106);
and UO_413 (O_413,N_18688,N_19004);
or UO_414 (O_414,N_19517,N_19207);
nand UO_415 (O_415,N_17784,N_16457);
and UO_416 (O_416,N_16528,N_17074);
and UO_417 (O_417,N_19383,N_16916);
xor UO_418 (O_418,N_18031,N_18213);
nor UO_419 (O_419,N_18430,N_18544);
or UO_420 (O_420,N_16246,N_16369);
nor UO_421 (O_421,N_19856,N_16047);
or UO_422 (O_422,N_19893,N_18870);
nor UO_423 (O_423,N_16774,N_19869);
and UO_424 (O_424,N_17431,N_17406);
xor UO_425 (O_425,N_17896,N_17916);
or UO_426 (O_426,N_16274,N_18339);
nand UO_427 (O_427,N_18586,N_18226);
nor UO_428 (O_428,N_19867,N_19648);
or UO_429 (O_429,N_18183,N_17468);
nand UO_430 (O_430,N_19134,N_19573);
and UO_431 (O_431,N_16642,N_18953);
nand UO_432 (O_432,N_17471,N_17942);
or UO_433 (O_433,N_17856,N_18865);
and UO_434 (O_434,N_16341,N_17931);
and UO_435 (O_435,N_19646,N_18711);
and UO_436 (O_436,N_19835,N_19827);
nand UO_437 (O_437,N_16596,N_16884);
or UO_438 (O_438,N_19273,N_18993);
or UO_439 (O_439,N_16220,N_17329);
or UO_440 (O_440,N_19831,N_16789);
nand UO_441 (O_441,N_19277,N_18721);
nand UO_442 (O_442,N_18490,N_16358);
nand UO_443 (O_443,N_18745,N_18782);
nand UO_444 (O_444,N_17443,N_19522);
nand UO_445 (O_445,N_18613,N_19372);
or UO_446 (O_446,N_16909,N_18513);
nor UO_447 (O_447,N_16719,N_19566);
and UO_448 (O_448,N_17973,N_17628);
nor UO_449 (O_449,N_17936,N_16943);
or UO_450 (O_450,N_19073,N_19745);
or UO_451 (O_451,N_16478,N_19114);
xor UO_452 (O_452,N_18075,N_18605);
nand UO_453 (O_453,N_18686,N_18411);
and UO_454 (O_454,N_19555,N_19786);
and UO_455 (O_455,N_16787,N_18532);
nor UO_456 (O_456,N_16071,N_18637);
nor UO_457 (O_457,N_16805,N_17535);
nor UO_458 (O_458,N_18203,N_16946);
and UO_459 (O_459,N_18791,N_18369);
xnor UO_460 (O_460,N_16822,N_18065);
xnor UO_461 (O_461,N_17181,N_18976);
nor UO_462 (O_462,N_18024,N_19395);
or UO_463 (O_463,N_17392,N_17609);
nor UO_464 (O_464,N_18932,N_17066);
nor UO_465 (O_465,N_19008,N_19228);
nor UO_466 (O_466,N_16417,N_16339);
nor UO_467 (O_467,N_18447,N_19758);
or UO_468 (O_468,N_19851,N_17064);
nand UO_469 (O_469,N_18184,N_17421);
nand UO_470 (O_470,N_16771,N_19082);
nand UO_471 (O_471,N_16604,N_16765);
xor UO_472 (O_472,N_17571,N_19666);
nor UO_473 (O_473,N_16832,N_17653);
or UO_474 (O_474,N_18064,N_18258);
nand UO_475 (O_475,N_17679,N_19017);
or UO_476 (O_476,N_18069,N_16888);
nand UO_477 (O_477,N_17147,N_19313);
nand UO_478 (O_478,N_17331,N_17387);
nand UO_479 (O_479,N_17813,N_16567);
and UO_480 (O_480,N_16737,N_19194);
nor UO_481 (O_481,N_16392,N_17893);
and UO_482 (O_482,N_18736,N_17918);
xor UO_483 (O_483,N_19037,N_17025);
and UO_484 (O_484,N_18785,N_16328);
nand UO_485 (O_485,N_18853,N_18841);
or UO_486 (O_486,N_17382,N_17447);
nand UO_487 (O_487,N_19357,N_18832);
or UO_488 (O_488,N_16602,N_17861);
nor UO_489 (O_489,N_19050,N_18762);
nand UO_490 (O_490,N_18360,N_18375);
nor UO_491 (O_491,N_17118,N_19934);
nand UO_492 (O_492,N_17582,N_16458);
nor UO_493 (O_493,N_19842,N_18905);
or UO_494 (O_494,N_18991,N_17473);
nor UO_495 (O_495,N_16521,N_19971);
xnor UO_496 (O_496,N_16187,N_18595);
and UO_497 (O_497,N_17932,N_17279);
or UO_498 (O_498,N_18723,N_18765);
nand UO_499 (O_499,N_18702,N_19965);
and UO_500 (O_500,N_19204,N_16772);
or UO_501 (O_501,N_17881,N_17970);
or UO_502 (O_502,N_18222,N_17094);
xor UO_503 (O_503,N_19060,N_19283);
and UO_504 (O_504,N_18128,N_19530);
and UO_505 (O_505,N_17858,N_17425);
nand UO_506 (O_506,N_16639,N_18440);
and UO_507 (O_507,N_18461,N_19707);
and UO_508 (O_508,N_19520,N_17894);
or UO_509 (O_509,N_19764,N_17393);
and UO_510 (O_510,N_18289,N_19880);
and UO_511 (O_511,N_16669,N_17057);
nand UO_512 (O_512,N_18657,N_17745);
and UO_513 (O_513,N_17612,N_18284);
nand UO_514 (O_514,N_19765,N_17000);
nand UO_515 (O_515,N_16814,N_17336);
nor UO_516 (O_516,N_19972,N_17318);
nand UO_517 (O_517,N_19892,N_16385);
and UO_518 (O_518,N_16940,N_17558);
nand UO_519 (O_519,N_18078,N_19647);
or UO_520 (O_520,N_16927,N_17594);
nand UO_521 (O_521,N_19931,N_18391);
or UO_522 (O_522,N_19168,N_17797);
nor UO_523 (O_523,N_17424,N_19435);
and UO_524 (O_524,N_18775,N_18296);
nand UO_525 (O_525,N_18623,N_17562);
nor UO_526 (O_526,N_16777,N_17237);
xnor UO_527 (O_527,N_18649,N_19382);
and UO_528 (O_528,N_17816,N_19780);
xor UO_529 (O_529,N_18385,N_19045);
xnor UO_530 (O_530,N_17543,N_16555);
and UO_531 (O_531,N_19361,N_18548);
nand UO_532 (O_532,N_17645,N_19538);
and UO_533 (O_533,N_18663,N_19913);
xnor UO_534 (O_534,N_17037,N_17863);
nor UO_535 (O_535,N_17158,N_18123);
nor UO_536 (O_536,N_16858,N_17154);
and UO_537 (O_537,N_19521,N_18541);
nor UO_538 (O_538,N_19635,N_17532);
or UO_539 (O_539,N_18020,N_19940);
nand UO_540 (O_540,N_17156,N_18852);
nand UO_541 (O_541,N_17885,N_17717);
or UO_542 (O_542,N_18856,N_16003);
nor UO_543 (O_543,N_17004,N_17142);
xnor UO_544 (O_544,N_19367,N_16160);
and UO_545 (O_545,N_16515,N_16756);
or UO_546 (O_546,N_19091,N_18547);
and UO_547 (O_547,N_16312,N_17067);
nor UO_548 (O_548,N_18189,N_16522);
nor UO_549 (O_549,N_19007,N_16232);
nor UO_550 (O_550,N_18813,N_17719);
or UO_551 (O_551,N_16728,N_19093);
xor UO_552 (O_552,N_16296,N_16088);
or UO_553 (O_553,N_17747,N_17155);
nand UO_554 (O_554,N_17464,N_16184);
nor UO_555 (O_555,N_17943,N_16055);
nand UO_556 (O_556,N_16114,N_16082);
and UO_557 (O_557,N_16325,N_16785);
nand UO_558 (O_558,N_17873,N_19876);
nand UO_559 (O_559,N_17231,N_16034);
xor UO_560 (O_560,N_18842,N_19346);
nand UO_561 (O_561,N_18802,N_19334);
or UO_562 (O_562,N_19042,N_18520);
xor UO_563 (O_563,N_17399,N_19792);
nand UO_564 (O_564,N_19553,N_17144);
nor UO_565 (O_565,N_18272,N_18436);
and UO_566 (O_566,N_19784,N_17347);
or UO_567 (O_567,N_17659,N_17343);
and UO_568 (O_568,N_18732,N_19531);
xnor UO_569 (O_569,N_16766,N_18484);
or UO_570 (O_570,N_16536,N_16293);
nand UO_571 (O_571,N_17991,N_17735);
and UO_572 (O_572,N_16623,N_17174);
nand UO_573 (O_573,N_17058,N_19153);
nor UO_574 (O_574,N_18304,N_17912);
nor UO_575 (O_575,N_17500,N_16481);
xnor UO_576 (O_576,N_17149,N_18770);
xnor UO_577 (O_577,N_16835,N_18354);
or UO_578 (O_578,N_16124,N_19420);
and UO_579 (O_579,N_18434,N_19611);
nand UO_580 (O_580,N_18215,N_16147);
nor UO_581 (O_581,N_18333,N_17766);
nor UO_582 (O_582,N_19322,N_19429);
xor UO_583 (O_583,N_19664,N_18254);
and UO_584 (O_584,N_18564,N_18502);
or UO_585 (O_585,N_18001,N_17960);
nand UO_586 (O_586,N_18689,N_18892);
nor UO_587 (O_587,N_18596,N_19027);
and UO_588 (O_588,N_17886,N_16242);
or UO_589 (O_589,N_18195,N_16076);
and UO_590 (O_590,N_17109,N_16550);
nor UO_591 (O_591,N_16295,N_16870);
and UO_592 (O_592,N_18172,N_16753);
and UO_593 (O_593,N_19770,N_17319);
nor UO_594 (O_594,N_16037,N_16613);
and UO_595 (O_595,N_17171,N_16353);
or UO_596 (O_596,N_18669,N_19062);
nor UO_597 (O_597,N_17827,N_17678);
or UO_598 (O_598,N_16072,N_19741);
nor UO_599 (O_599,N_16287,N_19964);
or UO_600 (O_600,N_18780,N_18526);
nand UO_601 (O_601,N_17049,N_18608);
or UO_602 (O_602,N_17754,N_17361);
nand UO_603 (O_603,N_16360,N_19550);
or UO_604 (O_604,N_18415,N_17161);
xnor UO_605 (O_605,N_16162,N_19676);
nor UO_606 (O_606,N_19980,N_18901);
xor UO_607 (O_607,N_17216,N_19278);
nand UO_608 (O_608,N_17234,N_16650);
xnor UO_609 (O_609,N_19504,N_17048);
nand UO_610 (O_610,N_19406,N_18713);
nand UO_611 (O_611,N_19229,N_16336);
nand UO_612 (O_612,N_16720,N_17548);
nand UO_613 (O_613,N_17951,N_16827);
nand UO_614 (O_614,N_18090,N_16222);
or UO_615 (O_615,N_18177,N_17162);
nand UO_616 (O_616,N_16169,N_18468);
or UO_617 (O_617,N_19926,N_18288);
or UO_618 (O_618,N_18630,N_19484);
xor UO_619 (O_619,N_17725,N_16680);
and UO_620 (O_620,N_16565,N_17095);
nor UO_621 (O_621,N_18598,N_18896);
or UO_622 (O_622,N_18557,N_17887);
xor UO_623 (O_623,N_16299,N_16570);
nand UO_624 (O_624,N_16193,N_18045);
nor UO_625 (O_625,N_19824,N_16896);
nor UO_626 (O_626,N_16767,N_19071);
nand UO_627 (O_627,N_17712,N_17517);
or UO_628 (O_628,N_19706,N_19492);
or UO_629 (O_629,N_17209,N_17513);
nand UO_630 (O_630,N_16671,N_16951);
or UO_631 (O_631,N_16627,N_16506);
or UO_632 (O_632,N_19101,N_18148);
and UO_633 (O_633,N_19390,N_16897);
and UO_634 (O_634,N_19302,N_16539);
and UO_635 (O_635,N_16501,N_16007);
or UO_636 (O_636,N_17619,N_18061);
and UO_637 (O_637,N_16183,N_18622);
nand UO_638 (O_638,N_17903,N_19748);
or UO_639 (O_639,N_16996,N_17435);
nand UO_640 (O_640,N_19920,N_17855);
and UO_641 (O_641,N_17160,N_16430);
xnor UO_642 (O_642,N_16340,N_18620);
xor UO_643 (O_643,N_18499,N_16572);
and UO_644 (O_644,N_18720,N_19184);
and UO_645 (O_645,N_17622,N_17242);
and UO_646 (O_646,N_18160,N_17565);
and UO_647 (O_647,N_17989,N_17923);
nor UO_648 (O_648,N_16375,N_18164);
and UO_649 (O_649,N_18470,N_17175);
nor UO_650 (O_650,N_17385,N_16640);
nand UO_651 (O_651,N_17005,N_16806);
and UO_652 (O_652,N_18467,N_17414);
and UO_653 (O_653,N_18287,N_18477);
or UO_654 (O_654,N_16855,N_18011);
and UO_655 (O_655,N_19655,N_17790);
and UO_656 (O_656,N_16241,N_18175);
nor UO_657 (O_657,N_18017,N_19673);
nand UO_658 (O_658,N_18458,N_17070);
or UO_659 (O_659,N_18741,N_19585);
or UO_660 (O_660,N_18550,N_16074);
and UO_661 (O_661,N_16017,N_19247);
and UO_662 (O_662,N_17574,N_17371);
and UO_663 (O_663,N_18796,N_17578);
xnor UO_664 (O_664,N_19499,N_19637);
nor UO_665 (O_665,N_18041,N_19266);
xnor UO_666 (O_666,N_19438,N_17283);
xor UO_667 (O_667,N_19046,N_16783);
and UO_668 (O_668,N_18413,N_19015);
or UO_669 (O_669,N_18960,N_17757);
nand UO_670 (O_670,N_19379,N_16384);
or UO_671 (O_671,N_18540,N_17301);
nor UO_672 (O_672,N_19130,N_18163);
and UO_673 (O_673,N_18790,N_16304);
or UO_674 (O_674,N_19546,N_17650);
nand UO_675 (O_675,N_19216,N_16693);
and UO_676 (O_676,N_17426,N_19584);
or UO_677 (O_677,N_17081,N_19021);
and UO_678 (O_678,N_16891,N_16933);
xnor UO_679 (O_679,N_19186,N_16021);
or UO_680 (O_680,N_16874,N_19541);
or UO_681 (O_681,N_18383,N_18179);
nand UO_682 (O_682,N_17201,N_16028);
nand UO_683 (O_683,N_17990,N_18274);
nand UO_684 (O_684,N_19187,N_17975);
and UO_685 (O_685,N_17129,N_16380);
nor UO_686 (O_686,N_18773,N_19496);
and UO_687 (O_687,N_19465,N_18743);
xor UO_688 (O_688,N_19234,N_18465);
and UO_689 (O_689,N_16422,N_18431);
nor UO_690 (O_690,N_16705,N_16804);
and UO_691 (O_691,N_19335,N_17980);
nor UO_692 (O_692,N_17883,N_19422);
or UO_693 (O_693,N_17405,N_18648);
and UO_694 (O_694,N_17206,N_18404);
nor UO_695 (O_695,N_19643,N_18329);
and UO_696 (O_696,N_19106,N_17652);
or UO_697 (O_697,N_16105,N_17502);
xor UO_698 (O_698,N_16988,N_17633);
xor UO_699 (O_699,N_18040,N_19214);
nand UO_700 (O_700,N_16957,N_19280);
nand UO_701 (O_701,N_17281,N_16255);
and UO_702 (O_702,N_17222,N_18578);
xnor UO_703 (O_703,N_18996,N_18894);
nor UO_704 (O_704,N_17312,N_17439);
nor UO_705 (O_705,N_18153,N_18948);
or UO_706 (O_706,N_16371,N_19866);
and UO_707 (O_707,N_16654,N_19859);
and UO_708 (O_708,N_19590,N_16906);
and UO_709 (O_709,N_16553,N_18571);
and UO_710 (O_710,N_17110,N_16167);
nor UO_711 (O_711,N_19989,N_16059);
and UO_712 (O_712,N_19337,N_18417);
or UO_713 (O_713,N_16614,N_16136);
xor UO_714 (O_714,N_19645,N_17900);
nand UO_715 (O_715,N_19882,N_19617);
or UO_716 (O_716,N_19375,N_17656);
xnor UO_717 (O_717,N_19269,N_16216);
nand UO_718 (O_718,N_19239,N_17020);
nand UO_719 (O_719,N_19807,N_16202);
or UO_720 (O_720,N_18893,N_18300);
or UO_721 (O_721,N_16992,N_18994);
or UO_722 (O_722,N_17608,N_17396);
and UO_723 (O_723,N_17810,N_16426);
nand UO_724 (O_724,N_18625,N_18965);
or UO_725 (O_725,N_18186,N_19806);
xnor UO_726 (O_726,N_18555,N_18982);
nor UO_727 (O_727,N_17386,N_18086);
nand UO_728 (O_728,N_19563,N_17522);
or UO_729 (O_729,N_18006,N_19448);
and UO_730 (O_730,N_17841,N_19172);
xor UO_731 (O_731,N_16402,N_18319);
nor UO_732 (O_732,N_16791,N_16205);
and UO_733 (O_733,N_17925,N_18820);
and UO_734 (O_734,N_18497,N_18698);
or UO_735 (O_735,N_16780,N_16537);
or UO_736 (O_736,N_18977,N_17189);
or UO_737 (O_737,N_19115,N_18561);
xor UO_738 (O_738,N_18811,N_17835);
nor UO_739 (O_739,N_16256,N_17974);
nand UO_740 (O_740,N_17898,N_18536);
and UO_741 (O_741,N_18019,N_18639);
xnor UO_742 (O_742,N_17809,N_18923);
and UO_743 (O_743,N_17508,N_16759);
and UO_744 (O_744,N_17223,N_18230);
nor UO_745 (O_745,N_18756,N_19321);
nor UO_746 (O_746,N_18904,N_18938);
nor UO_747 (O_747,N_18989,N_17309);
or UO_748 (O_748,N_19294,N_18915);
and UO_749 (O_749,N_16035,N_19787);
or UO_750 (O_750,N_17438,N_19425);
nand UO_751 (O_751,N_17030,N_17673);
nor UO_752 (O_752,N_18699,N_16036);
or UO_753 (O_753,N_17864,N_17758);
nand UO_754 (O_754,N_16424,N_17830);
and UO_755 (O_755,N_19715,N_17681);
nand UO_756 (O_756,N_16319,N_18972);
nor UO_757 (O_757,N_18580,N_16541);
or UO_758 (O_758,N_17584,N_17693);
or UO_759 (O_759,N_19581,N_19565);
or UO_760 (O_760,N_19414,N_16611);
or UO_761 (O_761,N_18317,N_16453);
nor UO_762 (O_762,N_19299,N_18134);
or UO_763 (O_763,N_17011,N_18421);
or UO_764 (O_764,N_18062,N_19692);
or UO_765 (O_765,N_18830,N_18933);
nor UO_766 (O_766,N_18519,N_17344);
nor UO_767 (O_767,N_17356,N_19132);
nand UO_768 (O_768,N_18767,N_19714);
nand UO_769 (O_769,N_19434,N_18341);
xor UO_770 (O_770,N_19738,N_18878);
nor UO_771 (O_771,N_18424,N_19393);
nor UO_772 (O_772,N_17831,N_16552);
or UO_773 (O_773,N_18925,N_19028);
and UO_774 (O_774,N_17906,N_16509);
and UO_775 (O_775,N_16967,N_17082);
nand UO_776 (O_776,N_18323,N_19303);
or UO_777 (O_777,N_18074,N_18907);
and UO_778 (O_778,N_16703,N_18542);
or UO_779 (O_779,N_16218,N_19547);
or UO_780 (O_780,N_19967,N_16508);
nor UO_781 (O_781,N_16127,N_16769);
xnor UO_782 (O_782,N_16199,N_16862);
or UO_783 (O_783,N_16533,N_18554);
and UO_784 (O_784,N_19768,N_18661);
or UO_785 (O_785,N_19057,N_18252);
or UO_786 (O_786,N_18951,N_19949);
nand UO_787 (O_787,N_16033,N_16354);
or UO_788 (O_788,N_16266,N_19529);
or UO_789 (O_789,N_16580,N_18133);
xor UO_790 (O_790,N_19574,N_19437);
nor UO_791 (O_791,N_17413,N_16311);
xnor UO_792 (O_792,N_18966,N_16045);
nor UO_793 (O_793,N_18682,N_17704);
nor UO_794 (O_794,N_16377,N_16708);
and UO_795 (O_795,N_17352,N_16990);
and UO_796 (O_796,N_16854,N_19255);
nor UO_797 (O_797,N_17778,N_19907);
and UO_798 (O_798,N_19314,N_17328);
or UO_799 (O_799,N_18435,N_16332);
nand UO_800 (O_800,N_16739,N_18646);
and UO_801 (O_801,N_19583,N_17465);
nand UO_802 (O_802,N_17964,N_16815);
xor UO_803 (O_803,N_19257,N_19456);
nor UO_804 (O_804,N_17376,N_16675);
nor UO_805 (O_805,N_18511,N_17429);
nand UO_806 (O_806,N_19262,N_19104);
nor UO_807 (O_807,N_18777,N_19596);
and UO_808 (O_808,N_16212,N_18312);
nand UO_809 (O_809,N_19791,N_17325);
and UO_810 (O_810,N_19458,N_17530);
or UO_811 (O_811,N_16523,N_16103);
nor UO_812 (O_812,N_16619,N_19809);
nor UO_813 (O_813,N_18995,N_17642);
or UO_814 (O_814,N_16583,N_17288);
or UO_815 (O_815,N_17178,N_18201);
and UO_816 (O_816,N_16730,N_17967);
and UO_817 (O_817,N_19779,N_19509);
nand UO_818 (O_818,N_17191,N_19737);
nand UO_819 (O_819,N_19493,N_16645);
and UO_820 (O_820,N_16163,N_16608);
and UO_821 (O_821,N_17478,N_17007);
xnor UO_822 (O_822,N_16830,N_18627);
nor UO_823 (O_823,N_18572,N_18217);
nand UO_824 (O_824,N_18863,N_18055);
nand UO_825 (O_825,N_16949,N_17232);
and UO_826 (O_826,N_17847,N_18072);
nand UO_827 (O_827,N_16085,N_16448);
or UO_828 (O_828,N_16168,N_18758);
nand UO_829 (O_829,N_19821,N_18060);
and UO_830 (O_830,N_18460,N_17832);
or UO_831 (O_831,N_17876,N_18221);
nand UO_832 (O_832,N_18621,N_16490);
and UO_833 (O_833,N_16833,N_19169);
xor UO_834 (O_834,N_19154,N_16364);
or UO_835 (O_835,N_16099,N_17572);
and UO_836 (O_836,N_18566,N_17734);
or UO_837 (O_837,N_17746,N_16600);
and UO_838 (O_838,N_16903,N_17270);
nor UO_839 (O_839,N_18235,N_16568);
and UO_840 (O_840,N_18315,N_17485);
or UO_841 (O_841,N_19570,N_19001);
nand UO_842 (O_842,N_18593,N_19930);
nor UO_843 (O_843,N_17306,N_19549);
nand UO_844 (O_844,N_17454,N_18283);
and UO_845 (O_845,N_17760,N_19067);
nor UO_846 (O_846,N_17627,N_17196);
nand UO_847 (O_847,N_16429,N_19995);
and UO_848 (O_848,N_17782,N_19215);
nand UO_849 (O_849,N_17499,N_16011);
nand UO_850 (O_850,N_19289,N_17786);
nand UO_851 (O_851,N_19022,N_17934);
xnor UO_852 (O_852,N_16321,N_16069);
nor UO_853 (O_853,N_17999,N_19656);
xor UO_854 (O_854,N_18748,N_18837);
nand UO_855 (O_855,N_19732,N_19199);
and UO_856 (O_856,N_16626,N_17409);
or UO_857 (O_857,N_16133,N_17976);
nor UO_858 (O_858,N_17330,N_16977);
and UO_859 (O_859,N_17568,N_16091);
or UO_860 (O_860,N_18356,N_19976);
or UO_861 (O_861,N_18964,N_19108);
nand UO_862 (O_862,N_18442,N_17879);
nand UO_863 (O_863,N_18692,N_17542);
and UO_864 (O_864,N_19568,N_18316);
xnor UO_865 (O_865,N_17604,N_19138);
xnor UO_866 (O_866,N_17069,N_18553);
and UO_867 (O_867,N_17372,N_16798);
and UO_868 (O_868,N_17762,N_19477);
and UO_869 (O_869,N_16505,N_17556);
nor UO_870 (O_870,N_18665,N_18267);
nor UO_871 (O_871,N_17432,N_17878);
and UO_872 (O_872,N_16947,N_19447);
or UO_873 (O_873,N_17034,N_18632);
xnor UO_874 (O_874,N_16337,N_18776);
or UO_875 (O_875,N_19122,N_19279);
or UO_876 (O_876,N_19888,N_16450);
nor UO_877 (O_877,N_18803,N_17640);
and UO_878 (O_878,N_18407,N_18968);
nor UO_879 (O_879,N_18108,N_18182);
and UO_880 (O_880,N_16966,N_18039);
or UO_881 (O_881,N_19161,N_17822);
nor UO_882 (O_882,N_19301,N_19619);
and UO_883 (O_883,N_18694,N_19542);
nor UO_884 (O_884,N_19620,N_18970);
or UO_885 (O_885,N_19952,N_17630);
nor UO_886 (O_886,N_18918,N_17078);
nand UO_887 (O_887,N_16662,N_18584);
xor UO_888 (O_888,N_16172,N_17339);
nor UO_889 (O_889,N_17910,N_17179);
nor UO_890 (O_890,N_19124,N_16540);
xor UO_891 (O_891,N_18503,N_17637);
and UO_892 (O_892,N_17987,N_19133);
xnor UO_893 (O_893,N_19185,N_19139);
nand UO_894 (O_894,N_19742,N_19911);
nand UO_895 (O_895,N_18828,N_19076);
and UO_896 (O_896,N_18835,N_19638);
nor UO_897 (O_897,N_17036,N_16923);
and UO_898 (O_898,N_17363,N_16146);
nand UO_899 (O_899,N_16433,N_18053);
xor UO_900 (O_900,N_19959,N_19081);
and UO_901 (O_901,N_19384,N_19353);
nand UO_902 (O_902,N_18280,N_18219);
nor UO_903 (O_903,N_16924,N_19672);
nand UO_904 (O_904,N_17451,N_16014);
and UO_905 (O_905,N_16224,N_18193);
or UO_906 (O_906,N_19511,N_18351);
and UO_907 (O_907,N_17278,N_18198);
or UO_908 (O_908,N_18610,N_17692);
and UO_909 (O_909,N_18107,N_16123);
xnor UO_910 (O_910,N_19513,N_17920);
or UO_911 (O_911,N_19958,N_18903);
and UO_912 (O_912,N_16504,N_17003);
nand UO_913 (O_913,N_17304,N_17559);
or UO_914 (O_914,N_17132,N_18528);
nor UO_915 (O_915,N_18935,N_16934);
nor UO_916 (O_916,N_16370,N_19525);
nor UO_917 (O_917,N_18718,N_18394);
or UO_918 (O_918,N_17199,N_19523);
nand UO_919 (O_919,N_17172,N_18927);
xor UO_920 (O_920,N_18763,N_19933);
nor UO_921 (O_921,N_18673,N_17844);
and UO_922 (O_922,N_19749,N_17402);
xor UO_923 (O_923,N_16589,N_17458);
nor UO_924 (O_924,N_16956,N_19460);
or UO_925 (O_925,N_18330,N_16044);
or UO_926 (O_926,N_19545,N_17261);
nor UO_927 (O_927,N_16204,N_16970);
or UO_928 (O_928,N_16225,N_18224);
nand UO_929 (O_929,N_18619,N_17217);
and UO_930 (O_930,N_16405,N_16594);
nor UO_931 (O_931,N_18671,N_18101);
or UO_932 (O_932,N_16080,N_19305);
or UO_933 (O_933,N_18310,N_16997);
and UO_934 (O_934,N_17836,N_16819);
nor UO_935 (O_935,N_18373,N_17730);
or UO_936 (O_936,N_19863,N_16455);
nor UO_937 (O_937,N_18752,N_18236);
or UO_938 (O_938,N_19973,N_17087);
or UO_939 (O_939,N_18212,N_16801);
or UO_940 (O_940,N_17362,N_17869);
or UO_941 (O_941,N_19603,N_19319);
and UO_942 (O_942,N_18344,N_17180);
and UO_943 (O_943,N_19642,N_18180);
xnor UO_944 (O_944,N_17721,N_17143);
nor UO_945 (O_945,N_17521,N_19955);
nor UO_946 (O_946,N_17567,N_17230);
nor UO_947 (O_947,N_18740,N_17840);
nand UO_948 (O_948,N_17908,N_18010);
nand UO_949 (O_949,N_19560,N_17498);
or UO_950 (O_950,N_18504,N_19065);
nand UO_951 (O_951,N_16688,N_19723);
and UO_952 (O_952,N_16179,N_19895);
nand UO_953 (O_953,N_19601,N_19196);
nor UO_954 (O_954,N_16135,N_17664);
nand UO_955 (O_955,N_16154,N_19798);
nand UO_956 (O_956,N_17272,N_18940);
nand UO_957 (O_957,N_16794,N_18766);
or UO_958 (O_958,N_19796,N_16155);
nor UO_959 (O_959,N_18886,N_17345);
or UO_960 (O_960,N_17922,N_19005);
nand UO_961 (O_961,N_17065,N_16562);
nand UO_962 (O_962,N_19968,N_17099);
nor UO_963 (O_963,N_19579,N_18706);
nand UO_964 (O_964,N_19084,N_18668);
nand UO_965 (O_965,N_18523,N_19236);
nor UO_966 (O_966,N_19948,N_19537);
or UO_967 (O_967,N_17616,N_17151);
xnor UO_968 (O_968,N_19686,N_19461);
or UO_969 (O_969,N_16416,N_19559);
nor UO_970 (O_970,N_17954,N_17256);
or UO_971 (O_971,N_17190,N_17240);
nor UO_972 (O_972,N_17245,N_17765);
and UO_973 (O_973,N_16886,N_16935);
xor UO_974 (O_974,N_19998,N_18023);
nor UO_975 (O_975,N_16408,N_17449);
and UO_976 (O_976,N_16419,N_16655);
nand UO_977 (O_977,N_16067,N_19709);
or UO_978 (O_978,N_17307,N_16065);
nand UO_979 (O_979,N_19681,N_17829);
or UO_980 (O_980,N_17295,N_17865);
xnor UO_981 (O_981,N_16616,N_19902);
xnor UO_982 (O_982,N_19908,N_18214);
nor UO_983 (O_983,N_16571,N_19453);
or UO_984 (O_984,N_19333,N_18138);
and UO_985 (O_985,N_19733,N_19848);
nand UO_986 (O_986,N_19272,N_18073);
or UO_987 (O_987,N_16659,N_19467);
or UO_988 (O_988,N_16132,N_17668);
nand UO_989 (O_989,N_19757,N_19370);
nor UO_990 (O_990,N_17450,N_19898);
and UO_991 (O_991,N_19632,N_18969);
nor UO_992 (O_992,N_16828,N_17860);
and UO_993 (O_993,N_19936,N_18859);
or UO_994 (O_994,N_19009,N_17412);
and UO_995 (O_995,N_18656,N_17969);
or UO_996 (O_996,N_18147,N_18371);
or UO_997 (O_997,N_18618,N_17736);
xnor UO_998 (O_998,N_18261,N_19072);
nor UO_999 (O_999,N_18054,N_17825);
and UO_1000 (O_1000,N_17705,N_16831);
or UO_1001 (O_1001,N_19855,N_18273);
and UO_1002 (O_1002,N_19659,N_17086);
nor UO_1003 (O_1003,N_18097,N_19079);
and UO_1004 (O_1004,N_19159,N_17401);
or UO_1005 (O_1005,N_16758,N_18112);
or UO_1006 (O_1006,N_18883,N_19471);
nand UO_1007 (O_1007,N_16489,N_16475);
nor UO_1008 (O_1008,N_17148,N_18459);
nor UO_1009 (O_1009,N_17848,N_19785);
or UO_1010 (O_1010,N_17843,N_19201);
and UO_1011 (O_1011,N_19986,N_16578);
nand UO_1012 (O_1012,N_19360,N_19562);
or UO_1013 (O_1013,N_19990,N_17434);
or UO_1014 (O_1014,N_16229,N_16599);
or UO_1015 (O_1015,N_19527,N_16150);
or UO_1016 (O_1016,N_18882,N_19144);
and UO_1017 (O_1017,N_16964,N_16912);
and UO_1018 (O_1018,N_18678,N_19343);
and UO_1019 (O_1019,N_19113,N_19739);
nand UO_1020 (O_1020,N_17203,N_18412);
or UO_1021 (O_1021,N_19281,N_16603);
or UO_1022 (O_1022,N_18794,N_19589);
nor UO_1023 (O_1023,N_17545,N_18855);
or UO_1024 (O_1024,N_19149,N_16920);
xnor UO_1025 (O_1025,N_17098,N_18514);
or UO_1026 (O_1026,N_19896,N_18361);
nor UO_1027 (O_1027,N_19623,N_16670);
nand UO_1028 (O_1028,N_16367,N_16259);
and UO_1029 (O_1029,N_16525,N_16318);
nand UO_1030 (O_1030,N_16344,N_18292);
xor UO_1031 (O_1031,N_18402,N_18082);
nand UO_1032 (O_1032,N_16390,N_18798);
nand UO_1033 (O_1033,N_19891,N_17313);
nand UO_1034 (O_1034,N_17246,N_16494);
or UO_1035 (O_1035,N_19249,N_19436);
nor UO_1036 (O_1036,N_16872,N_18888);
xor UO_1037 (O_1037,N_19442,N_19388);
nand UO_1038 (O_1038,N_18524,N_17163);
xnor UO_1039 (O_1039,N_19282,N_17648);
and UO_1040 (O_1040,N_17707,N_18464);
or UO_1041 (O_1041,N_19691,N_17124);
and UO_1042 (O_1042,N_17649,N_18727);
and UO_1043 (O_1043,N_16476,N_16030);
nor UO_1044 (O_1044,N_18173,N_18816);
and UO_1045 (O_1045,N_16400,N_16751);
and UO_1046 (O_1046,N_17023,N_19195);
xnor UO_1047 (O_1047,N_19010,N_19790);
nand UO_1048 (O_1048,N_19794,N_16258);
nor UO_1049 (O_1049,N_16376,N_17569);
or UO_1050 (O_1050,N_16629,N_19347);
and UO_1051 (O_1051,N_18930,N_16355);
or UO_1052 (O_1052,N_18868,N_19049);
xnor UO_1053 (O_1053,N_18052,N_19200);
nor UO_1054 (O_1054,N_19864,N_18286);
xnor UO_1055 (O_1055,N_18381,N_18473);
and UO_1056 (O_1056,N_18583,N_19812);
xor UO_1057 (O_1057,N_17953,N_19380);
and UO_1058 (O_1058,N_17598,N_16294);
or UO_1059 (O_1059,N_19924,N_16517);
and UO_1060 (O_1060,N_19469,N_16491);
xor UO_1061 (O_1061,N_17100,N_17337);
xnor UO_1062 (O_1062,N_16174,N_17890);
and UO_1063 (O_1063,N_18427,N_16895);
xor UO_1064 (O_1064,N_17416,N_19352);
nand UO_1065 (O_1065,N_18321,N_19166);
or UO_1066 (O_1066,N_19296,N_18898);
and UO_1067 (O_1067,N_18050,N_19212);
nor UO_1068 (O_1068,N_16213,N_16998);
nor UO_1069 (O_1069,N_19627,N_19315);
nor UO_1070 (O_1070,N_18003,N_16972);
nand UO_1071 (O_1071,N_19327,N_18753);
and UO_1072 (O_1072,N_19288,N_16524);
xnor UO_1073 (O_1073,N_16869,N_18227);
and UO_1074 (O_1074,N_16087,N_16010);
nor UO_1075 (O_1075,N_19376,N_17587);
xnor UO_1076 (O_1076,N_18228,N_18747);
and UO_1077 (O_1077,N_16887,N_17526);
nand UO_1078 (O_1078,N_18754,N_16284);
and UO_1079 (O_1079,N_18826,N_17411);
nor UO_1080 (O_1080,N_17088,N_16275);
nand UO_1081 (O_1081,N_17815,N_18860);
nor UO_1082 (O_1082,N_16727,N_16032);
or UO_1083 (O_1083,N_17404,N_17463);
and UO_1084 (O_1084,N_19957,N_19917);
nor UO_1085 (O_1085,N_17369,N_17510);
and UO_1086 (O_1086,N_17589,N_16733);
nor UO_1087 (O_1087,N_18066,N_17236);
and UO_1088 (O_1088,N_17317,N_17992);
and UO_1089 (O_1089,N_16697,N_19726);
nand UO_1090 (O_1090,N_19879,N_19455);
nand UO_1091 (O_1091,N_17303,N_19699);
nand UO_1092 (O_1092,N_18788,N_19978);
nor UO_1093 (O_1093,N_17017,N_19966);
and UO_1094 (O_1094,N_18985,N_16215);
nor UO_1095 (O_1095,N_16018,N_19873);
nand UO_1096 (O_1096,N_19497,N_16403);
nand UO_1097 (O_1097,N_19354,N_17197);
and UO_1098 (O_1098,N_19090,N_16983);
nor UO_1099 (O_1099,N_17186,N_16750);
or UO_1100 (O_1100,N_17053,N_19540);
xor UO_1101 (O_1101,N_19409,N_17357);
xor UO_1102 (O_1102,N_18581,N_16098);
or UO_1103 (O_1103,N_16876,N_17555);
nor UO_1104 (O_1104,N_18577,N_17491);
nor UO_1105 (O_1105,N_16451,N_17495);
and UO_1106 (O_1106,N_18127,N_19189);
xor UO_1107 (O_1107,N_17321,N_18824);
and UO_1108 (O_1108,N_17229,N_16747);
nor UO_1109 (O_1109,N_18887,N_17979);
xnor UO_1110 (O_1110,N_16890,N_19291);
and UO_1111 (O_1111,N_18349,N_18425);
or UO_1112 (O_1112,N_19092,N_16738);
nor UO_1113 (O_1113,N_19772,N_19043);
or UO_1114 (O_1114,N_18192,N_17601);
and UO_1115 (O_1115,N_16068,N_16226);
or UO_1116 (O_1116,N_18462,N_16348);
nor UO_1117 (O_1117,N_19928,N_17289);
or UO_1118 (O_1118,N_18615,N_18141);
and UO_1119 (O_1119,N_17277,N_19064);
xor UO_1120 (O_1120,N_17293,N_18185);
nand UO_1121 (O_1121,N_18303,N_16690);
or UO_1122 (O_1122,N_19981,N_16338);
and UO_1123 (O_1123,N_17533,N_17805);
nor UO_1124 (O_1124,N_17680,N_16379);
or UO_1125 (O_1125,N_16974,N_18866);
or UO_1126 (O_1126,N_18482,N_18115);
nand UO_1127 (O_1127,N_18691,N_19532);
xnor UO_1128 (O_1128,N_17117,N_16062);
nand UO_1129 (O_1129,N_18854,N_18981);
or UO_1130 (O_1130,N_19403,N_19328);
and UO_1131 (O_1131,N_16632,N_16333);
or UO_1132 (O_1132,N_17101,N_17824);
or UO_1133 (O_1133,N_16944,N_17316);
and UO_1134 (O_1134,N_17198,N_19066);
and UO_1135 (O_1135,N_18890,N_19954);
and UO_1136 (O_1136,N_18457,N_18545);
nor UO_1137 (O_1137,N_18599,N_16792);
or UO_1138 (O_1138,N_19400,N_16512);
nand UO_1139 (O_1139,N_17167,N_19674);
or UO_1140 (O_1140,N_16314,N_16841);
and UO_1141 (O_1141,N_19652,N_16461);
nor UO_1142 (O_1142,N_16118,N_16820);
xor UO_1143 (O_1143,N_17021,N_18120);
and UO_1144 (O_1144,N_19751,N_18257);
nor UO_1145 (O_1145,N_17291,N_16189);
nor UO_1146 (O_1146,N_18543,N_18934);
xor UO_1147 (O_1147,N_17764,N_17259);
nor UO_1148 (O_1148,N_17012,N_19284);
nand UO_1149 (O_1149,N_17935,N_17956);
and UO_1150 (O_1150,N_17636,N_17515);
nor UO_1151 (O_1151,N_19078,N_16529);
nor UO_1152 (O_1152,N_17807,N_18233);
nand UO_1153 (O_1153,N_18635,N_16962);
nand UO_1154 (O_1154,N_19286,N_16316);
nand UO_1155 (O_1155,N_19192,N_19231);
and UO_1156 (O_1156,N_18641,N_19783);
xor UO_1157 (O_1157,N_16856,N_19224);
nand UO_1158 (O_1158,N_16846,N_19991);
or UO_1159 (O_1159,N_17833,N_16356);
nor UO_1160 (O_1160,N_17706,N_16138);
xor UO_1161 (O_1161,N_19518,N_16320);
or UO_1162 (O_1162,N_17767,N_17826);
and UO_1163 (O_1163,N_18986,N_17505);
or UO_1164 (O_1164,N_19374,N_18190);
xor UO_1165 (O_1165,N_17251,N_19576);
nand UO_1166 (O_1166,N_19956,N_18038);
and UO_1167 (O_1167,N_18362,N_17803);
nor UO_1168 (O_1168,N_17275,N_18990);
nand UO_1169 (O_1169,N_18199,N_17591);
and UO_1170 (O_1170,N_17561,N_17709);
nand UO_1171 (O_1171,N_17603,N_17715);
or UO_1172 (O_1172,N_17346,N_17534);
nor UO_1173 (O_1173,N_17182,N_16866);
nand UO_1174 (O_1174,N_17427,N_18494);
xor UO_1175 (O_1175,N_18978,N_17055);
nand UO_1176 (O_1176,N_17949,N_17091);
nor UO_1177 (O_1177,N_19223,N_16729);
nor UO_1178 (O_1178,N_17751,N_16714);
nand UO_1179 (O_1179,N_19181,N_16093);
and UO_1180 (O_1180,N_18365,N_17137);
or UO_1181 (O_1181,N_18081,N_17877);
xnor UO_1182 (O_1182,N_16276,N_16239);
or UO_1183 (O_1183,N_19921,N_16297);
or UO_1184 (O_1184,N_16824,N_16350);
or UO_1185 (O_1185,N_17033,N_19238);
nor UO_1186 (O_1186,N_16095,N_17050);
or UO_1187 (O_1187,N_16006,N_18654);
nand UO_1188 (O_1188,N_18757,N_16667);
nor UO_1189 (O_1189,N_16107,N_19480);
nor UO_1190 (O_1190,N_18617,N_19510);
nor UO_1191 (O_1191,N_16958,N_18071);
nand UO_1192 (O_1192,N_19363,N_18493);
and UO_1193 (O_1193,N_17305,N_18366);
and UO_1194 (O_1194,N_18931,N_19728);
nand UO_1195 (O_1195,N_17061,N_19244);
and UO_1196 (O_1196,N_19662,N_18664);
or UO_1197 (O_1197,N_19650,N_19432);
and UO_1198 (O_1198,N_19755,N_17623);
or UO_1199 (O_1199,N_16586,N_17403);
nand UO_1200 (O_1200,N_18444,N_19754);
and UO_1201 (O_1201,N_19682,N_16585);
nand UO_1202 (O_1202,N_18576,N_18769);
or UO_1203 (O_1203,N_18446,N_17531);
nor UO_1204 (O_1204,N_18102,N_16991);
nor UO_1205 (O_1205,N_16039,N_17683);
or UO_1206 (O_1206,N_19320,N_16009);
nor UO_1207 (O_1207,N_19841,N_17027);
nor UO_1208 (O_1208,N_18963,N_19401);
nor UO_1209 (O_1209,N_18735,N_16883);
nor UO_1210 (O_1210,N_16365,N_17651);
or UO_1211 (O_1211,N_19610,N_16724);
and UO_1212 (O_1212,N_16203,N_19571);
nor UO_1213 (O_1213,N_18327,N_19494);
nand UO_1214 (O_1214,N_16075,N_16968);
and UO_1215 (O_1215,N_18902,N_16764);
nor UO_1216 (O_1216,N_19803,N_17670);
or UO_1217 (O_1217,N_19854,N_16802);
and UO_1218 (O_1218,N_19256,N_17791);
and UO_1219 (O_1219,N_17398,N_18980);
and UO_1220 (O_1220,N_19597,N_18962);
nor UO_1221 (O_1221,N_16591,N_16741);
or UO_1222 (O_1222,N_17812,N_19394);
nor UO_1223 (O_1223,N_16078,N_18420);
nand UO_1224 (O_1224,N_18014,N_17518);
nor UO_1225 (O_1225,N_17420,N_19047);
xnor UO_1226 (O_1226,N_17647,N_19095);
nor UO_1227 (O_1227,N_17308,N_17006);
nor UO_1228 (O_1228,N_19474,N_17823);
nand UO_1229 (O_1229,N_18048,N_16188);
nand UO_1230 (O_1230,N_19771,N_17460);
or UO_1231 (O_1231,N_19089,N_19142);
and UO_1232 (O_1232,N_16668,N_17062);
and UO_1233 (O_1233,N_17737,N_18337);
or UO_1234 (O_1234,N_17268,N_16712);
or UO_1235 (O_1235,N_19258,N_17950);
nand UO_1236 (O_1236,N_17119,N_19428);
and UO_1237 (O_1237,N_19271,N_19906);
nor UO_1238 (O_1238,N_19445,N_18681);
nand UO_1239 (O_1239,N_19316,N_18211);
and UO_1240 (O_1240,N_19267,N_19502);
nand UO_1241 (O_1241,N_19536,N_19128);
and UO_1242 (O_1242,N_18453,N_18379);
nor UO_1243 (O_1243,N_16829,N_19897);
or UO_1244 (O_1244,N_17965,N_19923);
or UO_1245 (O_1245,N_16394,N_18423);
and UO_1246 (O_1246,N_19815,N_19123);
or UO_1247 (O_1247,N_16151,N_19845);
or UO_1248 (O_1248,N_19068,N_17981);
and UO_1249 (O_1249,N_18487,N_18238);
and UO_1250 (O_1250,N_16706,N_16622);
nor UO_1251 (O_1251,N_17032,N_16575);
nor UO_1252 (O_1252,N_17282,N_17859);
or UO_1253 (O_1253,N_19308,N_18795);
nor UO_1254 (O_1254,N_19519,N_16439);
nor UO_1255 (O_1255,N_16140,N_16235);
nor UO_1256 (O_1256,N_16557,N_16847);
nand UO_1257 (O_1257,N_18872,N_16247);
xor UO_1258 (O_1258,N_17957,N_18733);
nor UO_1259 (O_1259,N_18843,N_19011);
xor UO_1260 (O_1260,N_17955,N_18645);
nand UO_1261 (O_1261,N_17408,N_19251);
nor UO_1262 (O_1262,N_17752,N_19592);
or UO_1263 (O_1263,N_16664,N_16894);
and UO_1264 (O_1264,N_17655,N_16648);
and UO_1265 (O_1265,N_17292,N_18376);
xor UO_1266 (O_1266,N_18094,N_17866);
nand UO_1267 (O_1267,N_16060,N_19938);
nor UO_1268 (O_1268,N_18650,N_16236);
or UO_1269 (O_1269,N_17126,N_17682);
and UO_1270 (O_1270,N_19860,N_18124);
nor UO_1271 (O_1271,N_19524,N_16252);
xor UO_1272 (O_1272,N_19947,N_18921);
nand UO_1273 (O_1273,N_19259,N_17768);
nor UO_1274 (O_1274,N_19969,N_19805);
nor UO_1275 (O_1275,N_19055,N_18251);
nand UO_1276 (O_1276,N_16042,N_18210);
and UO_1277 (O_1277,N_17090,N_17915);
xnor UO_1278 (O_1278,N_18340,N_17892);
nand UO_1279 (O_1279,N_16156,N_17501);
and UO_1280 (O_1280,N_17576,N_18285);
nand UO_1281 (O_1281,N_16464,N_17674);
or UO_1282 (O_1282,N_19107,N_18111);
xor UO_1283 (O_1283,N_19818,N_19992);
xnor UO_1284 (O_1284,N_19371,N_19736);
and UO_1285 (O_1285,N_19392,N_18026);
and UO_1286 (O_1286,N_16101,N_19035);
nor UO_1287 (O_1287,N_19443,N_16681);
and UO_1288 (O_1288,N_17701,N_19086);
and UO_1289 (O_1289,N_17241,N_19838);
nand UO_1290 (O_1290,N_19735,N_17929);
nor UO_1291 (O_1291,N_16373,N_19075);
nand UO_1292 (O_1292,N_18188,N_18129);
nor UO_1293 (O_1293,N_16324,N_16177);
nand UO_1294 (O_1294,N_16857,N_19756);
xnor UO_1295 (O_1295,N_18380,N_19318);
or UO_1296 (O_1296,N_16286,N_17266);
or UO_1297 (O_1297,N_16161,N_19718);
and UO_1298 (O_1298,N_19825,N_17122);
nand UO_1299 (O_1299,N_19117,N_19150);
and UO_1300 (O_1300,N_19366,N_17525);
nand UO_1301 (O_1301,N_19002,N_19997);
and UO_1302 (O_1302,N_16676,N_18947);
nand UO_1303 (O_1303,N_17958,N_16686);
nand UO_1304 (O_1304,N_19408,N_16556);
nand UO_1305 (O_1305,N_17225,N_16015);
nand UO_1306 (O_1306,N_19535,N_18471);
and UO_1307 (O_1307,N_17849,N_16026);
nor UO_1308 (O_1308,N_17732,N_19889);
nor UO_1309 (O_1309,N_16159,N_16907);
or UO_1310 (O_1310,N_17731,N_17671);
nand UO_1311 (O_1311,N_19713,N_16300);
or UO_1312 (O_1312,N_16208,N_17880);
nand UO_1313 (O_1313,N_16931,N_17107);
and UO_1314 (O_1314,N_18409,N_18428);
xnor UO_1315 (O_1315,N_16499,N_18945);
nand UO_1316 (O_1316,N_16227,N_18197);
nor UO_1317 (O_1317,N_18716,N_18849);
nand UO_1318 (O_1318,N_19454,N_16157);
nor UO_1319 (O_1319,N_16396,N_17248);
nand UO_1320 (O_1320,N_19740,N_16658);
or UO_1321 (O_1321,N_19671,N_18131);
or UO_1322 (O_1322,N_18044,N_17123);
nor UO_1323 (O_1323,N_18495,N_16473);
or UO_1324 (O_1324,N_18241,N_19500);
xnor UO_1325 (O_1325,N_17355,N_19904);
or UO_1326 (O_1326,N_16362,N_19103);
nand UO_1327 (O_1327,N_16366,N_18140);
or UO_1328 (O_1328,N_18844,N_17728);
and UO_1329 (O_1329,N_18396,N_19843);
or UO_1330 (O_1330,N_19489,N_19220);
nor UO_1331 (O_1331,N_18158,N_16308);
nand UO_1332 (O_1332,N_17699,N_16442);
nor UO_1333 (O_1333,N_16843,N_18737);
and UO_1334 (O_1334,N_17921,N_16813);
nor UO_1335 (O_1335,N_19309,N_19982);
nor UO_1336 (O_1336,N_17136,N_17787);
nand UO_1337 (O_1337,N_16982,N_16513);
or UO_1338 (O_1338,N_17102,N_19193);
or UO_1339 (O_1339,N_17497,N_19752);
nand UO_1340 (O_1340,N_19491,N_18559);
or UO_1341 (O_1341,N_17315,N_16414);
nor UO_1342 (O_1342,N_18121,N_18749);
or UO_1343 (O_1343,N_17607,N_18660);
xor UO_1344 (O_1344,N_17296,N_17727);
and UO_1345 (O_1345,N_16176,N_18771);
and UO_1346 (O_1346,N_16588,N_16285);
or UO_1347 (O_1347,N_17043,N_16559);
xor UO_1348 (O_1348,N_18937,N_17031);
nor UO_1349 (O_1349,N_17335,N_18364);
nand UO_1350 (O_1350,N_19143,N_16538);
and UO_1351 (O_1351,N_19939,N_16527);
or UO_1352 (O_1352,N_16721,N_16053);
nor UO_1353 (O_1353,N_16086,N_17410);
or UO_1354 (O_1354,N_19040,N_17469);
or UO_1355 (O_1355,N_18355,N_16269);
nand UO_1356 (O_1356,N_17152,N_16692);
and UO_1357 (O_1357,N_18510,N_19507);
nand UO_1358 (O_1358,N_19533,N_17982);
or UO_1359 (O_1359,N_18818,N_18695);
or UO_1360 (O_1360,N_19819,N_16351);
nor UO_1361 (O_1361,N_18829,N_19962);
nor UO_1362 (O_1362,N_16875,N_19085);
nor UO_1363 (O_1363,N_19242,N_17314);
and UO_1364 (O_1364,N_16795,N_16104);
xor UO_1365 (O_1365,N_19943,N_18772);
nor UO_1366 (O_1366,N_18522,N_16178);
or UO_1367 (O_1367,N_19711,N_16779);
and UO_1368 (O_1368,N_16707,N_17177);
or UO_1369 (O_1369,N_16881,N_17108);
nor UO_1370 (O_1370,N_17632,N_18043);
nor UO_1371 (O_1371,N_17573,N_16840);
nor UO_1372 (O_1372,N_19378,N_17799);
xnor UO_1373 (O_1373,N_18881,N_18700);
and UO_1374 (O_1374,N_17527,N_18246);
and UO_1375 (O_1375,N_18509,N_18314);
or UO_1376 (O_1376,N_19719,N_16310);
nor UO_1377 (O_1377,N_18988,N_16305);
xor UO_1378 (O_1378,N_16945,N_18202);
nand UO_1379 (O_1379,N_19639,N_18433);
nor UO_1380 (O_1380,N_18810,N_18492);
nand UO_1381 (O_1381,N_16811,N_19996);
or UO_1382 (O_1382,N_16551,N_16952);
and UO_1383 (O_1383,N_19977,N_18987);
nor UO_1384 (O_1384,N_18191,N_19439);
xor UO_1385 (O_1385,N_19685,N_16507);
nand UO_1386 (O_1386,N_19349,N_18744);
nand UO_1387 (O_1387,N_16331,N_19558);
or UO_1388 (O_1388,N_17986,N_19003);
and UO_1389 (O_1389,N_19501,N_17047);
or UO_1390 (O_1390,N_16928,N_16410);
nand UO_1391 (O_1391,N_18156,N_16470);
xnor UO_1392 (O_1392,N_16534,N_17635);
or UO_1393 (O_1393,N_16716,N_16590);
nor UO_1394 (O_1394,N_19162,N_19483);
or UO_1395 (O_1395,N_17018,N_17394);
xnor UO_1396 (O_1396,N_17818,N_19761);
nand UO_1397 (O_1397,N_18168,N_17800);
and UO_1398 (O_1398,N_19235,N_18552);
nand UO_1399 (O_1399,N_16306,N_16122);
nor UO_1400 (O_1400,N_19276,N_19131);
or UO_1401 (O_1401,N_16079,N_17333);
or UO_1402 (O_1402,N_17354,N_18232);
and UO_1403 (O_1403,N_16112,N_17441);
nor UO_1404 (O_1404,N_19416,N_18332);
nor UO_1405 (O_1405,N_19036,N_16190);
and UO_1406 (O_1406,N_17214,N_19802);
nor UO_1407 (O_1407,N_16412,N_19410);
and UO_1408 (O_1408,N_17265,N_18378);
nor UO_1409 (O_1409,N_16421,N_19202);
nor UO_1410 (O_1410,N_16443,N_17224);
and UO_1411 (O_1411,N_19613,N_16953);
or UO_1412 (O_1412,N_17792,N_19810);
nand UO_1413 (O_1413,N_16735,N_17643);
nand UO_1414 (O_1414,N_17052,N_18051);
nand UO_1415 (O_1415,N_19777,N_19988);
nand UO_1416 (O_1416,N_16409,N_17948);
and UO_1417 (O_1417,N_18588,N_17837);
nand UO_1418 (O_1418,N_17228,N_19430);
nor UO_1419 (O_1419,N_18920,N_16592);
nor UO_1420 (O_1420,N_16641,N_17722);
or UO_1421 (O_1421,N_19341,N_18913);
and UO_1422 (O_1422,N_19339,N_16211);
nand UO_1423 (O_1423,N_16700,N_16904);
nand UO_1424 (O_1424,N_16761,N_17258);
nand UO_1425 (O_1425,N_17624,N_19012);
nand UO_1426 (O_1426,N_18036,N_19961);
or UO_1427 (O_1427,N_18207,N_19651);
nor UO_1428 (O_1428,N_18722,N_18475);
or UO_1429 (O_1429,N_17482,N_17658);
and UO_1430 (O_1430,N_17474,N_18449);
and UO_1431 (O_1431,N_19487,N_16234);
or UO_1432 (O_1432,N_19922,N_18218);
or UO_1433 (O_1433,N_17042,N_19614);
or UO_1434 (O_1434,N_19963,N_19683);
nor UO_1435 (O_1435,N_17891,N_19526);
xnor UO_1436 (O_1436,N_16131,N_16980);
and UO_1437 (O_1437,N_16404,N_18600);
or UO_1438 (O_1438,N_16620,N_17575);
and UO_1439 (O_1439,N_18403,N_17400);
nand UO_1440 (O_1440,N_19506,N_19155);
nand UO_1441 (O_1441,N_19479,N_17927);
nand UO_1442 (O_1442,N_18033,N_17919);
nand UO_1443 (O_1443,N_18633,N_19548);
and UO_1444 (O_1444,N_17937,N_19098);
nand UO_1445 (O_1445,N_18463,N_16171);
nand UO_1446 (O_1446,N_19056,N_18974);
nor UO_1447 (O_1447,N_16445,N_16233);
or UO_1448 (O_1448,N_16717,N_17644);
or UO_1449 (O_1449,N_19795,N_19323);
nand UO_1450 (O_1450,N_16219,N_16861);
and UO_1451 (O_1451,N_18135,N_19629);
or UO_1452 (O_1452,N_16926,N_19210);
and UO_1453 (O_1453,N_17422,N_16635);
nand UO_1454 (O_1454,N_17875,N_17997);
nor UO_1455 (O_1455,N_17436,N_19910);
nor UO_1456 (O_1456,N_19020,N_16022);
or UO_1457 (O_1457,N_16715,N_18359);
xor UO_1458 (O_1458,N_18352,N_16548);
or UO_1459 (O_1459,N_16290,N_16029);
nor UO_1460 (O_1460,N_19631,N_17961);
or UO_1461 (O_1461,N_16682,N_17966);
and UO_1462 (O_1462,N_19753,N_18225);
nor UO_1463 (O_1463,N_17111,N_18644);
nor UO_1464 (O_1464,N_17723,N_17621);
nor UO_1465 (O_1465,N_16263,N_18512);
and UO_1466 (O_1466,N_17274,N_17952);
xor UO_1467 (O_1467,N_18809,N_17077);
nand UO_1468 (O_1468,N_17072,N_19858);
or UO_1469 (O_1469,N_18454,N_17541);
xnor UO_1470 (O_1470,N_19427,N_17613);
or UO_1471 (O_1471,N_18249,N_16057);
nor UO_1472 (O_1472,N_16986,N_19679);
nand UO_1473 (O_1473,N_18290,N_19616);
and UO_1474 (O_1474,N_19190,N_18117);
or UO_1475 (O_1475,N_19975,N_17595);
nor UO_1476 (O_1476,N_19464,N_18046);
nand UO_1477 (O_1477,N_19304,N_17364);
and UO_1478 (O_1478,N_19290,N_18909);
or UO_1479 (O_1479,N_18959,N_18631);
and UO_1480 (O_1480,N_18231,N_17016);
and UO_1481 (O_1481,N_18871,N_19822);
nand UO_1482 (O_1482,N_17093,N_18807);
nor UO_1483 (O_1483,N_17397,N_16260);
or UO_1484 (O_1484,N_17238,N_16695);
or UO_1485 (O_1485,N_16277,N_17418);
and UO_1486 (O_1486,N_16282,N_18395);
or UO_1487 (O_1487,N_17038,N_16612);
nor UO_1488 (O_1488,N_18480,N_17183);
and UO_1489 (O_1489,N_19687,N_17207);
nor UO_1490 (O_1490,N_17029,N_16164);
nor UO_1491 (O_1491,N_17606,N_17661);
nand UO_1492 (O_1492,N_19567,N_19942);
nor UO_1493 (O_1493,N_16579,N_19670);
and UO_1494 (O_1494,N_18432,N_16853);
nand UO_1495 (O_1495,N_18704,N_18919);
or UO_1496 (O_1496,N_16463,N_16217);
nor UO_1497 (O_1497,N_16969,N_16503);
nand UO_1498 (O_1498,N_16584,N_17994);
or UO_1499 (O_1499,N_16361,N_17748);
or UO_1500 (O_1500,N_17828,N_18426);
and UO_1501 (O_1501,N_17563,N_19330);
and UO_1502 (O_1502,N_19126,N_17480);
nor UO_1503 (O_1503,N_17290,N_17740);
and UO_1504 (O_1504,N_16510,N_16469);
and UO_1505 (O_1505,N_19399,N_18088);
nor UO_1506 (O_1506,N_18535,N_16950);
nand UO_1507 (O_1507,N_16808,N_18256);
nor UO_1508 (O_1508,N_18680,N_17041);
and UO_1509 (O_1509,N_18679,N_17611);
and UO_1510 (O_1510,N_19157,N_19350);
nand UO_1511 (O_1511,N_18500,N_17785);
and UO_1512 (O_1512,N_16782,N_18845);
or UO_1513 (O_1513,N_19512,N_18885);
or UO_1514 (O_1514,N_17596,N_17820);
or UO_1515 (O_1515,N_18485,N_18263);
and UO_1516 (O_1516,N_17368,N_19539);
nor UO_1517 (O_1517,N_16302,N_18009);
and UO_1518 (O_1518,N_17738,N_19459);
nand UO_1519 (O_1519,N_16743,N_18240);
or UO_1520 (O_1520,N_17695,N_18601);
xnor UO_1521 (O_1521,N_16939,N_16349);
nor UO_1522 (O_1522,N_16267,N_18234);
nand UO_1523 (O_1523,N_19878,N_16254);
and UO_1524 (O_1524,N_16660,N_18092);
and UO_1525 (O_1525,N_18336,N_19912);
nand UO_1526 (O_1526,N_17801,N_18187);
and UO_1527 (O_1527,N_17138,N_17794);
and UO_1528 (O_1528,N_19268,N_19254);
nor UO_1529 (O_1529,N_18573,N_16486);
nand UO_1530 (O_1530,N_18291,N_16900);
and UO_1531 (O_1531,N_16170,N_18455);
xnor UO_1532 (O_1532,N_16978,N_19336);
nor UO_1533 (O_1533,N_17433,N_19449);
nor UO_1534 (O_1534,N_16094,N_17772);
or UO_1535 (O_1535,N_18768,N_16673);
and UO_1536 (O_1536,N_16836,N_19048);
nor UO_1537 (O_1537,N_18099,N_16630);
nor UO_1538 (O_1538,N_19252,N_16984);
nor UO_1539 (O_1539,N_17665,N_19365);
and UO_1540 (O_1540,N_16755,N_19364);
nand UO_1541 (O_1541,N_19865,N_16844);
nor UO_1542 (O_1542,N_17930,N_18030);
and UO_1543 (O_1543,N_16651,N_18825);
nor UO_1544 (O_1544,N_17351,N_16257);
nand UO_1545 (O_1545,N_19441,N_19232);
nand UO_1546 (O_1546,N_18975,N_18840);
or UO_1547 (O_1547,N_19300,N_19750);
nor UO_1548 (O_1548,N_18353,N_19929);
or UO_1549 (O_1549,N_16148,N_18658);
xnor UO_1550 (O_1550,N_16905,N_17739);
nand UO_1551 (O_1551,N_16574,N_16210);
or UO_1552 (O_1552,N_17590,N_19237);
and UO_1553 (O_1553,N_18873,N_17054);
or UO_1554 (O_1554,N_16864,N_17646);
or UO_1555 (O_1555,N_19667,N_18984);
and UO_1556 (O_1556,N_19102,N_18674);
xor UO_1557 (O_1557,N_18248,N_18167);
nand UO_1558 (O_1558,N_19515,N_19849);
nor UO_1559 (O_1559,N_16937,N_18895);
and UO_1560 (O_1560,N_19951,N_18697);
xnor UO_1561 (O_1561,N_18083,N_16048);
or UO_1562 (O_1562,N_19696,N_16454);
or UO_1563 (O_1563,N_16689,N_16652);
xor UO_1564 (O_1564,N_16056,N_19413);
or UO_1565 (O_1565,N_17395,N_18450);
nor UO_1566 (O_1566,N_16081,N_16837);
or UO_1567 (O_1567,N_17391,N_17153);
and UO_1568 (O_1568,N_19173,N_18877);
xor UO_1569 (O_1569,N_17085,N_19782);
and UO_1570 (O_1570,N_16043,N_19481);
nor UO_1571 (O_1571,N_16480,N_17059);
nor UO_1572 (O_1572,N_19219,N_18418);
nand UO_1573 (O_1573,N_16467,N_19490);
nand UO_1574 (O_1574,N_16674,N_16482);
or UO_1575 (O_1575,N_17459,N_17780);
nand UO_1576 (O_1576,N_19731,N_17776);
and UO_1577 (O_1577,N_16520,N_19881);
or UO_1578 (O_1578,N_19111,N_18851);
nor UO_1579 (O_1579,N_17477,N_18908);
nor UO_1580 (O_1580,N_19253,N_17511);
or UO_1581 (O_1581,N_19720,N_19608);
xor UO_1582 (O_1582,N_18143,N_18171);
nand UO_1583 (O_1583,N_19440,N_19246);
xnor UO_1584 (O_1584,N_19452,N_19505);
nor UO_1585 (O_1585,N_17600,N_18701);
and UO_1586 (O_1586,N_19919,N_16607);
nor UO_1587 (O_1587,N_18539,N_16768);
nor UO_1588 (O_1588,N_16273,N_18912);
or UO_1589 (O_1589,N_19182,N_16474);
nor UO_1590 (O_1590,N_17552,N_16852);
and UO_1591 (O_1591,N_17244,N_16397);
nand UO_1592 (O_1592,N_17026,N_16301);
nand UO_1593 (O_1593,N_16420,N_19657);
nor UO_1594 (O_1594,N_16352,N_16223);
and UO_1595 (O_1595,N_17276,N_16702);
nand UO_1596 (O_1596,N_16317,N_18783);
nor UO_1597 (O_1597,N_18655,N_17332);
xnor UO_1598 (O_1598,N_17476,N_18155);
and UO_1599 (O_1599,N_17977,N_16342);
or UO_1600 (O_1600,N_17173,N_16960);
or UO_1601 (O_1601,N_17868,N_19274);
nand UO_1602 (O_1602,N_16192,N_19033);
and UO_1603 (O_1603,N_17184,N_18914);
nor UO_1604 (O_1604,N_18313,N_19874);
or UO_1605 (O_1605,N_16561,N_16796);
nand UO_1606 (O_1606,N_16547,N_18441);
or UO_1607 (O_1607,N_16391,N_19387);
nand UO_1608 (O_1608,N_16089,N_19677);
and UO_1609 (O_1609,N_19292,N_18683);
xor UO_1610 (O_1610,N_17538,N_17437);
and UO_1611 (O_1611,N_18000,N_18080);
and UO_1612 (O_1612,N_18479,N_19830);
and UO_1613 (O_1613,N_19766,N_16821);
and UO_1614 (O_1614,N_16845,N_16754);
xor UO_1615 (O_1615,N_17213,N_17917);
nand UO_1616 (O_1616,N_17264,N_17133);
and UO_1617 (O_1617,N_16110,N_17867);
nor UO_1618 (O_1618,N_18161,N_16879);
nor UO_1619 (O_1619,N_16382,N_16573);
and UO_1620 (O_1620,N_17145,N_19398);
nor UO_1621 (O_1621,N_18710,N_16460);
xnor UO_1622 (O_1622,N_17696,N_17170);
nand UO_1623 (O_1623,N_19109,N_16279);
nand UO_1624 (O_1624,N_16679,N_18157);
nand UO_1625 (O_1625,N_18817,N_18268);
and UO_1626 (O_1626,N_16793,N_19396);
and UO_1627 (O_1627,N_18388,N_17708);
or UO_1628 (O_1628,N_16423,N_16195);
and UO_1629 (O_1629,N_16389,N_18325);
or UO_1630 (O_1630,N_19119,N_16181);
nor UO_1631 (O_1631,N_17220,N_18439);
nor UO_1632 (O_1632,N_19211,N_17350);
nor UO_1633 (O_1633,N_18302,N_16447);
xor UO_1634 (O_1634,N_18264,N_17327);
nor UO_1635 (O_1635,N_16838,N_17597);
and UO_1636 (O_1636,N_18708,N_18137);
or UO_1637 (O_1637,N_16049,N_16418);
xor UO_1638 (O_1638,N_17697,N_18612);
and UO_1639 (O_1639,N_16244,N_17419);
nand UO_1640 (O_1640,N_16963,N_16401);
and UO_1641 (O_1641,N_19058,N_19206);
nand UO_1642 (O_1642,N_19953,N_19389);
or UO_1643 (O_1643,N_19069,N_16175);
or UO_1644 (O_1644,N_18452,N_16115);
or UO_1645 (O_1645,N_18847,N_17761);
nand UO_1646 (O_1646,N_19816,N_18142);
nor UO_1647 (O_1647,N_18734,N_18305);
xnor UO_1648 (O_1648,N_19708,N_17586);
or UO_1649 (O_1649,N_19914,N_17551);
or UO_1650 (O_1650,N_19944,N_19325);
nand UO_1651 (O_1651,N_19836,N_16902);
and UO_1652 (O_1652,N_16031,N_16699);
and UO_1653 (O_1653,N_17654,N_16867);
and UO_1654 (O_1654,N_16601,N_17483);
nor UO_1655 (O_1655,N_19861,N_16781);
nand UO_1656 (O_1656,N_19760,N_16558);
and UO_1657 (O_1657,N_16041,N_16250);
nor UO_1658 (O_1658,N_18739,N_18297);
xnor UO_1659 (O_1659,N_16116,N_17486);
or UO_1660 (O_1660,N_18093,N_16158);
nand UO_1661 (O_1661,N_18113,N_19070);
nand UO_1662 (O_1662,N_16001,N_17195);
nor UO_1663 (O_1663,N_17046,N_18259);
nand UO_1664 (O_1664,N_18755,N_16544);
and UO_1665 (O_1665,N_17667,N_16666);
and UO_1666 (O_1666,N_19950,N_17946);
or UO_1667 (O_1667,N_18149,N_16989);
and UO_1668 (O_1668,N_17549,N_19759);
nor UO_1669 (O_1669,N_19675,N_16638);
or UO_1670 (O_1670,N_18941,N_18200);
xor UO_1671 (O_1671,N_18746,N_18216);
or UO_1672 (O_1672,N_17806,N_16871);
nand UO_1673 (O_1673,N_18387,N_18357);
and UO_1674 (O_1674,N_18875,N_18438);
nor UO_1675 (O_1675,N_16309,N_19551);
and UO_1676 (O_1676,N_19668,N_16000);
nor UO_1677 (O_1677,N_17360,N_17779);
nor UO_1678 (O_1678,N_18831,N_19188);
and UO_1679 (O_1679,N_17821,N_16684);
nor UO_1680 (O_1680,N_19514,N_18879);
or UO_1681 (O_1681,N_16096,N_16270);
and UO_1682 (O_1682,N_18204,N_17781);
nor UO_1683 (O_1683,N_17928,N_16387);
nor UO_1684 (O_1684,N_16581,N_16672);
nor UO_1685 (O_1685,N_19178,N_16025);
nor UO_1686 (O_1686,N_16661,N_16637);
and UO_1687 (O_1687,N_19663,N_16678);
nor UO_1688 (O_1688,N_18861,N_19063);
or UO_1689 (O_1689,N_19960,N_16092);
and UO_1690 (O_1690,N_16477,N_19653);
or UO_1691 (O_1691,N_19916,N_16228);
nor UO_1692 (O_1692,N_16842,N_18266);
or UO_1693 (O_1693,N_17523,N_17150);
or UO_1694 (O_1694,N_19712,N_16271);
and UO_1695 (O_1695,N_19862,N_16797);
nor UO_1696 (O_1696,N_19886,N_16598);
xnor UO_1697 (O_1697,N_16327,N_16653);
nand UO_1698 (O_1698,N_19516,N_17257);
nand UO_1699 (O_1699,N_17341,N_17010);
nor UO_1700 (O_1700,N_19385,N_17379);
nand UO_1701 (O_1701,N_16994,N_18021);
nor UO_1702 (O_1702,N_17384,N_17560);
and UO_1703 (O_1703,N_19543,N_16788);
and UO_1704 (O_1704,N_19935,N_18812);
nor UO_1705 (O_1705,N_17724,N_16313);
xnor UO_1706 (O_1706,N_18363,N_17971);
nand UO_1707 (O_1707,N_18531,N_19230);
or UO_1708 (O_1708,N_18276,N_19808);
xnor UO_1709 (O_1709,N_18277,N_19203);
and UO_1710 (O_1710,N_18206,N_16810);
nand UO_1711 (O_1711,N_18939,N_19564);
xnor UO_1712 (O_1712,N_18801,N_19099);
nor UO_1713 (O_1713,N_19100,N_16061);
nand UO_1714 (O_1714,N_19344,N_16052);
or UO_1715 (O_1715,N_18223,N_18209);
nand UO_1716 (O_1716,N_18481,N_19205);
nor UO_1717 (O_1717,N_19306,N_17851);
or UO_1718 (O_1718,N_16691,N_17323);
and UO_1719 (O_1719,N_17698,N_18105);
nand UO_1720 (O_1720,N_18579,N_18527);
or UO_1721 (O_1721,N_17310,N_18575);
nand UO_1722 (O_1722,N_17689,N_18570);
and UO_1723 (O_1723,N_16546,N_17235);
or UO_1724 (O_1724,N_16129,N_17744);
and UO_1725 (O_1725,N_18880,N_17019);
and UO_1726 (O_1726,N_18659,N_18730);
nand UO_1727 (O_1727,N_19411,N_18946);
xnor UO_1728 (O_1728,N_19338,N_18521);
nand UO_1729 (O_1729,N_18370,N_17157);
nor UO_1730 (O_1730,N_16378,N_16848);
nor UO_1731 (O_1731,N_17788,N_17528);
nand UO_1732 (O_1732,N_19450,N_17131);
nand UO_1733 (O_1733,N_19588,N_17703);
nor UO_1734 (O_1734,N_16497,N_16145);
and UO_1735 (O_1735,N_18563,N_18281);
and UO_1736 (O_1736,N_16776,N_19871);
xnor UO_1737 (O_1737,N_18764,N_17811);
and UO_1738 (O_1738,N_16456,N_19226);
or UO_1739 (O_1739,N_19039,N_18602);
and UO_1740 (O_1740,N_16134,N_18483);
or UO_1741 (O_1741,N_18574,N_16437);
nand UO_1742 (O_1742,N_19034,N_17028);
and UO_1743 (O_1743,N_16483,N_18037);
nand UO_1744 (O_1744,N_17850,N_16459);
or UO_1745 (O_1745,N_17657,N_17286);
nor UO_1746 (O_1746,N_19351,N_16201);
and UO_1747 (O_1747,N_16877,N_19890);
nand UO_1748 (O_1748,N_19495,N_19265);
and UO_1749 (O_1749,N_18245,N_16166);
nor UO_1750 (O_1750,N_18125,N_18406);
xor UO_1751 (O_1751,N_17592,N_19877);
or UO_1752 (O_1752,N_16563,N_19684);
and UO_1753 (O_1753,N_18944,N_19482);
nand UO_1754 (O_1754,N_17862,N_17638);
and UO_1755 (O_1755,N_19180,N_17507);
or UO_1756 (O_1756,N_17580,N_16825);
or UO_1757 (O_1757,N_16395,N_16863);
or UO_1758 (O_1758,N_19580,N_19769);
nor UO_1759 (O_1759,N_19243,N_17759);
nand UO_1760 (O_1760,N_18307,N_19945);
or UO_1761 (O_1761,N_18408,N_16543);
xor UO_1762 (O_1762,N_17711,N_18002);
and UO_1763 (O_1763,N_16748,N_18999);
nor UO_1764 (O_1764,N_17349,N_18582);
and UO_1765 (O_1765,N_17570,N_18008);
nand UO_1766 (O_1766,N_16240,N_19421);
nand UO_1767 (O_1767,N_17895,N_19937);
nor UO_1768 (O_1768,N_19457,N_19811);
nor UO_1769 (O_1769,N_19198,N_16004);
nor UO_1770 (O_1770,N_16901,N_18358);
or UO_1771 (O_1771,N_17377,N_19356);
nor UO_1772 (O_1772,N_18146,N_19225);
nor UO_1773 (O_1773,N_19868,N_19797);
nor UO_1774 (O_1774,N_17529,N_16850);
nor UO_1775 (O_1775,N_17914,N_16704);
nor UO_1776 (O_1776,N_16298,N_17322);
nor UO_1777 (O_1777,N_19486,N_18850);
nor UO_1778 (O_1778,N_19006,N_19141);
nor UO_1779 (O_1779,N_16231,N_17423);
nand UO_1780 (O_1780,N_17445,N_19424);
nand UO_1781 (O_1781,N_16346,N_17210);
nand UO_1782 (O_1782,N_18491,N_19528);
and UO_1783 (O_1783,N_16649,N_18677);
nor UO_1784 (O_1784,N_19163,N_19023);
xor UO_1785 (O_1785,N_19355,N_16153);
or UO_1786 (O_1786,N_16070,N_18606);
nand UO_1787 (O_1787,N_19987,N_19941);
or UO_1788 (O_1788,N_16959,N_18956);
nor UO_1789 (O_1789,N_17804,N_19640);
or UO_1790 (O_1790,N_17015,N_18013);
nand UO_1791 (O_1791,N_16500,N_17554);
nand UO_1792 (O_1792,N_17675,N_17817);
and UO_1793 (O_1793,N_17390,N_18007);
xnor UO_1794 (O_1794,N_16722,N_16428);
nand UO_1795 (O_1795,N_18607,N_17297);
and UO_1796 (O_1796,N_18027,N_18822);
and UO_1797 (O_1797,N_17218,N_17536);
xnor UO_1798 (O_1798,N_16631,N_19094);
nand UO_1799 (O_1799,N_16008,N_18971);
and UO_1800 (O_1800,N_16566,N_16734);
or UO_1801 (O_1801,N_19575,N_19044);
and UO_1802 (O_1802,N_19470,N_17899);
nand UO_1803 (O_1803,N_18469,N_19600);
or UO_1804 (O_1804,N_19156,N_19694);
and UO_1805 (O_1805,N_16799,N_19097);
or UO_1806 (O_1806,N_16628,N_16152);
nand UO_1807 (O_1807,N_17985,N_19994);
nand UO_1808 (O_1808,N_16063,N_19171);
nor UO_1809 (O_1809,N_17539,N_17324);
nand UO_1810 (O_1810,N_19466,N_19402);
or UO_1811 (O_1811,N_17755,N_18466);
or UO_1812 (O_1812,N_17690,N_16736);
and UO_1813 (O_1813,N_19136,N_16411);
or UO_1814 (O_1814,N_19604,N_19077);
nor UO_1815 (O_1815,N_19660,N_18604);
or UO_1816 (O_1816,N_17884,N_18546);
and UO_1817 (O_1817,N_17808,N_17602);
nor UO_1818 (O_1818,N_16868,N_16593);
or UO_1819 (O_1819,N_18603,N_16432);
and UO_1820 (O_1820,N_18667,N_19112);
xor UO_1821 (O_1821,N_16763,N_17547);
nor UO_1822 (O_1822,N_19887,N_16024);
and UO_1823 (O_1823,N_17089,N_16013);
or UO_1824 (O_1824,N_19700,N_16760);
nor UO_1825 (O_1825,N_17512,N_17260);
nor UO_1826 (O_1826,N_16634,N_18611);
and UO_1827 (O_1827,N_17625,N_17493);
xor UO_1828 (O_1828,N_18833,N_17250);
and UO_1829 (O_1829,N_18196,N_19776);
or UO_1830 (O_1830,N_19250,N_18389);
and UO_1831 (O_1831,N_19636,N_16141);
nor UO_1832 (O_1832,N_18823,N_19488);
nand UO_1833 (O_1833,N_18136,N_18269);
and UO_1834 (O_1834,N_19473,N_17901);
and UO_1835 (O_1835,N_18016,N_17121);
nand UO_1836 (O_1836,N_19260,N_17358);
nor UO_1837 (O_1837,N_19644,N_18653);
nor UO_1838 (O_1838,N_16532,N_17710);
and UO_1839 (O_1839,N_16012,N_17599);
nand UO_1840 (O_1840,N_18910,N_19710);
nand UO_1841 (O_1841,N_16518,N_18750);
and UO_1842 (O_1842,N_19544,N_19324);
xor UO_1843 (O_1843,N_19368,N_18846);
nor UO_1844 (O_1844,N_16784,N_18057);
nand UO_1845 (O_1845,N_17001,N_19899);
and UO_1846 (O_1846,N_19625,N_18265);
or UO_1847 (O_1847,N_19582,N_16058);
nor UO_1848 (O_1848,N_19557,N_18651);
xnor UO_1849 (O_1849,N_19412,N_17462);
or UO_1850 (O_1850,N_19248,N_19734);
and UO_1851 (O_1851,N_17968,N_16554);
and UO_1852 (O_1852,N_16196,N_17686);
nor UO_1853 (O_1853,N_17271,N_16303);
nand UO_1854 (O_1854,N_16357,N_17593);
and UO_1855 (O_1855,N_18079,N_16778);
nor UO_1856 (O_1856,N_16981,N_18159);
or UO_1857 (O_1857,N_18592,N_16173);
nor UO_1858 (O_1858,N_19804,N_18565);
or UO_1859 (O_1859,N_18208,N_16656);
and UO_1860 (O_1860,N_18858,N_19297);
xor UO_1861 (O_1861,N_17557,N_16237);
or UO_1862 (O_1862,N_18515,N_16892);
nor UO_1863 (O_1863,N_17140,N_16665);
nor UO_1864 (O_1864,N_19725,N_18629);
nand UO_1865 (O_1865,N_19031,N_18194);
or UO_1866 (O_1866,N_16330,N_16381);
or UO_1867 (O_1867,N_19087,N_19724);
or UO_1868 (O_1868,N_19909,N_18719);
nand UO_1869 (O_1869,N_19615,N_17524);
or UO_1870 (O_1870,N_19240,N_18242);
or UO_1871 (O_1871,N_16498,N_19813);
or UO_1872 (O_1872,N_18869,N_17933);
nand UO_1873 (O_1873,N_19405,N_19847);
nand UO_1874 (O_1874,N_17793,N_16077);
nand UO_1875 (O_1875,N_16363,N_18174);
nand UO_1876 (O_1876,N_18145,N_17300);
or UO_1877 (O_1877,N_16773,N_17202);
xnor UO_1878 (O_1878,N_19026,N_16762);
nor UO_1879 (O_1879,N_18087,N_16329);
and UO_1880 (O_1880,N_17905,N_16685);
or UO_1881 (O_1881,N_18784,N_16723);
or UO_1882 (O_1882,N_16100,N_19721);
and UO_1883 (O_1883,N_19578,N_18476);
or UO_1884 (O_1884,N_18628,N_19833);
or UO_1885 (O_1885,N_16644,N_18144);
and UO_1886 (O_1886,N_17139,N_19386);
nand UO_1887 (O_1887,N_16531,N_18585);
nand UO_1888 (O_1888,N_17773,N_16936);
xor UO_1889 (O_1889,N_19468,N_16019);
nand UO_1890 (O_1890,N_17254,N_18705);
or UO_1891 (O_1891,N_16917,N_18726);
and UO_1892 (O_1892,N_18220,N_16230);
xnor UO_1893 (O_1893,N_16744,N_17802);
nor UO_1894 (O_1894,N_19762,N_19463);
nor UO_1895 (O_1895,N_18443,N_17193);
and UO_1896 (O_1896,N_17255,N_16431);
nand UO_1897 (O_1897,N_17466,N_17448);
nor UO_1898 (O_1898,N_18309,N_17084);
and UO_1899 (O_1899,N_16911,N_16484);
nand UO_1900 (O_1900,N_17962,N_16915);
nor UO_1901 (O_1901,N_18997,N_17839);
nand UO_1902 (O_1902,N_19624,N_17614);
or UO_1903 (O_1903,N_19014,N_19052);
nand UO_1904 (O_1904,N_19946,N_17819);
and UO_1905 (O_1905,N_16050,N_17993);
xor UO_1906 (O_1906,N_18386,N_18643);
nor UO_1907 (O_1907,N_18992,N_19915);
nor UO_1908 (O_1908,N_19342,N_19844);
or UO_1909 (O_1909,N_19840,N_17944);
nor UO_1910 (O_1910,N_18295,N_17114);
xnor UO_1911 (O_1911,N_19669,N_16194);
nor UO_1912 (O_1912,N_19870,N_18929);
or UO_1913 (O_1913,N_18326,N_16999);
xnor UO_1914 (O_1914,N_18032,N_16027);
or UO_1915 (O_1915,N_19970,N_17383);
and UO_1916 (O_1916,N_18472,N_19140);
and UO_1917 (O_1917,N_19918,N_18891);
nand UO_1918 (O_1918,N_19446,N_16292);
and UO_1919 (O_1919,N_18789,N_17904);
nand UO_1920 (O_1920,N_19038,N_18589);
and UO_1921 (O_1921,N_19105,N_18343);
nand UO_1922 (O_1922,N_17909,N_18399);
nand UO_1923 (O_1923,N_16197,N_16108);
and UO_1924 (O_1924,N_16930,N_17120);
and UO_1925 (O_1925,N_18114,N_18278);
nand UO_1926 (O_1926,N_17096,N_18374);
or UO_1927 (O_1927,N_16143,N_16083);
or UO_1928 (O_1928,N_18569,N_16595);
xor UO_1929 (O_1929,N_17660,N_16938);
or UO_1930 (O_1930,N_17470,N_18685);
and UO_1931 (O_1931,N_17299,N_18237);
nand UO_1932 (O_1932,N_18293,N_16307);
nor UO_1933 (O_1933,N_17115,N_17620);
xor UO_1934 (O_1934,N_18533,N_16064);
and UO_1935 (O_1935,N_19695,N_16633);
and UO_1936 (O_1936,N_16709,N_19183);
or UO_1937 (O_1937,N_18590,N_18922);
or UO_1938 (O_1938,N_17212,N_18696);
xnor UO_1939 (O_1939,N_17267,N_17373);
nor UO_1940 (O_1940,N_16731,N_18118);
and UO_1941 (O_1941,N_17453,N_17294);
nand UO_1942 (O_1942,N_18729,N_17185);
or UO_1943 (O_1943,N_16479,N_19191);
and UO_1944 (O_1944,N_19894,N_19630);
or UO_1945 (O_1945,N_18260,N_16545);
or UO_1946 (O_1946,N_17846,N_19217);
and UO_1947 (O_1947,N_19618,N_19606);
and UO_1948 (O_1948,N_18250,N_16914);
nor UO_1949 (O_1949,N_19984,N_19462);
nor UO_1950 (O_1950,N_16921,N_16186);
nand UO_1951 (O_1951,N_18299,N_18675);
xnor UO_1952 (O_1952,N_18076,N_18338);
nand UO_1953 (O_1953,N_18814,N_16137);
nor UO_1954 (O_1954,N_16809,N_16898);
nor UO_1955 (O_1955,N_18640,N_18320);
nand UO_1956 (O_1956,N_16406,N_19693);
nor UO_1957 (O_1957,N_18703,N_16882);
and UO_1958 (O_1958,N_19451,N_18808);
xnor UO_1959 (O_1959,N_16038,N_16386);
or UO_1960 (O_1960,N_16922,N_18936);
nand UO_1961 (O_1961,N_17298,N_19587);
xor UO_1962 (O_1962,N_17487,N_16511);
and UO_1963 (O_1963,N_16398,N_19688);
and UO_1964 (O_1964,N_19167,N_17022);
and UO_1965 (O_1965,N_19359,N_17467);
nor UO_1966 (O_1966,N_17677,N_18109);
nand UO_1967 (O_1967,N_16955,N_16427);
xor UO_1968 (O_1968,N_18666,N_18130);
or UO_1969 (O_1969,N_16322,N_19146);
nand UO_1970 (O_1970,N_16005,N_17166);
or UO_1971 (O_1971,N_17187,N_18549);
or UO_1972 (O_1972,N_16893,N_17902);
nand UO_1973 (O_1973,N_18942,N_17662);
xnor UO_1974 (O_1974,N_16097,N_19218);
or UO_1975 (O_1975,N_19852,N_18377);
or UO_1976 (O_1976,N_17367,N_18609);
nor UO_1977 (O_1977,N_19121,N_19417);
or UO_1978 (O_1978,N_18456,N_19554);
and UO_1979 (O_1979,N_16610,N_19016);
or UO_1980 (O_1980,N_16214,N_18900);
nand UO_1981 (O_1981,N_17417,N_17615);
nand UO_1982 (O_1982,N_16577,N_19391);
or UO_1983 (O_1983,N_18709,N_18398);
nor UO_1984 (O_1984,N_17200,N_17509);
or UO_1985 (O_1985,N_16182,N_18085);
nand UO_1986 (O_1986,N_18335,N_17720);
and UO_1987 (O_1987,N_16941,N_18821);
nor UO_1988 (O_1988,N_16807,N_18170);
nand UO_1989 (O_1989,N_16415,N_16393);
or UO_1990 (O_1990,N_17694,N_16516);
or UO_1991 (O_1991,N_19834,N_18392);
xnor UO_1992 (O_1992,N_18505,N_16549);
or UO_1993 (O_1993,N_19165,N_17285);
xnor UO_1994 (O_1994,N_18634,N_18839);
nor UO_1995 (O_1995,N_16248,N_18422);
xnor UO_1996 (O_1996,N_16200,N_19817);
nand UO_1997 (O_1997,N_17116,N_18015);
or UO_1998 (O_1998,N_19641,N_17475);
xor UO_1999 (O_1999,N_18178,N_16207);
and UO_2000 (O_2000,N_16975,N_19927);
and UO_2001 (O_2001,N_16789,N_19845);
and UO_2002 (O_2002,N_16368,N_17486);
or UO_2003 (O_2003,N_16842,N_18525);
and UO_2004 (O_2004,N_18533,N_17341);
nor UO_2005 (O_2005,N_18595,N_17259);
nand UO_2006 (O_2006,N_18254,N_19784);
or UO_2007 (O_2007,N_16990,N_19575);
and UO_2008 (O_2008,N_16870,N_17243);
nor UO_2009 (O_2009,N_18955,N_18231);
nand UO_2010 (O_2010,N_18792,N_19180);
nor UO_2011 (O_2011,N_17157,N_19232);
and UO_2012 (O_2012,N_19826,N_17574);
nor UO_2013 (O_2013,N_18069,N_19261);
nand UO_2014 (O_2014,N_17041,N_19324);
nor UO_2015 (O_2015,N_19211,N_16156);
nor UO_2016 (O_2016,N_16148,N_18815);
nand UO_2017 (O_2017,N_18767,N_18187);
or UO_2018 (O_2018,N_19217,N_19356);
and UO_2019 (O_2019,N_17868,N_18630);
nand UO_2020 (O_2020,N_18467,N_18318);
nor UO_2021 (O_2021,N_16103,N_19524);
and UO_2022 (O_2022,N_18255,N_17477);
or UO_2023 (O_2023,N_18694,N_19888);
nand UO_2024 (O_2024,N_17118,N_19630);
and UO_2025 (O_2025,N_17832,N_19395);
nand UO_2026 (O_2026,N_16917,N_16520);
and UO_2027 (O_2027,N_16128,N_19899);
nand UO_2028 (O_2028,N_17489,N_18907);
xnor UO_2029 (O_2029,N_19291,N_16897);
nand UO_2030 (O_2030,N_19220,N_17830);
or UO_2031 (O_2031,N_16254,N_16937);
and UO_2032 (O_2032,N_18852,N_18002);
or UO_2033 (O_2033,N_16037,N_19495);
nor UO_2034 (O_2034,N_16997,N_17252);
nand UO_2035 (O_2035,N_19372,N_18900);
nor UO_2036 (O_2036,N_16990,N_17064);
nand UO_2037 (O_2037,N_17980,N_18076);
xnor UO_2038 (O_2038,N_17857,N_16237);
xor UO_2039 (O_2039,N_18385,N_18215);
xor UO_2040 (O_2040,N_19263,N_18566);
or UO_2041 (O_2041,N_18115,N_19026);
nand UO_2042 (O_2042,N_18544,N_16282);
nor UO_2043 (O_2043,N_16079,N_17926);
or UO_2044 (O_2044,N_18807,N_19219);
and UO_2045 (O_2045,N_16726,N_17607);
xnor UO_2046 (O_2046,N_19717,N_16087);
and UO_2047 (O_2047,N_18641,N_16714);
or UO_2048 (O_2048,N_16930,N_19208);
or UO_2049 (O_2049,N_16489,N_16925);
nand UO_2050 (O_2050,N_17337,N_17591);
or UO_2051 (O_2051,N_17351,N_16709);
xor UO_2052 (O_2052,N_16140,N_18684);
xor UO_2053 (O_2053,N_18231,N_19213);
nor UO_2054 (O_2054,N_16071,N_18965);
nand UO_2055 (O_2055,N_18621,N_16434);
nand UO_2056 (O_2056,N_17081,N_18091);
nand UO_2057 (O_2057,N_17162,N_17432);
nand UO_2058 (O_2058,N_16749,N_17863);
xor UO_2059 (O_2059,N_19112,N_18976);
nor UO_2060 (O_2060,N_19071,N_18914);
or UO_2061 (O_2061,N_18058,N_18767);
or UO_2062 (O_2062,N_18081,N_16635);
nor UO_2063 (O_2063,N_18929,N_16339);
or UO_2064 (O_2064,N_17899,N_17794);
or UO_2065 (O_2065,N_19133,N_19675);
and UO_2066 (O_2066,N_16829,N_16261);
and UO_2067 (O_2067,N_19369,N_17412);
nand UO_2068 (O_2068,N_19043,N_16934);
or UO_2069 (O_2069,N_17144,N_17972);
and UO_2070 (O_2070,N_16002,N_16719);
and UO_2071 (O_2071,N_16539,N_18301);
and UO_2072 (O_2072,N_19147,N_18665);
xnor UO_2073 (O_2073,N_17961,N_16839);
and UO_2074 (O_2074,N_19864,N_18354);
and UO_2075 (O_2075,N_16128,N_16721);
nor UO_2076 (O_2076,N_18709,N_18108);
or UO_2077 (O_2077,N_19867,N_16277);
and UO_2078 (O_2078,N_17806,N_18190);
and UO_2079 (O_2079,N_19530,N_19658);
nor UO_2080 (O_2080,N_19220,N_18849);
or UO_2081 (O_2081,N_18014,N_18824);
and UO_2082 (O_2082,N_16896,N_17918);
nand UO_2083 (O_2083,N_18886,N_19683);
and UO_2084 (O_2084,N_18391,N_19585);
nor UO_2085 (O_2085,N_16684,N_17171);
and UO_2086 (O_2086,N_19416,N_16277);
or UO_2087 (O_2087,N_18321,N_17848);
nand UO_2088 (O_2088,N_18375,N_19205);
and UO_2089 (O_2089,N_16171,N_16761);
or UO_2090 (O_2090,N_18399,N_18179);
xnor UO_2091 (O_2091,N_18353,N_16826);
or UO_2092 (O_2092,N_18275,N_17011);
nand UO_2093 (O_2093,N_16011,N_17714);
nand UO_2094 (O_2094,N_17836,N_17245);
or UO_2095 (O_2095,N_16415,N_18025);
and UO_2096 (O_2096,N_17994,N_18498);
nand UO_2097 (O_2097,N_18750,N_18230);
and UO_2098 (O_2098,N_18958,N_18506);
or UO_2099 (O_2099,N_17739,N_19901);
and UO_2100 (O_2100,N_17616,N_19053);
and UO_2101 (O_2101,N_18490,N_16287);
and UO_2102 (O_2102,N_16010,N_17963);
nor UO_2103 (O_2103,N_19740,N_19034);
nand UO_2104 (O_2104,N_18334,N_18205);
or UO_2105 (O_2105,N_17278,N_18987);
and UO_2106 (O_2106,N_19081,N_19378);
xor UO_2107 (O_2107,N_19797,N_18004);
or UO_2108 (O_2108,N_16236,N_19335);
and UO_2109 (O_2109,N_19576,N_19741);
nand UO_2110 (O_2110,N_16787,N_19304);
or UO_2111 (O_2111,N_16084,N_19150);
nor UO_2112 (O_2112,N_16608,N_17982);
xnor UO_2113 (O_2113,N_19414,N_17368);
xor UO_2114 (O_2114,N_17345,N_18623);
nand UO_2115 (O_2115,N_17164,N_16125);
nor UO_2116 (O_2116,N_18006,N_16138);
or UO_2117 (O_2117,N_16804,N_17684);
or UO_2118 (O_2118,N_17479,N_17323);
xor UO_2119 (O_2119,N_16676,N_16587);
and UO_2120 (O_2120,N_18905,N_17485);
and UO_2121 (O_2121,N_19708,N_19953);
nand UO_2122 (O_2122,N_17855,N_18064);
or UO_2123 (O_2123,N_17999,N_19758);
nor UO_2124 (O_2124,N_18470,N_19118);
and UO_2125 (O_2125,N_17573,N_17925);
and UO_2126 (O_2126,N_18396,N_17120);
or UO_2127 (O_2127,N_16043,N_17917);
and UO_2128 (O_2128,N_18281,N_19111);
or UO_2129 (O_2129,N_16671,N_17487);
nand UO_2130 (O_2130,N_18829,N_16744);
and UO_2131 (O_2131,N_16753,N_18706);
xnor UO_2132 (O_2132,N_19807,N_19207);
or UO_2133 (O_2133,N_18628,N_16861);
and UO_2134 (O_2134,N_18918,N_19810);
and UO_2135 (O_2135,N_17154,N_18939);
nand UO_2136 (O_2136,N_16424,N_19747);
or UO_2137 (O_2137,N_17174,N_17577);
or UO_2138 (O_2138,N_16054,N_18053);
and UO_2139 (O_2139,N_19733,N_17188);
or UO_2140 (O_2140,N_19343,N_16862);
and UO_2141 (O_2141,N_19776,N_17317);
nand UO_2142 (O_2142,N_17610,N_17648);
nand UO_2143 (O_2143,N_17513,N_18833);
and UO_2144 (O_2144,N_18434,N_18898);
and UO_2145 (O_2145,N_19371,N_18054);
xor UO_2146 (O_2146,N_19571,N_17769);
nor UO_2147 (O_2147,N_16998,N_16505);
and UO_2148 (O_2148,N_19638,N_17046);
nor UO_2149 (O_2149,N_19015,N_19301);
and UO_2150 (O_2150,N_18563,N_17784);
xor UO_2151 (O_2151,N_17560,N_16623);
and UO_2152 (O_2152,N_16211,N_16715);
and UO_2153 (O_2153,N_17149,N_19621);
nand UO_2154 (O_2154,N_18597,N_17173);
nor UO_2155 (O_2155,N_16560,N_17837);
and UO_2156 (O_2156,N_18426,N_16532);
nor UO_2157 (O_2157,N_18489,N_18273);
nand UO_2158 (O_2158,N_18868,N_17023);
or UO_2159 (O_2159,N_18749,N_17726);
and UO_2160 (O_2160,N_19551,N_19937);
nand UO_2161 (O_2161,N_19232,N_17108);
and UO_2162 (O_2162,N_18318,N_19181);
nor UO_2163 (O_2163,N_17090,N_19919);
xor UO_2164 (O_2164,N_17603,N_18019);
nor UO_2165 (O_2165,N_19426,N_18720);
nand UO_2166 (O_2166,N_17774,N_16830);
nor UO_2167 (O_2167,N_18603,N_19793);
nor UO_2168 (O_2168,N_16458,N_19772);
nand UO_2169 (O_2169,N_17414,N_18971);
nand UO_2170 (O_2170,N_18070,N_17462);
nand UO_2171 (O_2171,N_18992,N_19913);
and UO_2172 (O_2172,N_17544,N_18820);
and UO_2173 (O_2173,N_16612,N_17144);
nor UO_2174 (O_2174,N_19538,N_18110);
or UO_2175 (O_2175,N_16548,N_16502);
and UO_2176 (O_2176,N_17047,N_18560);
nand UO_2177 (O_2177,N_17692,N_19609);
and UO_2178 (O_2178,N_19875,N_16962);
xor UO_2179 (O_2179,N_17220,N_19511);
and UO_2180 (O_2180,N_17869,N_18555);
nand UO_2181 (O_2181,N_18332,N_17091);
and UO_2182 (O_2182,N_17294,N_19565);
or UO_2183 (O_2183,N_18417,N_19155);
nand UO_2184 (O_2184,N_16719,N_16937);
nor UO_2185 (O_2185,N_18194,N_16638);
nor UO_2186 (O_2186,N_19260,N_16901);
nor UO_2187 (O_2187,N_17819,N_18597);
or UO_2188 (O_2188,N_18976,N_18249);
nand UO_2189 (O_2189,N_18961,N_19522);
nand UO_2190 (O_2190,N_19054,N_16745);
or UO_2191 (O_2191,N_18678,N_17162);
nand UO_2192 (O_2192,N_16358,N_19439);
and UO_2193 (O_2193,N_17493,N_19227);
nand UO_2194 (O_2194,N_19893,N_16457);
or UO_2195 (O_2195,N_18823,N_16162);
and UO_2196 (O_2196,N_17282,N_18908);
and UO_2197 (O_2197,N_16542,N_17823);
or UO_2198 (O_2198,N_16981,N_17780);
nand UO_2199 (O_2199,N_17161,N_16663);
or UO_2200 (O_2200,N_19016,N_19739);
nand UO_2201 (O_2201,N_18481,N_18049);
nand UO_2202 (O_2202,N_16804,N_16716);
or UO_2203 (O_2203,N_19145,N_19060);
or UO_2204 (O_2204,N_18716,N_17495);
or UO_2205 (O_2205,N_19021,N_17356);
nand UO_2206 (O_2206,N_17456,N_16907);
or UO_2207 (O_2207,N_18691,N_19292);
and UO_2208 (O_2208,N_19749,N_18710);
nand UO_2209 (O_2209,N_19068,N_17052);
xor UO_2210 (O_2210,N_16710,N_16550);
nor UO_2211 (O_2211,N_19701,N_18636);
and UO_2212 (O_2212,N_17482,N_16420);
or UO_2213 (O_2213,N_18845,N_17929);
nand UO_2214 (O_2214,N_18234,N_18241);
nand UO_2215 (O_2215,N_18598,N_16947);
xor UO_2216 (O_2216,N_18078,N_19826);
and UO_2217 (O_2217,N_16699,N_18202);
nand UO_2218 (O_2218,N_19852,N_17425);
nor UO_2219 (O_2219,N_17932,N_16287);
nor UO_2220 (O_2220,N_16422,N_17445);
and UO_2221 (O_2221,N_17679,N_17109);
nor UO_2222 (O_2222,N_19827,N_19717);
or UO_2223 (O_2223,N_18337,N_16029);
and UO_2224 (O_2224,N_18539,N_18039);
nor UO_2225 (O_2225,N_18105,N_18835);
nor UO_2226 (O_2226,N_18395,N_16299);
nand UO_2227 (O_2227,N_17654,N_17099);
and UO_2228 (O_2228,N_17611,N_19444);
nand UO_2229 (O_2229,N_16112,N_18417);
nand UO_2230 (O_2230,N_17279,N_19770);
nor UO_2231 (O_2231,N_18215,N_16575);
xnor UO_2232 (O_2232,N_19860,N_18608);
nand UO_2233 (O_2233,N_17905,N_18259);
nand UO_2234 (O_2234,N_18556,N_19464);
or UO_2235 (O_2235,N_17544,N_17877);
nor UO_2236 (O_2236,N_17938,N_19837);
and UO_2237 (O_2237,N_18452,N_18066);
and UO_2238 (O_2238,N_18878,N_17291);
or UO_2239 (O_2239,N_19657,N_19199);
xnor UO_2240 (O_2240,N_17988,N_17733);
nor UO_2241 (O_2241,N_16153,N_18555);
or UO_2242 (O_2242,N_17585,N_16477);
xnor UO_2243 (O_2243,N_16854,N_18442);
nand UO_2244 (O_2244,N_18121,N_18163);
and UO_2245 (O_2245,N_19660,N_19272);
and UO_2246 (O_2246,N_18681,N_18947);
or UO_2247 (O_2247,N_18698,N_19183);
nor UO_2248 (O_2248,N_17600,N_17839);
nand UO_2249 (O_2249,N_18389,N_17390);
or UO_2250 (O_2250,N_16498,N_18487);
or UO_2251 (O_2251,N_18326,N_18613);
nor UO_2252 (O_2252,N_19919,N_19471);
xnor UO_2253 (O_2253,N_16032,N_18960);
or UO_2254 (O_2254,N_16015,N_16395);
nand UO_2255 (O_2255,N_17324,N_18287);
and UO_2256 (O_2256,N_17758,N_17884);
or UO_2257 (O_2257,N_17086,N_16849);
nor UO_2258 (O_2258,N_19685,N_19206);
xor UO_2259 (O_2259,N_18267,N_19143);
and UO_2260 (O_2260,N_18875,N_19666);
nand UO_2261 (O_2261,N_18825,N_19623);
and UO_2262 (O_2262,N_16678,N_18131);
xnor UO_2263 (O_2263,N_16190,N_17937);
or UO_2264 (O_2264,N_18736,N_19807);
and UO_2265 (O_2265,N_16172,N_16515);
nor UO_2266 (O_2266,N_16847,N_18357);
nor UO_2267 (O_2267,N_18695,N_16994);
nand UO_2268 (O_2268,N_16311,N_17557);
nand UO_2269 (O_2269,N_18738,N_16837);
xnor UO_2270 (O_2270,N_16869,N_16148);
and UO_2271 (O_2271,N_17570,N_19366);
nor UO_2272 (O_2272,N_17879,N_19923);
nand UO_2273 (O_2273,N_19785,N_17791);
xnor UO_2274 (O_2274,N_16814,N_18718);
nand UO_2275 (O_2275,N_19833,N_19801);
nor UO_2276 (O_2276,N_18682,N_19932);
nand UO_2277 (O_2277,N_19790,N_17795);
and UO_2278 (O_2278,N_19648,N_17957);
nor UO_2279 (O_2279,N_18315,N_18707);
nand UO_2280 (O_2280,N_16797,N_18279);
nor UO_2281 (O_2281,N_17384,N_18261);
nand UO_2282 (O_2282,N_18212,N_18694);
nand UO_2283 (O_2283,N_16731,N_16689);
nand UO_2284 (O_2284,N_16174,N_17271);
xnor UO_2285 (O_2285,N_16418,N_18122);
xor UO_2286 (O_2286,N_17829,N_16156);
nand UO_2287 (O_2287,N_16846,N_16522);
or UO_2288 (O_2288,N_17125,N_17242);
and UO_2289 (O_2289,N_19145,N_17443);
nand UO_2290 (O_2290,N_19338,N_17896);
or UO_2291 (O_2291,N_18104,N_18563);
and UO_2292 (O_2292,N_18723,N_19023);
nand UO_2293 (O_2293,N_16046,N_19384);
or UO_2294 (O_2294,N_16214,N_19032);
nand UO_2295 (O_2295,N_17800,N_19405);
or UO_2296 (O_2296,N_16022,N_18216);
and UO_2297 (O_2297,N_16435,N_16152);
or UO_2298 (O_2298,N_17488,N_16872);
and UO_2299 (O_2299,N_17847,N_18496);
nand UO_2300 (O_2300,N_16328,N_16243);
and UO_2301 (O_2301,N_17881,N_17172);
nor UO_2302 (O_2302,N_16405,N_17255);
or UO_2303 (O_2303,N_17065,N_17881);
nor UO_2304 (O_2304,N_19001,N_19260);
nor UO_2305 (O_2305,N_16298,N_17804);
and UO_2306 (O_2306,N_19970,N_16019);
nand UO_2307 (O_2307,N_18067,N_18697);
xnor UO_2308 (O_2308,N_19689,N_17633);
xor UO_2309 (O_2309,N_17866,N_19617);
or UO_2310 (O_2310,N_17100,N_17378);
nor UO_2311 (O_2311,N_19868,N_17852);
or UO_2312 (O_2312,N_19879,N_18164);
and UO_2313 (O_2313,N_16825,N_16922);
nand UO_2314 (O_2314,N_19955,N_17286);
nand UO_2315 (O_2315,N_19327,N_17259);
nor UO_2316 (O_2316,N_19919,N_18127);
and UO_2317 (O_2317,N_19142,N_18305);
or UO_2318 (O_2318,N_19046,N_17718);
or UO_2319 (O_2319,N_18954,N_17640);
and UO_2320 (O_2320,N_19009,N_16019);
nand UO_2321 (O_2321,N_19715,N_19433);
nor UO_2322 (O_2322,N_18527,N_18904);
or UO_2323 (O_2323,N_18505,N_16947);
and UO_2324 (O_2324,N_16277,N_16335);
nor UO_2325 (O_2325,N_19289,N_17907);
or UO_2326 (O_2326,N_16610,N_16109);
nor UO_2327 (O_2327,N_19398,N_16703);
nor UO_2328 (O_2328,N_17412,N_18292);
xnor UO_2329 (O_2329,N_18031,N_17782);
xnor UO_2330 (O_2330,N_19566,N_18869);
nor UO_2331 (O_2331,N_18622,N_17047);
nor UO_2332 (O_2332,N_19742,N_18484);
nand UO_2333 (O_2333,N_19995,N_18116);
or UO_2334 (O_2334,N_16747,N_19030);
or UO_2335 (O_2335,N_17127,N_17949);
xor UO_2336 (O_2336,N_19284,N_17163);
or UO_2337 (O_2337,N_19613,N_19812);
nor UO_2338 (O_2338,N_18679,N_17159);
xnor UO_2339 (O_2339,N_19554,N_17305);
nand UO_2340 (O_2340,N_16110,N_19087);
xnor UO_2341 (O_2341,N_17675,N_16272);
and UO_2342 (O_2342,N_18165,N_17843);
and UO_2343 (O_2343,N_19975,N_16253);
and UO_2344 (O_2344,N_18473,N_19964);
and UO_2345 (O_2345,N_19821,N_19516);
or UO_2346 (O_2346,N_17446,N_19607);
nand UO_2347 (O_2347,N_17694,N_19495);
nor UO_2348 (O_2348,N_17539,N_18249);
or UO_2349 (O_2349,N_17131,N_16527);
nand UO_2350 (O_2350,N_16333,N_19589);
nor UO_2351 (O_2351,N_16535,N_19074);
nor UO_2352 (O_2352,N_19491,N_17829);
and UO_2353 (O_2353,N_19945,N_17735);
and UO_2354 (O_2354,N_17972,N_19760);
nor UO_2355 (O_2355,N_18521,N_18920);
nor UO_2356 (O_2356,N_18917,N_16928);
nand UO_2357 (O_2357,N_17747,N_19589);
xor UO_2358 (O_2358,N_18785,N_16004);
or UO_2359 (O_2359,N_17753,N_17289);
and UO_2360 (O_2360,N_19093,N_19282);
nand UO_2361 (O_2361,N_18513,N_16314);
or UO_2362 (O_2362,N_18283,N_17641);
nor UO_2363 (O_2363,N_17263,N_18455);
and UO_2364 (O_2364,N_19560,N_16286);
xor UO_2365 (O_2365,N_19958,N_19100);
or UO_2366 (O_2366,N_18843,N_18128);
nor UO_2367 (O_2367,N_17758,N_16312);
nor UO_2368 (O_2368,N_18258,N_16474);
nand UO_2369 (O_2369,N_16719,N_17950);
or UO_2370 (O_2370,N_17240,N_19754);
nor UO_2371 (O_2371,N_16121,N_17633);
xnor UO_2372 (O_2372,N_19263,N_19683);
nor UO_2373 (O_2373,N_17444,N_19242);
xnor UO_2374 (O_2374,N_18025,N_18651);
nand UO_2375 (O_2375,N_18884,N_19453);
nor UO_2376 (O_2376,N_17304,N_16818);
nand UO_2377 (O_2377,N_18876,N_16968);
nand UO_2378 (O_2378,N_19539,N_19832);
or UO_2379 (O_2379,N_18885,N_16138);
and UO_2380 (O_2380,N_18431,N_17934);
and UO_2381 (O_2381,N_17562,N_19422);
nor UO_2382 (O_2382,N_19990,N_16750);
and UO_2383 (O_2383,N_16198,N_19626);
nand UO_2384 (O_2384,N_19289,N_17181);
and UO_2385 (O_2385,N_19163,N_19963);
nand UO_2386 (O_2386,N_16445,N_17171);
nor UO_2387 (O_2387,N_18272,N_19268);
nand UO_2388 (O_2388,N_17864,N_18176);
or UO_2389 (O_2389,N_16246,N_17808);
and UO_2390 (O_2390,N_17110,N_17493);
nor UO_2391 (O_2391,N_19717,N_19260);
and UO_2392 (O_2392,N_17297,N_16569);
and UO_2393 (O_2393,N_16293,N_17650);
or UO_2394 (O_2394,N_17201,N_19525);
nand UO_2395 (O_2395,N_18919,N_19445);
nor UO_2396 (O_2396,N_19346,N_17381);
and UO_2397 (O_2397,N_18020,N_18904);
nor UO_2398 (O_2398,N_18031,N_16152);
nor UO_2399 (O_2399,N_18002,N_16009);
or UO_2400 (O_2400,N_16836,N_18232);
and UO_2401 (O_2401,N_19590,N_19626);
nand UO_2402 (O_2402,N_18237,N_16879);
and UO_2403 (O_2403,N_19196,N_19398);
nor UO_2404 (O_2404,N_19580,N_16006);
or UO_2405 (O_2405,N_19863,N_19538);
nor UO_2406 (O_2406,N_19270,N_17032);
or UO_2407 (O_2407,N_19761,N_16880);
nand UO_2408 (O_2408,N_19170,N_16572);
xor UO_2409 (O_2409,N_19270,N_18688);
or UO_2410 (O_2410,N_19485,N_19661);
and UO_2411 (O_2411,N_17045,N_16132);
nor UO_2412 (O_2412,N_17933,N_16488);
and UO_2413 (O_2413,N_18372,N_17101);
nor UO_2414 (O_2414,N_19153,N_17485);
or UO_2415 (O_2415,N_17979,N_18873);
or UO_2416 (O_2416,N_17536,N_16648);
nand UO_2417 (O_2417,N_17815,N_19856);
nor UO_2418 (O_2418,N_19512,N_19450);
nor UO_2419 (O_2419,N_17609,N_16846);
and UO_2420 (O_2420,N_19918,N_19084);
nand UO_2421 (O_2421,N_19956,N_16436);
xor UO_2422 (O_2422,N_16907,N_18540);
and UO_2423 (O_2423,N_19758,N_17158);
nand UO_2424 (O_2424,N_16110,N_18829);
nor UO_2425 (O_2425,N_17492,N_16255);
or UO_2426 (O_2426,N_17108,N_18898);
nand UO_2427 (O_2427,N_16381,N_19703);
nor UO_2428 (O_2428,N_19597,N_17688);
nor UO_2429 (O_2429,N_19506,N_16844);
and UO_2430 (O_2430,N_19583,N_17464);
nand UO_2431 (O_2431,N_18150,N_18417);
and UO_2432 (O_2432,N_18088,N_16841);
nor UO_2433 (O_2433,N_17330,N_18109);
or UO_2434 (O_2434,N_17210,N_16493);
xnor UO_2435 (O_2435,N_18777,N_19183);
or UO_2436 (O_2436,N_17806,N_16896);
and UO_2437 (O_2437,N_19393,N_18330);
nand UO_2438 (O_2438,N_19802,N_18230);
nor UO_2439 (O_2439,N_17190,N_16488);
nand UO_2440 (O_2440,N_18701,N_19653);
and UO_2441 (O_2441,N_18336,N_16448);
or UO_2442 (O_2442,N_16776,N_17309);
nor UO_2443 (O_2443,N_18473,N_17931);
nor UO_2444 (O_2444,N_17515,N_19527);
and UO_2445 (O_2445,N_16455,N_18271);
or UO_2446 (O_2446,N_18328,N_18555);
and UO_2447 (O_2447,N_19108,N_18973);
xnor UO_2448 (O_2448,N_19073,N_16011);
or UO_2449 (O_2449,N_16039,N_16848);
nor UO_2450 (O_2450,N_16311,N_19305);
and UO_2451 (O_2451,N_16868,N_16632);
nand UO_2452 (O_2452,N_19793,N_19949);
and UO_2453 (O_2453,N_16235,N_19319);
or UO_2454 (O_2454,N_19930,N_18939);
or UO_2455 (O_2455,N_19102,N_16586);
or UO_2456 (O_2456,N_18240,N_16997);
or UO_2457 (O_2457,N_17098,N_19687);
and UO_2458 (O_2458,N_16404,N_18859);
or UO_2459 (O_2459,N_16832,N_19082);
and UO_2460 (O_2460,N_19027,N_18116);
or UO_2461 (O_2461,N_19081,N_18008);
or UO_2462 (O_2462,N_17148,N_18405);
or UO_2463 (O_2463,N_19805,N_19280);
and UO_2464 (O_2464,N_19323,N_16024);
and UO_2465 (O_2465,N_16724,N_17840);
xnor UO_2466 (O_2466,N_18215,N_17443);
nand UO_2467 (O_2467,N_19217,N_19545);
xnor UO_2468 (O_2468,N_18709,N_19627);
or UO_2469 (O_2469,N_17498,N_17469);
nor UO_2470 (O_2470,N_17582,N_17347);
nand UO_2471 (O_2471,N_16819,N_16548);
xnor UO_2472 (O_2472,N_19272,N_19899);
and UO_2473 (O_2473,N_17974,N_19519);
nand UO_2474 (O_2474,N_16153,N_18028);
nor UO_2475 (O_2475,N_19082,N_16889);
and UO_2476 (O_2476,N_16309,N_18307);
or UO_2477 (O_2477,N_19967,N_16410);
xnor UO_2478 (O_2478,N_19562,N_16560);
and UO_2479 (O_2479,N_19642,N_17612);
or UO_2480 (O_2480,N_19396,N_16210);
nand UO_2481 (O_2481,N_16675,N_18747);
nand UO_2482 (O_2482,N_16583,N_18943);
xor UO_2483 (O_2483,N_16725,N_16313);
and UO_2484 (O_2484,N_18589,N_18210);
nand UO_2485 (O_2485,N_18447,N_16538);
and UO_2486 (O_2486,N_19681,N_19067);
nand UO_2487 (O_2487,N_16746,N_17173);
nor UO_2488 (O_2488,N_18274,N_19985);
or UO_2489 (O_2489,N_19487,N_19986);
nor UO_2490 (O_2490,N_17667,N_18060);
or UO_2491 (O_2491,N_17023,N_19375);
nand UO_2492 (O_2492,N_17093,N_16487);
nor UO_2493 (O_2493,N_16474,N_18317);
xnor UO_2494 (O_2494,N_18550,N_17720);
nor UO_2495 (O_2495,N_16036,N_17443);
or UO_2496 (O_2496,N_19893,N_19179);
xor UO_2497 (O_2497,N_19901,N_17526);
or UO_2498 (O_2498,N_17582,N_18062);
or UO_2499 (O_2499,N_16185,N_17871);
endmodule