module basic_1000_10000_1500_5_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
or U0 (N_0,In_778,In_591);
nand U1 (N_1,In_20,In_912);
nand U2 (N_2,In_586,In_397);
or U3 (N_3,In_109,In_982);
nor U4 (N_4,In_998,In_914);
or U5 (N_5,In_613,In_343);
nand U6 (N_6,In_913,In_240);
xnor U7 (N_7,In_715,In_774);
nand U8 (N_8,In_988,In_666);
nand U9 (N_9,In_130,In_156);
xor U10 (N_10,In_780,In_796);
xnor U11 (N_11,In_980,In_987);
nor U12 (N_12,In_274,In_733);
nand U13 (N_13,In_445,In_451);
nand U14 (N_14,In_436,In_635);
or U15 (N_15,In_937,In_55);
nor U16 (N_16,In_930,In_562);
xor U17 (N_17,In_655,In_814);
nor U18 (N_18,In_730,In_800);
and U19 (N_19,In_724,In_631);
xor U20 (N_20,In_720,In_753);
nand U21 (N_21,In_359,In_489);
nor U22 (N_22,In_381,In_515);
nor U23 (N_23,In_968,In_140);
nor U24 (N_24,In_483,In_79);
xor U25 (N_25,In_152,In_467);
or U26 (N_26,In_547,In_488);
nand U27 (N_27,In_554,In_447);
nor U28 (N_28,In_690,In_962);
nor U29 (N_29,In_16,In_194);
nand U30 (N_30,In_292,In_511);
xor U31 (N_31,In_165,In_854);
xor U32 (N_32,In_951,In_626);
or U33 (N_33,In_658,In_205);
or U34 (N_34,In_990,In_233);
or U35 (N_35,In_289,In_875);
nand U36 (N_36,In_97,In_934);
or U37 (N_37,In_563,In_369);
nor U38 (N_38,In_40,In_965);
xnor U39 (N_39,In_142,In_908);
or U40 (N_40,In_576,In_306);
nand U41 (N_41,In_199,In_475);
nand U42 (N_42,In_509,In_276);
nor U43 (N_43,In_559,In_405);
xor U44 (N_44,In_969,In_352);
xor U45 (N_45,In_1,In_820);
and U46 (N_46,In_776,In_763);
xor U47 (N_47,In_337,In_798);
nand U48 (N_48,In_593,In_725);
and U49 (N_49,In_261,In_956);
and U50 (N_50,In_13,In_944);
nor U51 (N_51,In_594,In_627);
or U52 (N_52,In_301,In_883);
nand U53 (N_53,In_450,In_887);
and U54 (N_54,In_510,In_967);
nand U55 (N_55,In_919,In_174);
or U56 (N_56,In_963,In_8);
xnor U57 (N_57,In_193,In_342);
xor U58 (N_58,In_191,In_374);
nand U59 (N_59,In_757,In_444);
or U60 (N_60,In_824,In_936);
and U61 (N_61,In_268,In_615);
and U62 (N_62,In_380,In_339);
or U63 (N_63,In_201,In_383);
and U64 (N_64,In_32,In_648);
and U65 (N_65,In_535,In_809);
and U66 (N_66,In_146,In_717);
and U67 (N_67,In_569,In_882);
nand U68 (N_68,In_611,In_411);
nand U69 (N_69,In_155,In_263);
nand U70 (N_70,In_441,In_65);
and U71 (N_71,In_435,In_151);
xnor U72 (N_72,In_417,In_42);
nand U73 (N_73,In_499,In_625);
or U74 (N_74,In_681,In_993);
and U75 (N_75,In_110,In_350);
nand U76 (N_76,In_644,In_366);
xnor U77 (N_77,In_66,In_312);
nand U78 (N_78,In_970,In_288);
nand U79 (N_79,In_362,In_822);
nand U80 (N_80,In_400,In_190);
nand U81 (N_81,In_920,In_685);
or U82 (N_82,In_552,In_196);
xor U83 (N_83,In_197,In_929);
nor U84 (N_84,In_797,In_222);
or U85 (N_85,In_113,In_791);
and U86 (N_86,In_863,In_885);
and U87 (N_87,In_916,In_154);
and U88 (N_88,In_884,In_255);
or U89 (N_89,In_293,In_57);
xnor U90 (N_90,In_888,In_474);
or U91 (N_91,In_587,In_530);
and U92 (N_92,In_748,In_759);
nand U93 (N_93,In_830,In_340);
nor U94 (N_94,In_101,In_957);
nand U95 (N_95,In_582,In_115);
and U96 (N_96,In_722,In_389);
and U97 (N_97,In_873,In_280);
nand U98 (N_98,In_198,In_786);
nand U99 (N_99,In_972,In_633);
xnor U100 (N_100,In_646,In_837);
xnor U101 (N_101,In_528,In_401);
nand U102 (N_102,In_418,In_758);
and U103 (N_103,In_950,In_899);
and U104 (N_104,In_567,In_457);
nor U105 (N_105,In_324,In_124);
nand U106 (N_106,In_501,In_213);
and U107 (N_107,In_247,In_54);
nor U108 (N_108,In_707,In_995);
xnor U109 (N_109,In_202,In_107);
or U110 (N_110,In_56,In_741);
xor U111 (N_111,In_895,In_902);
and U112 (N_112,In_866,In_727);
xor U113 (N_113,In_828,In_946);
nand U114 (N_114,In_807,In_241);
or U115 (N_115,In_657,In_82);
nand U116 (N_116,In_639,In_903);
or U117 (N_117,In_660,In_137);
nand U118 (N_118,In_461,In_938);
nand U119 (N_119,In_906,In_76);
xnor U120 (N_120,In_367,In_321);
and U121 (N_121,In_329,In_166);
xnor U122 (N_122,In_51,In_291);
or U123 (N_123,In_254,In_491);
nand U124 (N_124,In_439,In_48);
nand U125 (N_125,In_163,In_95);
or U126 (N_126,In_847,In_448);
or U127 (N_127,In_393,In_220);
nand U128 (N_128,In_585,In_67);
nand U129 (N_129,In_861,In_440);
xnor U130 (N_130,In_663,In_258);
nand U131 (N_131,In_710,In_355);
nand U132 (N_132,In_179,In_356);
or U133 (N_133,In_541,In_577);
nor U134 (N_134,In_652,In_465);
nor U135 (N_135,In_632,In_955);
nand U136 (N_136,In_766,In_572);
or U137 (N_137,In_556,In_286);
nor U138 (N_138,In_395,In_848);
or U139 (N_139,In_75,In_413);
and U140 (N_140,In_207,In_564);
and U141 (N_141,In_463,In_93);
xnor U142 (N_142,In_169,In_905);
or U143 (N_143,In_846,In_821);
nand U144 (N_144,In_573,In_159);
or U145 (N_145,In_309,In_87);
nand U146 (N_146,In_296,In_53);
nand U147 (N_147,In_9,In_102);
nor U148 (N_148,In_571,In_38);
nor U149 (N_149,In_894,In_546);
nor U150 (N_150,In_864,In_98);
or U151 (N_151,In_496,In_415);
or U152 (N_152,In_466,In_813);
or U153 (N_153,In_772,In_495);
or U154 (N_154,In_749,In_616);
xnor U155 (N_155,In_600,In_334);
and U156 (N_156,In_880,In_295);
xor U157 (N_157,In_227,In_624);
or U158 (N_158,In_376,In_925);
and U159 (N_159,In_224,In_214);
or U160 (N_160,In_302,In_328);
or U161 (N_161,In_867,In_699);
or U162 (N_162,In_71,In_891);
xnor U163 (N_163,In_520,In_674);
and U164 (N_164,In_898,In_747);
and U165 (N_165,In_331,In_931);
nand U166 (N_166,In_7,In_349);
xor U167 (N_167,In_206,In_519);
or U168 (N_168,In_384,In_935);
xnor U169 (N_169,In_117,In_294);
nor U170 (N_170,In_396,In_765);
and U171 (N_171,In_2,In_596);
nor U172 (N_172,In_271,In_503);
nand U173 (N_173,In_456,In_819);
nor U174 (N_174,In_915,In_428);
xnor U175 (N_175,In_618,In_529);
nand U176 (N_176,In_365,In_39);
and U177 (N_177,In_63,In_917);
and U178 (N_178,In_278,In_126);
and U179 (N_179,In_602,In_816);
nand U180 (N_180,In_574,In_852);
nand U181 (N_181,In_364,In_592);
or U182 (N_182,In_147,In_997);
nor U183 (N_183,In_645,In_422);
and U184 (N_184,In_740,In_752);
nor U185 (N_185,In_77,In_92);
or U186 (N_186,In_327,In_85);
or U187 (N_187,In_104,In_125);
nor U188 (N_188,In_948,In_728);
xnor U189 (N_189,In_120,In_354);
xnor U190 (N_190,In_810,In_595);
and U191 (N_191,In_210,In_536);
and U192 (N_192,In_277,In_811);
and U193 (N_193,In_701,In_881);
nor U194 (N_194,In_886,In_494);
or U195 (N_195,In_808,In_656);
nand U196 (N_196,In_285,In_392);
and U197 (N_197,In_253,In_832);
or U198 (N_198,In_472,In_344);
and U199 (N_199,In_675,In_314);
nand U200 (N_200,In_500,In_538);
xnor U201 (N_201,In_485,In_22);
nor U202 (N_202,In_187,In_838);
nor U203 (N_203,In_144,In_792);
nand U204 (N_204,In_942,In_234);
xnor U205 (N_205,In_802,In_532);
nor U206 (N_206,In_298,In_437);
nand U207 (N_207,In_490,In_922);
and U208 (N_208,In_901,In_839);
or U209 (N_209,In_88,In_226);
or U210 (N_210,In_818,In_319);
xor U211 (N_211,In_357,In_427);
and U212 (N_212,In_578,In_412);
nand U213 (N_213,In_70,In_527);
nand U214 (N_214,In_99,In_111);
nand U215 (N_215,In_696,In_406);
xor U216 (N_216,In_96,In_236);
and U217 (N_217,In_812,In_353);
xnor U218 (N_218,In_691,In_743);
or U219 (N_219,In_332,In_985);
and U220 (N_220,In_398,In_745);
xnor U221 (N_221,In_219,In_709);
or U222 (N_222,In_770,In_284);
and U223 (N_223,In_471,In_131);
and U224 (N_224,In_108,In_269);
and U225 (N_225,In_348,In_341);
nor U226 (N_226,In_148,In_548);
nand U227 (N_227,In_761,In_960);
nand U228 (N_228,In_735,In_24);
nand U229 (N_229,In_172,In_620);
nand U230 (N_230,In_26,In_473);
nand U231 (N_231,In_134,In_928);
xor U232 (N_232,In_505,In_50);
xnor U233 (N_233,In_686,In_958);
nor U234 (N_234,In_550,In_744);
nor U235 (N_235,In_370,In_647);
nor U236 (N_236,In_754,In_175);
xnor U237 (N_237,In_636,In_755);
nor U238 (N_238,In_638,In_713);
or U239 (N_239,In_23,In_316);
or U240 (N_240,In_221,In_333);
nand U241 (N_241,In_78,In_670);
and U242 (N_242,In_856,In_242);
nor U243 (N_243,In_539,In_927);
and U244 (N_244,In_892,In_94);
xor U245 (N_245,In_208,In_850);
nand U246 (N_246,In_617,In_414);
xnor U247 (N_247,In_588,In_464);
xnor U248 (N_248,In_843,In_878);
or U249 (N_249,In_599,In_363);
nand U250 (N_250,In_999,In_371);
nand U251 (N_251,In_751,In_317);
nor U252 (N_252,In_303,In_844);
and U253 (N_253,In_664,In_659);
nand U254 (N_254,In_143,In_229);
xor U255 (N_255,In_768,In_83);
nand U256 (N_256,In_662,In_653);
xor U257 (N_257,In_952,In_521);
and U258 (N_258,In_185,In_607);
nand U259 (N_259,In_61,In_114);
nand U260 (N_260,In_424,In_932);
or U261 (N_261,In_228,In_265);
and U262 (N_262,In_799,In_943);
or U263 (N_263,In_281,In_801);
or U264 (N_264,In_129,In_345);
and U265 (N_265,In_477,In_216);
and U266 (N_266,In_641,In_320);
xnor U267 (N_267,In_218,In_103);
nand U268 (N_268,In_35,In_589);
nand U269 (N_269,In_158,In_118);
or U270 (N_270,In_267,In_991);
xor U271 (N_271,In_795,In_37);
or U272 (N_272,In_983,In_391);
nor U273 (N_273,In_453,In_835);
nor U274 (N_274,In_608,In_27);
nor U275 (N_275,In_966,In_698);
nand U276 (N_276,In_858,In_30);
nor U277 (N_277,In_251,In_106);
and U278 (N_278,In_336,In_910);
nand U279 (N_279,In_697,In_257);
nand U280 (N_280,In_570,In_84);
and U281 (N_281,In_394,In_784);
or U282 (N_282,In_678,In_823);
nand U283 (N_283,In_700,In_432);
nand U284 (N_284,In_726,In_283);
nand U285 (N_285,In_29,In_523);
and U286 (N_286,In_89,In_311);
nand U287 (N_287,In_650,In_403);
nand U288 (N_288,In_971,In_868);
xnor U289 (N_289,In_734,In_679);
nand U290 (N_290,In_924,In_803);
nor U291 (N_291,In_454,In_918);
xor U292 (N_292,In_209,In_695);
nand U293 (N_293,In_513,In_731);
nand U294 (N_294,In_945,In_525);
and U295 (N_295,In_176,In_788);
xor U296 (N_296,In_44,In_273);
and U297 (N_297,In_954,In_211);
nor U298 (N_298,In_637,In_462);
nor U299 (N_299,In_430,In_45);
nor U300 (N_300,In_649,In_497);
nand U301 (N_301,In_794,In_90);
xnor U302 (N_302,In_323,In_634);
or U303 (N_303,In_272,In_180);
nor U304 (N_304,In_673,In_904);
nand U305 (N_305,In_192,In_58);
nand U306 (N_306,In_896,In_455);
xnor U307 (N_307,In_771,In_677);
nor U308 (N_308,In_718,In_590);
nand U309 (N_309,In_153,In_994);
and U310 (N_310,In_609,In_189);
and U311 (N_311,In_729,In_708);
xor U312 (N_312,In_669,In_979);
and U313 (N_313,In_874,In_390);
nand U314 (N_314,In_237,In_167);
and U315 (N_315,In_119,In_533);
or U316 (N_316,In_893,In_705);
nor U317 (N_317,In_420,In_12);
nand U318 (N_318,In_246,In_575);
xor U319 (N_319,In_826,In_584);
or U320 (N_320,In_122,In_672);
xor U321 (N_321,In_60,In_668);
or U322 (N_322,In_351,In_760);
nor U323 (N_323,In_890,In_978);
and U324 (N_324,In_325,In_827);
and U325 (N_325,In_643,In_28);
or U326 (N_326,In_642,In_481);
xor U327 (N_327,In_825,In_121);
nor U328 (N_328,In_235,In_361);
and U329 (N_329,In_502,In_157);
nor U330 (N_330,In_33,In_841);
or U331 (N_331,In_671,In_711);
or U332 (N_332,In_526,In_865);
nor U333 (N_333,In_326,In_851);
and U334 (N_334,In_68,In_31);
nand U335 (N_335,In_41,In_565);
xor U336 (N_336,In_833,In_19);
and U337 (N_337,In_81,In_248);
and U338 (N_338,In_429,In_750);
xor U339 (N_339,In_560,In_4);
or U340 (N_340,In_112,In_181);
xnor U341 (N_341,In_603,In_249);
and U342 (N_342,In_493,In_382);
and U343 (N_343,In_402,In_279);
xor U344 (N_344,In_716,In_540);
and U345 (N_345,In_168,In_46);
and U346 (N_346,In_80,In_133);
nor U347 (N_347,In_162,In_426);
xnor U348 (N_348,In_597,In_872);
and U349 (N_349,In_419,In_262);
and U350 (N_350,In_777,In_47);
xor U351 (N_351,In_178,In_375);
nand U352 (N_352,In_34,In_0);
or U353 (N_353,In_399,In_684);
or U354 (N_354,In_287,In_409);
nor U355 (N_355,In_787,In_225);
nor U356 (N_356,In_446,In_416);
xor U357 (N_357,In_25,In_64);
or U358 (N_358,In_531,In_443);
or U359 (N_359,In_223,In_598);
and U360 (N_360,In_621,In_388);
nor U361 (N_361,In_842,In_692);
xnor U362 (N_362,In_537,In_845);
xor U363 (N_363,In_857,In_512);
and U364 (N_364,In_407,In_186);
xnor U365 (N_365,In_996,In_762);
xor U366 (N_366,In_358,In_719);
xor U367 (N_367,In_315,In_171);
nand U368 (N_368,In_859,In_127);
or U369 (N_369,In_425,In_3);
xnor U370 (N_370,In_612,In_378);
or U371 (N_371,In_478,In_373);
and U372 (N_372,In_543,In_313);
or U373 (N_373,In_853,In_610);
and U374 (N_374,In_974,In_785);
and U375 (N_375,In_940,In_732);
and U376 (N_376,In_136,In_651);
and U377 (N_377,In_551,In_877);
xnor U378 (N_378,In_693,In_184);
nor U379 (N_379,In_712,In_738);
nor U380 (N_380,In_583,In_11);
nor U381 (N_381,In_486,In_69);
or U382 (N_382,In_909,In_561);
or U383 (N_383,In_230,In_487);
nor U384 (N_384,In_911,In_270);
and U385 (N_385,In_173,In_682);
or U386 (N_386,In_6,In_15);
xor U387 (N_387,In_300,In_264);
nor U388 (N_388,In_479,In_806);
and U389 (N_389,In_900,In_135);
or U390 (N_390,In_275,In_452);
and U391 (N_391,In_74,In_266);
or U392 (N_392,In_123,In_975);
nand U393 (N_393,In_683,In_132);
or U394 (N_394,In_204,In_542);
xnor U395 (N_395,In_177,In_150);
or U396 (N_396,In_601,In_756);
nand U397 (N_397,In_161,In_423);
or U398 (N_398,In_238,In_933);
xnor U399 (N_399,In_62,In_769);
xor U400 (N_400,In_862,In_976);
or U401 (N_401,In_630,In_897);
xor U402 (N_402,In_665,In_195);
and U403 (N_403,In_307,In_188);
and U404 (N_404,In_18,In_516);
xnor U405 (N_405,In_746,In_183);
nor U406 (N_406,In_484,In_459);
nand U407 (N_407,In_322,In_433);
xnor U408 (N_408,In_986,In_580);
or U409 (N_409,In_524,In_953);
or U410 (N_410,In_73,In_805);
or U411 (N_411,In_939,In_581);
and U412 (N_412,In_921,In_368);
nand U413 (N_413,In_470,In_386);
and U414 (N_414,In_245,In_579);
nand U415 (N_415,In_767,In_139);
and U416 (N_416,In_304,In_687);
nand U417 (N_417,In_605,In_779);
xnor U418 (N_418,In_310,In_517);
nand U419 (N_419,In_492,In_829);
and U420 (N_420,In_871,In_703);
or U421 (N_421,In_14,In_721);
xor U422 (N_422,In_318,In_989);
and U423 (N_423,In_654,In_566);
nand U424 (N_424,In_973,In_545);
xor U425 (N_425,In_105,In_256);
nand U426 (N_426,In_522,In_667);
or U427 (N_427,In_508,In_421);
nor U428 (N_428,In_141,In_387);
or U429 (N_429,In_804,In_714);
nor U430 (N_430,In_377,In_379);
or U431 (N_431,In_72,In_408);
nand U432 (N_432,In_568,In_476);
nand U433 (N_433,In_790,In_640);
or U434 (N_434,In_59,In_855);
or U435 (N_435,In_460,In_783);
or U436 (N_436,In_17,In_623);
and U437 (N_437,In_555,In_498);
xnor U438 (N_438,In_116,In_21);
and U439 (N_439,In_959,In_789);
or U440 (N_440,In_468,In_149);
xnor U441 (N_441,In_212,In_250);
or U442 (N_442,In_629,In_438);
nand U443 (N_443,In_434,In_145);
nand U444 (N_444,In_338,In_372);
nand U445 (N_445,In_518,In_614);
and U446 (N_446,In_290,In_5);
nand U447 (N_447,In_308,In_992);
or U448 (N_448,In_544,In_330);
nand U449 (N_449,In_817,In_764);
nor U450 (N_450,In_182,In_549);
or U451 (N_451,In_244,In_964);
xor U452 (N_452,In_680,In_782);
xor U453 (N_453,In_299,In_619);
or U454 (N_454,In_203,In_243);
nor U455 (N_455,In_981,In_217);
nand U456 (N_456,In_507,In_442);
or U457 (N_457,In_941,In_604);
and U458 (N_458,In_449,In_977);
or U459 (N_459,In_431,In_252);
xor U460 (N_460,In_360,In_160);
and U461 (N_461,In_949,In_534);
nor U462 (N_462,In_737,In_706);
nor U463 (N_463,In_773,In_704);
nand U464 (N_464,In_128,In_480);
and U465 (N_465,In_138,In_723);
or U466 (N_466,In_849,In_926);
and U467 (N_467,In_49,In_10);
nand U468 (N_468,In_907,In_781);
nor U469 (N_469,In_688,In_558);
nand U470 (N_470,In_834,In_506);
nand U471 (N_471,In_458,In_260);
nor U472 (N_472,In_231,In_876);
and U473 (N_473,In_482,In_504);
nand U474 (N_474,In_889,In_661);
nand U475 (N_475,In_742,In_239);
nor U476 (N_476,In_831,In_232);
nor U477 (N_477,In_689,In_385);
nand U478 (N_478,In_200,In_622);
and U479 (N_479,In_346,In_305);
nor U480 (N_480,In_694,In_86);
nor U481 (N_481,In_961,In_984);
nor U482 (N_482,In_793,In_947);
xor U483 (N_483,In_347,In_775);
nand U484 (N_484,In_282,In_739);
nor U485 (N_485,In_52,In_836);
nand U486 (N_486,In_170,In_469);
nand U487 (N_487,In_410,In_259);
nor U488 (N_488,In_676,In_36);
and U489 (N_489,In_702,In_164);
xor U490 (N_490,In_869,In_215);
and U491 (N_491,In_557,In_335);
or U492 (N_492,In_860,In_840);
and U493 (N_493,In_923,In_100);
or U494 (N_494,In_815,In_91);
xnor U495 (N_495,In_879,In_606);
or U496 (N_496,In_297,In_628);
or U497 (N_497,In_736,In_404);
xor U498 (N_498,In_553,In_870);
xor U499 (N_499,In_514,In_43);
and U500 (N_500,In_457,In_785);
xor U501 (N_501,In_585,In_309);
nor U502 (N_502,In_393,In_497);
nor U503 (N_503,In_157,In_868);
or U504 (N_504,In_543,In_408);
xnor U505 (N_505,In_513,In_785);
xnor U506 (N_506,In_113,In_249);
nor U507 (N_507,In_917,In_342);
nand U508 (N_508,In_692,In_105);
nand U509 (N_509,In_678,In_728);
xnor U510 (N_510,In_885,In_687);
xor U511 (N_511,In_661,In_121);
or U512 (N_512,In_90,In_150);
nor U513 (N_513,In_510,In_444);
and U514 (N_514,In_120,In_570);
and U515 (N_515,In_814,In_572);
and U516 (N_516,In_597,In_213);
xnor U517 (N_517,In_147,In_578);
xnor U518 (N_518,In_611,In_979);
or U519 (N_519,In_325,In_244);
nand U520 (N_520,In_123,In_557);
nor U521 (N_521,In_828,In_402);
nand U522 (N_522,In_194,In_297);
and U523 (N_523,In_52,In_834);
nand U524 (N_524,In_610,In_67);
nor U525 (N_525,In_909,In_395);
or U526 (N_526,In_654,In_202);
xnor U527 (N_527,In_860,In_129);
or U528 (N_528,In_489,In_532);
or U529 (N_529,In_180,In_945);
xnor U530 (N_530,In_220,In_208);
and U531 (N_531,In_53,In_61);
nand U532 (N_532,In_513,In_35);
xor U533 (N_533,In_437,In_287);
or U534 (N_534,In_840,In_859);
and U535 (N_535,In_618,In_563);
and U536 (N_536,In_637,In_474);
nand U537 (N_537,In_688,In_263);
or U538 (N_538,In_856,In_388);
or U539 (N_539,In_839,In_682);
or U540 (N_540,In_9,In_383);
and U541 (N_541,In_935,In_718);
and U542 (N_542,In_976,In_765);
or U543 (N_543,In_84,In_976);
or U544 (N_544,In_995,In_973);
or U545 (N_545,In_925,In_371);
and U546 (N_546,In_35,In_440);
nor U547 (N_547,In_515,In_206);
nor U548 (N_548,In_782,In_622);
and U549 (N_549,In_42,In_0);
nand U550 (N_550,In_517,In_868);
or U551 (N_551,In_496,In_180);
nor U552 (N_552,In_867,In_255);
xnor U553 (N_553,In_135,In_63);
xor U554 (N_554,In_175,In_893);
nor U555 (N_555,In_71,In_376);
nand U556 (N_556,In_619,In_122);
or U557 (N_557,In_741,In_995);
xor U558 (N_558,In_244,In_67);
or U559 (N_559,In_42,In_490);
or U560 (N_560,In_409,In_391);
nand U561 (N_561,In_73,In_750);
nor U562 (N_562,In_699,In_694);
or U563 (N_563,In_504,In_108);
or U564 (N_564,In_567,In_538);
or U565 (N_565,In_52,In_157);
or U566 (N_566,In_934,In_224);
and U567 (N_567,In_304,In_484);
or U568 (N_568,In_259,In_338);
and U569 (N_569,In_973,In_601);
and U570 (N_570,In_790,In_435);
nand U571 (N_571,In_766,In_498);
nand U572 (N_572,In_484,In_818);
xor U573 (N_573,In_169,In_27);
xor U574 (N_574,In_975,In_47);
nor U575 (N_575,In_611,In_213);
nor U576 (N_576,In_987,In_14);
and U577 (N_577,In_682,In_299);
and U578 (N_578,In_420,In_523);
nor U579 (N_579,In_633,In_534);
or U580 (N_580,In_800,In_476);
xnor U581 (N_581,In_261,In_966);
nor U582 (N_582,In_635,In_50);
and U583 (N_583,In_133,In_322);
and U584 (N_584,In_154,In_351);
xor U585 (N_585,In_73,In_644);
or U586 (N_586,In_767,In_93);
nand U587 (N_587,In_189,In_622);
nor U588 (N_588,In_699,In_14);
xnor U589 (N_589,In_333,In_159);
nor U590 (N_590,In_728,In_475);
and U591 (N_591,In_613,In_549);
nor U592 (N_592,In_409,In_374);
nand U593 (N_593,In_542,In_103);
and U594 (N_594,In_894,In_70);
or U595 (N_595,In_225,In_747);
nand U596 (N_596,In_71,In_123);
nand U597 (N_597,In_407,In_896);
xor U598 (N_598,In_388,In_252);
or U599 (N_599,In_876,In_460);
xnor U600 (N_600,In_178,In_587);
or U601 (N_601,In_448,In_864);
or U602 (N_602,In_750,In_673);
xor U603 (N_603,In_297,In_451);
nor U604 (N_604,In_596,In_293);
and U605 (N_605,In_642,In_774);
and U606 (N_606,In_795,In_248);
nand U607 (N_607,In_885,In_459);
or U608 (N_608,In_780,In_668);
xnor U609 (N_609,In_662,In_383);
xnor U610 (N_610,In_792,In_609);
nand U611 (N_611,In_599,In_844);
or U612 (N_612,In_288,In_863);
xnor U613 (N_613,In_644,In_72);
xor U614 (N_614,In_665,In_624);
nor U615 (N_615,In_467,In_715);
or U616 (N_616,In_954,In_352);
xor U617 (N_617,In_526,In_351);
nand U618 (N_618,In_724,In_313);
and U619 (N_619,In_787,In_702);
nor U620 (N_620,In_545,In_286);
xnor U621 (N_621,In_221,In_957);
xor U622 (N_622,In_502,In_455);
and U623 (N_623,In_3,In_292);
and U624 (N_624,In_200,In_746);
or U625 (N_625,In_682,In_69);
and U626 (N_626,In_660,In_383);
nor U627 (N_627,In_69,In_367);
nand U628 (N_628,In_944,In_561);
nand U629 (N_629,In_913,In_743);
and U630 (N_630,In_652,In_776);
or U631 (N_631,In_635,In_314);
or U632 (N_632,In_475,In_511);
nand U633 (N_633,In_906,In_818);
or U634 (N_634,In_649,In_443);
xnor U635 (N_635,In_257,In_468);
xnor U636 (N_636,In_714,In_92);
xnor U637 (N_637,In_458,In_917);
xor U638 (N_638,In_15,In_134);
nor U639 (N_639,In_325,In_360);
nand U640 (N_640,In_481,In_464);
or U641 (N_641,In_296,In_136);
nand U642 (N_642,In_49,In_878);
nand U643 (N_643,In_768,In_76);
xor U644 (N_644,In_755,In_98);
nand U645 (N_645,In_701,In_81);
nor U646 (N_646,In_439,In_871);
nor U647 (N_647,In_507,In_571);
or U648 (N_648,In_820,In_866);
nor U649 (N_649,In_126,In_855);
nor U650 (N_650,In_713,In_173);
and U651 (N_651,In_26,In_425);
xnor U652 (N_652,In_296,In_946);
nor U653 (N_653,In_650,In_247);
nand U654 (N_654,In_172,In_917);
or U655 (N_655,In_387,In_741);
xor U656 (N_656,In_264,In_734);
or U657 (N_657,In_718,In_449);
nor U658 (N_658,In_690,In_350);
xnor U659 (N_659,In_495,In_22);
xor U660 (N_660,In_48,In_549);
and U661 (N_661,In_437,In_480);
xnor U662 (N_662,In_352,In_754);
xnor U663 (N_663,In_286,In_734);
xor U664 (N_664,In_235,In_970);
xor U665 (N_665,In_482,In_869);
nand U666 (N_666,In_25,In_665);
xnor U667 (N_667,In_851,In_399);
or U668 (N_668,In_236,In_87);
and U669 (N_669,In_610,In_438);
xor U670 (N_670,In_926,In_834);
or U671 (N_671,In_930,In_546);
xor U672 (N_672,In_327,In_992);
xor U673 (N_673,In_488,In_371);
and U674 (N_674,In_763,In_13);
xor U675 (N_675,In_799,In_745);
nand U676 (N_676,In_498,In_285);
xor U677 (N_677,In_36,In_681);
nand U678 (N_678,In_440,In_536);
xor U679 (N_679,In_621,In_795);
nor U680 (N_680,In_384,In_821);
and U681 (N_681,In_675,In_519);
or U682 (N_682,In_35,In_361);
xnor U683 (N_683,In_776,In_625);
and U684 (N_684,In_898,In_124);
or U685 (N_685,In_301,In_455);
nand U686 (N_686,In_849,In_678);
nor U687 (N_687,In_875,In_741);
or U688 (N_688,In_653,In_397);
nor U689 (N_689,In_783,In_542);
xor U690 (N_690,In_728,In_411);
nand U691 (N_691,In_661,In_802);
or U692 (N_692,In_444,In_809);
and U693 (N_693,In_397,In_275);
xnor U694 (N_694,In_544,In_841);
nand U695 (N_695,In_504,In_587);
xor U696 (N_696,In_305,In_659);
xor U697 (N_697,In_80,In_355);
or U698 (N_698,In_984,In_788);
or U699 (N_699,In_584,In_141);
and U700 (N_700,In_999,In_35);
or U701 (N_701,In_298,In_945);
and U702 (N_702,In_798,In_458);
xor U703 (N_703,In_629,In_278);
xor U704 (N_704,In_429,In_571);
nand U705 (N_705,In_456,In_240);
xor U706 (N_706,In_664,In_916);
and U707 (N_707,In_912,In_358);
xnor U708 (N_708,In_529,In_917);
or U709 (N_709,In_24,In_355);
nor U710 (N_710,In_709,In_153);
xnor U711 (N_711,In_421,In_980);
nor U712 (N_712,In_214,In_555);
nor U713 (N_713,In_391,In_167);
xnor U714 (N_714,In_509,In_81);
nor U715 (N_715,In_738,In_209);
nor U716 (N_716,In_602,In_833);
and U717 (N_717,In_750,In_689);
nand U718 (N_718,In_11,In_471);
and U719 (N_719,In_958,In_656);
nor U720 (N_720,In_438,In_766);
nand U721 (N_721,In_439,In_211);
xor U722 (N_722,In_466,In_395);
or U723 (N_723,In_255,In_832);
and U724 (N_724,In_499,In_111);
and U725 (N_725,In_103,In_801);
nand U726 (N_726,In_332,In_66);
nand U727 (N_727,In_261,In_930);
nor U728 (N_728,In_866,In_444);
xor U729 (N_729,In_223,In_761);
xnor U730 (N_730,In_911,In_947);
nand U731 (N_731,In_241,In_866);
nand U732 (N_732,In_360,In_914);
nand U733 (N_733,In_705,In_689);
or U734 (N_734,In_548,In_221);
nand U735 (N_735,In_119,In_124);
nor U736 (N_736,In_545,In_554);
xnor U737 (N_737,In_623,In_683);
nor U738 (N_738,In_389,In_157);
nand U739 (N_739,In_100,In_639);
xnor U740 (N_740,In_311,In_749);
or U741 (N_741,In_622,In_68);
or U742 (N_742,In_683,In_300);
xor U743 (N_743,In_168,In_667);
xor U744 (N_744,In_151,In_757);
xor U745 (N_745,In_68,In_231);
and U746 (N_746,In_653,In_9);
nor U747 (N_747,In_589,In_931);
and U748 (N_748,In_237,In_343);
nor U749 (N_749,In_71,In_645);
xor U750 (N_750,In_456,In_121);
and U751 (N_751,In_169,In_855);
and U752 (N_752,In_998,In_888);
nand U753 (N_753,In_892,In_775);
or U754 (N_754,In_540,In_715);
or U755 (N_755,In_727,In_348);
nand U756 (N_756,In_402,In_696);
and U757 (N_757,In_199,In_735);
nand U758 (N_758,In_335,In_597);
nand U759 (N_759,In_483,In_97);
and U760 (N_760,In_384,In_408);
or U761 (N_761,In_598,In_674);
xnor U762 (N_762,In_768,In_893);
and U763 (N_763,In_969,In_974);
xnor U764 (N_764,In_486,In_532);
xnor U765 (N_765,In_696,In_412);
or U766 (N_766,In_805,In_752);
or U767 (N_767,In_236,In_591);
or U768 (N_768,In_495,In_350);
nand U769 (N_769,In_998,In_769);
and U770 (N_770,In_566,In_792);
nor U771 (N_771,In_325,In_395);
nor U772 (N_772,In_423,In_837);
and U773 (N_773,In_586,In_824);
nand U774 (N_774,In_522,In_81);
nor U775 (N_775,In_464,In_735);
or U776 (N_776,In_387,In_343);
or U777 (N_777,In_547,In_773);
nand U778 (N_778,In_248,In_198);
nor U779 (N_779,In_562,In_339);
nor U780 (N_780,In_809,In_327);
nand U781 (N_781,In_233,In_319);
xnor U782 (N_782,In_292,In_197);
and U783 (N_783,In_26,In_294);
xnor U784 (N_784,In_328,In_609);
and U785 (N_785,In_612,In_264);
and U786 (N_786,In_378,In_266);
and U787 (N_787,In_962,In_970);
nand U788 (N_788,In_527,In_558);
nand U789 (N_789,In_75,In_555);
nand U790 (N_790,In_165,In_135);
nand U791 (N_791,In_287,In_27);
or U792 (N_792,In_835,In_572);
xor U793 (N_793,In_672,In_779);
xor U794 (N_794,In_5,In_664);
and U795 (N_795,In_91,In_10);
or U796 (N_796,In_249,In_296);
nand U797 (N_797,In_149,In_540);
nand U798 (N_798,In_111,In_302);
and U799 (N_799,In_225,In_668);
nand U800 (N_800,In_438,In_88);
or U801 (N_801,In_502,In_870);
nand U802 (N_802,In_355,In_993);
nor U803 (N_803,In_166,In_588);
or U804 (N_804,In_355,In_9);
nand U805 (N_805,In_687,In_508);
nor U806 (N_806,In_581,In_158);
nor U807 (N_807,In_840,In_668);
and U808 (N_808,In_632,In_384);
nand U809 (N_809,In_77,In_645);
nor U810 (N_810,In_293,In_491);
nand U811 (N_811,In_349,In_459);
nor U812 (N_812,In_375,In_147);
nand U813 (N_813,In_37,In_513);
nand U814 (N_814,In_338,In_787);
nand U815 (N_815,In_579,In_800);
nor U816 (N_816,In_147,In_97);
and U817 (N_817,In_426,In_732);
xnor U818 (N_818,In_239,In_252);
and U819 (N_819,In_979,In_505);
xnor U820 (N_820,In_769,In_145);
xnor U821 (N_821,In_875,In_200);
nor U822 (N_822,In_5,In_950);
nand U823 (N_823,In_477,In_709);
or U824 (N_824,In_690,In_41);
nand U825 (N_825,In_932,In_631);
xnor U826 (N_826,In_408,In_639);
nor U827 (N_827,In_297,In_781);
and U828 (N_828,In_974,In_204);
nand U829 (N_829,In_452,In_29);
and U830 (N_830,In_74,In_272);
nand U831 (N_831,In_731,In_510);
and U832 (N_832,In_149,In_795);
xor U833 (N_833,In_731,In_566);
or U834 (N_834,In_518,In_125);
and U835 (N_835,In_943,In_279);
nor U836 (N_836,In_22,In_292);
nand U837 (N_837,In_358,In_804);
and U838 (N_838,In_69,In_300);
nor U839 (N_839,In_813,In_906);
or U840 (N_840,In_394,In_49);
or U841 (N_841,In_38,In_141);
or U842 (N_842,In_35,In_51);
nor U843 (N_843,In_821,In_337);
nor U844 (N_844,In_353,In_340);
xnor U845 (N_845,In_511,In_28);
or U846 (N_846,In_474,In_328);
xor U847 (N_847,In_781,In_498);
or U848 (N_848,In_606,In_151);
or U849 (N_849,In_702,In_695);
and U850 (N_850,In_410,In_285);
or U851 (N_851,In_803,In_42);
xor U852 (N_852,In_894,In_29);
xnor U853 (N_853,In_406,In_577);
xor U854 (N_854,In_995,In_897);
nor U855 (N_855,In_775,In_443);
nand U856 (N_856,In_67,In_186);
nand U857 (N_857,In_602,In_470);
or U858 (N_858,In_850,In_735);
xor U859 (N_859,In_529,In_777);
nor U860 (N_860,In_50,In_301);
or U861 (N_861,In_824,In_626);
nor U862 (N_862,In_993,In_525);
and U863 (N_863,In_509,In_586);
or U864 (N_864,In_390,In_831);
or U865 (N_865,In_432,In_521);
xnor U866 (N_866,In_363,In_101);
and U867 (N_867,In_345,In_980);
and U868 (N_868,In_592,In_309);
nor U869 (N_869,In_691,In_373);
and U870 (N_870,In_392,In_518);
xnor U871 (N_871,In_423,In_12);
xor U872 (N_872,In_636,In_98);
nor U873 (N_873,In_204,In_113);
nand U874 (N_874,In_54,In_845);
and U875 (N_875,In_57,In_556);
nor U876 (N_876,In_941,In_200);
xnor U877 (N_877,In_430,In_75);
and U878 (N_878,In_803,In_408);
xnor U879 (N_879,In_962,In_215);
xnor U880 (N_880,In_918,In_185);
nand U881 (N_881,In_686,In_620);
nand U882 (N_882,In_286,In_356);
and U883 (N_883,In_895,In_403);
and U884 (N_884,In_80,In_451);
nor U885 (N_885,In_883,In_881);
and U886 (N_886,In_540,In_589);
and U887 (N_887,In_364,In_331);
nand U888 (N_888,In_783,In_255);
or U889 (N_889,In_748,In_340);
nand U890 (N_890,In_696,In_673);
and U891 (N_891,In_622,In_255);
or U892 (N_892,In_106,In_790);
nand U893 (N_893,In_209,In_693);
or U894 (N_894,In_94,In_177);
or U895 (N_895,In_323,In_828);
and U896 (N_896,In_945,In_677);
xnor U897 (N_897,In_861,In_328);
or U898 (N_898,In_153,In_691);
or U899 (N_899,In_243,In_634);
nor U900 (N_900,In_89,In_751);
or U901 (N_901,In_241,In_921);
nand U902 (N_902,In_368,In_415);
xnor U903 (N_903,In_625,In_833);
and U904 (N_904,In_37,In_865);
or U905 (N_905,In_427,In_822);
nor U906 (N_906,In_401,In_650);
nor U907 (N_907,In_628,In_609);
nor U908 (N_908,In_976,In_27);
nor U909 (N_909,In_91,In_774);
nand U910 (N_910,In_685,In_35);
and U911 (N_911,In_846,In_969);
or U912 (N_912,In_800,In_749);
nor U913 (N_913,In_7,In_231);
xor U914 (N_914,In_239,In_23);
and U915 (N_915,In_75,In_783);
or U916 (N_916,In_99,In_799);
nand U917 (N_917,In_650,In_101);
or U918 (N_918,In_601,In_264);
xor U919 (N_919,In_841,In_779);
and U920 (N_920,In_573,In_633);
or U921 (N_921,In_786,In_526);
or U922 (N_922,In_352,In_325);
nand U923 (N_923,In_202,In_157);
or U924 (N_924,In_178,In_256);
xor U925 (N_925,In_891,In_235);
nor U926 (N_926,In_509,In_459);
xnor U927 (N_927,In_666,In_36);
or U928 (N_928,In_3,In_193);
nand U929 (N_929,In_2,In_595);
or U930 (N_930,In_444,In_134);
nand U931 (N_931,In_444,In_774);
xnor U932 (N_932,In_80,In_696);
nand U933 (N_933,In_115,In_362);
or U934 (N_934,In_501,In_976);
and U935 (N_935,In_936,In_105);
or U936 (N_936,In_96,In_664);
nand U937 (N_937,In_801,In_244);
nor U938 (N_938,In_613,In_806);
or U939 (N_939,In_543,In_201);
and U940 (N_940,In_923,In_102);
xnor U941 (N_941,In_296,In_843);
nor U942 (N_942,In_702,In_496);
or U943 (N_943,In_305,In_508);
nand U944 (N_944,In_418,In_55);
and U945 (N_945,In_903,In_829);
and U946 (N_946,In_746,In_240);
and U947 (N_947,In_300,In_32);
xor U948 (N_948,In_581,In_995);
nor U949 (N_949,In_393,In_584);
nand U950 (N_950,In_132,In_895);
and U951 (N_951,In_277,In_165);
nand U952 (N_952,In_554,In_880);
or U953 (N_953,In_532,In_872);
xnor U954 (N_954,In_166,In_389);
nor U955 (N_955,In_377,In_815);
xor U956 (N_956,In_439,In_328);
or U957 (N_957,In_476,In_463);
nor U958 (N_958,In_909,In_242);
and U959 (N_959,In_949,In_919);
nand U960 (N_960,In_937,In_313);
nand U961 (N_961,In_526,In_131);
and U962 (N_962,In_729,In_143);
xor U963 (N_963,In_359,In_41);
nor U964 (N_964,In_30,In_668);
nor U965 (N_965,In_472,In_787);
nand U966 (N_966,In_324,In_644);
or U967 (N_967,In_124,In_749);
and U968 (N_968,In_801,In_996);
nand U969 (N_969,In_517,In_707);
xnor U970 (N_970,In_707,In_74);
nand U971 (N_971,In_512,In_548);
nor U972 (N_972,In_782,In_625);
and U973 (N_973,In_317,In_262);
nand U974 (N_974,In_232,In_582);
xnor U975 (N_975,In_82,In_160);
nand U976 (N_976,In_761,In_460);
and U977 (N_977,In_372,In_976);
and U978 (N_978,In_395,In_701);
and U979 (N_979,In_388,In_29);
xor U980 (N_980,In_936,In_634);
xnor U981 (N_981,In_417,In_403);
nand U982 (N_982,In_856,In_466);
or U983 (N_983,In_781,In_997);
xor U984 (N_984,In_164,In_522);
and U985 (N_985,In_578,In_840);
or U986 (N_986,In_466,In_102);
and U987 (N_987,In_307,In_475);
nand U988 (N_988,In_673,In_726);
nor U989 (N_989,In_352,In_868);
nand U990 (N_990,In_672,In_266);
nand U991 (N_991,In_97,In_110);
xnor U992 (N_992,In_971,In_731);
nor U993 (N_993,In_51,In_982);
nand U994 (N_994,In_695,In_95);
nor U995 (N_995,In_408,In_772);
nand U996 (N_996,In_360,In_556);
or U997 (N_997,In_395,In_532);
nand U998 (N_998,In_405,In_867);
or U999 (N_999,In_317,In_287);
or U1000 (N_1000,In_658,In_379);
and U1001 (N_1001,In_798,In_856);
or U1002 (N_1002,In_87,In_552);
or U1003 (N_1003,In_459,In_492);
nand U1004 (N_1004,In_885,In_111);
xor U1005 (N_1005,In_767,In_319);
xnor U1006 (N_1006,In_275,In_708);
xor U1007 (N_1007,In_831,In_47);
or U1008 (N_1008,In_848,In_315);
xor U1009 (N_1009,In_566,In_733);
and U1010 (N_1010,In_522,In_985);
xor U1011 (N_1011,In_788,In_215);
xnor U1012 (N_1012,In_217,In_267);
xor U1013 (N_1013,In_135,In_964);
or U1014 (N_1014,In_837,In_148);
or U1015 (N_1015,In_942,In_895);
xor U1016 (N_1016,In_263,In_589);
nor U1017 (N_1017,In_170,In_145);
nand U1018 (N_1018,In_863,In_875);
or U1019 (N_1019,In_849,In_765);
and U1020 (N_1020,In_782,In_908);
and U1021 (N_1021,In_662,In_312);
and U1022 (N_1022,In_953,In_38);
or U1023 (N_1023,In_501,In_948);
xor U1024 (N_1024,In_766,In_69);
nor U1025 (N_1025,In_32,In_218);
nand U1026 (N_1026,In_536,In_866);
and U1027 (N_1027,In_416,In_625);
nor U1028 (N_1028,In_275,In_214);
nor U1029 (N_1029,In_84,In_793);
or U1030 (N_1030,In_283,In_478);
nor U1031 (N_1031,In_317,In_109);
and U1032 (N_1032,In_198,In_440);
xor U1033 (N_1033,In_887,In_788);
xnor U1034 (N_1034,In_758,In_156);
or U1035 (N_1035,In_488,In_498);
xor U1036 (N_1036,In_533,In_942);
nand U1037 (N_1037,In_470,In_606);
and U1038 (N_1038,In_852,In_421);
nor U1039 (N_1039,In_7,In_949);
xor U1040 (N_1040,In_72,In_425);
and U1041 (N_1041,In_251,In_882);
nor U1042 (N_1042,In_241,In_930);
or U1043 (N_1043,In_559,In_795);
and U1044 (N_1044,In_79,In_885);
xnor U1045 (N_1045,In_877,In_134);
nor U1046 (N_1046,In_154,In_202);
nor U1047 (N_1047,In_668,In_734);
nor U1048 (N_1048,In_665,In_865);
nand U1049 (N_1049,In_881,In_155);
and U1050 (N_1050,In_24,In_897);
nand U1051 (N_1051,In_59,In_471);
or U1052 (N_1052,In_364,In_471);
and U1053 (N_1053,In_172,In_648);
nor U1054 (N_1054,In_433,In_733);
xor U1055 (N_1055,In_526,In_932);
or U1056 (N_1056,In_503,In_590);
xnor U1057 (N_1057,In_703,In_299);
nor U1058 (N_1058,In_325,In_453);
or U1059 (N_1059,In_553,In_349);
and U1060 (N_1060,In_658,In_485);
or U1061 (N_1061,In_999,In_901);
or U1062 (N_1062,In_76,In_144);
nand U1063 (N_1063,In_634,In_533);
xor U1064 (N_1064,In_884,In_991);
xnor U1065 (N_1065,In_212,In_829);
or U1066 (N_1066,In_429,In_911);
xor U1067 (N_1067,In_406,In_931);
nand U1068 (N_1068,In_599,In_263);
or U1069 (N_1069,In_224,In_570);
or U1070 (N_1070,In_660,In_152);
xnor U1071 (N_1071,In_789,In_23);
nor U1072 (N_1072,In_475,In_419);
nand U1073 (N_1073,In_477,In_921);
and U1074 (N_1074,In_957,In_284);
nand U1075 (N_1075,In_912,In_511);
or U1076 (N_1076,In_54,In_158);
and U1077 (N_1077,In_402,In_239);
xnor U1078 (N_1078,In_133,In_202);
nand U1079 (N_1079,In_398,In_371);
or U1080 (N_1080,In_271,In_226);
xnor U1081 (N_1081,In_816,In_966);
nor U1082 (N_1082,In_877,In_503);
xor U1083 (N_1083,In_643,In_286);
or U1084 (N_1084,In_181,In_588);
or U1085 (N_1085,In_802,In_606);
nor U1086 (N_1086,In_660,In_919);
and U1087 (N_1087,In_569,In_643);
or U1088 (N_1088,In_380,In_554);
xor U1089 (N_1089,In_272,In_748);
nand U1090 (N_1090,In_83,In_182);
nor U1091 (N_1091,In_689,In_568);
or U1092 (N_1092,In_203,In_677);
nor U1093 (N_1093,In_466,In_145);
nand U1094 (N_1094,In_324,In_667);
xnor U1095 (N_1095,In_321,In_687);
xnor U1096 (N_1096,In_980,In_201);
or U1097 (N_1097,In_733,In_316);
nand U1098 (N_1098,In_453,In_163);
nor U1099 (N_1099,In_143,In_896);
xnor U1100 (N_1100,In_223,In_479);
and U1101 (N_1101,In_194,In_949);
and U1102 (N_1102,In_856,In_295);
and U1103 (N_1103,In_602,In_446);
nor U1104 (N_1104,In_784,In_170);
nand U1105 (N_1105,In_166,In_231);
and U1106 (N_1106,In_386,In_222);
nor U1107 (N_1107,In_891,In_53);
and U1108 (N_1108,In_636,In_579);
nand U1109 (N_1109,In_193,In_178);
nor U1110 (N_1110,In_795,In_467);
and U1111 (N_1111,In_459,In_632);
or U1112 (N_1112,In_286,In_352);
nand U1113 (N_1113,In_52,In_706);
nand U1114 (N_1114,In_647,In_601);
nand U1115 (N_1115,In_842,In_352);
and U1116 (N_1116,In_412,In_909);
nand U1117 (N_1117,In_772,In_194);
nor U1118 (N_1118,In_904,In_993);
and U1119 (N_1119,In_873,In_716);
nand U1120 (N_1120,In_156,In_93);
nor U1121 (N_1121,In_21,In_510);
or U1122 (N_1122,In_775,In_616);
and U1123 (N_1123,In_259,In_149);
or U1124 (N_1124,In_514,In_885);
or U1125 (N_1125,In_464,In_458);
xor U1126 (N_1126,In_557,In_30);
and U1127 (N_1127,In_862,In_41);
nand U1128 (N_1128,In_635,In_122);
and U1129 (N_1129,In_500,In_149);
and U1130 (N_1130,In_539,In_625);
nand U1131 (N_1131,In_485,In_513);
or U1132 (N_1132,In_418,In_676);
and U1133 (N_1133,In_134,In_942);
and U1134 (N_1134,In_685,In_549);
or U1135 (N_1135,In_814,In_377);
xnor U1136 (N_1136,In_826,In_334);
nor U1137 (N_1137,In_427,In_249);
or U1138 (N_1138,In_482,In_464);
and U1139 (N_1139,In_373,In_698);
nor U1140 (N_1140,In_289,In_743);
xor U1141 (N_1141,In_479,In_960);
and U1142 (N_1142,In_461,In_103);
or U1143 (N_1143,In_729,In_520);
nand U1144 (N_1144,In_594,In_654);
or U1145 (N_1145,In_982,In_508);
and U1146 (N_1146,In_934,In_261);
and U1147 (N_1147,In_592,In_46);
nand U1148 (N_1148,In_710,In_462);
and U1149 (N_1149,In_277,In_767);
nand U1150 (N_1150,In_806,In_848);
or U1151 (N_1151,In_366,In_459);
nand U1152 (N_1152,In_207,In_304);
nand U1153 (N_1153,In_746,In_1);
and U1154 (N_1154,In_323,In_357);
or U1155 (N_1155,In_495,In_625);
and U1156 (N_1156,In_74,In_522);
or U1157 (N_1157,In_20,In_864);
nand U1158 (N_1158,In_315,In_550);
and U1159 (N_1159,In_647,In_717);
or U1160 (N_1160,In_696,In_454);
nor U1161 (N_1161,In_557,In_524);
xnor U1162 (N_1162,In_691,In_54);
or U1163 (N_1163,In_423,In_584);
and U1164 (N_1164,In_207,In_109);
nand U1165 (N_1165,In_823,In_560);
nor U1166 (N_1166,In_488,In_230);
xnor U1167 (N_1167,In_812,In_119);
nor U1168 (N_1168,In_505,In_781);
xnor U1169 (N_1169,In_117,In_660);
and U1170 (N_1170,In_791,In_696);
xnor U1171 (N_1171,In_913,In_37);
nand U1172 (N_1172,In_587,In_938);
or U1173 (N_1173,In_626,In_285);
nand U1174 (N_1174,In_85,In_779);
nand U1175 (N_1175,In_549,In_277);
nand U1176 (N_1176,In_911,In_962);
nor U1177 (N_1177,In_827,In_92);
and U1178 (N_1178,In_47,In_326);
xor U1179 (N_1179,In_366,In_506);
nor U1180 (N_1180,In_737,In_334);
and U1181 (N_1181,In_784,In_679);
nor U1182 (N_1182,In_444,In_591);
xor U1183 (N_1183,In_622,In_799);
nor U1184 (N_1184,In_452,In_69);
nor U1185 (N_1185,In_847,In_88);
and U1186 (N_1186,In_803,In_402);
nor U1187 (N_1187,In_695,In_643);
and U1188 (N_1188,In_299,In_626);
xor U1189 (N_1189,In_918,In_458);
nor U1190 (N_1190,In_356,In_599);
xor U1191 (N_1191,In_250,In_137);
nand U1192 (N_1192,In_716,In_200);
xor U1193 (N_1193,In_693,In_779);
nor U1194 (N_1194,In_673,In_284);
xnor U1195 (N_1195,In_654,In_748);
or U1196 (N_1196,In_142,In_283);
or U1197 (N_1197,In_958,In_111);
xnor U1198 (N_1198,In_75,In_694);
nor U1199 (N_1199,In_730,In_611);
and U1200 (N_1200,In_14,In_184);
nor U1201 (N_1201,In_170,In_26);
xnor U1202 (N_1202,In_911,In_251);
nor U1203 (N_1203,In_521,In_227);
nor U1204 (N_1204,In_302,In_400);
or U1205 (N_1205,In_83,In_809);
nor U1206 (N_1206,In_422,In_442);
nand U1207 (N_1207,In_894,In_824);
nor U1208 (N_1208,In_746,In_772);
and U1209 (N_1209,In_980,In_928);
xnor U1210 (N_1210,In_136,In_535);
xor U1211 (N_1211,In_510,In_824);
nand U1212 (N_1212,In_198,In_725);
or U1213 (N_1213,In_523,In_958);
xnor U1214 (N_1214,In_109,In_742);
or U1215 (N_1215,In_420,In_247);
xor U1216 (N_1216,In_5,In_73);
nand U1217 (N_1217,In_706,In_171);
nand U1218 (N_1218,In_827,In_921);
nor U1219 (N_1219,In_110,In_836);
nor U1220 (N_1220,In_981,In_684);
xnor U1221 (N_1221,In_95,In_13);
or U1222 (N_1222,In_699,In_784);
nor U1223 (N_1223,In_166,In_875);
or U1224 (N_1224,In_521,In_885);
or U1225 (N_1225,In_559,In_873);
or U1226 (N_1226,In_922,In_895);
xor U1227 (N_1227,In_603,In_187);
nand U1228 (N_1228,In_477,In_520);
or U1229 (N_1229,In_653,In_616);
xnor U1230 (N_1230,In_770,In_295);
and U1231 (N_1231,In_324,In_660);
xnor U1232 (N_1232,In_233,In_105);
or U1233 (N_1233,In_610,In_433);
and U1234 (N_1234,In_225,In_54);
nor U1235 (N_1235,In_201,In_688);
nand U1236 (N_1236,In_523,In_321);
nand U1237 (N_1237,In_389,In_857);
and U1238 (N_1238,In_266,In_498);
and U1239 (N_1239,In_461,In_398);
or U1240 (N_1240,In_168,In_699);
xor U1241 (N_1241,In_516,In_281);
and U1242 (N_1242,In_963,In_410);
nor U1243 (N_1243,In_710,In_298);
nor U1244 (N_1244,In_918,In_349);
or U1245 (N_1245,In_404,In_268);
nand U1246 (N_1246,In_672,In_528);
nand U1247 (N_1247,In_81,In_278);
nand U1248 (N_1248,In_270,In_72);
nand U1249 (N_1249,In_34,In_341);
nor U1250 (N_1250,In_683,In_691);
and U1251 (N_1251,In_838,In_65);
xnor U1252 (N_1252,In_575,In_806);
or U1253 (N_1253,In_432,In_205);
and U1254 (N_1254,In_990,In_469);
nand U1255 (N_1255,In_41,In_674);
nor U1256 (N_1256,In_692,In_913);
xnor U1257 (N_1257,In_223,In_116);
or U1258 (N_1258,In_393,In_249);
nor U1259 (N_1259,In_758,In_91);
xnor U1260 (N_1260,In_211,In_801);
nand U1261 (N_1261,In_357,In_928);
nand U1262 (N_1262,In_200,In_937);
xnor U1263 (N_1263,In_994,In_114);
or U1264 (N_1264,In_819,In_898);
nor U1265 (N_1265,In_885,In_962);
xnor U1266 (N_1266,In_882,In_419);
and U1267 (N_1267,In_903,In_220);
xnor U1268 (N_1268,In_686,In_378);
nand U1269 (N_1269,In_672,In_353);
and U1270 (N_1270,In_50,In_974);
and U1271 (N_1271,In_544,In_22);
or U1272 (N_1272,In_395,In_991);
or U1273 (N_1273,In_746,In_20);
nand U1274 (N_1274,In_191,In_32);
nor U1275 (N_1275,In_544,In_55);
xnor U1276 (N_1276,In_868,In_475);
and U1277 (N_1277,In_208,In_346);
or U1278 (N_1278,In_146,In_901);
and U1279 (N_1279,In_478,In_764);
and U1280 (N_1280,In_452,In_166);
and U1281 (N_1281,In_27,In_898);
xnor U1282 (N_1282,In_941,In_353);
xnor U1283 (N_1283,In_268,In_353);
xor U1284 (N_1284,In_916,In_393);
or U1285 (N_1285,In_491,In_875);
nor U1286 (N_1286,In_794,In_342);
xnor U1287 (N_1287,In_808,In_508);
xnor U1288 (N_1288,In_983,In_672);
or U1289 (N_1289,In_741,In_832);
xnor U1290 (N_1290,In_826,In_112);
or U1291 (N_1291,In_578,In_497);
xnor U1292 (N_1292,In_155,In_713);
nor U1293 (N_1293,In_44,In_744);
nor U1294 (N_1294,In_367,In_100);
and U1295 (N_1295,In_768,In_706);
nand U1296 (N_1296,In_852,In_837);
xnor U1297 (N_1297,In_944,In_881);
nor U1298 (N_1298,In_356,In_13);
or U1299 (N_1299,In_278,In_714);
nand U1300 (N_1300,In_482,In_169);
and U1301 (N_1301,In_670,In_398);
and U1302 (N_1302,In_445,In_656);
or U1303 (N_1303,In_491,In_30);
and U1304 (N_1304,In_178,In_325);
and U1305 (N_1305,In_206,In_482);
nor U1306 (N_1306,In_387,In_514);
nand U1307 (N_1307,In_360,In_257);
xor U1308 (N_1308,In_841,In_906);
and U1309 (N_1309,In_261,In_225);
or U1310 (N_1310,In_874,In_612);
or U1311 (N_1311,In_701,In_9);
xor U1312 (N_1312,In_104,In_496);
nor U1313 (N_1313,In_340,In_311);
nor U1314 (N_1314,In_291,In_608);
or U1315 (N_1315,In_150,In_519);
or U1316 (N_1316,In_658,In_925);
or U1317 (N_1317,In_592,In_15);
and U1318 (N_1318,In_331,In_827);
nand U1319 (N_1319,In_46,In_641);
or U1320 (N_1320,In_89,In_948);
and U1321 (N_1321,In_185,In_852);
and U1322 (N_1322,In_431,In_331);
nand U1323 (N_1323,In_385,In_823);
and U1324 (N_1324,In_924,In_404);
and U1325 (N_1325,In_676,In_402);
and U1326 (N_1326,In_228,In_682);
nand U1327 (N_1327,In_639,In_690);
or U1328 (N_1328,In_466,In_213);
and U1329 (N_1329,In_503,In_146);
xnor U1330 (N_1330,In_289,In_659);
nor U1331 (N_1331,In_563,In_694);
or U1332 (N_1332,In_319,In_200);
xnor U1333 (N_1333,In_231,In_642);
nand U1334 (N_1334,In_651,In_727);
or U1335 (N_1335,In_866,In_811);
or U1336 (N_1336,In_979,In_485);
xnor U1337 (N_1337,In_315,In_566);
and U1338 (N_1338,In_280,In_38);
xnor U1339 (N_1339,In_447,In_817);
nor U1340 (N_1340,In_818,In_829);
and U1341 (N_1341,In_993,In_248);
nor U1342 (N_1342,In_938,In_293);
nand U1343 (N_1343,In_301,In_509);
nand U1344 (N_1344,In_71,In_391);
and U1345 (N_1345,In_650,In_115);
xor U1346 (N_1346,In_448,In_138);
or U1347 (N_1347,In_607,In_146);
or U1348 (N_1348,In_939,In_267);
and U1349 (N_1349,In_836,In_653);
nor U1350 (N_1350,In_734,In_363);
xnor U1351 (N_1351,In_225,In_337);
and U1352 (N_1352,In_862,In_141);
nor U1353 (N_1353,In_882,In_764);
xor U1354 (N_1354,In_303,In_672);
nor U1355 (N_1355,In_474,In_880);
nand U1356 (N_1356,In_291,In_427);
nor U1357 (N_1357,In_718,In_267);
xor U1358 (N_1358,In_6,In_927);
and U1359 (N_1359,In_852,In_872);
or U1360 (N_1360,In_788,In_433);
or U1361 (N_1361,In_579,In_949);
nand U1362 (N_1362,In_977,In_559);
or U1363 (N_1363,In_278,In_671);
or U1364 (N_1364,In_624,In_297);
xnor U1365 (N_1365,In_350,In_818);
nor U1366 (N_1366,In_108,In_796);
or U1367 (N_1367,In_330,In_838);
nor U1368 (N_1368,In_50,In_15);
xnor U1369 (N_1369,In_716,In_986);
xor U1370 (N_1370,In_71,In_878);
and U1371 (N_1371,In_529,In_531);
and U1372 (N_1372,In_207,In_844);
nor U1373 (N_1373,In_777,In_542);
or U1374 (N_1374,In_698,In_632);
nor U1375 (N_1375,In_528,In_148);
or U1376 (N_1376,In_991,In_101);
nand U1377 (N_1377,In_126,In_203);
nand U1378 (N_1378,In_260,In_357);
or U1379 (N_1379,In_524,In_482);
xnor U1380 (N_1380,In_689,In_259);
and U1381 (N_1381,In_218,In_493);
nand U1382 (N_1382,In_543,In_453);
and U1383 (N_1383,In_585,In_113);
nor U1384 (N_1384,In_378,In_459);
nor U1385 (N_1385,In_716,In_468);
xor U1386 (N_1386,In_20,In_508);
or U1387 (N_1387,In_397,In_261);
xor U1388 (N_1388,In_121,In_972);
nor U1389 (N_1389,In_229,In_868);
or U1390 (N_1390,In_439,In_896);
and U1391 (N_1391,In_889,In_180);
or U1392 (N_1392,In_67,In_90);
nor U1393 (N_1393,In_476,In_674);
and U1394 (N_1394,In_54,In_494);
nand U1395 (N_1395,In_590,In_399);
and U1396 (N_1396,In_28,In_947);
xnor U1397 (N_1397,In_445,In_464);
and U1398 (N_1398,In_950,In_850);
or U1399 (N_1399,In_640,In_727);
nand U1400 (N_1400,In_190,In_510);
and U1401 (N_1401,In_352,In_510);
or U1402 (N_1402,In_136,In_7);
or U1403 (N_1403,In_464,In_994);
and U1404 (N_1404,In_822,In_592);
xor U1405 (N_1405,In_298,In_350);
nand U1406 (N_1406,In_595,In_944);
xnor U1407 (N_1407,In_388,In_117);
and U1408 (N_1408,In_295,In_535);
nor U1409 (N_1409,In_846,In_168);
xor U1410 (N_1410,In_859,In_5);
and U1411 (N_1411,In_235,In_690);
and U1412 (N_1412,In_888,In_169);
nor U1413 (N_1413,In_26,In_184);
nand U1414 (N_1414,In_582,In_320);
nand U1415 (N_1415,In_614,In_543);
or U1416 (N_1416,In_88,In_898);
xor U1417 (N_1417,In_830,In_211);
or U1418 (N_1418,In_162,In_852);
xor U1419 (N_1419,In_150,In_657);
nand U1420 (N_1420,In_737,In_816);
nand U1421 (N_1421,In_417,In_662);
nand U1422 (N_1422,In_885,In_797);
nor U1423 (N_1423,In_194,In_108);
or U1424 (N_1424,In_753,In_588);
and U1425 (N_1425,In_486,In_832);
and U1426 (N_1426,In_152,In_330);
and U1427 (N_1427,In_716,In_458);
and U1428 (N_1428,In_180,In_685);
or U1429 (N_1429,In_990,In_462);
and U1430 (N_1430,In_583,In_366);
xnor U1431 (N_1431,In_247,In_383);
xor U1432 (N_1432,In_160,In_312);
and U1433 (N_1433,In_832,In_745);
nand U1434 (N_1434,In_576,In_688);
and U1435 (N_1435,In_283,In_379);
or U1436 (N_1436,In_371,In_979);
xnor U1437 (N_1437,In_150,In_958);
or U1438 (N_1438,In_607,In_737);
xor U1439 (N_1439,In_268,In_620);
xor U1440 (N_1440,In_589,In_184);
nand U1441 (N_1441,In_426,In_711);
nor U1442 (N_1442,In_227,In_186);
or U1443 (N_1443,In_540,In_672);
nor U1444 (N_1444,In_573,In_27);
and U1445 (N_1445,In_103,In_987);
xnor U1446 (N_1446,In_259,In_887);
xnor U1447 (N_1447,In_222,In_287);
and U1448 (N_1448,In_80,In_457);
nor U1449 (N_1449,In_663,In_169);
nand U1450 (N_1450,In_773,In_273);
nand U1451 (N_1451,In_963,In_623);
xor U1452 (N_1452,In_79,In_354);
xnor U1453 (N_1453,In_121,In_275);
or U1454 (N_1454,In_871,In_989);
nor U1455 (N_1455,In_362,In_556);
xnor U1456 (N_1456,In_602,In_198);
and U1457 (N_1457,In_644,In_38);
or U1458 (N_1458,In_101,In_484);
and U1459 (N_1459,In_557,In_999);
nand U1460 (N_1460,In_950,In_871);
or U1461 (N_1461,In_772,In_744);
nor U1462 (N_1462,In_770,In_303);
nor U1463 (N_1463,In_303,In_188);
nor U1464 (N_1464,In_80,In_741);
nand U1465 (N_1465,In_719,In_706);
nand U1466 (N_1466,In_202,In_429);
nand U1467 (N_1467,In_460,In_326);
or U1468 (N_1468,In_457,In_218);
and U1469 (N_1469,In_523,In_527);
or U1470 (N_1470,In_914,In_479);
and U1471 (N_1471,In_133,In_109);
xor U1472 (N_1472,In_672,In_990);
or U1473 (N_1473,In_798,In_218);
xor U1474 (N_1474,In_626,In_19);
nor U1475 (N_1475,In_534,In_425);
nand U1476 (N_1476,In_632,In_181);
and U1477 (N_1477,In_336,In_456);
or U1478 (N_1478,In_874,In_456);
and U1479 (N_1479,In_736,In_498);
nor U1480 (N_1480,In_96,In_519);
nand U1481 (N_1481,In_599,In_425);
and U1482 (N_1482,In_636,In_71);
nor U1483 (N_1483,In_138,In_740);
nor U1484 (N_1484,In_913,In_582);
and U1485 (N_1485,In_8,In_598);
and U1486 (N_1486,In_712,In_530);
xor U1487 (N_1487,In_783,In_545);
xor U1488 (N_1488,In_507,In_851);
nand U1489 (N_1489,In_954,In_590);
xnor U1490 (N_1490,In_910,In_41);
or U1491 (N_1491,In_780,In_737);
xor U1492 (N_1492,In_936,In_140);
nand U1493 (N_1493,In_190,In_90);
xor U1494 (N_1494,In_151,In_70);
nor U1495 (N_1495,In_304,In_276);
and U1496 (N_1496,In_358,In_961);
xnor U1497 (N_1497,In_976,In_516);
nand U1498 (N_1498,In_357,In_615);
and U1499 (N_1499,In_12,In_976);
and U1500 (N_1500,In_219,In_251);
and U1501 (N_1501,In_958,In_547);
nor U1502 (N_1502,In_144,In_784);
or U1503 (N_1503,In_989,In_334);
xor U1504 (N_1504,In_944,In_434);
and U1505 (N_1505,In_630,In_547);
nor U1506 (N_1506,In_616,In_550);
and U1507 (N_1507,In_760,In_311);
and U1508 (N_1508,In_941,In_431);
and U1509 (N_1509,In_993,In_233);
nand U1510 (N_1510,In_548,In_137);
nor U1511 (N_1511,In_444,In_255);
nand U1512 (N_1512,In_899,In_809);
and U1513 (N_1513,In_209,In_246);
and U1514 (N_1514,In_958,In_548);
xnor U1515 (N_1515,In_348,In_900);
or U1516 (N_1516,In_252,In_974);
nor U1517 (N_1517,In_13,In_567);
xor U1518 (N_1518,In_601,In_107);
nor U1519 (N_1519,In_711,In_254);
xor U1520 (N_1520,In_135,In_607);
or U1521 (N_1521,In_250,In_697);
and U1522 (N_1522,In_878,In_450);
nor U1523 (N_1523,In_355,In_96);
xor U1524 (N_1524,In_982,In_113);
or U1525 (N_1525,In_171,In_499);
nor U1526 (N_1526,In_718,In_445);
or U1527 (N_1527,In_31,In_912);
nor U1528 (N_1528,In_481,In_851);
nor U1529 (N_1529,In_143,In_999);
or U1530 (N_1530,In_259,In_469);
or U1531 (N_1531,In_505,In_846);
and U1532 (N_1532,In_33,In_352);
or U1533 (N_1533,In_799,In_141);
and U1534 (N_1534,In_756,In_337);
nor U1535 (N_1535,In_171,In_463);
and U1536 (N_1536,In_436,In_121);
or U1537 (N_1537,In_686,In_961);
nor U1538 (N_1538,In_210,In_451);
nor U1539 (N_1539,In_370,In_307);
or U1540 (N_1540,In_540,In_643);
nand U1541 (N_1541,In_222,In_478);
or U1542 (N_1542,In_79,In_622);
and U1543 (N_1543,In_820,In_88);
nor U1544 (N_1544,In_115,In_694);
or U1545 (N_1545,In_578,In_810);
nand U1546 (N_1546,In_97,In_505);
nand U1547 (N_1547,In_895,In_546);
nand U1548 (N_1548,In_930,In_451);
nor U1549 (N_1549,In_269,In_910);
or U1550 (N_1550,In_730,In_545);
and U1551 (N_1551,In_621,In_156);
nor U1552 (N_1552,In_472,In_143);
nand U1553 (N_1553,In_694,In_914);
and U1554 (N_1554,In_452,In_614);
nand U1555 (N_1555,In_369,In_414);
nor U1556 (N_1556,In_306,In_691);
xnor U1557 (N_1557,In_611,In_943);
or U1558 (N_1558,In_452,In_798);
xor U1559 (N_1559,In_361,In_622);
and U1560 (N_1560,In_609,In_692);
or U1561 (N_1561,In_108,In_731);
xnor U1562 (N_1562,In_534,In_407);
nor U1563 (N_1563,In_317,In_384);
nor U1564 (N_1564,In_845,In_163);
nor U1565 (N_1565,In_174,In_528);
xor U1566 (N_1566,In_158,In_809);
nand U1567 (N_1567,In_504,In_69);
nor U1568 (N_1568,In_937,In_123);
nand U1569 (N_1569,In_112,In_820);
nand U1570 (N_1570,In_494,In_448);
nor U1571 (N_1571,In_142,In_34);
and U1572 (N_1572,In_633,In_581);
nor U1573 (N_1573,In_99,In_20);
and U1574 (N_1574,In_265,In_216);
nand U1575 (N_1575,In_385,In_116);
xor U1576 (N_1576,In_199,In_6);
xnor U1577 (N_1577,In_455,In_456);
xnor U1578 (N_1578,In_193,In_409);
nand U1579 (N_1579,In_834,In_233);
and U1580 (N_1580,In_798,In_49);
nand U1581 (N_1581,In_688,In_215);
nand U1582 (N_1582,In_633,In_895);
or U1583 (N_1583,In_444,In_927);
nor U1584 (N_1584,In_960,In_309);
or U1585 (N_1585,In_816,In_473);
or U1586 (N_1586,In_492,In_138);
xor U1587 (N_1587,In_642,In_655);
xor U1588 (N_1588,In_623,In_914);
or U1589 (N_1589,In_363,In_518);
or U1590 (N_1590,In_830,In_10);
and U1591 (N_1591,In_214,In_156);
and U1592 (N_1592,In_400,In_786);
nand U1593 (N_1593,In_970,In_568);
nor U1594 (N_1594,In_7,In_590);
nor U1595 (N_1595,In_893,In_162);
nand U1596 (N_1596,In_643,In_190);
and U1597 (N_1597,In_755,In_289);
or U1598 (N_1598,In_884,In_794);
and U1599 (N_1599,In_724,In_201);
nor U1600 (N_1600,In_245,In_92);
nand U1601 (N_1601,In_800,In_426);
or U1602 (N_1602,In_378,In_24);
or U1603 (N_1603,In_267,In_844);
nand U1604 (N_1604,In_254,In_151);
xor U1605 (N_1605,In_124,In_435);
and U1606 (N_1606,In_527,In_590);
nor U1607 (N_1607,In_297,In_490);
and U1608 (N_1608,In_977,In_557);
nor U1609 (N_1609,In_838,In_895);
xor U1610 (N_1610,In_41,In_550);
nand U1611 (N_1611,In_648,In_957);
xor U1612 (N_1612,In_721,In_46);
or U1613 (N_1613,In_687,In_824);
nor U1614 (N_1614,In_230,In_451);
xor U1615 (N_1615,In_196,In_772);
xor U1616 (N_1616,In_175,In_979);
or U1617 (N_1617,In_784,In_132);
nor U1618 (N_1618,In_369,In_532);
xnor U1619 (N_1619,In_331,In_893);
and U1620 (N_1620,In_682,In_112);
xor U1621 (N_1621,In_620,In_210);
nor U1622 (N_1622,In_763,In_20);
nor U1623 (N_1623,In_375,In_815);
and U1624 (N_1624,In_888,In_858);
nand U1625 (N_1625,In_273,In_94);
nand U1626 (N_1626,In_361,In_244);
xor U1627 (N_1627,In_502,In_304);
and U1628 (N_1628,In_630,In_944);
or U1629 (N_1629,In_571,In_710);
nand U1630 (N_1630,In_577,In_985);
and U1631 (N_1631,In_85,In_349);
or U1632 (N_1632,In_225,In_266);
or U1633 (N_1633,In_638,In_32);
and U1634 (N_1634,In_118,In_192);
and U1635 (N_1635,In_822,In_974);
nor U1636 (N_1636,In_607,In_167);
or U1637 (N_1637,In_841,In_659);
and U1638 (N_1638,In_185,In_3);
and U1639 (N_1639,In_873,In_674);
or U1640 (N_1640,In_716,In_98);
xnor U1641 (N_1641,In_891,In_502);
nor U1642 (N_1642,In_499,In_551);
nand U1643 (N_1643,In_408,In_132);
and U1644 (N_1644,In_734,In_469);
nand U1645 (N_1645,In_996,In_815);
nand U1646 (N_1646,In_738,In_4);
and U1647 (N_1647,In_573,In_863);
nand U1648 (N_1648,In_375,In_961);
xor U1649 (N_1649,In_543,In_864);
nor U1650 (N_1650,In_594,In_895);
nor U1651 (N_1651,In_77,In_403);
xnor U1652 (N_1652,In_452,In_912);
nor U1653 (N_1653,In_138,In_626);
or U1654 (N_1654,In_115,In_843);
or U1655 (N_1655,In_973,In_32);
and U1656 (N_1656,In_75,In_73);
or U1657 (N_1657,In_494,In_372);
or U1658 (N_1658,In_880,In_0);
or U1659 (N_1659,In_16,In_427);
or U1660 (N_1660,In_895,In_436);
nand U1661 (N_1661,In_769,In_958);
or U1662 (N_1662,In_999,In_122);
xor U1663 (N_1663,In_41,In_614);
and U1664 (N_1664,In_657,In_500);
nor U1665 (N_1665,In_136,In_689);
or U1666 (N_1666,In_913,In_585);
xor U1667 (N_1667,In_112,In_715);
and U1668 (N_1668,In_246,In_412);
xnor U1669 (N_1669,In_673,In_618);
nand U1670 (N_1670,In_335,In_356);
nor U1671 (N_1671,In_320,In_104);
or U1672 (N_1672,In_563,In_783);
nor U1673 (N_1673,In_686,In_127);
and U1674 (N_1674,In_595,In_404);
nor U1675 (N_1675,In_211,In_23);
nor U1676 (N_1676,In_15,In_362);
xnor U1677 (N_1677,In_95,In_973);
nor U1678 (N_1678,In_189,In_965);
nor U1679 (N_1679,In_34,In_778);
or U1680 (N_1680,In_233,In_269);
or U1681 (N_1681,In_134,In_772);
or U1682 (N_1682,In_396,In_733);
nor U1683 (N_1683,In_954,In_666);
nand U1684 (N_1684,In_120,In_856);
xor U1685 (N_1685,In_969,In_788);
xor U1686 (N_1686,In_535,In_294);
nand U1687 (N_1687,In_363,In_853);
nor U1688 (N_1688,In_363,In_222);
and U1689 (N_1689,In_806,In_141);
and U1690 (N_1690,In_157,In_33);
and U1691 (N_1691,In_721,In_565);
nor U1692 (N_1692,In_125,In_666);
and U1693 (N_1693,In_592,In_811);
and U1694 (N_1694,In_376,In_286);
nor U1695 (N_1695,In_9,In_563);
xnor U1696 (N_1696,In_694,In_368);
nor U1697 (N_1697,In_674,In_402);
nand U1698 (N_1698,In_309,In_107);
xor U1699 (N_1699,In_569,In_962);
and U1700 (N_1700,In_642,In_353);
and U1701 (N_1701,In_862,In_282);
and U1702 (N_1702,In_698,In_31);
and U1703 (N_1703,In_77,In_9);
or U1704 (N_1704,In_166,In_349);
nand U1705 (N_1705,In_100,In_223);
or U1706 (N_1706,In_901,In_674);
nand U1707 (N_1707,In_992,In_647);
and U1708 (N_1708,In_491,In_37);
and U1709 (N_1709,In_678,In_395);
xnor U1710 (N_1710,In_652,In_478);
xnor U1711 (N_1711,In_199,In_372);
nor U1712 (N_1712,In_148,In_184);
nor U1713 (N_1713,In_563,In_827);
nand U1714 (N_1714,In_662,In_620);
nand U1715 (N_1715,In_307,In_190);
or U1716 (N_1716,In_361,In_545);
nor U1717 (N_1717,In_867,In_395);
xor U1718 (N_1718,In_676,In_125);
nor U1719 (N_1719,In_81,In_880);
or U1720 (N_1720,In_720,In_96);
xor U1721 (N_1721,In_423,In_967);
xor U1722 (N_1722,In_125,In_770);
and U1723 (N_1723,In_126,In_787);
xnor U1724 (N_1724,In_125,In_128);
nor U1725 (N_1725,In_418,In_741);
or U1726 (N_1726,In_360,In_925);
nand U1727 (N_1727,In_529,In_146);
nor U1728 (N_1728,In_16,In_62);
xor U1729 (N_1729,In_966,In_235);
nor U1730 (N_1730,In_383,In_919);
nor U1731 (N_1731,In_676,In_635);
nor U1732 (N_1732,In_331,In_815);
xnor U1733 (N_1733,In_788,In_687);
and U1734 (N_1734,In_301,In_342);
nor U1735 (N_1735,In_843,In_696);
xor U1736 (N_1736,In_179,In_13);
or U1737 (N_1737,In_694,In_567);
or U1738 (N_1738,In_747,In_211);
nor U1739 (N_1739,In_560,In_219);
xor U1740 (N_1740,In_932,In_732);
nand U1741 (N_1741,In_934,In_597);
nand U1742 (N_1742,In_845,In_807);
or U1743 (N_1743,In_262,In_257);
nand U1744 (N_1744,In_134,In_94);
and U1745 (N_1745,In_6,In_597);
or U1746 (N_1746,In_352,In_992);
nor U1747 (N_1747,In_733,In_126);
and U1748 (N_1748,In_19,In_214);
and U1749 (N_1749,In_661,In_655);
or U1750 (N_1750,In_545,In_727);
xnor U1751 (N_1751,In_539,In_306);
nand U1752 (N_1752,In_33,In_276);
nand U1753 (N_1753,In_76,In_253);
or U1754 (N_1754,In_131,In_858);
nor U1755 (N_1755,In_546,In_556);
or U1756 (N_1756,In_728,In_4);
xor U1757 (N_1757,In_652,In_258);
nand U1758 (N_1758,In_372,In_999);
or U1759 (N_1759,In_378,In_381);
and U1760 (N_1760,In_948,In_264);
or U1761 (N_1761,In_3,In_751);
or U1762 (N_1762,In_292,In_58);
and U1763 (N_1763,In_164,In_969);
and U1764 (N_1764,In_393,In_384);
nand U1765 (N_1765,In_738,In_638);
or U1766 (N_1766,In_223,In_753);
nor U1767 (N_1767,In_893,In_507);
xor U1768 (N_1768,In_799,In_119);
or U1769 (N_1769,In_187,In_79);
nor U1770 (N_1770,In_244,In_293);
and U1771 (N_1771,In_513,In_724);
nor U1772 (N_1772,In_932,In_988);
nand U1773 (N_1773,In_297,In_445);
xor U1774 (N_1774,In_441,In_147);
nand U1775 (N_1775,In_335,In_744);
xor U1776 (N_1776,In_525,In_657);
nand U1777 (N_1777,In_834,In_282);
xnor U1778 (N_1778,In_484,In_313);
nor U1779 (N_1779,In_556,In_625);
nand U1780 (N_1780,In_418,In_811);
and U1781 (N_1781,In_574,In_633);
nand U1782 (N_1782,In_727,In_608);
nor U1783 (N_1783,In_928,In_730);
nand U1784 (N_1784,In_684,In_78);
nor U1785 (N_1785,In_508,In_464);
nand U1786 (N_1786,In_536,In_898);
and U1787 (N_1787,In_421,In_476);
and U1788 (N_1788,In_435,In_916);
and U1789 (N_1789,In_3,In_15);
nor U1790 (N_1790,In_684,In_161);
nand U1791 (N_1791,In_931,In_804);
and U1792 (N_1792,In_742,In_997);
or U1793 (N_1793,In_866,In_253);
and U1794 (N_1794,In_892,In_201);
xnor U1795 (N_1795,In_719,In_703);
xor U1796 (N_1796,In_145,In_221);
and U1797 (N_1797,In_202,In_845);
and U1798 (N_1798,In_418,In_903);
or U1799 (N_1799,In_677,In_731);
and U1800 (N_1800,In_63,In_328);
xnor U1801 (N_1801,In_326,In_880);
nor U1802 (N_1802,In_594,In_521);
nor U1803 (N_1803,In_746,In_721);
nand U1804 (N_1804,In_963,In_137);
and U1805 (N_1805,In_371,In_282);
xor U1806 (N_1806,In_433,In_521);
xnor U1807 (N_1807,In_326,In_806);
and U1808 (N_1808,In_265,In_511);
nor U1809 (N_1809,In_677,In_913);
nor U1810 (N_1810,In_407,In_275);
and U1811 (N_1811,In_614,In_189);
nor U1812 (N_1812,In_641,In_248);
nand U1813 (N_1813,In_985,In_260);
and U1814 (N_1814,In_757,In_187);
nand U1815 (N_1815,In_501,In_109);
and U1816 (N_1816,In_819,In_710);
and U1817 (N_1817,In_574,In_370);
xor U1818 (N_1818,In_236,In_60);
xor U1819 (N_1819,In_840,In_438);
or U1820 (N_1820,In_901,In_602);
or U1821 (N_1821,In_725,In_391);
xnor U1822 (N_1822,In_958,In_204);
nor U1823 (N_1823,In_242,In_908);
nor U1824 (N_1824,In_870,In_934);
nor U1825 (N_1825,In_107,In_308);
and U1826 (N_1826,In_70,In_90);
nor U1827 (N_1827,In_414,In_263);
xor U1828 (N_1828,In_729,In_232);
or U1829 (N_1829,In_205,In_219);
nor U1830 (N_1830,In_861,In_47);
xor U1831 (N_1831,In_480,In_444);
or U1832 (N_1832,In_684,In_263);
and U1833 (N_1833,In_67,In_477);
or U1834 (N_1834,In_865,In_137);
nor U1835 (N_1835,In_389,In_122);
xnor U1836 (N_1836,In_768,In_797);
or U1837 (N_1837,In_474,In_193);
and U1838 (N_1838,In_264,In_72);
and U1839 (N_1839,In_568,In_876);
and U1840 (N_1840,In_292,In_196);
nand U1841 (N_1841,In_685,In_791);
nor U1842 (N_1842,In_220,In_156);
xor U1843 (N_1843,In_155,In_277);
or U1844 (N_1844,In_320,In_607);
nand U1845 (N_1845,In_548,In_651);
or U1846 (N_1846,In_880,In_890);
xnor U1847 (N_1847,In_155,In_606);
xor U1848 (N_1848,In_820,In_842);
nor U1849 (N_1849,In_894,In_411);
nor U1850 (N_1850,In_653,In_253);
xor U1851 (N_1851,In_851,In_649);
nand U1852 (N_1852,In_82,In_829);
or U1853 (N_1853,In_689,In_582);
nor U1854 (N_1854,In_383,In_246);
nor U1855 (N_1855,In_904,In_991);
xor U1856 (N_1856,In_198,In_322);
nor U1857 (N_1857,In_897,In_540);
and U1858 (N_1858,In_616,In_325);
xnor U1859 (N_1859,In_329,In_653);
xor U1860 (N_1860,In_971,In_930);
and U1861 (N_1861,In_24,In_20);
xnor U1862 (N_1862,In_304,In_59);
xnor U1863 (N_1863,In_229,In_924);
and U1864 (N_1864,In_80,In_462);
and U1865 (N_1865,In_993,In_828);
nor U1866 (N_1866,In_854,In_461);
and U1867 (N_1867,In_684,In_705);
or U1868 (N_1868,In_391,In_472);
nand U1869 (N_1869,In_973,In_54);
xnor U1870 (N_1870,In_792,In_719);
xor U1871 (N_1871,In_19,In_469);
or U1872 (N_1872,In_826,In_340);
and U1873 (N_1873,In_352,In_140);
nor U1874 (N_1874,In_9,In_171);
and U1875 (N_1875,In_197,In_471);
xor U1876 (N_1876,In_732,In_172);
or U1877 (N_1877,In_935,In_853);
xnor U1878 (N_1878,In_299,In_908);
nor U1879 (N_1879,In_513,In_406);
or U1880 (N_1880,In_76,In_800);
xnor U1881 (N_1881,In_832,In_61);
or U1882 (N_1882,In_743,In_140);
nor U1883 (N_1883,In_656,In_438);
nand U1884 (N_1884,In_406,In_917);
xnor U1885 (N_1885,In_379,In_665);
nand U1886 (N_1886,In_918,In_266);
and U1887 (N_1887,In_939,In_749);
and U1888 (N_1888,In_213,In_67);
xor U1889 (N_1889,In_536,In_129);
and U1890 (N_1890,In_823,In_272);
nand U1891 (N_1891,In_883,In_420);
nand U1892 (N_1892,In_118,In_924);
or U1893 (N_1893,In_733,In_38);
xor U1894 (N_1894,In_527,In_745);
and U1895 (N_1895,In_447,In_775);
nor U1896 (N_1896,In_565,In_942);
and U1897 (N_1897,In_23,In_113);
nor U1898 (N_1898,In_489,In_950);
and U1899 (N_1899,In_909,In_56);
and U1900 (N_1900,In_502,In_732);
nand U1901 (N_1901,In_370,In_245);
and U1902 (N_1902,In_685,In_904);
xnor U1903 (N_1903,In_735,In_976);
and U1904 (N_1904,In_395,In_359);
nor U1905 (N_1905,In_317,In_269);
nor U1906 (N_1906,In_509,In_911);
and U1907 (N_1907,In_103,In_48);
and U1908 (N_1908,In_249,In_234);
xor U1909 (N_1909,In_923,In_718);
nor U1910 (N_1910,In_565,In_657);
nand U1911 (N_1911,In_833,In_989);
nor U1912 (N_1912,In_390,In_868);
xor U1913 (N_1913,In_542,In_208);
nor U1914 (N_1914,In_609,In_911);
and U1915 (N_1915,In_404,In_947);
nand U1916 (N_1916,In_1,In_977);
xnor U1917 (N_1917,In_633,In_53);
nor U1918 (N_1918,In_923,In_459);
and U1919 (N_1919,In_852,In_183);
and U1920 (N_1920,In_458,In_591);
nor U1921 (N_1921,In_327,In_542);
nand U1922 (N_1922,In_35,In_257);
xor U1923 (N_1923,In_336,In_861);
or U1924 (N_1924,In_140,In_463);
or U1925 (N_1925,In_32,In_189);
xnor U1926 (N_1926,In_281,In_847);
or U1927 (N_1927,In_691,In_819);
xor U1928 (N_1928,In_851,In_123);
nand U1929 (N_1929,In_192,In_85);
and U1930 (N_1930,In_657,In_253);
xnor U1931 (N_1931,In_176,In_700);
and U1932 (N_1932,In_885,In_981);
nor U1933 (N_1933,In_129,In_329);
xnor U1934 (N_1934,In_5,In_580);
nand U1935 (N_1935,In_375,In_221);
xor U1936 (N_1936,In_752,In_468);
nand U1937 (N_1937,In_654,In_133);
nand U1938 (N_1938,In_776,In_566);
nor U1939 (N_1939,In_304,In_757);
and U1940 (N_1940,In_896,In_609);
xnor U1941 (N_1941,In_150,In_966);
nand U1942 (N_1942,In_385,In_984);
nand U1943 (N_1943,In_121,In_687);
xnor U1944 (N_1944,In_466,In_170);
or U1945 (N_1945,In_798,In_951);
or U1946 (N_1946,In_65,In_293);
or U1947 (N_1947,In_564,In_939);
or U1948 (N_1948,In_421,In_714);
nor U1949 (N_1949,In_827,In_373);
nor U1950 (N_1950,In_362,In_236);
and U1951 (N_1951,In_771,In_699);
nand U1952 (N_1952,In_561,In_301);
and U1953 (N_1953,In_62,In_758);
nand U1954 (N_1954,In_662,In_698);
nor U1955 (N_1955,In_312,In_191);
nor U1956 (N_1956,In_583,In_954);
nor U1957 (N_1957,In_725,In_418);
xnor U1958 (N_1958,In_634,In_807);
nand U1959 (N_1959,In_802,In_536);
xnor U1960 (N_1960,In_725,In_845);
or U1961 (N_1961,In_874,In_552);
nand U1962 (N_1962,In_258,In_269);
and U1963 (N_1963,In_375,In_928);
xnor U1964 (N_1964,In_250,In_151);
or U1965 (N_1965,In_36,In_768);
or U1966 (N_1966,In_300,In_611);
xnor U1967 (N_1967,In_517,In_225);
nor U1968 (N_1968,In_297,In_660);
nand U1969 (N_1969,In_431,In_646);
nand U1970 (N_1970,In_239,In_648);
or U1971 (N_1971,In_892,In_222);
or U1972 (N_1972,In_207,In_657);
nand U1973 (N_1973,In_465,In_733);
nand U1974 (N_1974,In_917,In_363);
and U1975 (N_1975,In_162,In_734);
or U1976 (N_1976,In_728,In_609);
nand U1977 (N_1977,In_102,In_584);
nor U1978 (N_1978,In_501,In_741);
xnor U1979 (N_1979,In_521,In_198);
or U1980 (N_1980,In_29,In_766);
and U1981 (N_1981,In_317,In_539);
nand U1982 (N_1982,In_389,In_509);
xnor U1983 (N_1983,In_128,In_514);
xnor U1984 (N_1984,In_630,In_347);
and U1985 (N_1985,In_913,In_888);
or U1986 (N_1986,In_963,In_79);
nor U1987 (N_1987,In_280,In_699);
or U1988 (N_1988,In_68,In_151);
nand U1989 (N_1989,In_274,In_706);
nor U1990 (N_1990,In_487,In_915);
nand U1991 (N_1991,In_773,In_972);
and U1992 (N_1992,In_36,In_38);
and U1993 (N_1993,In_432,In_282);
xor U1994 (N_1994,In_968,In_505);
or U1995 (N_1995,In_251,In_532);
and U1996 (N_1996,In_555,In_387);
and U1997 (N_1997,In_597,In_507);
or U1998 (N_1998,In_122,In_531);
nor U1999 (N_1999,In_753,In_688);
or U2000 (N_2000,N_471,N_746);
xor U2001 (N_2001,N_742,N_269);
xor U2002 (N_2002,N_1868,N_1339);
nor U2003 (N_2003,N_59,N_1264);
and U2004 (N_2004,N_854,N_34);
nand U2005 (N_2005,N_308,N_1401);
nand U2006 (N_2006,N_361,N_1886);
xnor U2007 (N_2007,N_999,N_1414);
and U2008 (N_2008,N_1581,N_727);
or U2009 (N_2009,N_522,N_1307);
xnor U2010 (N_2010,N_717,N_583);
nand U2011 (N_2011,N_1104,N_1603);
or U2012 (N_2012,N_1495,N_403);
and U2013 (N_2013,N_149,N_131);
nand U2014 (N_2014,N_1334,N_716);
xnor U2015 (N_2015,N_782,N_320);
and U2016 (N_2016,N_757,N_1745);
and U2017 (N_2017,N_1281,N_1828);
xor U2018 (N_2018,N_1150,N_133);
nand U2019 (N_2019,N_1650,N_1376);
and U2020 (N_2020,N_1137,N_409);
xnor U2021 (N_2021,N_951,N_381);
nand U2022 (N_2022,N_1017,N_137);
nor U2023 (N_2023,N_950,N_857);
and U2024 (N_2024,N_1683,N_1684);
or U2025 (N_2025,N_1527,N_922);
xor U2026 (N_2026,N_518,N_1557);
xor U2027 (N_2027,N_238,N_1440);
xor U2028 (N_2028,N_635,N_1083);
xor U2029 (N_2029,N_214,N_737);
or U2030 (N_2030,N_1275,N_1102);
nand U2031 (N_2031,N_976,N_1432);
or U2032 (N_2032,N_554,N_89);
nor U2033 (N_2033,N_249,N_1512);
xnor U2034 (N_2034,N_743,N_1464);
or U2035 (N_2035,N_1473,N_424);
and U2036 (N_2036,N_649,N_1192);
or U2037 (N_2037,N_1167,N_1630);
nand U2038 (N_2038,N_1299,N_1730);
nand U2039 (N_2039,N_1571,N_1114);
xnor U2040 (N_2040,N_1491,N_20);
nand U2041 (N_2041,N_970,N_392);
or U2042 (N_2042,N_1072,N_636);
or U2043 (N_2043,N_1795,N_711);
nand U2044 (N_2044,N_1695,N_929);
nor U2045 (N_2045,N_1981,N_1799);
or U2046 (N_2046,N_968,N_1907);
nor U2047 (N_2047,N_1615,N_1113);
nand U2048 (N_2048,N_1201,N_1621);
nor U2049 (N_2049,N_1126,N_433);
xor U2050 (N_2050,N_1124,N_945);
nand U2051 (N_2051,N_707,N_1593);
or U2052 (N_2052,N_973,N_612);
and U2053 (N_2053,N_106,N_1601);
nand U2054 (N_2054,N_1807,N_1225);
and U2055 (N_2055,N_524,N_419);
and U2056 (N_2056,N_1531,N_138);
or U2057 (N_2057,N_1858,N_58);
nand U2058 (N_2058,N_1353,N_1924);
xnor U2059 (N_2059,N_195,N_1012);
or U2060 (N_2060,N_1951,N_1677);
and U2061 (N_2061,N_573,N_1311);
xor U2062 (N_2062,N_1469,N_749);
xnor U2063 (N_2063,N_7,N_460);
xnor U2064 (N_2064,N_1285,N_302);
xor U2065 (N_2065,N_1529,N_1516);
and U2066 (N_2066,N_1091,N_348);
nor U2067 (N_2067,N_1266,N_157);
xnor U2068 (N_2068,N_1867,N_926);
nor U2069 (N_2069,N_700,N_179);
nand U2070 (N_2070,N_1324,N_74);
nor U2071 (N_2071,N_815,N_547);
and U2072 (N_2072,N_24,N_907);
nand U2073 (N_2073,N_1526,N_1530);
nor U2074 (N_2074,N_1269,N_5);
and U2075 (N_2075,N_108,N_1009);
xor U2076 (N_2076,N_1640,N_1826);
nor U2077 (N_2077,N_992,N_537);
and U2078 (N_2078,N_886,N_766);
nor U2079 (N_2079,N_294,N_1093);
xor U2080 (N_2080,N_834,N_1820);
xnor U2081 (N_2081,N_473,N_915);
and U2082 (N_2082,N_178,N_48);
nor U2083 (N_2083,N_299,N_1691);
and U2084 (N_2084,N_809,N_1866);
nor U2085 (N_2085,N_1653,N_1940);
and U2086 (N_2086,N_1336,N_1578);
nand U2087 (N_2087,N_344,N_738);
nand U2088 (N_2088,N_66,N_1437);
nor U2089 (N_2089,N_1520,N_523);
and U2090 (N_2090,N_695,N_1665);
nor U2091 (N_2091,N_847,N_1068);
nand U2092 (N_2092,N_1608,N_336);
nand U2093 (N_2093,N_1096,N_501);
or U2094 (N_2094,N_1233,N_197);
and U2095 (N_2095,N_1060,N_1561);
nand U2096 (N_2096,N_659,N_1628);
and U2097 (N_2097,N_1926,N_875);
nand U2098 (N_2098,N_677,N_1489);
nor U2099 (N_2099,N_1049,N_1818);
and U2100 (N_2100,N_375,N_1172);
or U2101 (N_2101,N_718,N_290);
and U2102 (N_2102,N_1084,N_1407);
xnor U2103 (N_2103,N_1367,N_1160);
nor U2104 (N_2104,N_693,N_648);
or U2105 (N_2105,N_698,N_446);
or U2106 (N_2106,N_1962,N_800);
or U2107 (N_2107,N_1816,N_1830);
xor U2108 (N_2108,N_1941,N_1917);
and U2109 (N_2109,N_1528,N_1077);
xnor U2110 (N_2110,N_1026,N_1203);
and U2111 (N_2111,N_1193,N_1323);
nand U2112 (N_2112,N_1610,N_1051);
nor U2113 (N_2113,N_350,N_241);
and U2114 (N_2114,N_856,N_1577);
nor U2115 (N_2115,N_1176,N_1788);
nand U2116 (N_2116,N_338,N_194);
nor U2117 (N_2117,N_1525,N_1048);
or U2118 (N_2118,N_1483,N_1293);
or U2119 (N_2119,N_1050,N_790);
nand U2120 (N_2120,N_1310,N_1344);
nor U2121 (N_2121,N_835,N_1613);
xor U2122 (N_2122,N_597,N_1287);
nor U2123 (N_2123,N_692,N_1993);
or U2124 (N_2124,N_644,N_980);
nor U2125 (N_2125,N_1257,N_882);
or U2126 (N_2126,N_223,N_461);
or U2127 (N_2127,N_1286,N_1121);
nor U2128 (N_2128,N_721,N_1800);
nand U2129 (N_2129,N_134,N_19);
and U2130 (N_2130,N_1064,N_1133);
nand U2131 (N_2131,N_1427,N_289);
and U2132 (N_2132,N_78,N_1261);
or U2133 (N_2133,N_1067,N_1181);
or U2134 (N_2134,N_1219,N_1802);
nand U2135 (N_2135,N_665,N_1115);
nor U2136 (N_2136,N_641,N_1002);
xor U2137 (N_2137,N_822,N_1063);
nand U2138 (N_2138,N_1547,N_953);
xor U2139 (N_2139,N_939,N_1622);
xor U2140 (N_2140,N_1715,N_203);
or U2141 (N_2141,N_1395,N_492);
or U2142 (N_2142,N_1027,N_795);
and U2143 (N_2143,N_511,N_1921);
nand U2144 (N_2144,N_53,N_971);
nand U2145 (N_2145,N_1862,N_1487);
or U2146 (N_2146,N_1748,N_65);
nand U2147 (N_2147,N_1726,N_1156);
and U2148 (N_2148,N_628,N_1689);
xor U2149 (N_2149,N_1216,N_1769);
nor U2150 (N_2150,N_569,N_921);
or U2151 (N_2151,N_832,N_1057);
or U2152 (N_2152,N_719,N_878);
xnor U2153 (N_2153,N_802,N_1108);
nor U2154 (N_2154,N_322,N_579);
and U2155 (N_2155,N_46,N_1517);
and U2156 (N_2156,N_586,N_1003);
xnor U2157 (N_2157,N_755,N_1345);
or U2158 (N_2158,N_243,N_1152);
or U2159 (N_2159,N_1479,N_352);
nor U2160 (N_2160,N_705,N_885);
or U2161 (N_2161,N_1641,N_1117);
xnor U2162 (N_2162,N_891,N_80);
nor U2163 (N_2163,N_1198,N_1869);
xor U2164 (N_2164,N_1348,N_825);
and U2165 (N_2165,N_188,N_591);
and U2166 (N_2166,N_829,N_725);
xor U2167 (N_2167,N_791,N_1184);
and U2168 (N_2168,N_867,N_587);
nand U2169 (N_2169,N_897,N_873);
nand U2170 (N_2170,N_1087,N_564);
and U2171 (N_2171,N_1379,N_812);
nor U2172 (N_2172,N_483,N_1758);
nor U2173 (N_2173,N_660,N_368);
nor U2174 (N_2174,N_1403,N_837);
or U2175 (N_2175,N_1729,N_1922);
nand U2176 (N_2176,N_342,N_803);
nand U2177 (N_2177,N_1971,N_1699);
nand U2178 (N_2178,N_1162,N_1036);
nor U2179 (N_2179,N_1980,N_1588);
and U2180 (N_2180,N_995,N_229);
nor U2181 (N_2181,N_1447,N_231);
and U2182 (N_2182,N_1189,N_874);
nor U2183 (N_2183,N_366,N_964);
nand U2184 (N_2184,N_1001,N_291);
nand U2185 (N_2185,N_396,N_672);
and U2186 (N_2186,N_696,N_836);
and U2187 (N_2187,N_470,N_516);
nor U2188 (N_2188,N_240,N_1296);
nand U2189 (N_2189,N_1766,N_192);
or U2190 (N_2190,N_566,N_1315);
xor U2191 (N_2191,N_175,N_1508);
nor U2192 (N_2192,N_437,N_1846);
or U2193 (N_2193,N_1082,N_817);
or U2194 (N_2194,N_706,N_1633);
and U2195 (N_2195,N_42,N_391);
and U2196 (N_2196,N_1902,N_1062);
nand U2197 (N_2197,N_373,N_1471);
nand U2198 (N_2198,N_627,N_855);
nor U2199 (N_2199,N_1270,N_1053);
or U2200 (N_2200,N_452,N_1654);
and U2201 (N_2201,N_216,N_1038);
nand U2202 (N_2202,N_590,N_578);
nor U2203 (N_2203,N_442,N_1331);
nand U2204 (N_2204,N_1870,N_1229);
xnor U2205 (N_2205,N_571,N_624);
xnor U2206 (N_2206,N_1493,N_270);
xor U2207 (N_2207,N_160,N_1812);
xor U2208 (N_2208,N_783,N_1058);
or U2209 (N_2209,N_625,N_1085);
and U2210 (N_2210,N_451,N_779);
or U2211 (N_2211,N_1194,N_1510);
xnor U2212 (N_2212,N_546,N_228);
nand U2213 (N_2213,N_1005,N_1514);
nand U2214 (N_2214,N_1207,N_986);
nor U2215 (N_2215,N_1943,N_588);
nor U2216 (N_2216,N_1488,N_101);
xnor U2217 (N_2217,N_475,N_543);
nand U2218 (N_2218,N_458,N_1777);
or U2219 (N_2219,N_703,N_1134);
or U2220 (N_2220,N_315,N_778);
xnor U2221 (N_2221,N_1366,N_1365);
nor U2222 (N_2222,N_193,N_887);
and U2223 (N_2223,N_1511,N_498);
nand U2224 (N_2224,N_1912,N_187);
and U2225 (N_2225,N_983,N_1056);
nand U2226 (N_2226,N_255,N_1765);
or U2227 (N_2227,N_64,N_1627);
and U2228 (N_2228,N_1556,N_337);
or U2229 (N_2229,N_1019,N_1438);
xnor U2230 (N_2230,N_1723,N_420);
xor U2231 (N_2231,N_1794,N_889);
xor U2232 (N_2232,N_467,N_1811);
xnor U2233 (N_2233,N_1781,N_892);
or U2234 (N_2234,N_1934,N_129);
nand U2235 (N_2235,N_1078,N_1475);
xor U2236 (N_2236,N_485,N_1532);
xnor U2237 (N_2237,N_1899,N_1059);
and U2238 (N_2238,N_949,N_1524);
or U2239 (N_2239,N_1635,N_77);
or U2240 (N_2240,N_1463,N_1970);
xor U2241 (N_2241,N_928,N_177);
and U2242 (N_2242,N_544,N_94);
nor U2243 (N_2243,N_1840,N_62);
nand U2244 (N_2244,N_152,N_1634);
xor U2245 (N_2245,N_1675,N_165);
nand U2246 (N_2246,N_865,N_557);
xor U2247 (N_2247,N_476,N_919);
nand U2248 (N_2248,N_1918,N_1923);
nor U2249 (N_2249,N_1791,N_455);
and U2250 (N_2250,N_1851,N_421);
or U2251 (N_2251,N_690,N_1406);
nor U2252 (N_2252,N_490,N_1140);
and U2253 (N_2253,N_1276,N_1265);
and U2254 (N_2254,N_923,N_1544);
xnor U2255 (N_2255,N_977,N_1171);
nand U2256 (N_2256,N_561,N_1982);
nor U2257 (N_2257,N_709,N_1537);
nor U2258 (N_2258,N_910,N_275);
nand U2259 (N_2259,N_917,N_1822);
nand U2260 (N_2260,N_345,N_390);
xnor U2261 (N_2261,N_4,N_503);
or U2262 (N_2262,N_1541,N_1903);
xnor U2263 (N_2263,N_1566,N_657);
nor U2264 (N_2264,N_1045,N_314);
and U2265 (N_2265,N_1564,N_1881);
nor U2266 (N_2266,N_43,N_793);
nor U2267 (N_2267,N_678,N_1245);
and U2268 (N_2268,N_1563,N_1289);
xor U2269 (N_2269,N_351,N_1901);
nand U2270 (N_2270,N_1103,N_1555);
and U2271 (N_2271,N_372,N_296);
nor U2272 (N_2272,N_1435,N_439);
xnor U2273 (N_2273,N_1241,N_1455);
and U2274 (N_2274,N_1377,N_1513);
xnor U2275 (N_2275,N_35,N_519);
xnor U2276 (N_2276,N_70,N_729);
nor U2277 (N_2277,N_981,N_1461);
and U2278 (N_2278,N_208,N_401);
and U2279 (N_2279,N_1280,N_1237);
nor U2280 (N_2280,N_634,N_1371);
nand U2281 (N_2281,N_1803,N_1070);
nor U2282 (N_2282,N_1277,N_1985);
and U2283 (N_2283,N_552,N_1255);
nor U2284 (N_2284,N_1094,N_714);
nand U2285 (N_2285,N_1480,N_1186);
nor U2286 (N_2286,N_158,N_1105);
nor U2287 (N_2287,N_549,N_371);
and U2288 (N_2288,N_472,N_1550);
nand U2289 (N_2289,N_667,N_423);
xnor U2290 (N_2290,N_602,N_1839);
and U2291 (N_2291,N_1925,N_772);
nand U2292 (N_2292,N_164,N_1211);
nor U2293 (N_2293,N_236,N_1753);
or U2294 (N_2294,N_144,N_204);
or U2295 (N_2295,N_828,N_510);
nor U2296 (N_2296,N_1243,N_227);
xor U2297 (N_2297,N_1873,N_1288);
nor U2298 (N_2298,N_1262,N_893);
and U2299 (N_2299,N_1565,N_1492);
or U2300 (N_2300,N_1118,N_1500);
or U2301 (N_2301,N_1232,N_1957);
or U2302 (N_2302,N_1597,N_1928);
and U2303 (N_2303,N_1725,N_162);
nor U2304 (N_2304,N_844,N_1533);
xnor U2305 (N_2305,N_380,N_944);
nand U2306 (N_2306,N_417,N_1953);
or U2307 (N_2307,N_934,N_1625);
nand U2308 (N_2308,N_1942,N_1761);
nand U2309 (N_2309,N_1031,N_1883);
nor U2310 (N_2310,N_1909,N_284);
and U2311 (N_2311,N_1195,N_978);
xnor U2312 (N_2312,N_1474,N_1877);
nor U2313 (N_2313,N_365,N_1039);
xor U2314 (N_2314,N_916,N_1430);
nand U2315 (N_2315,N_876,N_1560);
or U2316 (N_2316,N_261,N_57);
and U2317 (N_2317,N_1200,N_1385);
nand U2318 (N_2318,N_1671,N_1421);
nand U2319 (N_2319,N_1260,N_1099);
and U2320 (N_2320,N_1743,N_422);
nor U2321 (N_2321,N_898,N_210);
nand U2322 (N_2322,N_1596,N_1221);
xor U2323 (N_2323,N_768,N_997);
and U2324 (N_2324,N_1369,N_1620);
and U2325 (N_2325,N_689,N_1959);
or U2326 (N_2326,N_1485,N_1504);
or U2327 (N_2327,N_609,N_112);
or U2328 (N_2328,N_1010,N_1125);
xor U2329 (N_2329,N_1948,N_1111);
xnor U2330 (N_2330,N_1178,N_1518);
nand U2331 (N_2331,N_1011,N_147);
or U2332 (N_2332,N_1294,N_751);
nand U2333 (N_2333,N_140,N_1700);
nand U2334 (N_2334,N_237,N_715);
or U2335 (N_2335,N_76,N_1704);
xor U2336 (N_2336,N_1000,N_896);
or U2337 (N_2337,N_1484,N_356);
and U2338 (N_2338,N_87,N_379);
xnor U2339 (N_2339,N_1465,N_1810);
and U2340 (N_2340,N_124,N_1600);
nand U2341 (N_2341,N_479,N_226);
nand U2342 (N_2342,N_49,N_1894);
nor U2343 (N_2343,N_786,N_736);
or U2344 (N_2344,N_79,N_1789);
nor U2345 (N_2345,N_1747,N_1905);
or U2346 (N_2346,N_998,N_434);
nor U2347 (N_2347,N_697,N_1605);
or U2348 (N_2348,N_100,N_72);
nand U2349 (N_2349,N_1016,N_353);
xnor U2350 (N_2350,N_1204,N_1845);
nor U2351 (N_2351,N_1984,N_95);
or U2352 (N_2352,N_1764,N_153);
nand U2353 (N_2353,N_1383,N_254);
nand U2354 (N_2354,N_957,N_797);
and U2355 (N_2355,N_645,N_47);
nor U2356 (N_2356,N_1678,N_1013);
nand U2357 (N_2357,N_1545,N_572);
or U2358 (N_2358,N_913,N_448);
xnor U2359 (N_2359,N_1554,N_1988);
or U2360 (N_2360,N_1449,N_1669);
xor U2361 (N_2361,N_1263,N_185);
nand U2362 (N_2362,N_942,N_1703);
nand U2363 (N_2363,N_1954,N_413);
nand U2364 (N_2364,N_1817,N_1429);
and U2365 (N_2365,N_1770,N_1505);
nor U2366 (N_2366,N_1806,N_538);
nor U2367 (N_2367,N_151,N_1143);
or U2368 (N_2368,N_679,N_1249);
xor U2369 (N_2369,N_1169,N_1843);
xnor U2370 (N_2370,N_622,N_382);
or U2371 (N_2371,N_186,N_1833);
nand U2372 (N_2372,N_123,N_318);
nand U2373 (N_2373,N_506,N_1247);
xnor U2374 (N_2374,N_1579,N_107);
nand U2375 (N_2375,N_1874,N_947);
and U2376 (N_2376,N_600,N_1089);
and U2377 (N_2377,N_1419,N_1222);
nand U2378 (N_2378,N_385,N_346);
xnor U2379 (N_2379,N_1744,N_1977);
nand U2380 (N_2380,N_239,N_710);
xor U2381 (N_2381,N_1141,N_548);
and U2382 (N_2382,N_595,N_642);
xor U2383 (N_2383,N_935,N_1880);
nor U2384 (N_2384,N_1707,N_1428);
or U2385 (N_2385,N_861,N_621);
or U2386 (N_2386,N_267,N_903);
or U2387 (N_2387,N_1415,N_1022);
xnor U2388 (N_2388,N_1673,N_96);
and U2389 (N_2389,N_699,N_1693);
and U2390 (N_2390,N_1284,N_242);
nand U2391 (N_2391,N_606,N_769);
and U2392 (N_2392,N_1655,N_540);
nor U2393 (N_2393,N_713,N_456);
nand U2394 (N_2394,N_1737,N_1028);
or U2395 (N_2395,N_1997,N_765);
nor U2396 (N_2396,N_1210,N_1844);
and U2397 (N_2397,N_1523,N_325);
and U2398 (N_2398,N_1235,N_171);
or U2399 (N_2399,N_568,N_1963);
nand U2400 (N_2400,N_990,N_1303);
and U2401 (N_2401,N_507,N_1779);
nand U2402 (N_2402,N_445,N_1662);
and U2403 (N_2403,N_1944,N_1657);
xor U2404 (N_2404,N_1298,N_1047);
nor U2405 (N_2405,N_21,N_1842);
and U2406 (N_2406,N_438,N_1515);
and U2407 (N_2407,N_760,N_1130);
xor U2408 (N_2408,N_85,N_440);
nand U2409 (N_2409,N_1384,N_539);
xnor U2410 (N_2410,N_1969,N_494);
or U2411 (N_2411,N_858,N_1835);
or U2412 (N_2412,N_1496,N_545);
nor U2413 (N_2413,N_258,N_1920);
xor U2414 (N_2414,N_1127,N_1879);
nor U2415 (N_2415,N_1418,N_668);
xnor U2416 (N_2416,N_69,N_906);
or U2417 (N_2417,N_1044,N_1043);
nor U2418 (N_2418,N_1351,N_1754);
xor U2419 (N_2419,N_979,N_1180);
nand U2420 (N_2420,N_1785,N_1197);
nand U2421 (N_2421,N_1244,N_343);
and U2422 (N_2422,N_1895,N_638);
nand U2423 (N_2423,N_1041,N_1347);
xor U2424 (N_2424,N_1567,N_1268);
and U2425 (N_2425,N_1732,N_515);
xor U2426 (N_2426,N_202,N_222);
or U2427 (N_2427,N_491,N_16);
and U2428 (N_2428,N_1301,N_313);
or U2429 (N_2429,N_1606,N_257);
or U2430 (N_2430,N_816,N_170);
xnor U2431 (N_2431,N_724,N_444);
xnor U2432 (N_2432,N_1446,N_1205);
nand U2433 (N_2433,N_534,N_1123);
nor U2434 (N_2434,N_1340,N_307);
or U2435 (N_2435,N_63,N_754);
nor U2436 (N_2436,N_839,N_1538);
and U2437 (N_2437,N_1297,N_75);
and U2438 (N_2438,N_1904,N_787);
nor U2439 (N_2439,N_1431,N_555);
or U2440 (N_2440,N_1179,N_1402);
nand U2441 (N_2441,N_656,N_1898);
nand U2442 (N_2442,N_1034,N_1317);
xor U2443 (N_2443,N_477,N_266);
nor U2444 (N_2444,N_1604,N_528);
xor U2445 (N_2445,N_432,N_136);
or U2446 (N_2446,N_1652,N_367);
nor U2447 (N_2447,N_735,N_1424);
xnor U2448 (N_2448,N_1617,N_804);
or U2449 (N_2449,N_708,N_3);
and U2450 (N_2450,N_1486,N_418);
and U2451 (N_2451,N_1872,N_427);
or U2452 (N_2452,N_744,N_1226);
and U2453 (N_2453,N_1136,N_1539);
nand U2454 (N_2454,N_1476,N_1372);
and U2455 (N_2455,N_1316,N_468);
nor U2456 (N_2456,N_1937,N_673);
nand U2457 (N_2457,N_982,N_415);
nand U2458 (N_2458,N_1863,N_1052);
xnor U2459 (N_2459,N_1782,N_541);
nor U2460 (N_2460,N_376,N_1759);
and U2461 (N_2461,N_1956,N_559);
nand U2462 (N_2462,N_1787,N_1592);
nor U2463 (N_2463,N_1196,N_213);
and U2464 (N_2464,N_1456,N_1967);
nor U2465 (N_2465,N_400,N_1182);
and U2466 (N_2466,N_1570,N_1774);
or U2467 (N_2467,N_1815,N_527);
xor U2468 (N_2468,N_1423,N_1760);
nor U2469 (N_2469,N_142,N_1658);
or U2470 (N_2470,N_81,N_1054);
or U2471 (N_2471,N_680,N_1173);
nor U2472 (N_2472,N_675,N_395);
xor U2473 (N_2473,N_1636,N_311);
or U2474 (N_2474,N_1467,N_647);
nand U2475 (N_2475,N_1177,N_1014);
nor U2476 (N_2476,N_1408,N_480);
or U2477 (N_2477,N_463,N_1497);
nand U2478 (N_2478,N_762,N_181);
or U2479 (N_2479,N_1950,N_1021);
and U2480 (N_2480,N_1599,N_404);
nor U2481 (N_2481,N_334,N_1468);
and U2482 (N_2482,N_1792,N_862);
and U2483 (N_2483,N_39,N_1780);
nor U2484 (N_2484,N_30,N_1411);
xor U2485 (N_2485,N_1680,N_1046);
xnor U2486 (N_2486,N_1721,N_1460);
nor U2487 (N_2487,N_1559,N_1821);
or U2488 (N_2488,N_1661,N_792);
nand U2489 (N_2489,N_740,N_630);
or U2490 (N_2490,N_488,N_870);
nor U2491 (N_2491,N_652,N_1995);
nand U2492 (N_2492,N_1442,N_619);
or U2493 (N_2493,N_946,N_215);
and U2494 (N_2494,N_1676,N_1522);
nand U2495 (N_2495,N_1338,N_155);
or U2496 (N_2496,N_73,N_388);
nor U2497 (N_2497,N_894,N_758);
and U2498 (N_2498,N_987,N_1832);
nand U2499 (N_2499,N_97,N_701);
nand U2500 (N_2500,N_12,N_384);
nor U2501 (N_2501,N_38,N_196);
or U2502 (N_2502,N_1472,N_1801);
nor U2503 (N_2503,N_402,N_1343);
or U2504 (N_2504,N_848,N_1252);
xnor U2505 (N_2505,N_1300,N_932);
nand U2506 (N_2506,N_68,N_775);
or U2507 (N_2507,N_1035,N_1313);
or U2508 (N_2508,N_1163,N_1206);
and U2509 (N_2509,N_1309,N_172);
nor U2510 (N_2510,N_209,N_416);
or U2511 (N_2511,N_1887,N_224);
nand U2512 (N_2512,N_1109,N_1509);
xnor U2513 (N_2513,N_1931,N_925);
xnor U2514 (N_2514,N_1238,N_526);
and U2515 (N_2515,N_1100,N_1457);
and U2516 (N_2516,N_1400,N_317);
and U2517 (N_2517,N_259,N_1973);
nand U2518 (N_2518,N_1998,N_731);
nor U2519 (N_2519,N_1490,N_1482);
xor U2520 (N_2520,N_1081,N_1212);
nor U2521 (N_2521,N_1290,N_1306);
and U2522 (N_2522,N_486,N_796);
nor U2523 (N_2523,N_31,N_1534);
nand U2524 (N_2524,N_533,N_1018);
and U2525 (N_2525,N_1896,N_965);
nor U2526 (N_2526,N_33,N_788);
xnor U2527 (N_2527,N_1236,N_304);
and U2528 (N_2528,N_1733,N_620);
nand U2529 (N_2529,N_1332,N_605);
nor U2530 (N_2530,N_1521,N_377);
nor U2531 (N_2531,N_6,N_316);
nand U2532 (N_2532,N_1425,N_752);
and U2533 (N_2533,N_1352,N_1413);
nor U2534 (N_2534,N_14,N_341);
nor U2535 (N_2535,N_550,N_1337);
and U2536 (N_2536,N_1631,N_1572);
and U2537 (N_2537,N_22,N_1705);
nand U2538 (N_2538,N_128,N_1656);
nand U2539 (N_2539,N_952,N_774);
xor U2540 (N_2540,N_83,N_558);
nor U2541 (N_2541,N_121,N_669);
or U2542 (N_2542,N_1796,N_1139);
nand U2543 (N_2543,N_938,N_582);
nor U2544 (N_2544,N_247,N_739);
xor U2545 (N_2545,N_1763,N_1359);
nor U2546 (N_2546,N_1008,N_449);
xor U2547 (N_2547,N_1755,N_631);
nand U2548 (N_2548,N_278,N_1363);
xor U2549 (N_2549,N_1217,N_110);
or U2550 (N_2550,N_764,N_972);
and U2551 (N_2551,N_29,N_1499);
nand U2552 (N_2552,N_1623,N_1328);
nand U2553 (N_2553,N_1974,N_1246);
or U2554 (N_2554,N_1619,N_0);
or U2555 (N_2555,N_274,N_1850);
xor U2556 (N_2556,N_1146,N_937);
xnor U2557 (N_2557,N_309,N_1481);
or U2558 (N_2558,N_1914,N_148);
xnor U2559 (N_2559,N_508,N_653);
or U2560 (N_2560,N_1155,N_1387);
or U2561 (N_2561,N_996,N_1079);
nor U2562 (N_2562,N_285,N_109);
nor U2563 (N_2563,N_264,N_851);
and U2564 (N_2564,N_563,N_1396);
nand U2565 (N_2565,N_60,N_688);
and U2566 (N_2566,N_1302,N_598);
or U2567 (N_2567,N_1305,N_262);
nand U2568 (N_2568,N_1889,N_414);
or U2569 (N_2569,N_560,N_201);
nand U2570 (N_2570,N_1690,N_801);
nand U2571 (N_2571,N_1915,N_86);
and U2572 (N_2572,N_702,N_1930);
or U2573 (N_2573,N_813,N_819);
xor U2574 (N_2574,N_1731,N_643);
nand U2575 (N_2575,N_1295,N_1587);
nand U2576 (N_2576,N_1291,N_386);
and U2577 (N_2577,N_1335,N_674);
xnor U2578 (N_2578,N_1836,N_940);
nor U2579 (N_2579,N_1258,N_1107);
xor U2580 (N_2580,N_811,N_1314);
or U2581 (N_2581,N_1075,N_960);
nand U2582 (N_2582,N_105,N_1506);
nand U2583 (N_2583,N_849,N_1685);
and U2584 (N_2584,N_1553,N_1562);
or U2585 (N_2585,N_722,N_741);
nor U2586 (N_2586,N_1090,N_1042);
nand U2587 (N_2587,N_868,N_271);
nor U2588 (N_2588,N_363,N_1734);
or U2589 (N_2589,N_888,N_26);
xnor U2590 (N_2590,N_1390,N_502);
nand U2591 (N_2591,N_1853,N_1061);
or U2592 (N_2592,N_10,N_1738);
and U2593 (N_2593,N_1947,N_277);
xor U2594 (N_2594,N_1913,N_1996);
or U2595 (N_2595,N_1837,N_1852);
nand U2596 (N_2596,N_607,N_13);
and U2597 (N_2597,N_956,N_1961);
and U2598 (N_2598,N_1746,N_132);
xnor U2599 (N_2599,N_581,N_349);
or U2600 (N_2600,N_298,N_1955);
nor U2601 (N_2601,N_1098,N_530);
xnor U2602 (N_2602,N_126,N_1972);
xnor U2603 (N_2603,N_1712,N_1576);
nand U2604 (N_2604,N_1536,N_1242);
xor U2605 (N_2605,N_1370,N_1378);
nor U2606 (N_2606,N_18,N_1589);
xor U2607 (N_2607,N_1132,N_1535);
xnor U2608 (N_2608,N_1320,N_1586);
and U2609 (N_2609,N_1501,N_301);
nand U2610 (N_2610,N_1986,N_1416);
or U2611 (N_2611,N_1989,N_462);
nand U2612 (N_2612,N_1065,N_114);
nand U2613 (N_2613,N_1404,N_1071);
xor U2614 (N_2614,N_27,N_871);
nor U2615 (N_2615,N_912,N_1166);
xnor U2616 (N_2616,N_1202,N_1607);
and U2617 (N_2617,N_1020,N_576);
or U2618 (N_2618,N_640,N_36);
nand U2619 (N_2619,N_211,N_1936);
and U2620 (N_2620,N_1272,N_362);
and U2621 (N_2621,N_993,N_1569);
or U2622 (N_2622,N_975,N_777);
nand U2623 (N_2623,N_56,N_399);
nand U2624 (N_2624,N_1580,N_253);
nor U2625 (N_2625,N_633,N_1076);
or U2626 (N_2626,N_1271,N_1282);
and U2627 (N_2627,N_1742,N_103);
and U2628 (N_2628,N_1549,N_1354);
nand U2629 (N_2629,N_1398,N_273);
xor U2630 (N_2630,N_969,N_1187);
or U2631 (N_2631,N_664,N_616);
nor U2632 (N_2632,N_850,N_1097);
nand U2633 (N_2633,N_1426,N_1805);
nor U2634 (N_2634,N_899,N_726);
nand U2635 (N_2635,N_355,N_954);
or U2636 (N_2636,N_333,N_1834);
nand U2637 (N_2637,N_1088,N_1546);
or U2638 (N_2638,N_474,N_529);
nand U2639 (N_2639,N_119,N_525);
or U2640 (N_2640,N_1639,N_1120);
and U2641 (N_2641,N_601,N_1223);
or U2642 (N_2642,N_904,N_1389);
nor U2643 (N_2643,N_959,N_720);
nor U2644 (N_2644,N_205,N_1767);
nor U2645 (N_2645,N_1106,N_1386);
xor U2646 (N_2646,N_936,N_45);
xnor U2647 (N_2647,N_859,N_1);
nor U2648 (N_2648,N_963,N_1149);
xor U2649 (N_2649,N_1958,N_1900);
nor U2650 (N_2650,N_1735,N_500);
xor U2651 (N_2651,N_864,N_1023);
xor U2652 (N_2652,N_808,N_1185);
and U2653 (N_2653,N_1674,N_771);
nor U2654 (N_2654,N_872,N_1208);
xor U2655 (N_2655,N_1350,N_728);
xnor U2656 (N_2656,N_1848,N_1092);
or U2657 (N_2657,N_831,N_406);
nand U2658 (N_2658,N_323,N_1992);
or U2659 (N_2659,N_807,N_1004);
nor U2660 (N_2660,N_1254,N_1380);
xnor U2661 (N_2661,N_608,N_712);
or U2662 (N_2662,N_1624,N_1916);
or U2663 (N_2663,N_574,N_1584);
nand U2664 (N_2664,N_985,N_1714);
nand U2665 (N_2665,N_1702,N_1616);
nor U2666 (N_2666,N_232,N_1614);
nand U2667 (N_2667,N_1308,N_1025);
nand U2668 (N_2668,N_496,N_191);
or U2669 (N_2669,N_670,N_1319);
or U2670 (N_2670,N_1809,N_248);
nand U2671 (N_2671,N_339,N_682);
and U2672 (N_2672,N_50,N_453);
nand U2673 (N_2673,N_1772,N_1849);
xnor U2674 (N_2674,N_265,N_1583);
or U2675 (N_2675,N_1253,N_1585);
nor U2676 (N_2676,N_1643,N_1558);
xor U2677 (N_2677,N_784,N_1722);
or U2678 (N_2678,N_1720,N_1595);
nor U2679 (N_2679,N_1860,N_167);
or U2680 (N_2680,N_1329,N_1304);
nand U2681 (N_2681,N_1831,N_328);
nor U2682 (N_2682,N_176,N_1074);
xor U2683 (N_2683,N_1667,N_1405);
or U2684 (N_2684,N_1234,N_584);
nor U2685 (N_2685,N_310,N_268);
xor U2686 (N_2686,N_1644,N_331);
or U2687 (N_2687,N_637,N_908);
nand U2688 (N_2688,N_1341,N_509);
nor U2689 (N_2689,N_1283,N_1417);
and U2690 (N_2690,N_1910,N_1267);
nor U2691 (N_2691,N_948,N_481);
nand U2692 (N_2692,N_1462,N_658);
nor U2693 (N_2693,N_1990,N_1875);
or U2694 (N_2694,N_512,N_900);
and U2695 (N_2695,N_1736,N_359);
or U2696 (N_2696,N_1598,N_292);
nand U2697 (N_2697,N_671,N_1502);
nand U2698 (N_2698,N_1228,N_556);
nor U2699 (N_2699,N_1259,N_517);
or U2700 (N_2700,N_1548,N_1420);
nor U2701 (N_2701,N_694,N_1142);
and U2702 (N_2702,N_387,N_895);
nand U2703 (N_2703,N_429,N_1165);
nor U2704 (N_2704,N_890,N_1711);
xnor U2705 (N_2705,N_370,N_1751);
or U2706 (N_2706,N_833,N_1991);
nor U2707 (N_2707,N_430,N_378);
xor U2708 (N_2708,N_1322,N_798);
and U2709 (N_2709,N_1214,N_1666);
and U2710 (N_2710,N_28,N_1919);
nor U2711 (N_2711,N_330,N_853);
nand U2712 (N_2712,N_306,N_974);
nor U2713 (N_2713,N_1543,N_1368);
nand U2714 (N_2714,N_1888,N_1728);
and U2715 (N_2715,N_863,N_184);
nand U2716 (N_2716,N_272,N_1024);
and U2717 (N_2717,N_1632,N_1908);
nand U2718 (N_2718,N_881,N_773);
nor U2719 (N_2719,N_1670,N_759);
or U2720 (N_2720,N_1434,N_1507);
nor U2721 (N_2721,N_651,N_130);
or U2722 (N_2722,N_984,N_200);
and U2723 (N_2723,N_283,N_1356);
or U2724 (N_2724,N_190,N_161);
nor U2725 (N_2725,N_1191,N_37);
nand U2726 (N_2726,N_1679,N_1719);
xor U2727 (N_2727,N_593,N_877);
or U2728 (N_2728,N_1752,N_1412);
and U2729 (N_2729,N_329,N_410);
nor U2730 (N_2730,N_1122,N_1159);
or U2731 (N_2731,N_681,N_32);
nor U2732 (N_2732,N_905,N_666);
nor U2733 (N_2733,N_487,N_733);
and U2734 (N_2734,N_497,N_91);
xor U2735 (N_2735,N_408,N_122);
or U2736 (N_2736,N_88,N_1664);
nand U2737 (N_2737,N_2,N_1663);
or U2738 (N_2738,N_918,N_312);
xor U2739 (N_2739,N_596,N_1618);
and U2740 (N_2740,N_1648,N_763);
or U2741 (N_2741,N_360,N_821);
nand U2742 (N_2742,N_1865,N_1066);
xnor U2743 (N_2743,N_1575,N_233);
nand U2744 (N_2744,N_1709,N_1519);
and U2745 (N_2745,N_1101,N_482);
xor U2746 (N_2746,N_1073,N_1015);
xnor U2747 (N_2747,N_1360,N_398);
nor U2748 (N_2748,N_1927,N_623);
nand U2749 (N_2749,N_1741,N_189);
xor U2750 (N_2750,N_1854,N_852);
and U2751 (N_2751,N_745,N_1602);
xor U2752 (N_2752,N_1399,N_1771);
and U2753 (N_2753,N_1542,N_1983);
nor U2754 (N_2754,N_465,N_104);
and U2755 (N_2755,N_958,N_1827);
and U2756 (N_2756,N_988,N_1692);
nand U2757 (N_2757,N_962,N_1231);
nor U2758 (N_2758,N_1949,N_1220);
nand U2759 (N_2759,N_1706,N_288);
nor U2760 (N_2760,N_98,N_730);
xor U2761 (N_2761,N_1224,N_369);
and U2762 (N_2762,N_198,N_1422);
nand U2763 (N_2763,N_909,N_1727);
and U2764 (N_2764,N_1321,N_1778);
nor U2765 (N_2765,N_340,N_436);
or U2766 (N_2766,N_1775,N_1382);
or U2767 (N_2767,N_41,N_1450);
nor U2768 (N_2768,N_1444,N_1029);
nand U2769 (N_2769,N_450,N_838);
nor U2770 (N_2770,N_23,N_173);
and U2771 (N_2771,N_489,N_1864);
or U2772 (N_2772,N_686,N_901);
and U2773 (N_2773,N_55,N_141);
or U2774 (N_2774,N_245,N_553);
nor U2775 (N_2775,N_1965,N_260);
nor U2776 (N_2776,N_11,N_521);
or U2777 (N_2777,N_691,N_1933);
and U2778 (N_2778,N_321,N_626);
xor U2779 (N_2779,N_1776,N_326);
xor U2780 (N_2780,N_846,N_102);
xor U2781 (N_2781,N_676,N_484);
and U2782 (N_2782,N_1443,N_1147);
and U2783 (N_2783,N_1388,N_1138);
or U2784 (N_2784,N_113,N_943);
nor U2785 (N_2785,N_1797,N_1975);
nor U2786 (N_2786,N_1968,N_1696);
nand U2787 (N_2787,N_163,N_535);
nor U2788 (N_2788,N_407,N_684);
nand U2789 (N_2789,N_1498,N_1938);
nand U2790 (N_2790,N_1355,N_1668);
or U2791 (N_2791,N_770,N_44);
nor U2792 (N_2792,N_207,N_295);
and U2793 (N_2793,N_860,N_1740);
xor U2794 (N_2794,N_704,N_1813);
or U2795 (N_2795,N_1708,N_806);
nor U2796 (N_2796,N_256,N_206);
xnor U2797 (N_2797,N_1342,N_156);
nor U2798 (N_2798,N_1215,N_1032);
xnor U2799 (N_2799,N_1273,N_441);
nor U2800 (N_2800,N_1466,N_218);
nand U2801 (N_2801,N_1503,N_1161);
nand U2802 (N_2802,N_443,N_618);
nor U2803 (N_2803,N_466,N_1856);
and U2804 (N_2804,N_1478,N_1218);
and U2805 (N_2805,N_1540,N_1333);
xnor U2806 (N_2806,N_1590,N_880);
and U2807 (N_2807,N_234,N_1629);
nand U2808 (N_2808,N_1278,N_150);
and U2809 (N_2809,N_603,N_111);
or U2810 (N_2810,N_90,N_1213);
nand U2811 (N_2811,N_174,N_1312);
nor U2812 (N_2812,N_1274,N_459);
or U2813 (N_2813,N_1756,N_1151);
nor U2814 (N_2814,N_405,N_1932);
nor U2815 (N_2815,N_1394,N_1637);
xor U2816 (N_2816,N_1568,N_823);
nand U2817 (N_2817,N_1410,N_654);
and U2818 (N_2818,N_826,N_1451);
nor U2819 (N_2819,N_117,N_662);
xor U2820 (N_2820,N_1361,N_219);
nand U2821 (N_2821,N_1718,N_303);
and U2822 (N_2822,N_930,N_747);
or U2823 (N_2823,N_1688,N_454);
and U2824 (N_2824,N_499,N_287);
or U2825 (N_2825,N_159,N_1935);
or U2826 (N_2826,N_135,N_1594);
or U2827 (N_2827,N_305,N_924);
and U2828 (N_2828,N_599,N_748);
xnor U2829 (N_2829,N_282,N_1841);
nand U2830 (N_2830,N_1409,N_220);
nand U2831 (N_2831,N_1929,N_354);
nand U2832 (N_2832,N_580,N_1251);
xnor U2833 (N_2833,N_1183,N_879);
and U2834 (N_2834,N_383,N_1037);
nor U2835 (N_2835,N_562,N_639);
and U2836 (N_2836,N_1256,N_1349);
nand U2837 (N_2837,N_1128,N_1190);
nand U2838 (N_2838,N_961,N_1116);
and U2839 (N_2839,N_1144,N_794);
xnor U2840 (N_2840,N_263,N_1591);
or U2841 (N_2841,N_17,N_183);
xnor U2842 (N_2842,N_297,N_585);
and U2843 (N_2843,N_1876,N_1007);
or U2844 (N_2844,N_687,N_154);
and U2845 (N_2845,N_902,N_869);
nor U2846 (N_2846,N_1250,N_435);
xor U2847 (N_2847,N_1798,N_92);
nor U2848 (N_2848,N_276,N_824);
or U2849 (N_2849,N_663,N_8);
or U2850 (N_2850,N_1364,N_1227);
nand U2851 (N_2851,N_1859,N_567);
nand U2852 (N_2852,N_1154,N_1230);
and U2853 (N_2853,N_1978,N_394);
or U2854 (N_2854,N_182,N_1397);
or U2855 (N_2855,N_1790,N_221);
nor U2856 (N_2856,N_1381,N_551);
or U2857 (N_2857,N_1006,N_1724);
xor U2858 (N_2858,N_1891,N_613);
or U2859 (N_2859,N_252,N_1551);
or U2860 (N_2860,N_1454,N_25);
or U2861 (N_2861,N_883,N_1884);
nor U2862 (N_2862,N_810,N_611);
nor U2863 (N_2863,N_374,N_1892);
or U2864 (N_2864,N_1240,N_542);
or U2865 (N_2865,N_989,N_1847);
and U2866 (N_2866,N_1638,N_1439);
or U2867 (N_2867,N_1999,N_493);
or U2868 (N_2868,N_776,N_412);
xor U2869 (N_2869,N_1659,N_145);
nor U2870 (N_2870,N_1976,N_431);
and U2871 (N_2871,N_827,N_1199);
or U2872 (N_2872,N_753,N_447);
xor U2873 (N_2873,N_911,N_389);
nor U2874 (N_2874,N_1330,N_785);
and U2875 (N_2875,N_520,N_1452);
and U2876 (N_2876,N_1793,N_1681);
nand U2877 (N_2877,N_927,N_1749);
nor U2878 (N_2878,N_1814,N_683);
and U2879 (N_2879,N_532,N_1393);
xor U2880 (N_2880,N_1188,N_1964);
and U2881 (N_2881,N_143,N_1716);
nor U2882 (N_2882,N_1069,N_1838);
nand U2883 (N_2883,N_1878,N_1326);
and U2884 (N_2884,N_1642,N_1871);
nor U2885 (N_2885,N_1649,N_293);
and U2886 (N_2886,N_955,N_505);
and U2887 (N_2887,N_1952,N_118);
or U2888 (N_2888,N_127,N_1979);
nand U2889 (N_2889,N_830,N_1129);
nor U2890 (N_2890,N_1458,N_212);
or U2891 (N_2891,N_116,N_225);
and U2892 (N_2892,N_364,N_199);
xnor U2893 (N_2893,N_120,N_115);
or U2894 (N_2894,N_842,N_1651);
and U2895 (N_2895,N_250,N_1164);
or U2896 (N_2896,N_1392,N_300);
and U2897 (N_2897,N_1375,N_1325);
nand U2898 (N_2898,N_685,N_1327);
nand U2899 (N_2899,N_1448,N_1441);
or U2900 (N_2900,N_1170,N_1119);
nor U2901 (N_2901,N_1710,N_1612);
xor U2902 (N_2902,N_1080,N_866);
and U2903 (N_2903,N_457,N_1279);
nor U2904 (N_2904,N_1739,N_513);
and U2905 (N_2905,N_761,N_357);
xor U2906 (N_2906,N_332,N_1762);
nor U2907 (N_2907,N_1611,N_217);
or U2908 (N_2908,N_1694,N_1346);
xor U2909 (N_2909,N_1362,N_51);
nand U2910 (N_2910,N_15,N_411);
and U2911 (N_2911,N_358,N_324);
or U2912 (N_2912,N_650,N_1168);
nand U2913 (N_2913,N_280,N_1391);
xor U2914 (N_2914,N_425,N_629);
and U2915 (N_2915,N_841,N_565);
and U2916 (N_2916,N_495,N_1552);
nand U2917 (N_2917,N_1477,N_67);
xor U2918 (N_2918,N_393,N_920);
xnor U2919 (N_2919,N_1885,N_1808);
nand U2920 (N_2920,N_1040,N_967);
nor U2921 (N_2921,N_1784,N_244);
or U2922 (N_2922,N_1804,N_1701);
and U2923 (N_2923,N_723,N_780);
nand U2924 (N_2924,N_884,N_139);
nor U2925 (N_2925,N_933,N_428);
xor U2926 (N_2926,N_843,N_1647);
and U2927 (N_2927,N_1095,N_504);
nor U2928 (N_2928,N_146,N_93);
nand U2929 (N_2929,N_1318,N_820);
or U2930 (N_2930,N_1768,N_464);
and U2931 (N_2931,N_536,N_61);
nor U2932 (N_2932,N_1459,N_1358);
nor U2933 (N_2933,N_750,N_1939);
and U2934 (N_2934,N_994,N_1994);
or U2935 (N_2935,N_1987,N_166);
nand U2936 (N_2936,N_1783,N_1582);
and U2937 (N_2937,N_840,N_1819);
nor U2938 (N_2938,N_251,N_781);
nor U2939 (N_2939,N_1110,N_397);
or U2940 (N_2940,N_661,N_646);
nand U2941 (N_2941,N_615,N_1829);
or U2942 (N_2942,N_335,N_1175);
and U2943 (N_2943,N_1248,N_1373);
and U2944 (N_2944,N_1757,N_914);
nand U2945 (N_2945,N_478,N_1153);
nor U2946 (N_2946,N_54,N_426);
xor U2947 (N_2947,N_1470,N_589);
xnor U2948 (N_2948,N_1292,N_1609);
nor U2949 (N_2949,N_1946,N_1646);
or U2950 (N_2950,N_279,N_575);
nand U2951 (N_2951,N_1750,N_1209);
and U2952 (N_2952,N_991,N_1112);
and U2953 (N_2953,N_514,N_1966);
nand U2954 (N_2954,N_1897,N_1857);
and U2955 (N_2955,N_1030,N_1445);
and U2956 (N_2956,N_347,N_1148);
nor U2957 (N_2957,N_1686,N_1174);
or U2958 (N_2958,N_1698,N_1357);
nor U2959 (N_2959,N_1374,N_1773);
xnor U2960 (N_2960,N_592,N_1861);
and U2961 (N_2961,N_281,N_286);
and U2962 (N_2962,N_71,N_818);
nor U2963 (N_2963,N_1786,N_1157);
xnor U2964 (N_2964,N_931,N_1158);
xnor U2965 (N_2965,N_1911,N_1682);
nand U2966 (N_2966,N_570,N_40);
or U2967 (N_2967,N_577,N_941);
nor U2968 (N_2968,N_594,N_531);
nor U2969 (N_2969,N_1906,N_655);
or U2970 (N_2970,N_767,N_1239);
or U2971 (N_2971,N_52,N_1453);
nand U2972 (N_2972,N_469,N_1055);
nor U2973 (N_2973,N_235,N_614);
and U2974 (N_2974,N_1436,N_1890);
or U2975 (N_2975,N_1573,N_1823);
nor U2976 (N_2976,N_84,N_1960);
xor U2977 (N_2977,N_1717,N_246);
nor U2978 (N_2978,N_82,N_168);
nor U2979 (N_2979,N_732,N_327);
nand U2980 (N_2980,N_1855,N_1131);
and U2981 (N_2981,N_99,N_1086);
or U2982 (N_2982,N_734,N_1945);
nor U2983 (N_2983,N_756,N_789);
nor U2984 (N_2984,N_966,N_1645);
xor U2985 (N_2985,N_1574,N_805);
nand U2986 (N_2986,N_1713,N_604);
xnor U2987 (N_2987,N_1033,N_1135);
nor U2988 (N_2988,N_180,N_9);
and U2989 (N_2989,N_1672,N_845);
nor U2990 (N_2990,N_814,N_1433);
or U2991 (N_2991,N_1626,N_1697);
xnor U2992 (N_2992,N_1824,N_632);
nor U2993 (N_2993,N_319,N_1494);
nand U2994 (N_2994,N_1882,N_617);
and U2995 (N_2995,N_169,N_1825);
or U2996 (N_2996,N_230,N_799);
nand U2997 (N_2997,N_1660,N_610);
or U2998 (N_2998,N_1893,N_1687);
xnor U2999 (N_2999,N_125,N_1145);
nor U3000 (N_3000,N_391,N_859);
xnor U3001 (N_3001,N_1727,N_639);
or U3002 (N_3002,N_1954,N_470);
or U3003 (N_3003,N_865,N_1817);
nand U3004 (N_3004,N_1768,N_1539);
nor U3005 (N_3005,N_1033,N_1952);
or U3006 (N_3006,N_348,N_268);
nor U3007 (N_3007,N_895,N_1906);
xor U3008 (N_3008,N_1343,N_1223);
nand U3009 (N_3009,N_1014,N_1214);
or U3010 (N_3010,N_1030,N_209);
xor U3011 (N_3011,N_1553,N_531);
xnor U3012 (N_3012,N_1391,N_1506);
and U3013 (N_3013,N_1685,N_1339);
nand U3014 (N_3014,N_818,N_291);
nand U3015 (N_3015,N_620,N_1082);
and U3016 (N_3016,N_1226,N_591);
nand U3017 (N_3017,N_865,N_1081);
nor U3018 (N_3018,N_1224,N_1029);
xor U3019 (N_3019,N_1441,N_1226);
xor U3020 (N_3020,N_773,N_1427);
xor U3021 (N_3021,N_169,N_601);
nand U3022 (N_3022,N_1515,N_1616);
xor U3023 (N_3023,N_1380,N_671);
and U3024 (N_3024,N_1700,N_566);
nand U3025 (N_3025,N_1636,N_1536);
or U3026 (N_3026,N_1106,N_944);
or U3027 (N_3027,N_370,N_651);
nor U3028 (N_3028,N_1375,N_1532);
nor U3029 (N_3029,N_812,N_1159);
nand U3030 (N_3030,N_621,N_1892);
xor U3031 (N_3031,N_998,N_373);
xnor U3032 (N_3032,N_558,N_1322);
nand U3033 (N_3033,N_1371,N_659);
nand U3034 (N_3034,N_1816,N_1202);
nand U3035 (N_3035,N_1577,N_1836);
nand U3036 (N_3036,N_1580,N_134);
nor U3037 (N_3037,N_1565,N_735);
xor U3038 (N_3038,N_1545,N_1605);
nor U3039 (N_3039,N_1431,N_512);
or U3040 (N_3040,N_332,N_1405);
xor U3041 (N_3041,N_1285,N_376);
nor U3042 (N_3042,N_1092,N_1078);
nand U3043 (N_3043,N_1099,N_23);
and U3044 (N_3044,N_331,N_380);
nor U3045 (N_3045,N_1519,N_1834);
nand U3046 (N_3046,N_1131,N_1301);
nor U3047 (N_3047,N_973,N_1093);
nor U3048 (N_3048,N_11,N_1627);
or U3049 (N_3049,N_561,N_568);
nor U3050 (N_3050,N_1240,N_1506);
or U3051 (N_3051,N_1544,N_1165);
nor U3052 (N_3052,N_1207,N_1123);
or U3053 (N_3053,N_1959,N_76);
xor U3054 (N_3054,N_764,N_1548);
nand U3055 (N_3055,N_579,N_1890);
nand U3056 (N_3056,N_1451,N_1249);
or U3057 (N_3057,N_726,N_1323);
nand U3058 (N_3058,N_200,N_1069);
and U3059 (N_3059,N_1167,N_365);
nand U3060 (N_3060,N_620,N_1533);
nand U3061 (N_3061,N_367,N_204);
nor U3062 (N_3062,N_658,N_1293);
nor U3063 (N_3063,N_823,N_1059);
or U3064 (N_3064,N_148,N_79);
nand U3065 (N_3065,N_1784,N_1390);
and U3066 (N_3066,N_128,N_238);
or U3067 (N_3067,N_272,N_1074);
and U3068 (N_3068,N_360,N_409);
nor U3069 (N_3069,N_3,N_1656);
or U3070 (N_3070,N_224,N_455);
nor U3071 (N_3071,N_31,N_1449);
nor U3072 (N_3072,N_1938,N_187);
nand U3073 (N_3073,N_1829,N_608);
nand U3074 (N_3074,N_740,N_1310);
xor U3075 (N_3075,N_1514,N_655);
nor U3076 (N_3076,N_703,N_593);
nand U3077 (N_3077,N_1824,N_1994);
xnor U3078 (N_3078,N_200,N_1903);
nand U3079 (N_3079,N_1646,N_343);
and U3080 (N_3080,N_109,N_1565);
nand U3081 (N_3081,N_828,N_1917);
and U3082 (N_3082,N_976,N_1652);
nand U3083 (N_3083,N_377,N_1257);
and U3084 (N_3084,N_1693,N_1592);
xor U3085 (N_3085,N_233,N_596);
nor U3086 (N_3086,N_991,N_1038);
nor U3087 (N_3087,N_586,N_472);
nand U3088 (N_3088,N_1601,N_1151);
xnor U3089 (N_3089,N_1395,N_1785);
nand U3090 (N_3090,N_917,N_650);
nand U3091 (N_3091,N_1164,N_158);
nor U3092 (N_3092,N_1506,N_1501);
xnor U3093 (N_3093,N_940,N_1850);
nand U3094 (N_3094,N_938,N_1475);
nor U3095 (N_3095,N_460,N_41);
and U3096 (N_3096,N_1224,N_513);
and U3097 (N_3097,N_1312,N_1035);
or U3098 (N_3098,N_1230,N_1066);
nor U3099 (N_3099,N_615,N_1387);
or U3100 (N_3100,N_1622,N_921);
or U3101 (N_3101,N_1838,N_1462);
or U3102 (N_3102,N_127,N_1303);
and U3103 (N_3103,N_1927,N_1040);
and U3104 (N_3104,N_1796,N_1786);
or U3105 (N_3105,N_1400,N_793);
nor U3106 (N_3106,N_1834,N_1529);
nand U3107 (N_3107,N_405,N_274);
xnor U3108 (N_3108,N_379,N_750);
xor U3109 (N_3109,N_1561,N_731);
and U3110 (N_3110,N_1800,N_133);
nand U3111 (N_3111,N_273,N_569);
nor U3112 (N_3112,N_491,N_633);
or U3113 (N_3113,N_167,N_1404);
xor U3114 (N_3114,N_1222,N_769);
xor U3115 (N_3115,N_18,N_576);
and U3116 (N_3116,N_482,N_1036);
or U3117 (N_3117,N_865,N_1902);
nor U3118 (N_3118,N_1877,N_313);
or U3119 (N_3119,N_1590,N_437);
nand U3120 (N_3120,N_10,N_1968);
and U3121 (N_3121,N_769,N_1618);
xor U3122 (N_3122,N_711,N_1284);
and U3123 (N_3123,N_55,N_969);
or U3124 (N_3124,N_393,N_1311);
or U3125 (N_3125,N_1979,N_836);
nand U3126 (N_3126,N_1540,N_334);
nor U3127 (N_3127,N_1314,N_134);
xor U3128 (N_3128,N_148,N_1474);
nor U3129 (N_3129,N_841,N_1946);
or U3130 (N_3130,N_362,N_30);
xnor U3131 (N_3131,N_1568,N_1421);
xor U3132 (N_3132,N_1527,N_466);
and U3133 (N_3133,N_1847,N_1283);
nand U3134 (N_3134,N_59,N_249);
and U3135 (N_3135,N_1023,N_1551);
xnor U3136 (N_3136,N_1792,N_845);
and U3137 (N_3137,N_363,N_1467);
or U3138 (N_3138,N_371,N_1538);
nor U3139 (N_3139,N_1599,N_1068);
and U3140 (N_3140,N_630,N_737);
xor U3141 (N_3141,N_1712,N_1427);
and U3142 (N_3142,N_1026,N_1147);
xor U3143 (N_3143,N_861,N_614);
nor U3144 (N_3144,N_723,N_1529);
xnor U3145 (N_3145,N_1413,N_288);
or U3146 (N_3146,N_426,N_1673);
xor U3147 (N_3147,N_1671,N_999);
nor U3148 (N_3148,N_238,N_1178);
and U3149 (N_3149,N_284,N_1473);
nand U3150 (N_3150,N_1869,N_929);
nor U3151 (N_3151,N_88,N_564);
or U3152 (N_3152,N_176,N_1929);
nand U3153 (N_3153,N_1745,N_1967);
or U3154 (N_3154,N_524,N_1422);
nor U3155 (N_3155,N_1856,N_1702);
nand U3156 (N_3156,N_645,N_128);
and U3157 (N_3157,N_698,N_1180);
nand U3158 (N_3158,N_959,N_72);
or U3159 (N_3159,N_1043,N_711);
xnor U3160 (N_3160,N_1265,N_1601);
xnor U3161 (N_3161,N_1790,N_644);
and U3162 (N_3162,N_1667,N_317);
nor U3163 (N_3163,N_537,N_569);
nand U3164 (N_3164,N_1746,N_232);
nor U3165 (N_3165,N_1730,N_1685);
nor U3166 (N_3166,N_1819,N_558);
and U3167 (N_3167,N_553,N_1250);
or U3168 (N_3168,N_1486,N_1210);
and U3169 (N_3169,N_599,N_511);
and U3170 (N_3170,N_1582,N_1194);
xnor U3171 (N_3171,N_1018,N_954);
nand U3172 (N_3172,N_1695,N_1981);
xor U3173 (N_3173,N_1982,N_1745);
xnor U3174 (N_3174,N_260,N_1411);
or U3175 (N_3175,N_1912,N_1377);
nand U3176 (N_3176,N_174,N_1494);
nor U3177 (N_3177,N_1796,N_1691);
and U3178 (N_3178,N_1654,N_1919);
nor U3179 (N_3179,N_669,N_1003);
nor U3180 (N_3180,N_1821,N_296);
or U3181 (N_3181,N_86,N_99);
or U3182 (N_3182,N_1982,N_1886);
and U3183 (N_3183,N_1524,N_1067);
xor U3184 (N_3184,N_468,N_502);
nor U3185 (N_3185,N_1357,N_1489);
nor U3186 (N_3186,N_1476,N_1677);
xor U3187 (N_3187,N_390,N_1146);
and U3188 (N_3188,N_1781,N_1503);
or U3189 (N_3189,N_1201,N_1996);
and U3190 (N_3190,N_584,N_871);
nand U3191 (N_3191,N_147,N_1139);
or U3192 (N_3192,N_1118,N_838);
xnor U3193 (N_3193,N_1006,N_1398);
and U3194 (N_3194,N_1797,N_1980);
xnor U3195 (N_3195,N_1985,N_956);
or U3196 (N_3196,N_765,N_1271);
xor U3197 (N_3197,N_1849,N_1887);
nand U3198 (N_3198,N_970,N_128);
nor U3199 (N_3199,N_742,N_716);
nand U3200 (N_3200,N_1921,N_1718);
and U3201 (N_3201,N_1809,N_949);
and U3202 (N_3202,N_1973,N_161);
xnor U3203 (N_3203,N_1114,N_1989);
or U3204 (N_3204,N_809,N_1212);
xnor U3205 (N_3205,N_1386,N_359);
and U3206 (N_3206,N_1520,N_1333);
and U3207 (N_3207,N_935,N_1892);
or U3208 (N_3208,N_1074,N_1771);
xor U3209 (N_3209,N_1978,N_820);
and U3210 (N_3210,N_962,N_1816);
nand U3211 (N_3211,N_1218,N_177);
and U3212 (N_3212,N_1454,N_620);
and U3213 (N_3213,N_1444,N_602);
and U3214 (N_3214,N_1845,N_1142);
or U3215 (N_3215,N_42,N_176);
nor U3216 (N_3216,N_1039,N_765);
nor U3217 (N_3217,N_227,N_1046);
or U3218 (N_3218,N_715,N_1012);
xor U3219 (N_3219,N_771,N_1828);
and U3220 (N_3220,N_1402,N_166);
and U3221 (N_3221,N_949,N_415);
xor U3222 (N_3222,N_1401,N_1048);
xor U3223 (N_3223,N_242,N_1765);
nand U3224 (N_3224,N_712,N_1290);
and U3225 (N_3225,N_323,N_1138);
xor U3226 (N_3226,N_1914,N_51);
nand U3227 (N_3227,N_1542,N_1777);
nand U3228 (N_3228,N_469,N_191);
nor U3229 (N_3229,N_1364,N_14);
xnor U3230 (N_3230,N_463,N_1106);
xnor U3231 (N_3231,N_1407,N_1090);
and U3232 (N_3232,N_338,N_684);
and U3233 (N_3233,N_1240,N_1662);
or U3234 (N_3234,N_837,N_609);
and U3235 (N_3235,N_653,N_169);
nor U3236 (N_3236,N_1644,N_1943);
nor U3237 (N_3237,N_762,N_117);
nand U3238 (N_3238,N_1210,N_801);
and U3239 (N_3239,N_1338,N_1082);
or U3240 (N_3240,N_1709,N_497);
and U3241 (N_3241,N_578,N_130);
and U3242 (N_3242,N_749,N_624);
nand U3243 (N_3243,N_678,N_1742);
nand U3244 (N_3244,N_1932,N_1907);
nand U3245 (N_3245,N_357,N_1963);
nand U3246 (N_3246,N_63,N_896);
and U3247 (N_3247,N_1137,N_335);
nor U3248 (N_3248,N_1128,N_1044);
and U3249 (N_3249,N_1666,N_1111);
nor U3250 (N_3250,N_135,N_1180);
and U3251 (N_3251,N_165,N_1539);
nor U3252 (N_3252,N_1788,N_1049);
nand U3253 (N_3253,N_1048,N_1434);
or U3254 (N_3254,N_1376,N_1893);
and U3255 (N_3255,N_1935,N_1409);
and U3256 (N_3256,N_1620,N_1846);
nand U3257 (N_3257,N_1421,N_1442);
nand U3258 (N_3258,N_961,N_1811);
nor U3259 (N_3259,N_1831,N_1707);
nor U3260 (N_3260,N_850,N_576);
nor U3261 (N_3261,N_201,N_1758);
nand U3262 (N_3262,N_1183,N_254);
nor U3263 (N_3263,N_300,N_1685);
and U3264 (N_3264,N_990,N_683);
or U3265 (N_3265,N_1426,N_87);
xnor U3266 (N_3266,N_1209,N_1700);
xor U3267 (N_3267,N_389,N_1378);
or U3268 (N_3268,N_1242,N_540);
nand U3269 (N_3269,N_1236,N_640);
nand U3270 (N_3270,N_646,N_1705);
and U3271 (N_3271,N_1662,N_38);
xnor U3272 (N_3272,N_1664,N_1688);
and U3273 (N_3273,N_1313,N_1252);
nand U3274 (N_3274,N_1137,N_939);
nor U3275 (N_3275,N_1746,N_1382);
xnor U3276 (N_3276,N_881,N_1581);
or U3277 (N_3277,N_1726,N_1198);
or U3278 (N_3278,N_71,N_285);
nor U3279 (N_3279,N_1786,N_1695);
xnor U3280 (N_3280,N_394,N_823);
or U3281 (N_3281,N_275,N_1029);
xnor U3282 (N_3282,N_1516,N_1466);
or U3283 (N_3283,N_1877,N_212);
nor U3284 (N_3284,N_1181,N_726);
and U3285 (N_3285,N_54,N_347);
xnor U3286 (N_3286,N_1711,N_1840);
and U3287 (N_3287,N_329,N_1885);
and U3288 (N_3288,N_792,N_115);
or U3289 (N_3289,N_1031,N_1176);
nor U3290 (N_3290,N_1458,N_1648);
nor U3291 (N_3291,N_1044,N_1046);
nor U3292 (N_3292,N_1146,N_794);
nor U3293 (N_3293,N_349,N_625);
nand U3294 (N_3294,N_664,N_1577);
nor U3295 (N_3295,N_552,N_1828);
and U3296 (N_3296,N_233,N_377);
xnor U3297 (N_3297,N_1528,N_778);
and U3298 (N_3298,N_1752,N_118);
and U3299 (N_3299,N_501,N_1164);
or U3300 (N_3300,N_1078,N_665);
and U3301 (N_3301,N_372,N_1827);
nor U3302 (N_3302,N_1043,N_1311);
xor U3303 (N_3303,N_1178,N_1316);
nand U3304 (N_3304,N_1022,N_731);
nor U3305 (N_3305,N_238,N_466);
nand U3306 (N_3306,N_1180,N_1301);
or U3307 (N_3307,N_1248,N_1222);
nor U3308 (N_3308,N_864,N_126);
and U3309 (N_3309,N_1377,N_277);
nor U3310 (N_3310,N_53,N_177);
and U3311 (N_3311,N_1261,N_889);
xor U3312 (N_3312,N_865,N_901);
and U3313 (N_3313,N_276,N_624);
nor U3314 (N_3314,N_1255,N_1924);
xnor U3315 (N_3315,N_239,N_1265);
and U3316 (N_3316,N_1276,N_805);
and U3317 (N_3317,N_1032,N_988);
xor U3318 (N_3318,N_180,N_1312);
nand U3319 (N_3319,N_1890,N_207);
nand U3320 (N_3320,N_228,N_771);
nor U3321 (N_3321,N_408,N_1389);
nand U3322 (N_3322,N_907,N_294);
xnor U3323 (N_3323,N_964,N_1554);
xor U3324 (N_3324,N_1735,N_1048);
xor U3325 (N_3325,N_667,N_1552);
xor U3326 (N_3326,N_1732,N_860);
nor U3327 (N_3327,N_1752,N_644);
or U3328 (N_3328,N_882,N_552);
or U3329 (N_3329,N_1069,N_1825);
or U3330 (N_3330,N_863,N_1954);
and U3331 (N_3331,N_1438,N_263);
nor U3332 (N_3332,N_749,N_20);
or U3333 (N_3333,N_916,N_1268);
and U3334 (N_3334,N_997,N_1652);
xnor U3335 (N_3335,N_1087,N_483);
nand U3336 (N_3336,N_131,N_931);
and U3337 (N_3337,N_414,N_522);
or U3338 (N_3338,N_626,N_577);
and U3339 (N_3339,N_1489,N_779);
nand U3340 (N_3340,N_1307,N_1965);
and U3341 (N_3341,N_1055,N_1155);
or U3342 (N_3342,N_978,N_1402);
or U3343 (N_3343,N_909,N_1638);
xor U3344 (N_3344,N_931,N_130);
and U3345 (N_3345,N_1477,N_1932);
and U3346 (N_3346,N_381,N_699);
xnor U3347 (N_3347,N_256,N_1806);
nand U3348 (N_3348,N_1862,N_1329);
or U3349 (N_3349,N_1415,N_1409);
or U3350 (N_3350,N_505,N_1735);
or U3351 (N_3351,N_1759,N_1803);
xor U3352 (N_3352,N_1783,N_1549);
nand U3353 (N_3353,N_585,N_1458);
xor U3354 (N_3354,N_1347,N_385);
or U3355 (N_3355,N_546,N_1608);
nor U3356 (N_3356,N_1145,N_700);
and U3357 (N_3357,N_1131,N_1223);
nor U3358 (N_3358,N_1585,N_468);
nand U3359 (N_3359,N_1113,N_1627);
nand U3360 (N_3360,N_1177,N_1460);
xor U3361 (N_3361,N_1421,N_1369);
and U3362 (N_3362,N_1402,N_615);
and U3363 (N_3363,N_190,N_1190);
xor U3364 (N_3364,N_1101,N_1596);
nor U3365 (N_3365,N_929,N_1906);
nor U3366 (N_3366,N_1467,N_962);
nor U3367 (N_3367,N_1428,N_389);
xor U3368 (N_3368,N_589,N_1193);
nor U3369 (N_3369,N_1495,N_1018);
xor U3370 (N_3370,N_155,N_663);
and U3371 (N_3371,N_1499,N_1122);
nor U3372 (N_3372,N_1993,N_963);
nor U3373 (N_3373,N_1367,N_979);
nor U3374 (N_3374,N_1516,N_127);
nand U3375 (N_3375,N_693,N_1551);
or U3376 (N_3376,N_992,N_1887);
nor U3377 (N_3377,N_1219,N_1421);
xnor U3378 (N_3378,N_895,N_345);
or U3379 (N_3379,N_675,N_1667);
nand U3380 (N_3380,N_1475,N_1894);
or U3381 (N_3381,N_1292,N_1513);
nand U3382 (N_3382,N_1115,N_255);
xnor U3383 (N_3383,N_339,N_1120);
and U3384 (N_3384,N_393,N_813);
nand U3385 (N_3385,N_1975,N_1241);
and U3386 (N_3386,N_323,N_10);
nand U3387 (N_3387,N_1823,N_1458);
nor U3388 (N_3388,N_1762,N_1359);
nor U3389 (N_3389,N_301,N_460);
xor U3390 (N_3390,N_1625,N_790);
nand U3391 (N_3391,N_91,N_1196);
nor U3392 (N_3392,N_1121,N_1225);
nand U3393 (N_3393,N_1333,N_511);
nor U3394 (N_3394,N_282,N_45);
and U3395 (N_3395,N_1966,N_990);
xor U3396 (N_3396,N_1318,N_1693);
xor U3397 (N_3397,N_1624,N_1113);
xor U3398 (N_3398,N_684,N_1266);
nor U3399 (N_3399,N_1107,N_673);
and U3400 (N_3400,N_1,N_593);
or U3401 (N_3401,N_928,N_1579);
and U3402 (N_3402,N_1335,N_1647);
nand U3403 (N_3403,N_511,N_1729);
nand U3404 (N_3404,N_890,N_1293);
and U3405 (N_3405,N_1135,N_243);
nand U3406 (N_3406,N_1845,N_846);
nand U3407 (N_3407,N_210,N_1854);
xnor U3408 (N_3408,N_608,N_555);
xnor U3409 (N_3409,N_1561,N_1802);
nand U3410 (N_3410,N_1824,N_836);
and U3411 (N_3411,N_1357,N_1146);
nand U3412 (N_3412,N_745,N_533);
and U3413 (N_3413,N_1871,N_1724);
and U3414 (N_3414,N_185,N_1944);
nand U3415 (N_3415,N_863,N_256);
nand U3416 (N_3416,N_1191,N_1030);
nor U3417 (N_3417,N_504,N_55);
nand U3418 (N_3418,N_1593,N_1342);
nor U3419 (N_3419,N_1350,N_198);
and U3420 (N_3420,N_868,N_235);
or U3421 (N_3421,N_1208,N_554);
nor U3422 (N_3422,N_223,N_701);
nand U3423 (N_3423,N_1406,N_287);
nor U3424 (N_3424,N_1940,N_225);
or U3425 (N_3425,N_1904,N_1199);
nand U3426 (N_3426,N_1145,N_751);
and U3427 (N_3427,N_1860,N_329);
xor U3428 (N_3428,N_686,N_636);
xor U3429 (N_3429,N_305,N_1653);
xnor U3430 (N_3430,N_1257,N_523);
nor U3431 (N_3431,N_57,N_1456);
nand U3432 (N_3432,N_988,N_684);
xnor U3433 (N_3433,N_827,N_145);
and U3434 (N_3434,N_218,N_963);
nand U3435 (N_3435,N_1620,N_323);
nand U3436 (N_3436,N_1087,N_1748);
xnor U3437 (N_3437,N_1322,N_964);
nor U3438 (N_3438,N_869,N_443);
or U3439 (N_3439,N_1933,N_1164);
nor U3440 (N_3440,N_1019,N_1728);
and U3441 (N_3441,N_1085,N_416);
xor U3442 (N_3442,N_1719,N_1851);
nand U3443 (N_3443,N_1202,N_674);
xnor U3444 (N_3444,N_1537,N_1762);
and U3445 (N_3445,N_1897,N_696);
and U3446 (N_3446,N_682,N_698);
or U3447 (N_3447,N_577,N_853);
nor U3448 (N_3448,N_167,N_1973);
nand U3449 (N_3449,N_1271,N_1926);
xnor U3450 (N_3450,N_1480,N_308);
and U3451 (N_3451,N_829,N_887);
or U3452 (N_3452,N_1177,N_1984);
or U3453 (N_3453,N_229,N_293);
or U3454 (N_3454,N_713,N_231);
xor U3455 (N_3455,N_1849,N_1596);
xnor U3456 (N_3456,N_13,N_1115);
nand U3457 (N_3457,N_913,N_189);
xnor U3458 (N_3458,N_787,N_1741);
or U3459 (N_3459,N_1304,N_837);
and U3460 (N_3460,N_387,N_34);
xnor U3461 (N_3461,N_1129,N_917);
or U3462 (N_3462,N_667,N_375);
xnor U3463 (N_3463,N_430,N_384);
nor U3464 (N_3464,N_717,N_1284);
xor U3465 (N_3465,N_1825,N_768);
or U3466 (N_3466,N_1364,N_759);
xor U3467 (N_3467,N_1116,N_1712);
and U3468 (N_3468,N_1634,N_828);
nand U3469 (N_3469,N_1785,N_843);
and U3470 (N_3470,N_248,N_1970);
and U3471 (N_3471,N_1230,N_1745);
and U3472 (N_3472,N_1989,N_1442);
nor U3473 (N_3473,N_1898,N_981);
or U3474 (N_3474,N_1377,N_1094);
nor U3475 (N_3475,N_1956,N_1918);
or U3476 (N_3476,N_1097,N_596);
and U3477 (N_3477,N_641,N_1717);
xnor U3478 (N_3478,N_192,N_1461);
and U3479 (N_3479,N_1129,N_1821);
nor U3480 (N_3480,N_248,N_743);
or U3481 (N_3481,N_1809,N_310);
or U3482 (N_3482,N_794,N_110);
nor U3483 (N_3483,N_361,N_690);
nand U3484 (N_3484,N_1607,N_1888);
nand U3485 (N_3485,N_1974,N_636);
or U3486 (N_3486,N_809,N_446);
and U3487 (N_3487,N_787,N_336);
nand U3488 (N_3488,N_393,N_1837);
or U3489 (N_3489,N_869,N_233);
xnor U3490 (N_3490,N_163,N_1716);
nand U3491 (N_3491,N_1922,N_1465);
or U3492 (N_3492,N_79,N_835);
or U3493 (N_3493,N_1997,N_1280);
nand U3494 (N_3494,N_1665,N_648);
nor U3495 (N_3495,N_1238,N_377);
nor U3496 (N_3496,N_310,N_274);
xor U3497 (N_3497,N_1279,N_673);
and U3498 (N_3498,N_1559,N_1457);
nand U3499 (N_3499,N_1731,N_839);
nand U3500 (N_3500,N_1108,N_1644);
xor U3501 (N_3501,N_554,N_920);
nor U3502 (N_3502,N_1792,N_1797);
nand U3503 (N_3503,N_1070,N_1756);
nand U3504 (N_3504,N_1900,N_1654);
and U3505 (N_3505,N_219,N_451);
nor U3506 (N_3506,N_66,N_960);
and U3507 (N_3507,N_1872,N_1193);
nand U3508 (N_3508,N_1837,N_1637);
or U3509 (N_3509,N_1584,N_746);
and U3510 (N_3510,N_1212,N_1589);
nand U3511 (N_3511,N_165,N_1613);
xnor U3512 (N_3512,N_1275,N_883);
or U3513 (N_3513,N_1724,N_595);
xnor U3514 (N_3514,N_1829,N_1503);
and U3515 (N_3515,N_1842,N_716);
or U3516 (N_3516,N_955,N_137);
nand U3517 (N_3517,N_390,N_285);
nand U3518 (N_3518,N_1817,N_21);
xor U3519 (N_3519,N_1528,N_1293);
or U3520 (N_3520,N_610,N_1738);
nand U3521 (N_3521,N_1217,N_1428);
and U3522 (N_3522,N_1367,N_367);
nand U3523 (N_3523,N_1339,N_957);
or U3524 (N_3524,N_1116,N_1122);
and U3525 (N_3525,N_239,N_277);
or U3526 (N_3526,N_244,N_1649);
and U3527 (N_3527,N_1507,N_1089);
and U3528 (N_3528,N_1851,N_1564);
nand U3529 (N_3529,N_738,N_390);
nor U3530 (N_3530,N_279,N_715);
nor U3531 (N_3531,N_985,N_1019);
nor U3532 (N_3532,N_185,N_1352);
nand U3533 (N_3533,N_1010,N_1685);
or U3534 (N_3534,N_621,N_1160);
or U3535 (N_3535,N_871,N_1133);
nand U3536 (N_3536,N_1573,N_718);
nor U3537 (N_3537,N_1856,N_1700);
and U3538 (N_3538,N_193,N_1750);
nor U3539 (N_3539,N_446,N_673);
and U3540 (N_3540,N_390,N_481);
or U3541 (N_3541,N_287,N_1935);
or U3542 (N_3542,N_400,N_1767);
or U3543 (N_3543,N_328,N_75);
nor U3544 (N_3544,N_968,N_348);
nand U3545 (N_3545,N_1374,N_1919);
nor U3546 (N_3546,N_1371,N_1464);
and U3547 (N_3547,N_1621,N_1924);
or U3548 (N_3548,N_1727,N_282);
nor U3549 (N_3549,N_394,N_1194);
nor U3550 (N_3550,N_341,N_1756);
and U3551 (N_3551,N_614,N_456);
or U3552 (N_3552,N_1885,N_777);
and U3553 (N_3553,N_1974,N_1498);
nand U3554 (N_3554,N_778,N_1803);
xnor U3555 (N_3555,N_1778,N_545);
and U3556 (N_3556,N_1163,N_1753);
nand U3557 (N_3557,N_1165,N_1338);
nor U3558 (N_3558,N_62,N_1658);
and U3559 (N_3559,N_1132,N_1522);
nor U3560 (N_3560,N_1007,N_1891);
or U3561 (N_3561,N_956,N_195);
nand U3562 (N_3562,N_1056,N_298);
or U3563 (N_3563,N_1736,N_638);
nor U3564 (N_3564,N_1306,N_1791);
xnor U3565 (N_3565,N_227,N_1356);
xnor U3566 (N_3566,N_1805,N_617);
xnor U3567 (N_3567,N_722,N_975);
and U3568 (N_3568,N_236,N_1683);
or U3569 (N_3569,N_43,N_1231);
xor U3570 (N_3570,N_362,N_47);
or U3571 (N_3571,N_644,N_5);
nand U3572 (N_3572,N_322,N_1814);
nor U3573 (N_3573,N_888,N_905);
nand U3574 (N_3574,N_1110,N_987);
nor U3575 (N_3575,N_191,N_156);
nand U3576 (N_3576,N_187,N_1736);
or U3577 (N_3577,N_1341,N_1801);
nor U3578 (N_3578,N_961,N_1411);
nand U3579 (N_3579,N_1466,N_1728);
nand U3580 (N_3580,N_1351,N_472);
nor U3581 (N_3581,N_200,N_1103);
nor U3582 (N_3582,N_223,N_1890);
and U3583 (N_3583,N_1865,N_1023);
and U3584 (N_3584,N_918,N_795);
xor U3585 (N_3585,N_984,N_718);
or U3586 (N_3586,N_1171,N_1469);
or U3587 (N_3587,N_1024,N_1974);
xnor U3588 (N_3588,N_792,N_699);
xor U3589 (N_3589,N_997,N_1968);
nand U3590 (N_3590,N_1281,N_171);
and U3591 (N_3591,N_1865,N_786);
or U3592 (N_3592,N_1412,N_641);
nand U3593 (N_3593,N_963,N_1628);
nand U3594 (N_3594,N_1350,N_1843);
nand U3595 (N_3595,N_1725,N_1549);
nand U3596 (N_3596,N_1302,N_234);
and U3597 (N_3597,N_774,N_719);
xnor U3598 (N_3598,N_1065,N_1184);
xnor U3599 (N_3599,N_959,N_1770);
or U3600 (N_3600,N_1032,N_1264);
xor U3601 (N_3601,N_1183,N_1269);
nand U3602 (N_3602,N_1661,N_295);
nand U3603 (N_3603,N_661,N_1090);
nor U3604 (N_3604,N_1356,N_1879);
and U3605 (N_3605,N_526,N_1164);
and U3606 (N_3606,N_494,N_990);
nor U3607 (N_3607,N_1155,N_935);
nand U3608 (N_3608,N_283,N_386);
and U3609 (N_3609,N_1064,N_644);
or U3610 (N_3610,N_221,N_1743);
or U3611 (N_3611,N_452,N_529);
nor U3612 (N_3612,N_921,N_181);
nand U3613 (N_3613,N_1814,N_336);
and U3614 (N_3614,N_999,N_427);
or U3615 (N_3615,N_662,N_1803);
xor U3616 (N_3616,N_1153,N_393);
xnor U3617 (N_3617,N_77,N_942);
or U3618 (N_3618,N_923,N_1519);
or U3619 (N_3619,N_853,N_1889);
or U3620 (N_3620,N_1796,N_407);
and U3621 (N_3621,N_460,N_1074);
nor U3622 (N_3622,N_580,N_511);
or U3623 (N_3623,N_1991,N_632);
xnor U3624 (N_3624,N_1217,N_1676);
or U3625 (N_3625,N_1840,N_421);
xor U3626 (N_3626,N_1468,N_1095);
nor U3627 (N_3627,N_1787,N_464);
xor U3628 (N_3628,N_135,N_189);
xnor U3629 (N_3629,N_383,N_1527);
nand U3630 (N_3630,N_356,N_1199);
nand U3631 (N_3631,N_1403,N_1884);
and U3632 (N_3632,N_726,N_1411);
or U3633 (N_3633,N_1958,N_1307);
or U3634 (N_3634,N_139,N_1691);
and U3635 (N_3635,N_1710,N_1731);
and U3636 (N_3636,N_1338,N_432);
or U3637 (N_3637,N_1664,N_1404);
xor U3638 (N_3638,N_1262,N_1383);
nand U3639 (N_3639,N_213,N_167);
or U3640 (N_3640,N_1622,N_265);
and U3641 (N_3641,N_984,N_179);
or U3642 (N_3642,N_1972,N_1289);
and U3643 (N_3643,N_602,N_236);
nand U3644 (N_3644,N_1157,N_1745);
xnor U3645 (N_3645,N_339,N_1339);
and U3646 (N_3646,N_1019,N_1061);
or U3647 (N_3647,N_320,N_1142);
nand U3648 (N_3648,N_1288,N_1960);
nor U3649 (N_3649,N_1818,N_1720);
xor U3650 (N_3650,N_253,N_971);
or U3651 (N_3651,N_1980,N_1596);
and U3652 (N_3652,N_1036,N_923);
or U3653 (N_3653,N_1941,N_965);
and U3654 (N_3654,N_623,N_787);
nor U3655 (N_3655,N_1,N_1334);
and U3656 (N_3656,N_978,N_338);
or U3657 (N_3657,N_969,N_1972);
xnor U3658 (N_3658,N_1637,N_831);
or U3659 (N_3659,N_1592,N_1691);
and U3660 (N_3660,N_780,N_835);
xor U3661 (N_3661,N_363,N_1071);
nand U3662 (N_3662,N_221,N_846);
or U3663 (N_3663,N_37,N_111);
nor U3664 (N_3664,N_1884,N_1432);
nor U3665 (N_3665,N_128,N_1536);
nand U3666 (N_3666,N_1080,N_274);
and U3667 (N_3667,N_1982,N_994);
nand U3668 (N_3668,N_1071,N_835);
and U3669 (N_3669,N_430,N_1209);
nor U3670 (N_3670,N_796,N_472);
and U3671 (N_3671,N_619,N_640);
xnor U3672 (N_3672,N_465,N_611);
or U3673 (N_3673,N_1110,N_405);
nand U3674 (N_3674,N_668,N_1122);
nor U3675 (N_3675,N_1847,N_48);
xnor U3676 (N_3676,N_403,N_1171);
xor U3677 (N_3677,N_1901,N_876);
nor U3678 (N_3678,N_1674,N_1633);
and U3679 (N_3679,N_774,N_938);
nand U3680 (N_3680,N_800,N_1254);
or U3681 (N_3681,N_1227,N_1412);
and U3682 (N_3682,N_618,N_943);
xnor U3683 (N_3683,N_1791,N_495);
or U3684 (N_3684,N_1474,N_527);
or U3685 (N_3685,N_1711,N_711);
xnor U3686 (N_3686,N_283,N_1468);
or U3687 (N_3687,N_809,N_1317);
nand U3688 (N_3688,N_1189,N_309);
and U3689 (N_3689,N_1666,N_1384);
or U3690 (N_3690,N_885,N_1740);
nor U3691 (N_3691,N_1720,N_694);
nand U3692 (N_3692,N_181,N_1940);
and U3693 (N_3693,N_1454,N_1239);
xnor U3694 (N_3694,N_190,N_1767);
and U3695 (N_3695,N_1937,N_1818);
or U3696 (N_3696,N_1064,N_50);
xnor U3697 (N_3697,N_685,N_378);
xnor U3698 (N_3698,N_422,N_1067);
xnor U3699 (N_3699,N_1915,N_164);
xor U3700 (N_3700,N_769,N_1499);
nor U3701 (N_3701,N_1368,N_533);
and U3702 (N_3702,N_885,N_1446);
xnor U3703 (N_3703,N_1542,N_294);
nand U3704 (N_3704,N_1177,N_1379);
xor U3705 (N_3705,N_237,N_1162);
or U3706 (N_3706,N_979,N_1221);
nor U3707 (N_3707,N_1149,N_1483);
xor U3708 (N_3708,N_1458,N_550);
and U3709 (N_3709,N_1509,N_597);
and U3710 (N_3710,N_445,N_1887);
and U3711 (N_3711,N_1808,N_817);
or U3712 (N_3712,N_1630,N_1810);
xnor U3713 (N_3713,N_359,N_498);
and U3714 (N_3714,N_883,N_10);
and U3715 (N_3715,N_400,N_611);
nor U3716 (N_3716,N_1378,N_1816);
nand U3717 (N_3717,N_1164,N_780);
xnor U3718 (N_3718,N_248,N_393);
and U3719 (N_3719,N_518,N_1783);
and U3720 (N_3720,N_1311,N_544);
nand U3721 (N_3721,N_905,N_1523);
nor U3722 (N_3722,N_303,N_4);
xnor U3723 (N_3723,N_1124,N_1781);
nor U3724 (N_3724,N_675,N_1571);
or U3725 (N_3725,N_1049,N_1315);
xor U3726 (N_3726,N_950,N_1002);
and U3727 (N_3727,N_625,N_623);
nor U3728 (N_3728,N_405,N_1221);
xnor U3729 (N_3729,N_1985,N_1943);
nand U3730 (N_3730,N_500,N_1380);
nor U3731 (N_3731,N_311,N_1031);
nand U3732 (N_3732,N_1323,N_459);
or U3733 (N_3733,N_1198,N_680);
nand U3734 (N_3734,N_1326,N_1987);
or U3735 (N_3735,N_624,N_717);
nand U3736 (N_3736,N_1259,N_1369);
and U3737 (N_3737,N_1670,N_337);
nor U3738 (N_3738,N_775,N_478);
nor U3739 (N_3739,N_1516,N_878);
nand U3740 (N_3740,N_1032,N_936);
nor U3741 (N_3741,N_465,N_232);
or U3742 (N_3742,N_804,N_1100);
nor U3743 (N_3743,N_533,N_1798);
xor U3744 (N_3744,N_383,N_387);
or U3745 (N_3745,N_791,N_1070);
nor U3746 (N_3746,N_588,N_94);
and U3747 (N_3747,N_279,N_1483);
nand U3748 (N_3748,N_1763,N_1224);
or U3749 (N_3749,N_1849,N_1769);
nand U3750 (N_3750,N_795,N_617);
or U3751 (N_3751,N_1865,N_390);
or U3752 (N_3752,N_1748,N_1881);
and U3753 (N_3753,N_1543,N_724);
nand U3754 (N_3754,N_720,N_1266);
or U3755 (N_3755,N_1828,N_810);
nor U3756 (N_3756,N_1488,N_981);
nand U3757 (N_3757,N_964,N_172);
or U3758 (N_3758,N_195,N_1042);
nand U3759 (N_3759,N_1685,N_166);
or U3760 (N_3760,N_958,N_868);
and U3761 (N_3761,N_18,N_1831);
xor U3762 (N_3762,N_1189,N_513);
nor U3763 (N_3763,N_1197,N_586);
and U3764 (N_3764,N_1151,N_91);
nor U3765 (N_3765,N_1843,N_845);
or U3766 (N_3766,N_1850,N_700);
nand U3767 (N_3767,N_1868,N_798);
or U3768 (N_3768,N_698,N_61);
nor U3769 (N_3769,N_1928,N_332);
nand U3770 (N_3770,N_360,N_1962);
or U3771 (N_3771,N_493,N_155);
xor U3772 (N_3772,N_361,N_1194);
nand U3773 (N_3773,N_1634,N_1364);
nor U3774 (N_3774,N_1104,N_635);
and U3775 (N_3775,N_1632,N_1692);
nand U3776 (N_3776,N_1694,N_761);
nor U3777 (N_3777,N_756,N_450);
nor U3778 (N_3778,N_738,N_922);
nand U3779 (N_3779,N_1281,N_1956);
nand U3780 (N_3780,N_180,N_1988);
nor U3781 (N_3781,N_1217,N_1264);
xor U3782 (N_3782,N_760,N_87);
nor U3783 (N_3783,N_1798,N_834);
nand U3784 (N_3784,N_827,N_399);
nand U3785 (N_3785,N_1740,N_604);
xor U3786 (N_3786,N_1889,N_1699);
or U3787 (N_3787,N_1888,N_1268);
or U3788 (N_3788,N_270,N_1286);
nand U3789 (N_3789,N_983,N_298);
nor U3790 (N_3790,N_1676,N_1406);
and U3791 (N_3791,N_1864,N_102);
or U3792 (N_3792,N_204,N_1545);
nand U3793 (N_3793,N_791,N_175);
nor U3794 (N_3794,N_1859,N_349);
nand U3795 (N_3795,N_1699,N_933);
nor U3796 (N_3796,N_1671,N_754);
xnor U3797 (N_3797,N_1331,N_360);
nand U3798 (N_3798,N_1958,N_1112);
nand U3799 (N_3799,N_339,N_1444);
nor U3800 (N_3800,N_54,N_1375);
xnor U3801 (N_3801,N_634,N_235);
and U3802 (N_3802,N_1912,N_1014);
nor U3803 (N_3803,N_1028,N_753);
and U3804 (N_3804,N_783,N_685);
or U3805 (N_3805,N_1708,N_873);
or U3806 (N_3806,N_1041,N_1763);
xor U3807 (N_3807,N_1921,N_1165);
nand U3808 (N_3808,N_1767,N_958);
nand U3809 (N_3809,N_551,N_535);
nand U3810 (N_3810,N_1440,N_1024);
and U3811 (N_3811,N_814,N_109);
and U3812 (N_3812,N_1716,N_1834);
xor U3813 (N_3813,N_493,N_868);
nor U3814 (N_3814,N_1300,N_504);
xor U3815 (N_3815,N_1195,N_19);
and U3816 (N_3816,N_303,N_1421);
xnor U3817 (N_3817,N_1381,N_61);
and U3818 (N_3818,N_1719,N_1309);
and U3819 (N_3819,N_1678,N_645);
nor U3820 (N_3820,N_1851,N_1428);
xnor U3821 (N_3821,N_1071,N_1055);
xnor U3822 (N_3822,N_1732,N_673);
nand U3823 (N_3823,N_266,N_598);
nand U3824 (N_3824,N_850,N_200);
and U3825 (N_3825,N_1417,N_1896);
xor U3826 (N_3826,N_1090,N_1202);
xnor U3827 (N_3827,N_509,N_1116);
and U3828 (N_3828,N_1130,N_626);
or U3829 (N_3829,N_677,N_1275);
nand U3830 (N_3830,N_382,N_1594);
xnor U3831 (N_3831,N_1068,N_87);
nor U3832 (N_3832,N_770,N_521);
xnor U3833 (N_3833,N_1844,N_841);
xnor U3834 (N_3834,N_386,N_1119);
nand U3835 (N_3835,N_1887,N_1859);
xnor U3836 (N_3836,N_1327,N_956);
nor U3837 (N_3837,N_176,N_1147);
nor U3838 (N_3838,N_645,N_916);
or U3839 (N_3839,N_1543,N_472);
nand U3840 (N_3840,N_1653,N_1229);
nor U3841 (N_3841,N_1091,N_1083);
or U3842 (N_3842,N_37,N_257);
and U3843 (N_3843,N_512,N_918);
and U3844 (N_3844,N_1097,N_658);
or U3845 (N_3845,N_1819,N_330);
nor U3846 (N_3846,N_1543,N_953);
xor U3847 (N_3847,N_728,N_509);
xor U3848 (N_3848,N_986,N_1469);
and U3849 (N_3849,N_1202,N_1938);
and U3850 (N_3850,N_798,N_1280);
and U3851 (N_3851,N_1053,N_1973);
or U3852 (N_3852,N_930,N_1836);
xnor U3853 (N_3853,N_1709,N_180);
nor U3854 (N_3854,N_358,N_1005);
and U3855 (N_3855,N_9,N_1373);
or U3856 (N_3856,N_1097,N_1210);
xor U3857 (N_3857,N_139,N_1289);
xnor U3858 (N_3858,N_1906,N_969);
xor U3859 (N_3859,N_1271,N_218);
or U3860 (N_3860,N_970,N_59);
xor U3861 (N_3861,N_1013,N_972);
nand U3862 (N_3862,N_1572,N_569);
nand U3863 (N_3863,N_1953,N_1444);
xnor U3864 (N_3864,N_31,N_121);
and U3865 (N_3865,N_979,N_88);
nand U3866 (N_3866,N_494,N_274);
or U3867 (N_3867,N_503,N_612);
nor U3868 (N_3868,N_637,N_74);
nor U3869 (N_3869,N_592,N_1568);
or U3870 (N_3870,N_108,N_1925);
nand U3871 (N_3871,N_1627,N_957);
nand U3872 (N_3872,N_1966,N_350);
nor U3873 (N_3873,N_1865,N_934);
and U3874 (N_3874,N_1730,N_131);
and U3875 (N_3875,N_1891,N_478);
nor U3876 (N_3876,N_1775,N_561);
and U3877 (N_3877,N_17,N_568);
or U3878 (N_3878,N_1983,N_1631);
nand U3879 (N_3879,N_1176,N_978);
xor U3880 (N_3880,N_1837,N_865);
xor U3881 (N_3881,N_1980,N_885);
nand U3882 (N_3882,N_1741,N_1502);
or U3883 (N_3883,N_554,N_239);
or U3884 (N_3884,N_869,N_476);
or U3885 (N_3885,N_1318,N_698);
nand U3886 (N_3886,N_633,N_1995);
xnor U3887 (N_3887,N_452,N_607);
or U3888 (N_3888,N_101,N_603);
nor U3889 (N_3889,N_954,N_970);
and U3890 (N_3890,N_1021,N_1907);
and U3891 (N_3891,N_123,N_220);
or U3892 (N_3892,N_123,N_1973);
or U3893 (N_3893,N_1856,N_387);
or U3894 (N_3894,N_309,N_1622);
nor U3895 (N_3895,N_282,N_940);
or U3896 (N_3896,N_1376,N_1830);
nand U3897 (N_3897,N_1043,N_1559);
xor U3898 (N_3898,N_1707,N_686);
and U3899 (N_3899,N_1664,N_1888);
xor U3900 (N_3900,N_591,N_544);
nor U3901 (N_3901,N_339,N_1055);
and U3902 (N_3902,N_1362,N_106);
or U3903 (N_3903,N_1154,N_413);
or U3904 (N_3904,N_199,N_295);
and U3905 (N_3905,N_1693,N_1507);
or U3906 (N_3906,N_366,N_304);
xnor U3907 (N_3907,N_1037,N_502);
xnor U3908 (N_3908,N_1250,N_813);
nor U3909 (N_3909,N_641,N_727);
or U3910 (N_3910,N_1038,N_1121);
xor U3911 (N_3911,N_1974,N_1796);
and U3912 (N_3912,N_1314,N_306);
nand U3913 (N_3913,N_1898,N_1044);
nand U3914 (N_3914,N_1197,N_1199);
and U3915 (N_3915,N_215,N_804);
nor U3916 (N_3916,N_654,N_398);
nand U3917 (N_3917,N_86,N_1988);
nor U3918 (N_3918,N_202,N_418);
and U3919 (N_3919,N_1859,N_324);
nand U3920 (N_3920,N_1566,N_847);
nor U3921 (N_3921,N_341,N_1056);
xnor U3922 (N_3922,N_1192,N_360);
or U3923 (N_3923,N_923,N_146);
xnor U3924 (N_3924,N_424,N_890);
nand U3925 (N_3925,N_1189,N_625);
and U3926 (N_3926,N_911,N_544);
xor U3927 (N_3927,N_194,N_1268);
nor U3928 (N_3928,N_1530,N_1618);
nor U3929 (N_3929,N_802,N_1323);
nand U3930 (N_3930,N_1547,N_1293);
or U3931 (N_3931,N_176,N_1130);
nor U3932 (N_3932,N_1851,N_1380);
nand U3933 (N_3933,N_1532,N_409);
xnor U3934 (N_3934,N_723,N_144);
nand U3935 (N_3935,N_909,N_1352);
and U3936 (N_3936,N_1064,N_1003);
nand U3937 (N_3937,N_602,N_327);
xor U3938 (N_3938,N_740,N_1361);
and U3939 (N_3939,N_996,N_1568);
and U3940 (N_3940,N_1418,N_508);
or U3941 (N_3941,N_1227,N_1922);
and U3942 (N_3942,N_876,N_1432);
nor U3943 (N_3943,N_1806,N_204);
xnor U3944 (N_3944,N_850,N_1988);
nor U3945 (N_3945,N_803,N_166);
nand U3946 (N_3946,N_261,N_1415);
and U3947 (N_3947,N_1400,N_608);
xnor U3948 (N_3948,N_1591,N_731);
xnor U3949 (N_3949,N_1238,N_996);
and U3950 (N_3950,N_805,N_1525);
or U3951 (N_3951,N_653,N_1226);
xnor U3952 (N_3952,N_1645,N_1463);
nor U3953 (N_3953,N_566,N_1343);
or U3954 (N_3954,N_1164,N_1191);
nand U3955 (N_3955,N_555,N_1415);
xnor U3956 (N_3956,N_546,N_1622);
xor U3957 (N_3957,N_714,N_1750);
and U3958 (N_3958,N_1695,N_312);
xnor U3959 (N_3959,N_820,N_1755);
or U3960 (N_3960,N_389,N_1562);
nand U3961 (N_3961,N_463,N_1965);
nor U3962 (N_3962,N_98,N_540);
or U3963 (N_3963,N_392,N_995);
nand U3964 (N_3964,N_52,N_709);
nand U3965 (N_3965,N_1465,N_573);
and U3966 (N_3966,N_1262,N_794);
or U3967 (N_3967,N_144,N_1608);
nor U3968 (N_3968,N_135,N_1094);
nand U3969 (N_3969,N_1233,N_997);
and U3970 (N_3970,N_1208,N_287);
nand U3971 (N_3971,N_884,N_1858);
nor U3972 (N_3972,N_1536,N_549);
nand U3973 (N_3973,N_698,N_1808);
nor U3974 (N_3974,N_1042,N_1185);
or U3975 (N_3975,N_1031,N_767);
nand U3976 (N_3976,N_1572,N_576);
xor U3977 (N_3977,N_1235,N_263);
nor U3978 (N_3978,N_525,N_1065);
nand U3979 (N_3979,N_1752,N_1673);
or U3980 (N_3980,N_1841,N_422);
xnor U3981 (N_3981,N_206,N_211);
and U3982 (N_3982,N_935,N_1363);
or U3983 (N_3983,N_1771,N_1943);
or U3984 (N_3984,N_906,N_1141);
nor U3985 (N_3985,N_83,N_251);
or U3986 (N_3986,N_765,N_431);
and U3987 (N_3987,N_13,N_741);
xor U3988 (N_3988,N_835,N_1044);
and U3989 (N_3989,N_81,N_155);
or U3990 (N_3990,N_731,N_1606);
nor U3991 (N_3991,N_1524,N_909);
xor U3992 (N_3992,N_71,N_598);
and U3993 (N_3993,N_721,N_288);
xor U3994 (N_3994,N_1072,N_170);
and U3995 (N_3995,N_389,N_1794);
or U3996 (N_3996,N_1736,N_734);
xnor U3997 (N_3997,N_1016,N_690);
nand U3998 (N_3998,N_1903,N_1008);
nand U3999 (N_3999,N_902,N_1012);
or U4000 (N_4000,N_2682,N_3785);
and U4001 (N_4001,N_2753,N_2595);
nor U4002 (N_4002,N_3514,N_2407);
and U4003 (N_4003,N_3116,N_2176);
or U4004 (N_4004,N_3253,N_2388);
and U4005 (N_4005,N_3029,N_2013);
nor U4006 (N_4006,N_2646,N_2174);
xor U4007 (N_4007,N_2270,N_3999);
nor U4008 (N_4008,N_3538,N_3343);
xor U4009 (N_4009,N_2996,N_2980);
nand U4010 (N_4010,N_3789,N_2153);
nor U4011 (N_4011,N_3455,N_3685);
xnor U4012 (N_4012,N_2701,N_2846);
and U4013 (N_4013,N_3496,N_2396);
nor U4014 (N_4014,N_2289,N_2030);
or U4015 (N_4015,N_3268,N_2401);
and U4016 (N_4016,N_3681,N_3009);
nor U4017 (N_4017,N_3095,N_2042);
xnor U4018 (N_4018,N_3290,N_3796);
nand U4019 (N_4019,N_2895,N_3650);
or U4020 (N_4020,N_2878,N_3421);
xnor U4021 (N_4021,N_3655,N_2347);
nand U4022 (N_4022,N_3977,N_3443);
or U4023 (N_4023,N_3083,N_2080);
or U4024 (N_4024,N_3915,N_3028);
or U4025 (N_4025,N_2776,N_2015);
nand U4026 (N_4026,N_3300,N_2377);
nand U4027 (N_4027,N_3480,N_2265);
xor U4028 (N_4028,N_2920,N_3053);
nor U4029 (N_4029,N_2715,N_3407);
nor U4030 (N_4030,N_3213,N_2236);
nand U4031 (N_4031,N_3939,N_3146);
nand U4032 (N_4032,N_2184,N_3833);
nor U4033 (N_4033,N_2827,N_3241);
or U4034 (N_4034,N_2464,N_3805);
nand U4035 (N_4035,N_3822,N_2819);
xnor U4036 (N_4036,N_2198,N_3621);
nor U4037 (N_4037,N_3084,N_3026);
or U4038 (N_4038,N_2951,N_2580);
nand U4039 (N_4039,N_3882,N_3064);
xor U4040 (N_4040,N_2249,N_3248);
and U4041 (N_4041,N_3740,N_3405);
and U4042 (N_4042,N_3784,N_3778);
nand U4043 (N_4043,N_3824,N_2476);
or U4044 (N_4044,N_3288,N_3412);
nand U4045 (N_4045,N_2297,N_2736);
and U4046 (N_4046,N_2750,N_2922);
xnor U4047 (N_4047,N_3942,N_2143);
nand U4048 (N_4048,N_3045,N_2586);
nand U4049 (N_4049,N_3806,N_2752);
and U4050 (N_4050,N_2582,N_3724);
or U4051 (N_4051,N_2982,N_3555);
nand U4052 (N_4052,N_3467,N_2315);
nand U4053 (N_4053,N_3828,N_2933);
nand U4054 (N_4054,N_2572,N_2731);
or U4055 (N_4055,N_3326,N_2062);
or U4056 (N_4056,N_2535,N_2034);
and U4057 (N_4057,N_2303,N_2380);
or U4058 (N_4058,N_2037,N_2500);
or U4059 (N_4059,N_3834,N_2805);
nor U4060 (N_4060,N_2223,N_2378);
and U4061 (N_4061,N_3979,N_3088);
nand U4062 (N_4062,N_2311,N_3917);
or U4063 (N_4063,N_3101,N_2362);
and U4064 (N_4064,N_2240,N_3082);
or U4065 (N_4065,N_2219,N_3861);
nand U4066 (N_4066,N_3250,N_3551);
and U4067 (N_4067,N_2339,N_3245);
xnor U4068 (N_4068,N_2431,N_2438);
or U4069 (N_4069,N_2745,N_3646);
nor U4070 (N_4070,N_3588,N_3328);
nor U4071 (N_4071,N_3475,N_3281);
and U4072 (N_4072,N_3743,N_3878);
xnor U4073 (N_4073,N_3951,N_3956);
or U4074 (N_4074,N_2550,N_3821);
and U4075 (N_4075,N_2772,N_3903);
and U4076 (N_4076,N_3534,N_3441);
or U4077 (N_4077,N_2331,N_3715);
xor U4078 (N_4078,N_2204,N_3227);
or U4079 (N_4079,N_2697,N_3911);
and U4080 (N_4080,N_2931,N_2106);
and U4081 (N_4081,N_3141,N_2721);
or U4082 (N_4082,N_2995,N_2602);
or U4083 (N_4083,N_2127,N_3560);
xnor U4084 (N_4084,N_2093,N_3908);
nor U4085 (N_4085,N_2357,N_2038);
or U4086 (N_4086,N_3312,N_3945);
or U4087 (N_4087,N_3408,N_2248);
xor U4088 (N_4088,N_3868,N_3559);
nor U4089 (N_4089,N_3222,N_3234);
nand U4090 (N_4090,N_3390,N_2139);
and U4091 (N_4091,N_3447,N_2053);
nand U4092 (N_4092,N_3558,N_3949);
or U4093 (N_4093,N_3629,N_3633);
and U4094 (N_4094,N_2092,N_2228);
or U4095 (N_4095,N_3849,N_3684);
and U4096 (N_4096,N_2629,N_2145);
xnor U4097 (N_4097,N_2364,N_2436);
and U4098 (N_4098,N_2205,N_3072);
and U4099 (N_4099,N_3557,N_3089);
xnor U4100 (N_4100,N_3366,N_2040);
nand U4101 (N_4101,N_2829,N_3765);
nand U4102 (N_4102,N_3620,N_3719);
or U4103 (N_4103,N_3679,N_2094);
and U4104 (N_4104,N_2463,N_3004);
and U4105 (N_4105,N_2230,N_3733);
xnor U4106 (N_4106,N_2677,N_3205);
and U4107 (N_4107,N_3960,N_2381);
nand U4108 (N_4108,N_3183,N_2063);
and U4109 (N_4109,N_2314,N_2932);
nor U4110 (N_4110,N_3606,N_3372);
nand U4111 (N_4111,N_2087,N_3823);
nor U4112 (N_4112,N_3401,N_3152);
and U4113 (N_4113,N_3546,N_3973);
nor U4114 (N_4114,N_2972,N_3274);
and U4115 (N_4115,N_2402,N_3788);
nand U4116 (N_4116,N_2163,N_3449);
nand U4117 (N_4117,N_2345,N_2416);
nor U4118 (N_4118,N_3351,N_3065);
nor U4119 (N_4119,N_3611,N_3519);
nor U4120 (N_4120,N_3756,N_2432);
nor U4121 (N_4121,N_2564,N_2141);
and U4122 (N_4122,N_2644,N_3955);
and U4123 (N_4123,N_2823,N_3739);
nor U4124 (N_4124,N_2004,N_3052);
xnor U4125 (N_4125,N_3500,N_3427);
or U4126 (N_4126,N_2298,N_2927);
nor U4127 (N_4127,N_3148,N_3660);
or U4128 (N_4128,N_3110,N_2170);
nand U4129 (N_4129,N_3653,N_3483);
or U4130 (N_4130,N_2243,N_2001);
xor U4131 (N_4131,N_2625,N_2478);
or U4132 (N_4132,N_2511,N_2825);
nand U4133 (N_4133,N_2209,N_3658);
xor U4134 (N_4134,N_2130,N_2090);
and U4135 (N_4135,N_2964,N_3846);
and U4136 (N_4136,N_3835,N_2348);
and U4137 (N_4137,N_2585,N_2164);
nor U4138 (N_4138,N_3884,N_2957);
nand U4139 (N_4139,N_2142,N_3499);
nand U4140 (N_4140,N_3378,N_3905);
nor U4141 (N_4141,N_2253,N_3504);
nand U4142 (N_4142,N_3283,N_3392);
or U4143 (N_4143,N_3628,N_3505);
nand U4144 (N_4144,N_2909,N_3093);
xor U4145 (N_4145,N_2410,N_3215);
nor U4146 (N_4146,N_2672,N_2915);
and U4147 (N_4147,N_2747,N_2645);
or U4148 (N_4148,N_2764,N_2065);
nand U4149 (N_4149,N_2581,N_3194);
nand U4150 (N_4150,N_3022,N_3721);
nand U4151 (N_4151,N_3079,N_3744);
nand U4152 (N_4152,N_2941,N_2537);
nor U4153 (N_4153,N_3356,N_3576);
and U4154 (N_4154,N_2400,N_3921);
or U4155 (N_4155,N_2624,N_2016);
xor U4156 (N_4156,N_2523,N_3174);
xnor U4157 (N_4157,N_2733,N_2481);
and U4158 (N_4158,N_2981,N_2195);
or U4159 (N_4159,N_3510,N_2700);
nand U4160 (N_4160,N_3109,N_3466);
xnor U4161 (N_4161,N_3157,N_2556);
nand U4162 (N_4162,N_3114,N_2128);
nand U4163 (N_4163,N_2725,N_3767);
or U4164 (N_4164,N_3374,N_2443);
or U4165 (N_4165,N_2199,N_3035);
nor U4166 (N_4166,N_3568,N_2201);
nand U4167 (N_4167,N_3073,N_2883);
xor U4168 (N_4168,N_2826,N_2842);
nor U4169 (N_4169,N_2548,N_2849);
nand U4170 (N_4170,N_3542,N_2891);
and U4171 (N_4171,N_3857,N_2071);
xor U4172 (N_4172,N_3471,N_3107);
or U4173 (N_4173,N_3547,N_3468);
or U4174 (N_4174,N_2019,N_3860);
or U4175 (N_4175,N_3544,N_2858);
and U4176 (N_4176,N_2288,N_3316);
and U4177 (N_4177,N_2961,N_2674);
or U4178 (N_4178,N_2226,N_2074);
nand U4179 (N_4179,N_2816,N_3406);
nor U4180 (N_4180,N_2593,N_2947);
nor U4181 (N_4181,N_2992,N_3668);
nand U4182 (N_4182,N_3714,N_3501);
xor U4183 (N_4183,N_3923,N_3815);
nor U4184 (N_4184,N_2975,N_2856);
and U4185 (N_4185,N_2977,N_3612);
or U4186 (N_4186,N_2422,N_2706);
nand U4187 (N_4187,N_3790,N_2763);
and U4188 (N_4188,N_2872,N_2609);
nand U4189 (N_4189,N_2623,N_2335);
nand U4190 (N_4190,N_3780,N_3813);
or U4191 (N_4191,N_3413,N_3961);
xor U4192 (N_4192,N_3040,N_3380);
and U4193 (N_4193,N_3354,N_2177);
and U4194 (N_4194,N_2525,N_2104);
xor U4195 (N_4195,N_3456,N_3948);
and U4196 (N_4196,N_3676,N_3800);
nand U4197 (N_4197,N_2191,N_2620);
nand U4198 (N_4198,N_2867,N_3153);
or U4199 (N_4199,N_3391,N_3595);
nand U4200 (N_4200,N_3994,N_3880);
and U4201 (N_4201,N_3794,N_3386);
nand U4202 (N_4202,N_3062,N_3779);
and U4203 (N_4203,N_2954,N_2549);
or U4204 (N_4204,N_3803,N_3304);
nand U4205 (N_4205,N_2877,N_2108);
and U4206 (N_4206,N_2185,N_2167);
nor U4207 (N_4207,N_2699,N_2638);
xor U4208 (N_4208,N_2007,N_2359);
and U4209 (N_4209,N_3327,N_3970);
and U4210 (N_4210,N_2663,N_2262);
or U4211 (N_4211,N_2570,N_3043);
xor U4212 (N_4212,N_3985,N_2865);
xor U4213 (N_4213,N_2813,N_2719);
nand U4214 (N_4214,N_2383,N_3564);
and U4215 (N_4215,N_2113,N_3705);
and U4216 (N_4216,N_2073,N_2779);
xnor U4217 (N_4217,N_3171,N_2290);
nand U4218 (N_4218,N_3169,N_3424);
and U4219 (N_4219,N_3757,N_3397);
and U4220 (N_4220,N_2091,N_3840);
or U4221 (N_4221,N_2144,N_2134);
nor U4222 (N_4222,N_3862,N_2978);
nor U4223 (N_4223,N_2614,N_2146);
and U4224 (N_4224,N_2450,N_2250);
nor U4225 (N_4225,N_3000,N_2969);
xor U4226 (N_4226,N_2862,N_3047);
or U4227 (N_4227,N_3170,N_2350);
and U4228 (N_4228,N_3554,N_3003);
and U4229 (N_4229,N_2574,N_3596);
nor U4230 (N_4230,N_3229,N_2647);
xnor U4231 (N_4231,N_2387,N_3792);
nor U4232 (N_4232,N_3331,N_3609);
xor U4233 (N_4233,N_3753,N_3195);
nor U4234 (N_4234,N_2659,N_3549);
nor U4235 (N_4235,N_2434,N_2714);
or U4236 (N_4236,N_3420,N_3856);
or U4237 (N_4237,N_3113,N_2773);
nor U4238 (N_4238,N_2605,N_2423);
or U4239 (N_4239,N_3798,N_3820);
and U4240 (N_4240,N_3207,N_2890);
xor U4241 (N_4241,N_2168,N_3232);
nor U4242 (N_4242,N_3462,N_2882);
nand U4243 (N_4243,N_2923,N_2121);
nand U4244 (N_4244,N_2902,N_3048);
xor U4245 (N_4245,N_3147,N_2708);
and U4246 (N_4246,N_3002,N_3938);
nand U4247 (N_4247,N_2002,N_2538);
or U4248 (N_4248,N_3570,N_2384);
nor U4249 (N_4249,N_3126,N_2751);
or U4250 (N_4250,N_3603,N_3652);
nor U4251 (N_4251,N_2366,N_2488);
xor U4252 (N_4252,N_2547,N_2974);
or U4253 (N_4253,N_2894,N_3012);
xnor U4254 (N_4254,N_3452,N_2178);
and U4255 (N_4255,N_2258,N_2006);
nor U4256 (N_4256,N_2081,N_2797);
and U4257 (N_4257,N_2943,N_3690);
and U4258 (N_4258,N_2788,N_2305);
xnor U4259 (N_4259,N_3847,N_2122);
xnor U4260 (N_4260,N_2000,N_2551);
nand U4261 (N_4261,N_3099,N_3112);
or U4262 (N_4262,N_3654,N_3996);
nand U4263 (N_4263,N_3434,N_2782);
nand U4264 (N_4264,N_3341,N_3111);
xor U4265 (N_4265,N_3533,N_3329);
nand U4266 (N_4266,N_2403,N_3541);
or U4267 (N_4267,N_2958,N_2575);
nand U4268 (N_4268,N_2208,N_2010);
xor U4269 (N_4269,N_3158,N_3179);
nand U4270 (N_4270,N_3284,N_3428);
or U4271 (N_4271,N_3272,N_3269);
nand U4272 (N_4272,N_3370,N_2354);
nand U4273 (N_4273,N_2910,N_3843);
and U4274 (N_4274,N_2916,N_3937);
and U4275 (N_4275,N_2193,N_3314);
xor U4276 (N_4276,N_2160,N_3276);
nand U4277 (N_4277,N_2439,N_3663);
nor U4278 (N_4278,N_3931,N_3423);
nand U4279 (N_4279,N_2940,N_3478);
nand U4280 (N_4280,N_3075,N_3177);
nor U4281 (N_4281,N_3991,N_2031);
nor U4282 (N_4282,N_2477,N_3895);
xor U4283 (N_4283,N_3894,N_2847);
nor U4284 (N_4284,N_3348,N_3226);
nor U4285 (N_4285,N_3238,N_2800);
and U4286 (N_4286,N_3486,N_2351);
and U4287 (N_4287,N_2993,N_2541);
nand U4288 (N_4288,N_3918,N_2442);
and U4289 (N_4289,N_3339,N_2987);
and U4290 (N_4290,N_3287,N_2363);
nand U4291 (N_4291,N_2521,N_2202);
xnor U4292 (N_4292,N_2522,N_2504);
xnor U4293 (N_4293,N_2928,N_3747);
nor U4294 (N_4294,N_3574,N_3850);
nor U4295 (N_4295,N_3267,N_3662);
xor U4296 (N_4296,N_2785,N_3103);
or U4297 (N_4297,N_2341,N_2369);
or U4298 (N_4298,N_3254,N_3763);
nand U4299 (N_4299,N_3875,N_3742);
nor U4300 (N_4300,N_2101,N_2792);
nand U4301 (N_4301,N_2798,N_2194);
nand U4302 (N_4302,N_3873,N_2660);
or U4303 (N_4303,N_3271,N_2684);
and U4304 (N_4304,N_3362,N_3758);
or U4305 (N_4305,N_3635,N_3142);
nand U4306 (N_4306,N_2970,N_3930);
nand U4307 (N_4307,N_3617,N_2517);
xnor U4308 (N_4308,N_2405,N_2469);
or U4309 (N_4309,N_3122,N_2412);
and U4310 (N_4310,N_3307,N_2617);
nand U4311 (N_4311,N_3429,N_3968);
and U4312 (N_4312,N_3812,N_3165);
or U4313 (N_4313,N_2367,N_2386);
and U4314 (N_4314,N_2761,N_3829);
nand U4315 (N_4315,N_3333,N_2035);
and U4316 (N_4316,N_3459,N_3573);
nor U4317 (N_4317,N_3769,N_3605);
xnor U4318 (N_4318,N_2028,N_2633);
and U4319 (N_4319,N_2332,N_3602);
nand U4320 (N_4320,N_3978,N_3289);
xnor U4321 (N_4321,N_2310,N_2349);
nand U4322 (N_4322,N_2762,N_2713);
nor U4323 (N_4323,N_2085,N_2003);
and U4324 (N_4324,N_2246,N_2855);
xor U4325 (N_4325,N_3342,N_2132);
xnor U4326 (N_4326,N_3709,N_3776);
and U4327 (N_4327,N_3916,N_3046);
xnor U4328 (N_4328,N_3764,N_3502);
or U4329 (N_4329,N_3993,N_2277);
and U4330 (N_4330,N_3350,N_2151);
xor U4331 (N_4331,N_2634,N_3264);
and U4332 (N_4332,N_2681,N_2485);
nor U4333 (N_4333,N_3184,N_2186);
nand U4334 (N_4334,N_3220,N_3674);
xor U4335 (N_4335,N_3759,N_3360);
xor U4336 (N_4336,N_2861,N_2738);
xnor U4337 (N_4337,N_2118,N_2937);
and U4338 (N_4338,N_3683,N_2579);
nor U4339 (N_4339,N_2414,N_2919);
xor U4340 (N_4340,N_3485,N_2685);
nand U4341 (N_4341,N_2592,N_3006);
xnor U4342 (N_4342,N_3722,N_3393);
nand U4343 (N_4343,N_2115,N_2218);
nand U4344 (N_4344,N_2183,N_3347);
xor U4345 (N_4345,N_3597,N_2691);
nor U4346 (N_4346,N_3031,N_3197);
nand U4347 (N_4347,N_2278,N_3859);
nor U4348 (N_4348,N_2260,N_2415);
or U4349 (N_4349,N_2534,N_2527);
xnor U4350 (N_4350,N_3749,N_3732);
nor U4351 (N_4351,N_3433,N_2190);
nand U4352 (N_4352,N_2172,N_3256);
or U4353 (N_4353,N_2502,N_3200);
nor U4354 (N_4354,N_3149,N_3432);
and U4355 (N_4355,N_2734,N_3582);
or U4356 (N_4356,N_3487,N_2059);
or U4357 (N_4357,N_3367,N_2507);
xor U4358 (N_4358,N_2394,N_3318);
nor U4359 (N_4359,N_2207,N_3217);
and U4360 (N_4360,N_3419,N_2885);
and U4361 (N_4361,N_2705,N_2077);
nor U4362 (N_4362,N_2588,N_3458);
or U4363 (N_4363,N_2508,N_3801);
or U4364 (N_4364,N_2887,N_2320);
nor U4365 (N_4365,N_3521,N_3520);
xnor U4366 (N_4366,N_3581,N_3592);
nand U4367 (N_4367,N_2116,N_2326);
nand U4368 (N_4368,N_3578,N_2889);
or U4369 (N_4369,N_3061,N_3572);
xnor U4370 (N_4370,N_2656,N_3139);
or U4371 (N_4371,N_3212,N_2948);
nor U4372 (N_4372,N_2287,N_3155);
nand U4373 (N_4373,N_3493,N_2465);
xnor U4374 (N_4374,N_3926,N_3020);
xnor U4375 (N_4375,N_2470,N_3667);
nor U4376 (N_4376,N_3730,N_2355);
nor U4377 (N_4377,N_3713,N_3355);
and U4378 (N_4378,N_2675,N_2784);
xor U4379 (N_4379,N_3736,N_3365);
xor U4380 (N_4380,N_3565,N_3914);
xor U4381 (N_4381,N_3252,N_2487);
or U4382 (N_4382,N_3680,N_2642);
xnor U4383 (N_4383,N_3198,N_2991);
nand U4384 (N_4384,N_2033,N_3634);
nand U4385 (N_4385,N_2555,N_3497);
nor U4386 (N_4386,N_2942,N_3242);
or U4387 (N_4387,N_3553,N_3377);
or U4388 (N_4388,N_3422,N_3460);
xnor U4389 (N_4389,N_3296,N_2968);
xnor U4390 (N_4390,N_2227,N_2017);
xnor U4391 (N_4391,N_3618,N_3087);
or U4392 (N_4392,N_3876,N_2737);
and U4393 (N_4393,N_3168,N_2133);
and U4394 (N_4394,N_3913,N_2906);
and U4395 (N_4395,N_3933,N_3078);
nand U4396 (N_4396,N_2206,N_3748);
nor U4397 (N_4397,N_2222,N_3855);
nor U4398 (N_4398,N_3755,N_3610);
nor U4399 (N_4399,N_3368,N_2812);
nand U4400 (N_4400,N_3414,N_3998);
nor U4401 (N_4401,N_2173,N_3513);
xor U4402 (N_4402,N_2471,N_2859);
xnor U4403 (N_4403,N_3349,N_3224);
nand U4404 (N_4404,N_2009,N_3526);
xor U4405 (N_4405,N_3954,N_3866);
and U4406 (N_4406,N_2989,N_2950);
nand U4407 (N_4407,N_2055,N_3404);
xor U4408 (N_4408,N_2678,N_2409);
or U4409 (N_4409,N_2292,N_2576);
xnor U4410 (N_4410,N_2857,N_2622);
and U4411 (N_4411,N_3438,N_2333);
nor U4412 (N_4412,N_3844,N_3092);
nor U4413 (N_4413,N_2791,N_3886);
and U4414 (N_4414,N_2449,N_3928);
or U4415 (N_4415,N_3398,N_3745);
xnor U4416 (N_4416,N_2024,N_2196);
nand U4417 (N_4417,N_2323,N_2793);
xor U4418 (N_4418,N_2261,N_3874);
nor U4419 (N_4419,N_3137,N_3645);
and U4420 (N_4420,N_2162,N_3594);
and U4421 (N_4421,N_2371,N_3782);
or U4422 (N_4422,N_2293,N_3481);
nor U4423 (N_4423,N_2848,N_3545);
or U4424 (N_4424,N_2925,N_3670);
or U4425 (N_4425,N_3997,N_3591);
nand U4426 (N_4426,N_2528,N_3172);
xnor U4427 (N_4427,N_3664,N_2573);
and U4428 (N_4428,N_3540,N_2756);
nand U4429 (N_4429,N_3014,N_2854);
xor U4430 (N_4430,N_2393,N_2526);
nand U4431 (N_4431,N_2781,N_2382);
and U4432 (N_4432,N_3741,N_2631);
nand U4433 (N_4433,N_3058,N_3762);
or U4434 (N_4434,N_3057,N_2917);
xnor U4435 (N_4435,N_3166,N_3352);
xor U4436 (N_4436,N_3975,N_2879);
and U4437 (N_4437,N_2913,N_2011);
nand U4438 (N_4438,N_3892,N_2740);
nand U4439 (N_4439,N_2707,N_3221);
xor U4440 (N_4440,N_3297,N_3482);
or U4441 (N_4441,N_2985,N_2598);
nor U4442 (N_4442,N_3925,N_2529);
and U4443 (N_4443,N_2180,N_3185);
and U4444 (N_4444,N_3963,N_3989);
and U4445 (N_4445,N_2480,N_3131);
nand U4446 (N_4446,N_3959,N_2869);
nor U4447 (N_4447,N_3463,N_2759);
nand U4448 (N_4448,N_2389,N_3971);
nand U4449 (N_4449,N_2905,N_3774);
nand U4450 (N_4450,N_2497,N_3282);
xor U4451 (N_4451,N_2997,N_2467);
xor U4452 (N_4452,N_2900,N_3076);
xor U4453 (N_4453,N_2524,N_3865);
nor U4454 (N_4454,N_2235,N_2956);
nor U4455 (N_4455,N_3495,N_2078);
nand U4456 (N_4456,N_2828,N_3616);
nor U4457 (N_4457,N_3952,N_3522);
nor U4458 (N_4458,N_2129,N_2864);
xnor U4459 (N_4459,N_3947,N_2421);
and U4460 (N_4460,N_2637,N_2567);
xor U4461 (N_4461,N_3537,N_3100);
nand U4462 (N_4462,N_2365,N_3399);
xnor U4463 (N_4463,N_2741,N_2971);
or U4464 (N_4464,N_2216,N_3189);
nand U4465 (N_4465,N_2871,N_3251);
nand U4466 (N_4466,N_3509,N_2767);
nor U4467 (N_4467,N_2084,N_3912);
or U4468 (N_4468,N_3425,N_3783);
and U4469 (N_4469,N_3879,N_3607);
and U4470 (N_4470,N_2375,N_2503);
and U4471 (N_4471,N_3630,N_3145);
or U4472 (N_4472,N_2533,N_2232);
and U4473 (N_4473,N_2893,N_3472);
or U4474 (N_4474,N_3827,N_2337);
or U4475 (N_4475,N_2938,N_3070);
or U4476 (N_4476,N_3154,N_2221);
or U4477 (N_4477,N_3127,N_3190);
or U4478 (N_4478,N_3891,N_2693);
nand U4479 (N_4479,N_2903,N_3358);
nor U4480 (N_4480,N_2835,N_2182);
and U4481 (N_4481,N_3007,N_3067);
xor U4482 (N_4482,N_2896,N_3707);
and U4483 (N_4483,N_2664,N_2257);
and U4484 (N_4484,N_3243,N_3507);
nand U4485 (N_4485,N_2356,N_2043);
or U4486 (N_4486,N_3697,N_3144);
xnor U4487 (N_4487,N_2898,N_3086);
or U4488 (N_4488,N_3074,N_2051);
and U4489 (N_4489,N_2851,N_2911);
xor U4490 (N_4490,N_2192,N_3511);
and U4491 (N_4491,N_2291,N_3902);
xor U4492 (N_4492,N_2914,N_3228);
nor U4493 (N_4493,N_2999,N_2026);
or U4494 (N_4494,N_3702,N_2612);
xor U4495 (N_4495,N_2282,N_2994);
and U4496 (N_4496,N_2689,N_3257);
and U4497 (N_4497,N_3625,N_2735);
or U4498 (N_4498,N_3943,N_3647);
nand U4499 (N_4499,N_3426,N_2748);
and U4500 (N_4500,N_3017,N_3345);
nand U4501 (N_4501,N_3446,N_2952);
or U4502 (N_4502,N_2283,N_2520);
and U4503 (N_4503,N_2352,N_2770);
and U4504 (N_4504,N_3336,N_3718);
xor U4505 (N_4505,N_3966,N_2569);
or U4506 (N_4506,N_3286,N_2330);
xnor U4507 (N_4507,N_2850,N_2665);
nor U4508 (N_4508,N_2716,N_2743);
and U4509 (N_4509,N_2553,N_2641);
xor U4510 (N_4510,N_2309,N_2739);
and U4511 (N_4511,N_3121,N_3877);
or U4512 (N_4512,N_2098,N_3384);
nand U4513 (N_4513,N_2140,N_2072);
or U4514 (N_4514,N_2284,N_2874);
nor U4515 (N_4515,N_3944,N_3180);
and U4516 (N_4516,N_2694,N_2304);
nor U4517 (N_4517,N_2251,N_3208);
or U4518 (N_4518,N_2445,N_2824);
xor U4519 (N_4519,N_2760,N_3839);
nand U4520 (N_4520,N_3695,N_2054);
nor U4521 (N_4521,N_3319,N_3196);
xor U4522 (N_4522,N_3308,N_2984);
or U4523 (N_4523,N_2930,N_2881);
or U4524 (N_4524,N_2621,N_3870);
or U4525 (N_4525,N_2484,N_2607);
and U4526 (N_4526,N_3642,N_3830);
or U4527 (N_4527,N_2056,N_2908);
xnor U4528 (N_4528,N_3324,N_3291);
nor U4529 (N_4529,N_3448,N_3648);
and U4530 (N_4530,N_2138,N_3361);
xnor U4531 (N_4531,N_2008,N_2710);
nor U4532 (N_4532,N_3337,N_2424);
nand U4533 (N_4533,N_2018,N_2285);
xnor U4534 (N_4534,N_3761,N_2673);
nand U4535 (N_4535,N_2654,N_3159);
nand U4536 (N_4536,N_3303,N_3623);
nor U4537 (N_4537,N_3292,N_3808);
nor U4538 (N_4538,N_2299,N_3402);
xor U4539 (N_4539,N_2308,N_3863);
or U4540 (N_4540,N_2322,N_2703);
nand U4541 (N_4541,N_2670,N_3396);
or U4542 (N_4542,N_3786,N_2324);
or U4543 (N_4543,N_3136,N_2655);
or U4544 (N_4544,N_2317,N_3675);
nand U4545 (N_4545,N_3731,N_2473);
xor U4546 (N_4546,N_3474,N_3294);
nand U4547 (N_4547,N_3204,N_2267);
or U4548 (N_4548,N_3524,N_2109);
nor U4549 (N_4549,N_3301,N_2661);
xnor U4550 (N_4550,N_2212,N_2440);
or U4551 (N_4551,N_2532,N_3964);
nand U4552 (N_4552,N_2457,N_3832);
xor U4553 (N_4553,N_2821,N_3435);
or U4554 (N_4554,N_2247,N_2616);
and U4555 (N_4555,N_3305,N_3897);
or U4556 (N_4556,N_3081,N_2775);
nand U4557 (N_4557,N_3548,N_2047);
xor U4558 (N_4558,N_2912,N_3010);
nor U4559 (N_4559,N_3627,N_3953);
xor U4560 (N_4560,N_3699,N_2242);
and U4561 (N_4561,N_2934,N_3716);
xnor U4562 (N_4562,N_3117,N_3125);
nand U4563 (N_4563,N_2286,N_3787);
and U4564 (N_4564,N_3566,N_2604);
nand U4565 (N_4565,N_2413,N_3054);
nand U4566 (N_4566,N_3858,N_3793);
and U4567 (N_4567,N_3900,N_2046);
nor U4568 (N_4568,N_2712,N_2686);
or U4569 (N_4569,N_2462,N_2272);
xnor U4570 (N_4570,N_2565,N_3656);
xor U4571 (N_4571,N_3752,N_2430);
and U4572 (N_4572,N_3810,N_2768);
nand U4573 (N_4573,N_3962,N_2136);
xor U4574 (N_4574,N_2451,N_2029);
nand U4575 (N_4575,N_3363,N_2161);
xor U4576 (N_4576,N_2296,N_2446);
and U4577 (N_4577,N_3130,N_2068);
and U4578 (N_4578,N_2597,N_2123);
or U4579 (N_4579,N_2787,N_3907);
and U4580 (N_4580,N_3071,N_3920);
xor U4581 (N_4581,N_2610,N_3728);
or U4582 (N_4582,N_2039,N_3357);
nand U4583 (N_4583,N_3922,N_2965);
nand U4584 (N_4584,N_2513,N_3119);
nor U4585 (N_4585,N_2695,N_3278);
and U4586 (N_4586,N_3624,N_3854);
nor U4587 (N_4587,N_3373,N_3608);
nor U4588 (N_4588,N_3313,N_3016);
nand U4589 (N_4589,N_2509,N_3332);
and U4590 (N_4590,N_2408,N_2437);
or U4591 (N_4591,N_3027,N_3451);
nor U4592 (N_4592,N_3906,N_2590);
xor U4593 (N_4593,N_2474,N_3974);
or U4594 (N_4594,N_3836,N_3108);
xnor U4595 (N_4595,N_2578,N_3115);
nor U4596 (N_4596,N_2175,N_2188);
nand U4597 (N_4597,N_3104,N_3580);
nor U4598 (N_4598,N_3001,N_2269);
or U4599 (N_4599,N_2454,N_2546);
xnor U4600 (N_4600,N_3041,N_2810);
nand U4601 (N_4601,N_2853,N_3233);
and U4602 (N_4602,N_3682,N_3567);
or U4603 (N_4603,N_3871,N_3161);
and U4604 (N_4604,N_2096,N_2651);
nand U4605 (N_4605,N_3249,N_2374);
and U4606 (N_4606,N_3335,N_3231);
xor U4607 (N_4607,N_3881,N_2704);
nor U4608 (N_4608,N_2754,N_3376);
nor U4609 (N_4609,N_3935,N_3364);
and U4610 (N_4610,N_3015,N_2327);
or U4611 (N_4611,N_2876,N_2771);
nand U4612 (N_4612,N_2515,N_2530);
or U4613 (N_4613,N_2496,N_2147);
xnor U4614 (N_4614,N_2758,N_3816);
xor U4615 (N_4615,N_2559,N_2801);
and U4616 (N_4616,N_3600,N_2475);
xnor U4617 (N_4617,N_2099,N_2983);
nand U4618 (N_4618,N_3191,N_2492);
or U4619 (N_4619,N_3491,N_3613);
nand U4620 (N_4620,N_3295,N_2866);
nor U4621 (N_4621,N_2884,N_2543);
nor U4622 (N_4622,N_3476,N_3211);
xnor U4623 (N_4623,N_2924,N_2458);
and U4624 (N_4624,N_3178,N_2254);
nor U4625 (N_4625,N_2545,N_3631);
nor U4626 (N_4626,N_3410,N_2328);
xnor U4627 (N_4627,N_2486,N_2159);
xor U4628 (N_4628,N_3503,N_3842);
or U4629 (N_4629,N_3751,N_3643);
xnor U4630 (N_4630,N_2329,N_2483);
and U4631 (N_4631,N_2717,N_2599);
xnor U4632 (N_4632,N_3394,N_2131);
nand U4633 (N_4633,N_2976,N_2489);
xnor U4634 (N_4634,N_2360,N_3096);
and U4635 (N_4635,N_3193,N_3202);
nor U4636 (N_4636,N_2472,N_2953);
xor U4637 (N_4637,N_2005,N_3106);
or U4638 (N_4638,N_3201,N_2557);
xnor U4639 (N_4639,N_2840,N_2334);
and U4640 (N_4640,N_3388,N_2398);
nand U4641 (N_4641,N_3929,N_3910);
nor U4642 (N_4642,N_2390,N_3069);
and U4643 (N_4643,N_3693,N_2650);
nor U4644 (N_4644,N_3049,N_2100);
and U4645 (N_4645,N_3454,N_3330);
and U4646 (N_4646,N_3457,N_3123);
nor U4647 (N_4647,N_3235,N_3720);
nor U4648 (N_4648,N_2114,N_2817);
or U4649 (N_4649,N_2709,N_3008);
nand U4650 (N_4650,N_2732,N_2373);
or U4651 (N_4651,N_2692,N_2935);
nor U4652 (N_4652,N_2536,N_3889);
nor U4653 (N_4653,N_2873,N_2803);
xor U4654 (N_4654,N_2841,N_2233);
xor U4655 (N_4655,N_2544,N_2125);
and U4656 (N_4656,N_2340,N_2799);
and U4657 (N_4657,N_3203,N_2336);
or U4658 (N_4658,N_2584,N_2057);
and U4659 (N_4659,N_2720,N_2358);
and U4660 (N_4660,N_3431,N_2804);
or U4661 (N_4661,N_3704,N_3869);
and U4662 (N_4662,N_2279,N_2795);
or U4663 (N_4663,N_3638,N_2690);
and U4664 (N_4664,N_3883,N_3710);
nor U4665 (N_4665,N_3273,N_2636);
and U4666 (N_4666,N_3156,N_2224);
and U4667 (N_4667,N_3461,N_2124);
or U4668 (N_4668,N_3583,N_2820);
nor U4669 (N_4669,N_2676,N_3530);
and U4670 (N_4670,N_3706,N_2838);
or U4671 (N_4671,N_2516,N_2032);
or U4672 (N_4672,N_2506,N_2724);
nor U4673 (N_4673,N_3689,N_2263);
nand U4674 (N_4674,N_3671,N_3531);
nor U4675 (N_4675,N_2231,N_2833);
xor U4676 (N_4676,N_3430,N_3465);
nor U4677 (N_4677,N_3585,N_2036);
and U4678 (N_4678,N_2834,N_3085);
nand U4679 (N_4679,N_2766,N_2653);
or U4680 (N_4680,N_2082,N_2307);
nand U4681 (N_4681,N_2722,N_3992);
or U4682 (N_4682,N_3599,N_2306);
or U4683 (N_4683,N_2271,N_2126);
nand U4684 (N_4684,N_3050,N_3969);
xnor U4685 (N_4685,N_2425,N_3615);
nor U4686 (N_4686,N_2822,N_2558);
or U4687 (N_4687,N_3389,N_2482);
nand U4688 (N_4688,N_3379,N_2157);
xor U4689 (N_4689,N_2107,N_3306);
nand U4690 (N_4690,N_2765,N_2203);
and U4691 (N_4691,N_3244,N_3265);
xor U4692 (N_4692,N_2519,N_2777);
nand U4693 (N_4693,N_3677,N_2589);
nand U4694 (N_4694,N_2152,N_3619);
or U4695 (N_4695,N_3781,N_2729);
xor U4696 (N_4696,N_3601,N_3164);
or U4697 (N_4697,N_2962,N_3799);
or U4698 (N_4698,N_3771,N_3528);
and U4699 (N_4699,N_3770,N_2888);
nor U4700 (N_4700,N_3976,N_2229);
nor U4701 (N_4701,N_2769,N_3517);
xnor U4702 (N_4702,N_3411,N_3344);
nor U4703 (N_4703,N_3255,N_3772);
nor U4704 (N_4704,N_2863,N_2783);
nand U4705 (N_4705,N_2453,N_2596);
or U4706 (N_4706,N_2696,N_2459);
nor U4707 (N_4707,N_2619,N_3841);
and U4708 (N_4708,N_2171,N_3773);
or U4709 (N_4709,N_3132,N_3571);
and U4710 (N_4710,N_3896,N_2346);
nor U4711 (N_4711,N_3037,N_3135);
or U4712 (N_4712,N_2241,N_3005);
or U4713 (N_4713,N_3687,N_3199);
nor U4714 (N_4714,N_2234,N_2448);
nand U4715 (N_4715,N_2048,N_3506);
nor U4716 (N_4716,N_3831,N_2255);
xnor U4717 (N_4717,N_3192,N_2461);
nand U4718 (N_4718,N_3967,N_3021);
nand U4719 (N_4719,N_2067,N_3838);
nor U4720 (N_4720,N_2945,N_3315);
xnor U4721 (N_4721,N_3299,N_3280);
xnor U4722 (N_4722,N_2560,N_3077);
nor U4723 (N_4723,N_3409,N_2213);
nand U4724 (N_4724,N_2273,N_2566);
nor U4725 (N_4725,N_2211,N_2967);
xor U4726 (N_4726,N_3890,N_2811);
xnor U4727 (N_4727,N_2276,N_3760);
and U4728 (N_4728,N_3661,N_2963);
nand U4729 (N_4729,N_3225,N_2730);
nor U4730 (N_4730,N_2014,N_2657);
or U4731 (N_4731,N_3852,N_3321);
or U4732 (N_4732,N_3899,N_2926);
or U4733 (N_4733,N_3649,N_3802);
and U4734 (N_4734,N_2755,N_2907);
or U4735 (N_4735,N_2639,N_3160);
nand U4736 (N_4736,N_2680,N_3489);
and U4737 (N_4737,N_2698,N_3236);
nand U4738 (N_4738,N_3369,N_3323);
nand U4739 (N_4739,N_3266,N_3893);
nor U4740 (N_4740,N_3098,N_2514);
xnor U4741 (N_4741,N_3814,N_3766);
xor U4742 (N_4742,N_3262,N_3775);
and U4743 (N_4743,N_3128,N_2683);
nand U4744 (N_4744,N_3143,N_2112);
nor U4745 (N_4745,N_3686,N_2630);
nand U4746 (N_4746,N_2295,N_3637);
and U4747 (N_4747,N_2837,N_3277);
nand U4748 (N_4748,N_3091,N_3492);
nand U4749 (N_4749,N_2554,N_2076);
or U4750 (N_4750,N_2929,N_2154);
xor U4751 (N_4751,N_2256,N_2435);
and U4752 (N_4752,N_2892,N_2959);
nor U4753 (N_4753,N_2022,N_3359);
or U4754 (N_4754,N_3691,N_3066);
or U4755 (N_4755,N_2294,N_2615);
xnor U4756 (N_4756,N_3569,N_2300);
nor U4757 (N_4757,N_2606,N_3826);
xnor U4758 (N_4758,N_3317,N_2012);
or U4759 (N_4759,N_3490,N_2944);
nand U4760 (N_4760,N_2742,N_3575);
or U4761 (N_4761,N_2319,N_2103);
nand U4762 (N_4762,N_2749,N_3322);
xor U4763 (N_4763,N_2197,N_2746);
xor U4764 (N_4764,N_2649,N_3672);
nand U4765 (N_4765,N_3904,N_3735);
nand U4766 (N_4766,N_3809,N_3550);
nor U4767 (N_4767,N_3484,N_2025);
nor U4768 (N_4768,N_2069,N_3311);
nand U4769 (N_4769,N_2688,N_3584);
or U4770 (N_4770,N_3984,N_2095);
or U4771 (N_4771,N_2023,N_3727);
nor U4772 (N_4772,N_3263,N_3563);
xnor U4773 (N_4773,N_3590,N_2044);
xor U4774 (N_4774,N_3529,N_2148);
nor U4775 (N_4775,N_3182,N_3102);
nor U4776 (N_4776,N_3186,N_2045);
and U4777 (N_4777,N_2986,N_3279);
nor U4778 (N_4778,N_3381,N_3712);
and U4779 (N_4779,N_3415,N_2648);
nand U4780 (N_4780,N_3346,N_3777);
nor U4781 (N_4781,N_2137,N_2426);
or U4782 (N_4782,N_3247,N_2368);
or U4783 (N_4783,N_2456,N_3982);
xnor U4784 (N_4784,N_2831,N_3539);
and U4785 (N_4785,N_3586,N_3450);
or U4786 (N_4786,N_3039,N_3403);
xnor U4787 (N_4787,N_3941,N_2936);
nor U4788 (N_4788,N_3768,N_2563);
or U4789 (N_4789,N_2603,N_2921);
xnor U4790 (N_4790,N_2613,N_3579);
xor U4791 (N_4791,N_3651,N_2210);
and U4792 (N_4792,N_3614,N_3444);
or U4793 (N_4793,N_2268,N_3237);
nor U4794 (N_4794,N_3535,N_3442);
or U4795 (N_4795,N_2158,N_2608);
and U4796 (N_4796,N_2662,N_3025);
nand U4797 (N_4797,N_3400,N_3120);
and U4798 (N_4798,N_3791,N_2666);
and U4799 (N_4799,N_2744,N_2949);
nor U4800 (N_4800,N_2150,N_3163);
or U4801 (N_4801,N_3888,N_3097);
nand U4802 (N_4802,N_3940,N_3105);
xor U4803 (N_4803,N_2064,N_2667);
or U4804 (N_4804,N_2786,N_3957);
nand U4805 (N_4805,N_3665,N_2518);
nor U4806 (N_4806,N_2264,N_3024);
nand U4807 (N_4807,N_2418,N_3094);
nand U4808 (N_4808,N_2845,N_3223);
nand U4809 (N_4809,N_2061,N_3440);
or U4810 (N_4810,N_2512,N_2643);
xor U4811 (N_4811,N_2618,N_2561);
xnor U4812 (N_4812,N_3508,N_3068);
xor U4813 (N_4813,N_3817,N_3375);
or U4814 (N_4814,N_2790,N_2568);
and U4815 (N_4815,N_3972,N_2839);
nor U4816 (N_4816,N_3898,N_2217);
xor U4817 (N_4817,N_2789,N_3488);
nor U4818 (N_4818,N_3059,N_2832);
xnor U4819 (N_4819,N_3703,N_2411);
xor U4820 (N_4820,N_3060,N_2419);
nor U4821 (N_4821,N_2727,N_3436);
nor U4822 (N_4822,N_2156,N_2325);
or U4823 (N_4823,N_3848,N_2499);
xnor U4824 (N_4824,N_2189,N_2539);
xnor U4825 (N_4825,N_3033,N_2635);
nor U4826 (N_4826,N_3230,N_2301);
and U4827 (N_4827,N_3275,N_2600);
or U4828 (N_4828,N_3293,N_2244);
and U4829 (N_4829,N_2583,N_3167);
or U4830 (N_4830,N_2632,N_3383);
nor U4831 (N_4831,N_3924,N_3418);
xor U4832 (N_4832,N_2843,N_2404);
and U4833 (N_4833,N_2671,N_2119);
or U4834 (N_4834,N_2627,N_2342);
or U4835 (N_4835,N_3754,N_3604);
nor U4836 (N_4836,N_2252,N_3729);
xnor U4837 (N_4837,N_2302,N_2809);
xnor U4838 (N_4838,N_3309,N_3995);
xor U4839 (N_4839,N_2441,N_3417);
xor U4840 (N_4840,N_2379,N_3818);
nand U4841 (N_4841,N_3240,N_3118);
or U4842 (N_4842,N_3587,N_3851);
nor U4843 (N_4843,N_2215,N_2343);
or U4844 (N_4844,N_3919,N_2105);
or U4845 (N_4845,N_3395,N_3034);
and U4846 (N_4846,N_3063,N_3188);
or U4847 (N_4847,N_3927,N_2998);
and U4848 (N_4848,N_3717,N_2447);
and U4849 (N_4849,N_2111,N_2120);
and U4850 (N_4850,N_3218,N_3932);
nand U4851 (N_4851,N_2806,N_3845);
or U4852 (N_4852,N_3825,N_2179);
and U4853 (N_4853,N_3036,N_2966);
xnor U4854 (N_4854,N_3562,N_2318);
nor U4855 (N_4855,N_3819,N_3853);
nor U4856 (N_4856,N_2652,N_3965);
nor U4857 (N_4857,N_3990,N_3239);
and U4858 (N_4858,N_2239,N_2433);
nor U4859 (N_4859,N_2808,N_3988);
or U4860 (N_4860,N_2280,N_2155);
or U4861 (N_4861,N_3210,N_2397);
and U4862 (N_4862,N_3216,N_3525);
xnor U4863 (N_4863,N_2870,N_2542);
and U4864 (N_4864,N_2702,N_2939);
nand U4865 (N_4865,N_3804,N_3090);
nor U4866 (N_4866,N_2110,N_2711);
nor U4867 (N_4867,N_3516,N_2531);
xnor U4868 (N_4868,N_2562,N_3340);
nor U4869 (N_4869,N_2169,N_2391);
xnor U4870 (N_4870,N_3698,N_2050);
or U4871 (N_4871,N_3556,N_3134);
nand U4872 (N_4872,N_2658,N_3986);
and U4873 (N_4873,N_3151,N_2417);
nor U4874 (N_4874,N_2868,N_2918);
or U4875 (N_4875,N_2494,N_2200);
xor U4876 (N_4876,N_2135,N_3909);
nand U4877 (N_4877,N_2245,N_2904);
xnor U4878 (N_4878,N_3498,N_3181);
xor U4879 (N_4879,N_3692,N_3725);
xor U4880 (N_4880,N_2852,N_2097);
or U4881 (N_4881,N_2220,N_3325);
or U4882 (N_4882,N_3737,N_2058);
nor U4883 (N_4883,N_2640,N_2814);
xor U4884 (N_4884,N_3479,N_3353);
nor U4885 (N_4885,N_2468,N_3593);
xor U4886 (N_4886,N_3552,N_2495);
xnor U4887 (N_4887,N_2079,N_2338);
nand U4888 (N_4888,N_3536,N_3055);
nand U4889 (N_4889,N_3867,N_2875);
xnor U4890 (N_4890,N_3980,N_3285);
nor U4891 (N_4891,N_3887,N_2955);
xor U4892 (N_4892,N_2052,N_2728);
nor U4893 (N_4893,N_2490,N_3688);
xnor U4894 (N_4894,N_2901,N_3577);
or U4895 (N_4895,N_3946,N_2281);
xor U4896 (N_4896,N_3270,N_2066);
nand U4897 (N_4897,N_2466,N_2669);
nand U4898 (N_4898,N_2321,N_2611);
xor U4899 (N_4899,N_2540,N_2021);
and U4900 (N_4900,N_3416,N_3626);
nand U4901 (N_4901,N_2406,N_3561);
nor U4902 (N_4902,N_2679,N_3512);
nor U4903 (N_4903,N_2238,N_2376);
or U4904 (N_4904,N_3246,N_3811);
or U4905 (N_4905,N_2353,N_2399);
nor U4906 (N_4906,N_3807,N_2086);
nand U4907 (N_4907,N_3032,N_2880);
nand U4908 (N_4908,N_3302,N_3018);
nand U4909 (N_4909,N_3030,N_3708);
and U4910 (N_4910,N_2117,N_3527);
or U4911 (N_4911,N_3864,N_3644);
xor U4912 (N_4912,N_3598,N_2723);
or U4913 (N_4913,N_2960,N_3950);
and U4914 (N_4914,N_2427,N_3140);
nor U4915 (N_4915,N_3334,N_2149);
nor U4916 (N_4916,N_2577,N_3936);
nand U4917 (N_4917,N_2313,N_2225);
xor U4918 (N_4918,N_2165,N_3795);
or U4919 (N_4919,N_2316,N_3696);
xnor U4920 (N_4920,N_3666,N_2089);
and U4921 (N_4921,N_3259,N_2444);
xor U4922 (N_4922,N_3260,N_3044);
and U4923 (N_4923,N_2102,N_3701);
nor U4924 (N_4924,N_2266,N_2392);
nand U4925 (N_4925,N_2796,N_3470);
and U4926 (N_4926,N_2552,N_3669);
nand U4927 (N_4927,N_3532,N_2372);
and U4928 (N_4928,N_3371,N_3901);
and U4929 (N_4929,N_3622,N_2070);
or U4930 (N_4930,N_3310,N_3726);
nor U4931 (N_4931,N_2505,N_3872);
nor U4932 (N_4932,N_3673,N_3013);
and U4933 (N_4933,N_2344,N_2973);
and U4934 (N_4934,N_3723,N_2027);
xnor U4935 (N_4935,N_3543,N_3298);
xnor U4936 (N_4936,N_2830,N_3133);
xnor U4937 (N_4937,N_2780,N_3469);
or U4938 (N_4938,N_3473,N_3038);
nand U4939 (N_4939,N_3641,N_3150);
or U4940 (N_4940,N_3711,N_3837);
nor U4941 (N_4941,N_3439,N_3042);
nand U4942 (N_4942,N_3162,N_2899);
and U4943 (N_4943,N_3214,N_3445);
or U4944 (N_4944,N_2237,N_3124);
nor U4945 (N_4945,N_3173,N_2455);
nor U4946 (N_4946,N_3056,N_2794);
nor U4947 (N_4947,N_2312,N_3746);
nor U4948 (N_4948,N_3981,N_3453);
and U4949 (N_4949,N_3175,N_2594);
nand U4950 (N_4950,N_2587,N_2718);
nor U4951 (N_4951,N_3659,N_3639);
or U4952 (N_4952,N_3437,N_3385);
or U4953 (N_4953,N_2807,N_3477);
nor U4954 (N_4954,N_3632,N_2687);
xnor U4955 (N_4955,N_2836,N_3219);
or U4956 (N_4956,N_2187,N_3382);
or U4957 (N_4957,N_3518,N_3987);
or U4958 (N_4958,N_2946,N_2510);
nand U4959 (N_4959,N_2429,N_2214);
nand U4960 (N_4960,N_2075,N_3738);
xnor U4961 (N_4961,N_2668,N_2815);
nand U4962 (N_4962,N_3640,N_3338);
nor U4963 (N_4963,N_2361,N_3023);
nand U4964 (N_4964,N_3494,N_3885);
nand U4965 (N_4965,N_2275,N_2591);
xnor U4966 (N_4966,N_2493,N_2802);
nor U4967 (N_4967,N_3750,N_3797);
nand U4968 (N_4968,N_2452,N_3700);
nand U4969 (N_4969,N_3176,N_3657);
nand U4970 (N_4970,N_3678,N_3051);
nor U4971 (N_4971,N_3011,N_2979);
or U4972 (N_4972,N_2395,N_2259);
xnor U4973 (N_4973,N_2060,N_2166);
nor U4974 (N_4974,N_2428,N_3734);
nand U4975 (N_4975,N_2420,N_2626);
nor U4976 (N_4976,N_2774,N_2385);
or U4977 (N_4977,N_3958,N_2370);
xor U4978 (N_4978,N_3261,N_3515);
nor U4979 (N_4979,N_3320,N_3523);
nor U4980 (N_4980,N_2990,N_2860);
or U4981 (N_4981,N_3694,N_2181);
and U4982 (N_4982,N_3934,N_2274);
nor U4983 (N_4983,N_2571,N_2049);
or U4984 (N_4984,N_3080,N_2988);
or U4985 (N_4985,N_3019,N_2897);
xnor U4986 (N_4986,N_2020,N_3636);
or U4987 (N_4987,N_3983,N_2726);
xnor U4988 (N_4988,N_2601,N_3464);
xor U4989 (N_4989,N_3258,N_3589);
nor U4990 (N_4990,N_2479,N_2498);
nand U4991 (N_4991,N_2844,N_2818);
nor U4992 (N_4992,N_2041,N_3187);
nand U4993 (N_4993,N_3387,N_2460);
nand U4994 (N_4994,N_3129,N_3138);
and U4995 (N_4995,N_2088,N_2491);
xnor U4996 (N_4996,N_3206,N_2083);
xnor U4997 (N_4997,N_2757,N_3209);
nand U4998 (N_4998,N_2886,N_2778);
xnor U4999 (N_4999,N_2501,N_2628);
and U5000 (N_5000,N_3808,N_3108);
nor U5001 (N_5001,N_2162,N_3567);
or U5002 (N_5002,N_3777,N_2064);
nand U5003 (N_5003,N_3840,N_3032);
and U5004 (N_5004,N_2827,N_3713);
nand U5005 (N_5005,N_3251,N_3777);
and U5006 (N_5006,N_3697,N_3142);
nand U5007 (N_5007,N_2747,N_3916);
or U5008 (N_5008,N_3792,N_2761);
nand U5009 (N_5009,N_3566,N_2923);
nor U5010 (N_5010,N_2118,N_3350);
nor U5011 (N_5011,N_3499,N_2104);
or U5012 (N_5012,N_3923,N_2828);
or U5013 (N_5013,N_2270,N_3833);
and U5014 (N_5014,N_2301,N_3506);
xnor U5015 (N_5015,N_2298,N_3691);
xor U5016 (N_5016,N_2036,N_2486);
xnor U5017 (N_5017,N_3566,N_2663);
or U5018 (N_5018,N_3893,N_2647);
nor U5019 (N_5019,N_2963,N_2180);
or U5020 (N_5020,N_3823,N_3340);
xnor U5021 (N_5021,N_2512,N_2145);
xor U5022 (N_5022,N_2652,N_3902);
nor U5023 (N_5023,N_2544,N_3307);
and U5024 (N_5024,N_2910,N_3011);
nand U5025 (N_5025,N_2483,N_3510);
nand U5026 (N_5026,N_2171,N_3431);
nor U5027 (N_5027,N_2019,N_2568);
xor U5028 (N_5028,N_3342,N_3506);
or U5029 (N_5029,N_3226,N_2315);
nor U5030 (N_5030,N_3997,N_3959);
and U5031 (N_5031,N_3078,N_3176);
and U5032 (N_5032,N_3741,N_2378);
xnor U5033 (N_5033,N_2467,N_3334);
nor U5034 (N_5034,N_3182,N_3124);
or U5035 (N_5035,N_2059,N_3903);
xnor U5036 (N_5036,N_2446,N_3593);
xnor U5037 (N_5037,N_2100,N_2708);
xnor U5038 (N_5038,N_2371,N_2918);
nor U5039 (N_5039,N_3974,N_2216);
and U5040 (N_5040,N_2780,N_3093);
and U5041 (N_5041,N_3405,N_2181);
xor U5042 (N_5042,N_2917,N_2835);
xor U5043 (N_5043,N_3929,N_2522);
nand U5044 (N_5044,N_3750,N_2360);
and U5045 (N_5045,N_3009,N_2165);
or U5046 (N_5046,N_2081,N_3836);
nor U5047 (N_5047,N_3050,N_2500);
or U5048 (N_5048,N_2835,N_2043);
nand U5049 (N_5049,N_2813,N_2912);
or U5050 (N_5050,N_3416,N_3515);
and U5051 (N_5051,N_3752,N_3957);
nor U5052 (N_5052,N_2860,N_3272);
and U5053 (N_5053,N_3164,N_3085);
and U5054 (N_5054,N_2788,N_3198);
nand U5055 (N_5055,N_3870,N_2835);
and U5056 (N_5056,N_2661,N_3888);
nand U5057 (N_5057,N_2344,N_2076);
nor U5058 (N_5058,N_2248,N_3755);
or U5059 (N_5059,N_2673,N_2746);
nor U5060 (N_5060,N_2278,N_3565);
xnor U5061 (N_5061,N_3026,N_3560);
and U5062 (N_5062,N_2761,N_2989);
nor U5063 (N_5063,N_2207,N_2864);
or U5064 (N_5064,N_2505,N_3276);
nand U5065 (N_5065,N_3310,N_3982);
or U5066 (N_5066,N_3146,N_2019);
xor U5067 (N_5067,N_2542,N_2468);
nand U5068 (N_5068,N_2044,N_3655);
and U5069 (N_5069,N_2415,N_2715);
xor U5070 (N_5070,N_3612,N_3398);
or U5071 (N_5071,N_2786,N_2957);
nor U5072 (N_5072,N_3064,N_2293);
nand U5073 (N_5073,N_3445,N_2186);
and U5074 (N_5074,N_3121,N_3606);
or U5075 (N_5075,N_2569,N_2717);
nor U5076 (N_5076,N_3120,N_2650);
and U5077 (N_5077,N_2651,N_2094);
xor U5078 (N_5078,N_2776,N_2445);
nand U5079 (N_5079,N_3820,N_2545);
xnor U5080 (N_5080,N_2966,N_2340);
and U5081 (N_5081,N_3256,N_3214);
xor U5082 (N_5082,N_2610,N_2242);
and U5083 (N_5083,N_2399,N_2935);
or U5084 (N_5084,N_3762,N_3622);
and U5085 (N_5085,N_3031,N_2524);
or U5086 (N_5086,N_3436,N_2636);
and U5087 (N_5087,N_3421,N_3104);
nand U5088 (N_5088,N_2986,N_3648);
nor U5089 (N_5089,N_3492,N_3774);
nor U5090 (N_5090,N_3424,N_2413);
nor U5091 (N_5091,N_3145,N_2801);
nor U5092 (N_5092,N_2862,N_2289);
and U5093 (N_5093,N_3319,N_3223);
xor U5094 (N_5094,N_2020,N_3064);
nor U5095 (N_5095,N_2385,N_3713);
or U5096 (N_5096,N_2836,N_2252);
or U5097 (N_5097,N_2325,N_2125);
nand U5098 (N_5098,N_3219,N_2475);
xor U5099 (N_5099,N_2910,N_3734);
xnor U5100 (N_5100,N_2273,N_2419);
nand U5101 (N_5101,N_3250,N_2296);
nand U5102 (N_5102,N_3473,N_2488);
or U5103 (N_5103,N_2581,N_3498);
and U5104 (N_5104,N_3547,N_3663);
xor U5105 (N_5105,N_2918,N_3939);
or U5106 (N_5106,N_3569,N_3277);
nor U5107 (N_5107,N_2181,N_3253);
and U5108 (N_5108,N_2559,N_2348);
nor U5109 (N_5109,N_2475,N_2529);
xnor U5110 (N_5110,N_3612,N_2940);
xnor U5111 (N_5111,N_3116,N_3027);
and U5112 (N_5112,N_3364,N_2008);
nand U5113 (N_5113,N_2854,N_2292);
xnor U5114 (N_5114,N_3170,N_3132);
nor U5115 (N_5115,N_2866,N_2776);
nor U5116 (N_5116,N_2435,N_3401);
or U5117 (N_5117,N_2308,N_2786);
nand U5118 (N_5118,N_2486,N_2432);
nand U5119 (N_5119,N_3072,N_3061);
xnor U5120 (N_5120,N_3987,N_2705);
xor U5121 (N_5121,N_2978,N_2525);
or U5122 (N_5122,N_2401,N_3025);
and U5123 (N_5123,N_3138,N_3472);
and U5124 (N_5124,N_3632,N_3139);
nor U5125 (N_5125,N_2926,N_3485);
nor U5126 (N_5126,N_2246,N_2721);
nor U5127 (N_5127,N_2077,N_2290);
and U5128 (N_5128,N_3310,N_2400);
nand U5129 (N_5129,N_3654,N_3072);
nor U5130 (N_5130,N_2720,N_3272);
nand U5131 (N_5131,N_2498,N_2618);
nand U5132 (N_5132,N_3120,N_3621);
nand U5133 (N_5133,N_3014,N_3784);
xor U5134 (N_5134,N_3710,N_3036);
nand U5135 (N_5135,N_3067,N_3453);
and U5136 (N_5136,N_3824,N_3003);
and U5137 (N_5137,N_3873,N_3543);
and U5138 (N_5138,N_3164,N_3396);
nand U5139 (N_5139,N_3905,N_3902);
nand U5140 (N_5140,N_2843,N_2957);
nor U5141 (N_5141,N_2703,N_3497);
nand U5142 (N_5142,N_3610,N_3151);
and U5143 (N_5143,N_2891,N_2575);
and U5144 (N_5144,N_3685,N_3853);
and U5145 (N_5145,N_3829,N_2210);
nand U5146 (N_5146,N_2429,N_2818);
nand U5147 (N_5147,N_3246,N_3916);
xor U5148 (N_5148,N_3198,N_2533);
and U5149 (N_5149,N_2182,N_3184);
nor U5150 (N_5150,N_3650,N_2978);
xor U5151 (N_5151,N_3905,N_3393);
and U5152 (N_5152,N_2771,N_2487);
nor U5153 (N_5153,N_3624,N_2678);
nand U5154 (N_5154,N_3330,N_2867);
xnor U5155 (N_5155,N_2469,N_3995);
nand U5156 (N_5156,N_3241,N_3820);
xnor U5157 (N_5157,N_2549,N_3792);
xnor U5158 (N_5158,N_2050,N_2994);
and U5159 (N_5159,N_2062,N_2953);
and U5160 (N_5160,N_2850,N_2815);
nor U5161 (N_5161,N_3248,N_2889);
nor U5162 (N_5162,N_3320,N_3197);
and U5163 (N_5163,N_3758,N_2766);
xnor U5164 (N_5164,N_3707,N_2816);
or U5165 (N_5165,N_2753,N_3139);
or U5166 (N_5166,N_2783,N_2988);
xnor U5167 (N_5167,N_2432,N_3333);
or U5168 (N_5168,N_3327,N_3950);
or U5169 (N_5169,N_3879,N_3727);
and U5170 (N_5170,N_2664,N_2906);
nand U5171 (N_5171,N_2200,N_2812);
nand U5172 (N_5172,N_3045,N_2343);
nand U5173 (N_5173,N_3072,N_3998);
and U5174 (N_5174,N_3649,N_2888);
or U5175 (N_5175,N_2583,N_2756);
nand U5176 (N_5176,N_2202,N_2530);
or U5177 (N_5177,N_3967,N_3080);
and U5178 (N_5178,N_3974,N_3635);
or U5179 (N_5179,N_3903,N_2259);
xnor U5180 (N_5180,N_2357,N_2209);
xnor U5181 (N_5181,N_3532,N_3986);
or U5182 (N_5182,N_2668,N_2418);
nand U5183 (N_5183,N_3212,N_3368);
or U5184 (N_5184,N_3034,N_2812);
xnor U5185 (N_5185,N_2210,N_2613);
xor U5186 (N_5186,N_2483,N_2420);
nor U5187 (N_5187,N_2723,N_3440);
xnor U5188 (N_5188,N_2123,N_2877);
nor U5189 (N_5189,N_3782,N_3482);
or U5190 (N_5190,N_3077,N_3200);
nor U5191 (N_5191,N_3495,N_2647);
and U5192 (N_5192,N_3425,N_3171);
and U5193 (N_5193,N_3797,N_3654);
nor U5194 (N_5194,N_3122,N_2170);
and U5195 (N_5195,N_2059,N_2733);
nor U5196 (N_5196,N_2997,N_2789);
and U5197 (N_5197,N_2084,N_2304);
nand U5198 (N_5198,N_2877,N_2589);
nand U5199 (N_5199,N_2409,N_2449);
or U5200 (N_5200,N_2367,N_3707);
and U5201 (N_5201,N_2500,N_3952);
nor U5202 (N_5202,N_2709,N_3068);
or U5203 (N_5203,N_2411,N_2235);
nand U5204 (N_5204,N_2789,N_3292);
nand U5205 (N_5205,N_3142,N_3552);
or U5206 (N_5206,N_2693,N_2689);
nor U5207 (N_5207,N_2430,N_2757);
or U5208 (N_5208,N_2561,N_3804);
nand U5209 (N_5209,N_2937,N_2279);
or U5210 (N_5210,N_3688,N_3874);
xnor U5211 (N_5211,N_2927,N_2757);
and U5212 (N_5212,N_3466,N_2757);
and U5213 (N_5213,N_3025,N_3382);
nor U5214 (N_5214,N_2718,N_3935);
nand U5215 (N_5215,N_2998,N_3013);
xnor U5216 (N_5216,N_2510,N_2089);
and U5217 (N_5217,N_2498,N_3030);
nor U5218 (N_5218,N_3140,N_3165);
or U5219 (N_5219,N_3814,N_3238);
and U5220 (N_5220,N_2561,N_2476);
nor U5221 (N_5221,N_3971,N_2197);
or U5222 (N_5222,N_3394,N_3321);
and U5223 (N_5223,N_2652,N_2823);
and U5224 (N_5224,N_3968,N_2927);
and U5225 (N_5225,N_2280,N_3663);
nand U5226 (N_5226,N_3099,N_3903);
or U5227 (N_5227,N_2487,N_2843);
and U5228 (N_5228,N_2053,N_2555);
or U5229 (N_5229,N_2073,N_2812);
and U5230 (N_5230,N_2578,N_3171);
xnor U5231 (N_5231,N_3290,N_2286);
nand U5232 (N_5232,N_3220,N_3839);
nand U5233 (N_5233,N_3479,N_2802);
xnor U5234 (N_5234,N_2795,N_2380);
xnor U5235 (N_5235,N_2194,N_2874);
nand U5236 (N_5236,N_2586,N_3033);
or U5237 (N_5237,N_3739,N_3125);
xnor U5238 (N_5238,N_3503,N_2945);
nor U5239 (N_5239,N_3360,N_2903);
and U5240 (N_5240,N_2467,N_2736);
nor U5241 (N_5241,N_3969,N_2140);
nand U5242 (N_5242,N_3910,N_2884);
nor U5243 (N_5243,N_3181,N_3748);
nand U5244 (N_5244,N_2321,N_2859);
xor U5245 (N_5245,N_3939,N_2205);
xor U5246 (N_5246,N_2365,N_2080);
nor U5247 (N_5247,N_2554,N_2206);
xnor U5248 (N_5248,N_3560,N_2085);
xnor U5249 (N_5249,N_2411,N_3658);
xnor U5250 (N_5250,N_3630,N_2146);
xnor U5251 (N_5251,N_2779,N_2500);
nand U5252 (N_5252,N_2990,N_3282);
nand U5253 (N_5253,N_2135,N_3253);
nand U5254 (N_5254,N_3516,N_2621);
nor U5255 (N_5255,N_3252,N_2288);
and U5256 (N_5256,N_3851,N_3476);
and U5257 (N_5257,N_2908,N_2831);
nand U5258 (N_5258,N_2821,N_3648);
or U5259 (N_5259,N_2897,N_2232);
or U5260 (N_5260,N_3585,N_2998);
xnor U5261 (N_5261,N_2858,N_2351);
nand U5262 (N_5262,N_3875,N_3671);
xor U5263 (N_5263,N_3661,N_2526);
xor U5264 (N_5264,N_2723,N_3857);
nor U5265 (N_5265,N_2967,N_3048);
nand U5266 (N_5266,N_3283,N_3443);
or U5267 (N_5267,N_2437,N_2642);
and U5268 (N_5268,N_3156,N_3779);
nand U5269 (N_5269,N_2214,N_2176);
and U5270 (N_5270,N_3334,N_3142);
and U5271 (N_5271,N_3864,N_2765);
nor U5272 (N_5272,N_2316,N_3065);
xnor U5273 (N_5273,N_2349,N_3018);
or U5274 (N_5274,N_3925,N_3220);
nand U5275 (N_5275,N_3456,N_3881);
nor U5276 (N_5276,N_2605,N_2032);
or U5277 (N_5277,N_3673,N_3895);
nand U5278 (N_5278,N_3838,N_3103);
nor U5279 (N_5279,N_3651,N_2684);
nand U5280 (N_5280,N_3305,N_3995);
or U5281 (N_5281,N_2976,N_3000);
and U5282 (N_5282,N_2511,N_2282);
nor U5283 (N_5283,N_3855,N_3108);
nor U5284 (N_5284,N_2894,N_3770);
and U5285 (N_5285,N_2780,N_2991);
or U5286 (N_5286,N_3513,N_3503);
or U5287 (N_5287,N_3587,N_2187);
xnor U5288 (N_5288,N_3314,N_3919);
nor U5289 (N_5289,N_3492,N_3953);
xor U5290 (N_5290,N_2399,N_3598);
nand U5291 (N_5291,N_3522,N_3861);
nand U5292 (N_5292,N_3453,N_2350);
nand U5293 (N_5293,N_3079,N_2921);
and U5294 (N_5294,N_2200,N_3380);
or U5295 (N_5295,N_3656,N_2642);
xnor U5296 (N_5296,N_2099,N_3596);
or U5297 (N_5297,N_2863,N_2504);
xor U5298 (N_5298,N_2850,N_2353);
xor U5299 (N_5299,N_3457,N_3227);
nand U5300 (N_5300,N_2457,N_3209);
or U5301 (N_5301,N_3639,N_3398);
or U5302 (N_5302,N_3177,N_3441);
nor U5303 (N_5303,N_3059,N_3442);
or U5304 (N_5304,N_2682,N_3320);
nor U5305 (N_5305,N_3528,N_2057);
xnor U5306 (N_5306,N_2056,N_2561);
and U5307 (N_5307,N_2156,N_2327);
xnor U5308 (N_5308,N_2071,N_3712);
and U5309 (N_5309,N_2800,N_2938);
and U5310 (N_5310,N_2074,N_3711);
xor U5311 (N_5311,N_3839,N_3670);
and U5312 (N_5312,N_3702,N_2271);
nand U5313 (N_5313,N_3644,N_2739);
nor U5314 (N_5314,N_2044,N_2035);
and U5315 (N_5315,N_3415,N_3398);
or U5316 (N_5316,N_3019,N_2869);
and U5317 (N_5317,N_2357,N_2085);
nand U5318 (N_5318,N_2412,N_3626);
xor U5319 (N_5319,N_2298,N_2182);
nand U5320 (N_5320,N_2525,N_2826);
xnor U5321 (N_5321,N_2537,N_3758);
and U5322 (N_5322,N_2140,N_2584);
and U5323 (N_5323,N_2023,N_2321);
and U5324 (N_5324,N_3453,N_2046);
nand U5325 (N_5325,N_3281,N_3655);
and U5326 (N_5326,N_3122,N_2606);
and U5327 (N_5327,N_3023,N_2061);
xnor U5328 (N_5328,N_3868,N_3953);
and U5329 (N_5329,N_3805,N_2281);
and U5330 (N_5330,N_2291,N_2123);
nand U5331 (N_5331,N_2880,N_3209);
and U5332 (N_5332,N_3809,N_2816);
nand U5333 (N_5333,N_2948,N_3026);
and U5334 (N_5334,N_3422,N_3472);
xor U5335 (N_5335,N_3800,N_3132);
xnor U5336 (N_5336,N_3456,N_2720);
xor U5337 (N_5337,N_3985,N_3340);
or U5338 (N_5338,N_2900,N_2409);
or U5339 (N_5339,N_3199,N_3140);
nor U5340 (N_5340,N_2753,N_2613);
nor U5341 (N_5341,N_2211,N_2582);
and U5342 (N_5342,N_2250,N_2547);
nor U5343 (N_5343,N_2723,N_3930);
xnor U5344 (N_5344,N_3550,N_2040);
nand U5345 (N_5345,N_3092,N_2673);
or U5346 (N_5346,N_3582,N_2705);
nand U5347 (N_5347,N_3779,N_3965);
nand U5348 (N_5348,N_2668,N_2667);
nand U5349 (N_5349,N_2379,N_3685);
xor U5350 (N_5350,N_2577,N_3971);
nor U5351 (N_5351,N_3245,N_2786);
or U5352 (N_5352,N_2721,N_3808);
nand U5353 (N_5353,N_2136,N_3670);
xor U5354 (N_5354,N_2957,N_2148);
nor U5355 (N_5355,N_3558,N_3589);
nor U5356 (N_5356,N_3194,N_2199);
xnor U5357 (N_5357,N_2311,N_2844);
nor U5358 (N_5358,N_3122,N_3363);
nor U5359 (N_5359,N_2605,N_2277);
or U5360 (N_5360,N_3835,N_3301);
nor U5361 (N_5361,N_2149,N_2392);
or U5362 (N_5362,N_3754,N_2599);
nand U5363 (N_5363,N_3172,N_3951);
nand U5364 (N_5364,N_2354,N_3209);
and U5365 (N_5365,N_3514,N_2465);
nor U5366 (N_5366,N_3231,N_2872);
nand U5367 (N_5367,N_2262,N_2347);
nand U5368 (N_5368,N_2274,N_3505);
xor U5369 (N_5369,N_3965,N_2637);
nand U5370 (N_5370,N_3977,N_2953);
xnor U5371 (N_5371,N_3631,N_3439);
xor U5372 (N_5372,N_3479,N_3107);
nand U5373 (N_5373,N_2463,N_3591);
or U5374 (N_5374,N_2645,N_2963);
xnor U5375 (N_5375,N_3154,N_3959);
nor U5376 (N_5376,N_3468,N_3622);
nand U5377 (N_5377,N_3272,N_3596);
xor U5378 (N_5378,N_2667,N_2698);
nor U5379 (N_5379,N_3614,N_3903);
nor U5380 (N_5380,N_3105,N_2304);
and U5381 (N_5381,N_3013,N_3719);
xor U5382 (N_5382,N_3408,N_2282);
nor U5383 (N_5383,N_2926,N_3158);
nand U5384 (N_5384,N_2930,N_2587);
nor U5385 (N_5385,N_3465,N_3786);
nor U5386 (N_5386,N_2524,N_2450);
nor U5387 (N_5387,N_3718,N_3375);
nand U5388 (N_5388,N_2275,N_3460);
xnor U5389 (N_5389,N_2796,N_3465);
nand U5390 (N_5390,N_3996,N_2920);
nand U5391 (N_5391,N_3573,N_3206);
or U5392 (N_5392,N_3849,N_3510);
or U5393 (N_5393,N_3635,N_2946);
and U5394 (N_5394,N_3767,N_3216);
and U5395 (N_5395,N_2274,N_2839);
nor U5396 (N_5396,N_2040,N_2163);
and U5397 (N_5397,N_3511,N_2722);
xor U5398 (N_5398,N_2777,N_2302);
and U5399 (N_5399,N_2227,N_3617);
or U5400 (N_5400,N_2223,N_2399);
and U5401 (N_5401,N_3107,N_2944);
or U5402 (N_5402,N_3405,N_3083);
nand U5403 (N_5403,N_2952,N_3374);
nor U5404 (N_5404,N_3650,N_3906);
or U5405 (N_5405,N_2980,N_3309);
and U5406 (N_5406,N_3266,N_3441);
nor U5407 (N_5407,N_2865,N_2060);
nand U5408 (N_5408,N_3445,N_3494);
or U5409 (N_5409,N_2005,N_3598);
nand U5410 (N_5410,N_2356,N_3859);
or U5411 (N_5411,N_2434,N_3584);
nor U5412 (N_5412,N_3511,N_2283);
nor U5413 (N_5413,N_2688,N_3024);
nand U5414 (N_5414,N_2732,N_3478);
or U5415 (N_5415,N_2887,N_2222);
or U5416 (N_5416,N_2628,N_3089);
nand U5417 (N_5417,N_2596,N_3530);
nor U5418 (N_5418,N_2898,N_2893);
nor U5419 (N_5419,N_3505,N_2765);
nor U5420 (N_5420,N_3373,N_2964);
or U5421 (N_5421,N_2731,N_3964);
and U5422 (N_5422,N_2807,N_3417);
or U5423 (N_5423,N_3449,N_3442);
and U5424 (N_5424,N_2133,N_2663);
and U5425 (N_5425,N_3687,N_2800);
nand U5426 (N_5426,N_2201,N_3171);
nor U5427 (N_5427,N_3550,N_3767);
nand U5428 (N_5428,N_3095,N_3164);
and U5429 (N_5429,N_2850,N_3200);
nor U5430 (N_5430,N_3304,N_3474);
and U5431 (N_5431,N_2772,N_3709);
and U5432 (N_5432,N_3222,N_2738);
nor U5433 (N_5433,N_2631,N_3202);
or U5434 (N_5434,N_3752,N_2010);
nand U5435 (N_5435,N_3879,N_2737);
nand U5436 (N_5436,N_3335,N_2207);
and U5437 (N_5437,N_3051,N_2202);
or U5438 (N_5438,N_3880,N_3330);
xnor U5439 (N_5439,N_3344,N_2121);
and U5440 (N_5440,N_2987,N_3696);
nand U5441 (N_5441,N_2802,N_3292);
xnor U5442 (N_5442,N_2401,N_3009);
xor U5443 (N_5443,N_3103,N_2114);
nand U5444 (N_5444,N_3777,N_3357);
and U5445 (N_5445,N_3915,N_3937);
or U5446 (N_5446,N_3089,N_2741);
and U5447 (N_5447,N_2242,N_2248);
or U5448 (N_5448,N_2005,N_3675);
xnor U5449 (N_5449,N_2497,N_3704);
xnor U5450 (N_5450,N_3661,N_2220);
and U5451 (N_5451,N_2018,N_3454);
and U5452 (N_5452,N_3160,N_2714);
and U5453 (N_5453,N_2494,N_3375);
nand U5454 (N_5454,N_2486,N_2997);
nor U5455 (N_5455,N_3316,N_2252);
nor U5456 (N_5456,N_2971,N_2323);
xnor U5457 (N_5457,N_3396,N_3567);
nor U5458 (N_5458,N_3026,N_2047);
or U5459 (N_5459,N_3065,N_3625);
nand U5460 (N_5460,N_3832,N_3909);
or U5461 (N_5461,N_2766,N_3868);
and U5462 (N_5462,N_3405,N_3221);
and U5463 (N_5463,N_3169,N_2943);
nand U5464 (N_5464,N_3148,N_3501);
nor U5465 (N_5465,N_2436,N_2779);
and U5466 (N_5466,N_2143,N_3100);
nand U5467 (N_5467,N_2564,N_2871);
and U5468 (N_5468,N_2608,N_2174);
nand U5469 (N_5469,N_2821,N_2958);
nor U5470 (N_5470,N_2181,N_3634);
nand U5471 (N_5471,N_2394,N_3860);
nand U5472 (N_5472,N_3936,N_2716);
and U5473 (N_5473,N_2971,N_2212);
xor U5474 (N_5474,N_2421,N_3644);
nor U5475 (N_5475,N_3740,N_2926);
and U5476 (N_5476,N_2184,N_2698);
nor U5477 (N_5477,N_3202,N_2123);
nand U5478 (N_5478,N_2752,N_2265);
and U5479 (N_5479,N_2504,N_3419);
nand U5480 (N_5480,N_2027,N_3740);
xor U5481 (N_5481,N_3247,N_2716);
nand U5482 (N_5482,N_2935,N_2088);
nand U5483 (N_5483,N_3924,N_2534);
nor U5484 (N_5484,N_2881,N_2296);
nand U5485 (N_5485,N_3763,N_3426);
xnor U5486 (N_5486,N_3627,N_2644);
nand U5487 (N_5487,N_2822,N_2588);
or U5488 (N_5488,N_2860,N_2177);
and U5489 (N_5489,N_3230,N_3309);
xor U5490 (N_5490,N_3176,N_2593);
and U5491 (N_5491,N_3529,N_3892);
nand U5492 (N_5492,N_2395,N_3545);
nor U5493 (N_5493,N_2646,N_2556);
nor U5494 (N_5494,N_3845,N_3932);
xor U5495 (N_5495,N_2211,N_3722);
xnor U5496 (N_5496,N_3121,N_3590);
xnor U5497 (N_5497,N_2528,N_2167);
or U5498 (N_5498,N_3082,N_3214);
and U5499 (N_5499,N_3552,N_3325);
xnor U5500 (N_5500,N_3663,N_3177);
xnor U5501 (N_5501,N_2135,N_2025);
nor U5502 (N_5502,N_2077,N_2205);
xor U5503 (N_5503,N_2883,N_2876);
or U5504 (N_5504,N_2668,N_2270);
or U5505 (N_5505,N_3855,N_3901);
or U5506 (N_5506,N_2088,N_2339);
and U5507 (N_5507,N_2313,N_2146);
or U5508 (N_5508,N_3064,N_3501);
nand U5509 (N_5509,N_3008,N_2631);
xor U5510 (N_5510,N_2053,N_2141);
or U5511 (N_5511,N_3885,N_3340);
or U5512 (N_5512,N_2673,N_3783);
nand U5513 (N_5513,N_2071,N_2723);
nor U5514 (N_5514,N_3755,N_2783);
nor U5515 (N_5515,N_2728,N_2760);
nor U5516 (N_5516,N_2873,N_2065);
xnor U5517 (N_5517,N_3021,N_2046);
or U5518 (N_5518,N_2794,N_2740);
nand U5519 (N_5519,N_3942,N_2479);
and U5520 (N_5520,N_2239,N_3938);
or U5521 (N_5521,N_3902,N_2856);
nand U5522 (N_5522,N_3470,N_3015);
or U5523 (N_5523,N_2614,N_2947);
and U5524 (N_5524,N_2371,N_2111);
or U5525 (N_5525,N_2123,N_2183);
and U5526 (N_5526,N_3512,N_3606);
xor U5527 (N_5527,N_2892,N_3956);
and U5528 (N_5528,N_3194,N_2837);
nor U5529 (N_5529,N_2338,N_3034);
xor U5530 (N_5530,N_2224,N_2949);
or U5531 (N_5531,N_2634,N_3749);
or U5532 (N_5532,N_2768,N_2535);
nor U5533 (N_5533,N_3363,N_3877);
nand U5534 (N_5534,N_3359,N_3672);
nor U5535 (N_5535,N_2065,N_2059);
nor U5536 (N_5536,N_2982,N_3098);
xor U5537 (N_5537,N_3492,N_3389);
nand U5538 (N_5538,N_2819,N_3598);
and U5539 (N_5539,N_3582,N_3231);
xnor U5540 (N_5540,N_2207,N_3489);
xor U5541 (N_5541,N_2389,N_2928);
xor U5542 (N_5542,N_3488,N_3926);
xor U5543 (N_5543,N_2865,N_3387);
nand U5544 (N_5544,N_2155,N_3138);
xnor U5545 (N_5545,N_2125,N_3927);
and U5546 (N_5546,N_2395,N_2166);
xor U5547 (N_5547,N_3381,N_2380);
and U5548 (N_5548,N_2789,N_3682);
nor U5549 (N_5549,N_3818,N_2109);
or U5550 (N_5550,N_3229,N_2946);
or U5551 (N_5551,N_3793,N_3285);
nand U5552 (N_5552,N_2935,N_3688);
nor U5553 (N_5553,N_2737,N_3591);
xor U5554 (N_5554,N_3952,N_3717);
nand U5555 (N_5555,N_2696,N_2005);
or U5556 (N_5556,N_3650,N_2923);
or U5557 (N_5557,N_2470,N_2743);
nor U5558 (N_5558,N_3299,N_2055);
nand U5559 (N_5559,N_2924,N_3340);
nor U5560 (N_5560,N_3487,N_3218);
nand U5561 (N_5561,N_3117,N_3671);
or U5562 (N_5562,N_3768,N_2554);
xor U5563 (N_5563,N_3760,N_2424);
and U5564 (N_5564,N_3684,N_3425);
or U5565 (N_5565,N_3746,N_3932);
and U5566 (N_5566,N_3682,N_3766);
xnor U5567 (N_5567,N_3404,N_2301);
nor U5568 (N_5568,N_2428,N_3195);
nor U5569 (N_5569,N_2680,N_3180);
xor U5570 (N_5570,N_2254,N_3470);
or U5571 (N_5571,N_3252,N_3319);
and U5572 (N_5572,N_3854,N_2250);
nand U5573 (N_5573,N_2990,N_2296);
nand U5574 (N_5574,N_3121,N_3214);
or U5575 (N_5575,N_3888,N_2790);
or U5576 (N_5576,N_3649,N_2007);
nor U5577 (N_5577,N_2726,N_3450);
nor U5578 (N_5578,N_3709,N_2691);
xor U5579 (N_5579,N_3495,N_2813);
or U5580 (N_5580,N_3916,N_3872);
xnor U5581 (N_5581,N_2069,N_3705);
nor U5582 (N_5582,N_2952,N_3721);
or U5583 (N_5583,N_2321,N_3204);
nor U5584 (N_5584,N_3882,N_2850);
xor U5585 (N_5585,N_3238,N_3166);
xor U5586 (N_5586,N_2075,N_3894);
xnor U5587 (N_5587,N_2579,N_3145);
and U5588 (N_5588,N_3457,N_2480);
xnor U5589 (N_5589,N_2269,N_2156);
nor U5590 (N_5590,N_3766,N_2710);
nand U5591 (N_5591,N_2855,N_2135);
nor U5592 (N_5592,N_3352,N_2277);
or U5593 (N_5593,N_3841,N_2190);
nand U5594 (N_5594,N_2927,N_3728);
or U5595 (N_5595,N_2598,N_3092);
and U5596 (N_5596,N_2339,N_3781);
nor U5597 (N_5597,N_3481,N_3989);
xor U5598 (N_5598,N_2065,N_2908);
and U5599 (N_5599,N_2182,N_3797);
xor U5600 (N_5600,N_2565,N_2163);
nor U5601 (N_5601,N_2883,N_2556);
or U5602 (N_5602,N_2467,N_2877);
nor U5603 (N_5603,N_3577,N_3963);
nand U5604 (N_5604,N_3958,N_3609);
and U5605 (N_5605,N_3365,N_2315);
or U5606 (N_5606,N_3825,N_3669);
or U5607 (N_5607,N_2083,N_2495);
nor U5608 (N_5608,N_2374,N_3055);
xnor U5609 (N_5609,N_3080,N_3297);
nor U5610 (N_5610,N_2989,N_3009);
nor U5611 (N_5611,N_3060,N_2846);
nor U5612 (N_5612,N_2682,N_3163);
or U5613 (N_5613,N_2390,N_2366);
nand U5614 (N_5614,N_3074,N_2031);
and U5615 (N_5615,N_3643,N_2914);
or U5616 (N_5616,N_3915,N_3935);
nor U5617 (N_5617,N_3010,N_3039);
nand U5618 (N_5618,N_2325,N_2087);
nand U5619 (N_5619,N_3731,N_3870);
nor U5620 (N_5620,N_3119,N_2994);
or U5621 (N_5621,N_2541,N_3193);
xor U5622 (N_5622,N_2920,N_3260);
nor U5623 (N_5623,N_2818,N_3309);
and U5624 (N_5624,N_3818,N_2274);
nor U5625 (N_5625,N_2767,N_3789);
xnor U5626 (N_5626,N_2297,N_3634);
nor U5627 (N_5627,N_3481,N_3124);
nor U5628 (N_5628,N_3616,N_2610);
or U5629 (N_5629,N_2683,N_3778);
nand U5630 (N_5630,N_2036,N_2661);
nand U5631 (N_5631,N_3316,N_2941);
and U5632 (N_5632,N_2974,N_3022);
xnor U5633 (N_5633,N_3560,N_2239);
nor U5634 (N_5634,N_2097,N_2475);
and U5635 (N_5635,N_2526,N_3191);
nor U5636 (N_5636,N_3484,N_2175);
nor U5637 (N_5637,N_3174,N_2729);
nand U5638 (N_5638,N_3332,N_3113);
nand U5639 (N_5639,N_3546,N_2995);
nand U5640 (N_5640,N_3066,N_3456);
nand U5641 (N_5641,N_3322,N_3752);
or U5642 (N_5642,N_3640,N_2083);
xnor U5643 (N_5643,N_2067,N_3444);
nor U5644 (N_5644,N_2281,N_3993);
and U5645 (N_5645,N_2400,N_3854);
xor U5646 (N_5646,N_2426,N_3153);
or U5647 (N_5647,N_2850,N_3725);
nor U5648 (N_5648,N_3731,N_2188);
and U5649 (N_5649,N_3085,N_3842);
nor U5650 (N_5650,N_3679,N_2850);
nand U5651 (N_5651,N_3879,N_3676);
xor U5652 (N_5652,N_3419,N_2907);
xnor U5653 (N_5653,N_3737,N_2446);
or U5654 (N_5654,N_2884,N_3614);
nand U5655 (N_5655,N_3211,N_2250);
or U5656 (N_5656,N_2248,N_2285);
and U5657 (N_5657,N_3594,N_3646);
xnor U5658 (N_5658,N_3339,N_3376);
nand U5659 (N_5659,N_2558,N_3053);
nor U5660 (N_5660,N_2918,N_3797);
xor U5661 (N_5661,N_3478,N_3278);
nand U5662 (N_5662,N_2782,N_3413);
xor U5663 (N_5663,N_2784,N_3220);
and U5664 (N_5664,N_2106,N_2336);
or U5665 (N_5665,N_2830,N_2285);
and U5666 (N_5666,N_3716,N_3254);
and U5667 (N_5667,N_2232,N_3496);
or U5668 (N_5668,N_3616,N_3031);
nand U5669 (N_5669,N_3520,N_2104);
and U5670 (N_5670,N_2747,N_3838);
nor U5671 (N_5671,N_2192,N_3910);
or U5672 (N_5672,N_3906,N_2467);
and U5673 (N_5673,N_3004,N_2232);
xor U5674 (N_5674,N_2496,N_2777);
xor U5675 (N_5675,N_3047,N_3251);
or U5676 (N_5676,N_3526,N_2719);
or U5677 (N_5677,N_3398,N_3250);
nand U5678 (N_5678,N_2058,N_3699);
xnor U5679 (N_5679,N_2418,N_2141);
nor U5680 (N_5680,N_3609,N_3205);
nand U5681 (N_5681,N_3017,N_3249);
xnor U5682 (N_5682,N_2689,N_2534);
xnor U5683 (N_5683,N_2646,N_3480);
xnor U5684 (N_5684,N_2515,N_3423);
and U5685 (N_5685,N_2929,N_3981);
nor U5686 (N_5686,N_2747,N_2841);
or U5687 (N_5687,N_3554,N_3236);
and U5688 (N_5688,N_3429,N_2768);
nor U5689 (N_5689,N_2720,N_3222);
nand U5690 (N_5690,N_3096,N_2631);
nor U5691 (N_5691,N_2567,N_2225);
nor U5692 (N_5692,N_3907,N_2547);
xor U5693 (N_5693,N_2740,N_3567);
nand U5694 (N_5694,N_2095,N_2447);
nand U5695 (N_5695,N_3476,N_2820);
xor U5696 (N_5696,N_2028,N_3312);
and U5697 (N_5697,N_3639,N_3303);
or U5698 (N_5698,N_3006,N_2965);
nor U5699 (N_5699,N_2807,N_2824);
and U5700 (N_5700,N_2966,N_3295);
xor U5701 (N_5701,N_2097,N_3390);
nand U5702 (N_5702,N_3931,N_3954);
or U5703 (N_5703,N_2589,N_3918);
xnor U5704 (N_5704,N_3254,N_2789);
or U5705 (N_5705,N_2195,N_2164);
nor U5706 (N_5706,N_3725,N_2992);
nand U5707 (N_5707,N_2517,N_3867);
xor U5708 (N_5708,N_2617,N_2852);
nand U5709 (N_5709,N_2796,N_2176);
nor U5710 (N_5710,N_3864,N_2664);
or U5711 (N_5711,N_3073,N_2962);
nor U5712 (N_5712,N_3431,N_2012);
or U5713 (N_5713,N_3480,N_3733);
xor U5714 (N_5714,N_2721,N_3066);
nand U5715 (N_5715,N_3060,N_3147);
and U5716 (N_5716,N_3151,N_3451);
and U5717 (N_5717,N_3289,N_2163);
or U5718 (N_5718,N_3346,N_2094);
nand U5719 (N_5719,N_3068,N_3308);
and U5720 (N_5720,N_3634,N_2626);
nor U5721 (N_5721,N_3314,N_2045);
nand U5722 (N_5722,N_2224,N_3966);
or U5723 (N_5723,N_2055,N_2123);
nand U5724 (N_5724,N_3672,N_2079);
nand U5725 (N_5725,N_2265,N_3765);
nand U5726 (N_5726,N_2388,N_3185);
or U5727 (N_5727,N_2378,N_2882);
xnor U5728 (N_5728,N_2260,N_2130);
xor U5729 (N_5729,N_3859,N_3721);
and U5730 (N_5730,N_3870,N_3920);
xnor U5731 (N_5731,N_2576,N_2227);
or U5732 (N_5732,N_2893,N_3683);
or U5733 (N_5733,N_2753,N_2115);
or U5734 (N_5734,N_2091,N_2067);
nand U5735 (N_5735,N_2818,N_2756);
xor U5736 (N_5736,N_3012,N_3133);
xor U5737 (N_5737,N_2691,N_3125);
and U5738 (N_5738,N_3384,N_2374);
or U5739 (N_5739,N_3455,N_2863);
nand U5740 (N_5740,N_3135,N_3905);
or U5741 (N_5741,N_2188,N_3134);
xnor U5742 (N_5742,N_2429,N_2909);
nor U5743 (N_5743,N_2467,N_2603);
and U5744 (N_5744,N_2563,N_2333);
and U5745 (N_5745,N_2556,N_2607);
or U5746 (N_5746,N_2875,N_2425);
xor U5747 (N_5747,N_3367,N_2836);
and U5748 (N_5748,N_3681,N_2089);
or U5749 (N_5749,N_3723,N_2999);
nor U5750 (N_5750,N_3179,N_3762);
nor U5751 (N_5751,N_2928,N_3266);
and U5752 (N_5752,N_3084,N_3592);
or U5753 (N_5753,N_3701,N_3955);
nand U5754 (N_5754,N_3929,N_3384);
xor U5755 (N_5755,N_3452,N_2669);
and U5756 (N_5756,N_3119,N_2007);
nand U5757 (N_5757,N_2818,N_2237);
and U5758 (N_5758,N_3338,N_2401);
and U5759 (N_5759,N_3449,N_3797);
or U5760 (N_5760,N_2738,N_3836);
nor U5761 (N_5761,N_2666,N_3507);
and U5762 (N_5762,N_3676,N_3413);
nor U5763 (N_5763,N_3684,N_3717);
xnor U5764 (N_5764,N_2422,N_3204);
and U5765 (N_5765,N_3841,N_2859);
xnor U5766 (N_5766,N_2495,N_2561);
nor U5767 (N_5767,N_3791,N_3010);
xnor U5768 (N_5768,N_2639,N_2833);
xnor U5769 (N_5769,N_2888,N_3091);
nor U5770 (N_5770,N_2666,N_2719);
xnor U5771 (N_5771,N_3287,N_3823);
xor U5772 (N_5772,N_3670,N_2516);
and U5773 (N_5773,N_3677,N_3401);
or U5774 (N_5774,N_3307,N_2164);
and U5775 (N_5775,N_3434,N_2077);
or U5776 (N_5776,N_2249,N_2039);
nand U5777 (N_5777,N_3396,N_3478);
nand U5778 (N_5778,N_2897,N_3575);
xor U5779 (N_5779,N_2859,N_2128);
nand U5780 (N_5780,N_2785,N_3852);
or U5781 (N_5781,N_3186,N_3961);
xor U5782 (N_5782,N_3682,N_2359);
nor U5783 (N_5783,N_2703,N_2764);
nand U5784 (N_5784,N_3124,N_2419);
and U5785 (N_5785,N_3460,N_2883);
and U5786 (N_5786,N_3398,N_3101);
nand U5787 (N_5787,N_2716,N_3519);
xnor U5788 (N_5788,N_2985,N_3535);
and U5789 (N_5789,N_2740,N_2081);
and U5790 (N_5790,N_3365,N_3487);
xor U5791 (N_5791,N_3962,N_3507);
nor U5792 (N_5792,N_3879,N_3896);
and U5793 (N_5793,N_2730,N_3973);
nand U5794 (N_5794,N_2363,N_3564);
xor U5795 (N_5795,N_2901,N_2302);
nor U5796 (N_5796,N_2803,N_3425);
nand U5797 (N_5797,N_2385,N_3237);
xnor U5798 (N_5798,N_3939,N_2056);
and U5799 (N_5799,N_2655,N_2764);
nand U5800 (N_5800,N_3664,N_2731);
and U5801 (N_5801,N_3018,N_3148);
and U5802 (N_5802,N_2482,N_3798);
nor U5803 (N_5803,N_2693,N_2713);
nor U5804 (N_5804,N_2547,N_2278);
or U5805 (N_5805,N_2937,N_3799);
nor U5806 (N_5806,N_3827,N_3926);
or U5807 (N_5807,N_2300,N_3516);
nand U5808 (N_5808,N_3524,N_3451);
or U5809 (N_5809,N_3690,N_2981);
nor U5810 (N_5810,N_3673,N_3283);
xor U5811 (N_5811,N_3534,N_3742);
xnor U5812 (N_5812,N_2059,N_3231);
or U5813 (N_5813,N_3978,N_3613);
xnor U5814 (N_5814,N_2273,N_2633);
or U5815 (N_5815,N_3138,N_3207);
or U5816 (N_5816,N_3879,N_2027);
and U5817 (N_5817,N_2146,N_2743);
xor U5818 (N_5818,N_3033,N_2165);
nand U5819 (N_5819,N_3837,N_2233);
and U5820 (N_5820,N_3708,N_3382);
nor U5821 (N_5821,N_3388,N_2158);
nor U5822 (N_5822,N_3781,N_3040);
xor U5823 (N_5823,N_2156,N_3866);
nor U5824 (N_5824,N_3185,N_2959);
nand U5825 (N_5825,N_2342,N_3947);
or U5826 (N_5826,N_2573,N_2485);
nor U5827 (N_5827,N_2566,N_3570);
xor U5828 (N_5828,N_3053,N_2674);
nand U5829 (N_5829,N_3727,N_2060);
or U5830 (N_5830,N_3863,N_2056);
or U5831 (N_5831,N_3081,N_2983);
or U5832 (N_5832,N_3393,N_2592);
nor U5833 (N_5833,N_2017,N_2608);
nor U5834 (N_5834,N_2679,N_3183);
nand U5835 (N_5835,N_2034,N_3955);
or U5836 (N_5836,N_2869,N_2098);
and U5837 (N_5837,N_2092,N_3958);
or U5838 (N_5838,N_3618,N_2704);
xor U5839 (N_5839,N_2011,N_3033);
nand U5840 (N_5840,N_3870,N_3136);
nand U5841 (N_5841,N_2354,N_2766);
xor U5842 (N_5842,N_2532,N_2189);
nor U5843 (N_5843,N_2352,N_2511);
xor U5844 (N_5844,N_3955,N_3049);
or U5845 (N_5845,N_2343,N_3521);
nor U5846 (N_5846,N_2430,N_3400);
nand U5847 (N_5847,N_3966,N_2115);
nor U5848 (N_5848,N_3504,N_2998);
nor U5849 (N_5849,N_2229,N_2349);
xor U5850 (N_5850,N_2840,N_3348);
xor U5851 (N_5851,N_3929,N_2916);
nor U5852 (N_5852,N_3507,N_2453);
or U5853 (N_5853,N_3650,N_3959);
and U5854 (N_5854,N_2731,N_3146);
nor U5855 (N_5855,N_3730,N_2668);
xnor U5856 (N_5856,N_2152,N_3240);
xnor U5857 (N_5857,N_3382,N_3004);
nor U5858 (N_5858,N_3820,N_3520);
or U5859 (N_5859,N_3953,N_2626);
nor U5860 (N_5860,N_3896,N_3080);
or U5861 (N_5861,N_2891,N_3689);
nand U5862 (N_5862,N_3823,N_3857);
nand U5863 (N_5863,N_3072,N_2597);
or U5864 (N_5864,N_3673,N_2991);
nor U5865 (N_5865,N_3766,N_3801);
or U5866 (N_5866,N_3836,N_3809);
xor U5867 (N_5867,N_3166,N_3840);
or U5868 (N_5868,N_2641,N_2628);
xnor U5869 (N_5869,N_3101,N_3676);
or U5870 (N_5870,N_2830,N_2408);
nand U5871 (N_5871,N_2256,N_2482);
or U5872 (N_5872,N_2317,N_2556);
and U5873 (N_5873,N_2053,N_3522);
and U5874 (N_5874,N_2019,N_2389);
xnor U5875 (N_5875,N_3240,N_3671);
xnor U5876 (N_5876,N_2999,N_2573);
xnor U5877 (N_5877,N_3604,N_2854);
or U5878 (N_5878,N_2440,N_2848);
xnor U5879 (N_5879,N_2896,N_3110);
and U5880 (N_5880,N_2724,N_3171);
nand U5881 (N_5881,N_2684,N_2200);
nor U5882 (N_5882,N_2249,N_2709);
or U5883 (N_5883,N_2605,N_3291);
nor U5884 (N_5884,N_3936,N_3621);
nor U5885 (N_5885,N_2369,N_3092);
or U5886 (N_5886,N_2735,N_2504);
nor U5887 (N_5887,N_3655,N_2184);
or U5888 (N_5888,N_3737,N_3065);
xor U5889 (N_5889,N_3722,N_3678);
and U5890 (N_5890,N_3258,N_3941);
nand U5891 (N_5891,N_2321,N_2194);
and U5892 (N_5892,N_3460,N_3256);
xnor U5893 (N_5893,N_2567,N_2747);
xor U5894 (N_5894,N_3292,N_2447);
xor U5895 (N_5895,N_3310,N_3300);
or U5896 (N_5896,N_3549,N_3161);
nand U5897 (N_5897,N_3139,N_2122);
nand U5898 (N_5898,N_2959,N_3292);
and U5899 (N_5899,N_2906,N_3590);
nor U5900 (N_5900,N_2189,N_3582);
xnor U5901 (N_5901,N_3446,N_3823);
nor U5902 (N_5902,N_3865,N_2677);
or U5903 (N_5903,N_2676,N_2379);
or U5904 (N_5904,N_2007,N_3491);
or U5905 (N_5905,N_3589,N_2463);
or U5906 (N_5906,N_2882,N_3252);
xor U5907 (N_5907,N_3592,N_2535);
or U5908 (N_5908,N_3864,N_2657);
nor U5909 (N_5909,N_3425,N_2432);
nand U5910 (N_5910,N_3758,N_2073);
or U5911 (N_5911,N_2538,N_2877);
and U5912 (N_5912,N_3854,N_2901);
and U5913 (N_5913,N_3168,N_2854);
nor U5914 (N_5914,N_2854,N_3522);
nand U5915 (N_5915,N_3071,N_3928);
nor U5916 (N_5916,N_2205,N_3520);
or U5917 (N_5917,N_3071,N_2653);
and U5918 (N_5918,N_2792,N_2004);
or U5919 (N_5919,N_3484,N_2110);
or U5920 (N_5920,N_3273,N_2274);
nand U5921 (N_5921,N_3518,N_3425);
xor U5922 (N_5922,N_2042,N_3737);
nand U5923 (N_5923,N_2111,N_2594);
and U5924 (N_5924,N_3608,N_2361);
or U5925 (N_5925,N_3227,N_3250);
xnor U5926 (N_5926,N_2830,N_2689);
nand U5927 (N_5927,N_2426,N_3985);
xor U5928 (N_5928,N_2323,N_2283);
xnor U5929 (N_5929,N_2471,N_3137);
nor U5930 (N_5930,N_3107,N_2209);
nand U5931 (N_5931,N_2711,N_2152);
nor U5932 (N_5932,N_2483,N_2717);
xor U5933 (N_5933,N_2838,N_3525);
and U5934 (N_5934,N_2766,N_2914);
and U5935 (N_5935,N_3130,N_3461);
xnor U5936 (N_5936,N_2696,N_3101);
nor U5937 (N_5937,N_2672,N_3562);
or U5938 (N_5938,N_3865,N_3348);
or U5939 (N_5939,N_2226,N_3833);
xor U5940 (N_5940,N_2755,N_3030);
or U5941 (N_5941,N_2511,N_2985);
nand U5942 (N_5942,N_2313,N_2874);
xor U5943 (N_5943,N_2058,N_2836);
xor U5944 (N_5944,N_2431,N_3117);
xnor U5945 (N_5945,N_2335,N_2072);
nand U5946 (N_5946,N_2333,N_3638);
or U5947 (N_5947,N_2447,N_3481);
nand U5948 (N_5948,N_2441,N_2350);
and U5949 (N_5949,N_3481,N_2449);
xnor U5950 (N_5950,N_2607,N_2889);
nand U5951 (N_5951,N_3324,N_2042);
xor U5952 (N_5952,N_3375,N_3122);
xnor U5953 (N_5953,N_3292,N_2594);
and U5954 (N_5954,N_3377,N_2749);
and U5955 (N_5955,N_3019,N_3504);
and U5956 (N_5956,N_3090,N_2851);
or U5957 (N_5957,N_2207,N_3620);
xnor U5958 (N_5958,N_3516,N_2891);
nor U5959 (N_5959,N_2643,N_2670);
nand U5960 (N_5960,N_3891,N_3559);
xor U5961 (N_5961,N_3743,N_2137);
nand U5962 (N_5962,N_2409,N_3888);
nor U5963 (N_5963,N_3468,N_3913);
nor U5964 (N_5964,N_3665,N_3273);
xnor U5965 (N_5965,N_3538,N_2771);
and U5966 (N_5966,N_3840,N_3588);
nor U5967 (N_5967,N_3326,N_3750);
nor U5968 (N_5968,N_2626,N_3823);
nor U5969 (N_5969,N_2640,N_3393);
nand U5970 (N_5970,N_2669,N_2797);
and U5971 (N_5971,N_2302,N_3335);
and U5972 (N_5972,N_2443,N_2559);
and U5973 (N_5973,N_2530,N_2481);
nand U5974 (N_5974,N_2904,N_3528);
xnor U5975 (N_5975,N_3325,N_2565);
xnor U5976 (N_5976,N_3454,N_3322);
xnor U5977 (N_5977,N_3124,N_3955);
nand U5978 (N_5978,N_3565,N_3986);
nor U5979 (N_5979,N_2218,N_2705);
xor U5980 (N_5980,N_3625,N_2859);
and U5981 (N_5981,N_2893,N_2496);
and U5982 (N_5982,N_2150,N_3958);
and U5983 (N_5983,N_3704,N_3592);
and U5984 (N_5984,N_2982,N_3745);
and U5985 (N_5985,N_2932,N_2031);
nand U5986 (N_5986,N_3605,N_2869);
xor U5987 (N_5987,N_3143,N_3579);
or U5988 (N_5988,N_2988,N_2194);
or U5989 (N_5989,N_3885,N_2368);
xor U5990 (N_5990,N_2282,N_2482);
and U5991 (N_5991,N_3150,N_3923);
xnor U5992 (N_5992,N_3891,N_3597);
nand U5993 (N_5993,N_2755,N_3839);
or U5994 (N_5994,N_2472,N_3571);
nand U5995 (N_5995,N_3610,N_3945);
or U5996 (N_5996,N_3676,N_2877);
nand U5997 (N_5997,N_2328,N_2384);
and U5998 (N_5998,N_2664,N_2726);
nor U5999 (N_5999,N_3871,N_3651);
and U6000 (N_6000,N_5730,N_5128);
nor U6001 (N_6001,N_4878,N_5957);
nand U6002 (N_6002,N_4879,N_5211);
xor U6003 (N_6003,N_4714,N_5398);
or U6004 (N_6004,N_4024,N_4884);
and U6005 (N_6005,N_5636,N_5772);
or U6006 (N_6006,N_5980,N_5659);
xnor U6007 (N_6007,N_5131,N_4314);
nor U6008 (N_6008,N_4982,N_5439);
nand U6009 (N_6009,N_5074,N_4711);
nor U6010 (N_6010,N_4703,N_5991);
or U6011 (N_6011,N_4874,N_5195);
and U6012 (N_6012,N_4926,N_4281);
nor U6013 (N_6013,N_5129,N_5606);
xnor U6014 (N_6014,N_4981,N_4073);
nor U6015 (N_6015,N_5075,N_4306);
nor U6016 (N_6016,N_5565,N_4352);
nand U6017 (N_6017,N_5603,N_5831);
or U6018 (N_6018,N_4244,N_4038);
xnor U6019 (N_6019,N_4691,N_5599);
nand U6020 (N_6020,N_4374,N_5043);
nor U6021 (N_6021,N_5276,N_4030);
nand U6022 (N_6022,N_4622,N_5016);
or U6023 (N_6023,N_5001,N_5975);
or U6024 (N_6024,N_4354,N_4415);
nor U6025 (N_6025,N_5178,N_4147);
or U6026 (N_6026,N_5568,N_5271);
nor U6027 (N_6027,N_5623,N_5548);
xnor U6028 (N_6028,N_4126,N_4284);
nand U6029 (N_6029,N_5572,N_4364);
nand U6030 (N_6030,N_5589,N_5169);
nand U6031 (N_6031,N_5620,N_4905);
nor U6032 (N_6032,N_4370,N_4097);
xnor U6033 (N_6033,N_4846,N_4280);
or U6034 (N_6034,N_4270,N_4952);
or U6035 (N_6035,N_5146,N_4810);
xnor U6036 (N_6036,N_5172,N_5305);
nand U6037 (N_6037,N_5929,N_5750);
or U6038 (N_6038,N_5301,N_4074);
and U6039 (N_6039,N_4474,N_4532);
nor U6040 (N_6040,N_4588,N_4529);
nor U6041 (N_6041,N_5449,N_5539);
or U6042 (N_6042,N_5463,N_5840);
or U6043 (N_6043,N_4423,N_4004);
or U6044 (N_6044,N_5933,N_5186);
or U6045 (N_6045,N_4720,N_5518);
or U6046 (N_6046,N_5820,N_5564);
and U6047 (N_6047,N_5291,N_5734);
or U6048 (N_6048,N_5235,N_5685);
and U6049 (N_6049,N_4402,N_4142);
and U6050 (N_6050,N_5934,N_4484);
and U6051 (N_6051,N_5000,N_4184);
or U6052 (N_6052,N_5237,N_5132);
and U6053 (N_6053,N_5837,N_5220);
and U6054 (N_6054,N_4885,N_4632);
or U6055 (N_6055,N_4642,N_5756);
xnor U6056 (N_6056,N_5344,N_4022);
nor U6057 (N_6057,N_5771,N_4338);
xor U6058 (N_6058,N_4158,N_5650);
or U6059 (N_6059,N_5407,N_5731);
nand U6060 (N_6060,N_4688,N_4823);
or U6061 (N_6061,N_4076,N_5893);
xor U6062 (N_6062,N_5749,N_4503);
and U6063 (N_6063,N_4334,N_4646);
nor U6064 (N_6064,N_5338,N_5020);
xor U6065 (N_6065,N_4072,N_4429);
nor U6066 (N_6066,N_4021,N_5445);
xor U6067 (N_6067,N_5616,N_4909);
nand U6068 (N_6068,N_5224,N_4790);
xor U6069 (N_6069,N_4295,N_4150);
or U6070 (N_6070,N_4335,N_5268);
nor U6071 (N_6071,N_4692,N_5414);
nor U6072 (N_6072,N_4591,N_5423);
xor U6073 (N_6073,N_5948,N_4726);
or U6074 (N_6074,N_4485,N_4685);
nor U6075 (N_6075,N_4657,N_5847);
xor U6076 (N_6076,N_4040,N_5661);
xnor U6077 (N_6077,N_5160,N_4548);
nor U6078 (N_6078,N_5150,N_5262);
and U6079 (N_6079,N_4710,N_4459);
nand U6080 (N_6080,N_4255,N_4820);
xnor U6081 (N_6081,N_5610,N_5144);
xor U6082 (N_6082,N_4995,N_4351);
nor U6083 (N_6083,N_4340,N_5736);
nor U6084 (N_6084,N_5964,N_5993);
nand U6085 (N_6085,N_5508,N_5118);
xnor U6086 (N_6086,N_4294,N_4590);
xor U6087 (N_6087,N_4378,N_4218);
xnor U6088 (N_6088,N_4203,N_5708);
and U6089 (N_6089,N_5514,N_4207);
xor U6090 (N_6090,N_4424,N_4077);
or U6091 (N_6091,N_4835,N_5763);
nand U6092 (N_6092,N_5827,N_4464);
or U6093 (N_6093,N_4491,N_4029);
xnor U6094 (N_6094,N_4736,N_5180);
xnor U6095 (N_6095,N_5381,N_4227);
nor U6096 (N_6096,N_4966,N_5509);
nand U6097 (N_6097,N_4365,N_4265);
xor U6098 (N_6098,N_4621,N_5039);
nand U6099 (N_6099,N_4282,N_4181);
and U6100 (N_6100,N_4213,N_5258);
nand U6101 (N_6101,N_4221,N_5857);
or U6102 (N_6102,N_5096,N_4543);
nor U6103 (N_6103,N_4933,N_4100);
xor U6104 (N_6104,N_5063,N_4141);
and U6105 (N_6105,N_4961,N_5139);
and U6106 (N_6106,N_4858,N_5808);
nor U6107 (N_6107,N_4807,N_4816);
and U6108 (N_6108,N_4558,N_4027);
nand U6109 (N_6109,N_4009,N_5491);
xor U6110 (N_6110,N_5851,N_4974);
and U6111 (N_6111,N_4683,N_4135);
and U6112 (N_6112,N_5212,N_4896);
and U6113 (N_6113,N_4323,N_4036);
nand U6114 (N_6114,N_4535,N_4919);
nand U6115 (N_6115,N_5900,N_5162);
and U6116 (N_6116,N_5037,N_4967);
xor U6117 (N_6117,N_4717,N_5982);
or U6118 (N_6118,N_5351,N_4845);
or U6119 (N_6119,N_5867,N_4048);
xnor U6120 (N_6120,N_5451,N_5115);
nand U6121 (N_6121,N_4894,N_4214);
and U6122 (N_6122,N_5870,N_4388);
nor U6123 (N_6123,N_4748,N_4245);
or U6124 (N_6124,N_5813,N_5773);
nor U6125 (N_6125,N_5926,N_5370);
nand U6126 (N_6126,N_5283,N_4902);
xnor U6127 (N_6127,N_4589,N_5494);
xnor U6128 (N_6128,N_5033,N_4643);
nand U6129 (N_6129,N_4687,N_5322);
xor U6130 (N_6130,N_4507,N_4864);
nor U6131 (N_6131,N_4387,N_4478);
nor U6132 (N_6132,N_4153,N_4442);
xor U6133 (N_6133,N_5923,N_4644);
xor U6134 (N_6134,N_5284,N_5937);
nand U6135 (N_6135,N_4680,N_5009);
and U6136 (N_6136,N_4787,N_4738);
nand U6137 (N_6137,N_4003,N_5368);
nor U6138 (N_6138,N_5595,N_5824);
nand U6139 (N_6139,N_5081,N_5768);
and U6140 (N_6140,N_5170,N_5223);
nand U6141 (N_6141,N_4877,N_4922);
nand U6142 (N_6142,N_5393,N_5350);
xor U6143 (N_6143,N_5878,N_4447);
xor U6144 (N_6144,N_5054,N_5404);
and U6145 (N_6145,N_4479,N_5645);
nand U6146 (N_6146,N_4463,N_5134);
and U6147 (N_6147,N_5739,N_4851);
and U6148 (N_6148,N_4185,N_4421);
nor U6149 (N_6149,N_4121,N_5713);
nor U6150 (N_6150,N_5303,N_4599);
or U6151 (N_6151,N_4825,N_4962);
and U6152 (N_6152,N_5287,N_5727);
nor U6153 (N_6153,N_5361,N_4771);
or U6154 (N_6154,N_4718,N_4705);
and U6155 (N_6155,N_4605,N_4292);
and U6156 (N_6156,N_4530,N_4565);
nor U6157 (N_6157,N_5758,N_4273);
and U6158 (N_6158,N_4347,N_5440);
nand U6159 (N_6159,N_5068,N_4663);
xnor U6160 (N_6160,N_5873,N_5458);
xor U6161 (N_6161,N_4086,N_5903);
xor U6162 (N_6162,N_4899,N_4749);
xnor U6163 (N_6163,N_5688,N_5123);
or U6164 (N_6164,N_5138,N_4192);
and U6165 (N_6165,N_5670,N_5587);
xnor U6166 (N_6166,N_4345,N_4095);
and U6167 (N_6167,N_5437,N_5493);
or U6168 (N_6168,N_5364,N_4719);
and U6169 (N_6169,N_5969,N_5041);
xnor U6170 (N_6170,N_4536,N_5087);
or U6171 (N_6171,N_5108,N_5578);
nand U6172 (N_6172,N_4986,N_5097);
nor U6173 (N_6173,N_4330,N_5540);
or U6174 (N_6174,N_5047,N_5053);
xor U6175 (N_6175,N_5639,N_5002);
or U6176 (N_6176,N_4942,N_4968);
nor U6177 (N_6177,N_5515,N_4163);
and U6178 (N_6178,N_5882,N_5859);
nor U6179 (N_6179,N_5862,N_5183);
xnor U6180 (N_6180,N_4159,N_5455);
and U6181 (N_6181,N_4113,N_5299);
nor U6182 (N_6182,N_4665,N_5298);
nand U6183 (N_6183,N_4827,N_4861);
nor U6184 (N_6184,N_5928,N_5663);
nand U6185 (N_6185,N_4260,N_5924);
xnor U6186 (N_6186,N_5916,N_5409);
or U6187 (N_6187,N_4346,N_4137);
xnor U6188 (N_6188,N_4585,N_4007);
nor U6189 (N_6189,N_4118,N_5692);
nand U6190 (N_6190,N_4540,N_4627);
nor U6191 (N_6191,N_5120,N_4519);
xor U6192 (N_6192,N_5545,N_4993);
or U6193 (N_6193,N_5495,N_5537);
nand U6194 (N_6194,N_5310,N_5532);
nand U6195 (N_6195,N_4286,N_5358);
nor U6196 (N_6196,N_4235,N_4018);
or U6197 (N_6197,N_4015,N_5967);
and U6198 (N_6198,N_4239,N_5754);
nand U6199 (N_6199,N_5861,N_4283);
nand U6200 (N_6200,N_4495,N_4327);
and U6201 (N_6201,N_5555,N_5872);
xor U6202 (N_6202,N_5743,N_4489);
nor U6203 (N_6203,N_4678,N_4984);
nand U6204 (N_6204,N_5046,N_4624);
or U6205 (N_6205,N_4947,N_5959);
nand U6206 (N_6206,N_5216,N_5091);
or U6207 (N_6207,N_5105,N_5441);
nor U6208 (N_6208,N_5275,N_5696);
nand U6209 (N_6209,N_4145,N_5018);
nand U6210 (N_6210,N_4689,N_4668);
and U6211 (N_6211,N_5601,N_5446);
nand U6212 (N_6212,N_5856,N_5420);
nor U6213 (N_6213,N_5333,N_4871);
nor U6214 (N_6214,N_5821,N_5617);
and U6215 (N_6215,N_5678,N_5524);
nor U6216 (N_6216,N_4716,N_4050);
and U6217 (N_6217,N_5148,N_4586);
nor U6218 (N_6218,N_4553,N_5832);
xor U6219 (N_6219,N_4462,N_4840);
nor U6220 (N_6220,N_5230,N_5686);
xor U6221 (N_6221,N_5523,N_5668);
and U6222 (N_6222,N_4037,N_4108);
xor U6223 (N_6223,N_5366,N_4882);
nand U6224 (N_6224,N_5726,N_5811);
xnor U6225 (N_6225,N_4659,N_4469);
or U6226 (N_6226,N_5462,N_5428);
nand U6227 (N_6227,N_4672,N_5533);
and U6228 (N_6228,N_5239,N_4715);
nor U6229 (N_6229,N_5529,N_5931);
nor U6230 (N_6230,N_4602,N_4950);
xnor U6231 (N_6231,N_5411,N_5113);
nand U6232 (N_6232,N_4795,N_5992);
and U6233 (N_6233,N_5839,N_4941);
nor U6234 (N_6234,N_4853,N_5683);
and U6235 (N_6235,N_4082,N_4641);
nor U6236 (N_6236,N_4238,N_5667);
and U6237 (N_6237,N_4348,N_4202);
or U6238 (N_6238,N_4060,N_5644);
nand U6239 (N_6239,N_4729,N_5863);
and U6240 (N_6240,N_4408,N_4569);
nand U6241 (N_6241,N_5430,N_5825);
or U6242 (N_6242,N_5391,N_5191);
nand U6243 (N_6243,N_5202,N_5621);
nor U6244 (N_6244,N_4708,N_4104);
xor U6245 (N_6245,N_4811,N_5674);
nor U6246 (N_6246,N_5835,N_4232);
nor U6247 (N_6247,N_4413,N_5765);
xor U6248 (N_6248,N_5904,N_4985);
and U6249 (N_6249,N_5076,N_4443);
and U6250 (N_6250,N_5100,N_5700);
and U6251 (N_6251,N_5422,N_4386);
xnor U6252 (N_6252,N_4410,N_5340);
xor U6253 (N_6253,N_4005,N_4293);
nand U6254 (N_6254,N_4881,N_4913);
or U6255 (N_6255,N_5226,N_4200);
nand U6256 (N_6256,N_5712,N_4655);
and U6257 (N_6257,N_5999,N_5040);
and U6258 (N_6258,N_4236,N_5316);
and U6259 (N_6259,N_4833,N_4712);
nor U6260 (N_6260,N_5345,N_5550);
or U6261 (N_6261,N_4817,N_4722);
nor U6262 (N_6262,N_4721,N_5014);
or U6263 (N_6263,N_5531,N_4697);
nor U6264 (N_6264,N_5764,N_4128);
or U6265 (N_6265,N_4531,N_5206);
and U6266 (N_6266,N_4092,N_4862);
and U6267 (N_6267,N_5311,N_4106);
nor U6268 (N_6268,N_5522,N_5173);
or U6269 (N_6269,N_5588,N_4626);
nand U6270 (N_6270,N_5112,N_5329);
xor U6271 (N_6271,N_5244,N_5476);
nor U6272 (N_6272,N_5774,N_5828);
and U6273 (N_6273,N_5106,N_5653);
and U6274 (N_6274,N_4998,N_4026);
xnor U6275 (N_6275,N_5279,N_4144);
and U6276 (N_6276,N_5849,N_4932);
or U6277 (N_6277,N_4287,N_5798);
xnor U6278 (N_6278,N_5103,N_4978);
or U6279 (N_6279,N_4547,N_4724);
nand U6280 (N_6280,N_4971,N_5387);
nor U6281 (N_6281,N_5919,N_5921);
or U6282 (N_6282,N_5164,N_5791);
or U6283 (N_6283,N_5334,N_4580);
nor U6284 (N_6284,N_5786,N_4915);
or U6285 (N_6285,N_5630,N_5519);
nor U6286 (N_6286,N_4400,N_4369);
nand U6287 (N_6287,N_4326,N_5152);
xnor U6288 (N_6288,N_5400,N_4956);
or U6289 (N_6289,N_5552,N_4361);
or U6290 (N_6290,N_5662,N_4911);
xor U6291 (N_6291,N_5070,N_4465);
nand U6292 (N_6292,N_5360,N_5023);
nand U6293 (N_6293,N_5675,N_5841);
or U6294 (N_6294,N_4631,N_5952);
xnor U6295 (N_6295,N_4759,N_4813);
and U6296 (N_6296,N_4337,N_4785);
nor U6297 (N_6297,N_5289,N_4700);
or U6298 (N_6298,N_4473,N_4633);
and U6299 (N_6299,N_4120,N_4803);
xor U6300 (N_6300,N_5945,N_4240);
and U6301 (N_6301,N_5829,N_5892);
and U6302 (N_6302,N_5499,N_5879);
xnor U6303 (N_6303,N_4544,N_5673);
nand U6304 (N_6304,N_4069,N_4176);
nand U6305 (N_6305,N_4615,N_4903);
or U6306 (N_6306,N_5871,N_5910);
nand U6307 (N_6307,N_5107,N_5048);
and U6308 (N_6308,N_5011,N_5938);
and U6309 (N_6309,N_4635,N_4737);
nor U6310 (N_6310,N_4904,N_4454);
or U6311 (N_6311,N_4333,N_4233);
nand U6312 (N_6312,N_5032,N_5542);
nor U6313 (N_6313,N_4557,N_4772);
xor U6314 (N_6314,N_5543,N_4943);
nor U6315 (N_6315,N_4197,N_5012);
nor U6316 (N_6316,N_5573,N_5954);
and U6317 (N_6317,N_5464,N_5779);
nor U6318 (N_6318,N_5489,N_5019);
nor U6319 (N_6319,N_4883,N_4847);
nand U6320 (N_6320,N_4582,N_4654);
or U6321 (N_6321,N_4774,N_4796);
and U6322 (N_6322,N_4533,N_4850);
and U6323 (N_6323,N_5907,N_5228);
nor U6324 (N_6324,N_5325,N_5693);
nor U6325 (N_6325,N_4047,N_4570);
or U6326 (N_6326,N_5988,N_4814);
or U6327 (N_6327,N_5868,N_5718);
xnor U6328 (N_6328,N_5243,N_5317);
or U6329 (N_6329,N_4760,N_5177);
and U6330 (N_6330,N_5922,N_5044);
xnor U6331 (N_6331,N_4776,N_5735);
nand U6332 (N_6332,N_5719,N_4205);
nor U6333 (N_6333,N_4806,N_4357);
or U6334 (N_6334,N_4893,N_4545);
or U6335 (N_6335,N_5784,N_5137);
nor U6336 (N_6336,N_5456,N_4449);
and U6337 (N_6337,N_5003,N_5836);
nor U6338 (N_6338,N_4559,N_4763);
or U6339 (N_6339,N_4384,N_5450);
or U6340 (N_6340,N_4516,N_4766);
xor U6341 (N_6341,N_4980,N_4561);
or U6342 (N_6342,N_4499,N_5465);
nand U6343 (N_6343,N_4250,N_4241);
or U6344 (N_6344,N_5030,N_4867);
and U6345 (N_6345,N_4897,N_5278);
and U6346 (N_6346,N_5260,N_4648);
nand U6347 (N_6347,N_5891,N_4910);
nor U6348 (N_6348,N_5527,N_4953);
xnor U6349 (N_6349,N_5082,N_4187);
xnor U6350 (N_6350,N_4812,N_4681);
xor U6351 (N_6351,N_5810,N_5241);
and U6352 (N_6352,N_5042,N_5308);
or U6353 (N_6353,N_5008,N_5013);
xor U6354 (N_6354,N_4204,N_4527);
xor U6355 (N_6355,N_4380,N_5869);
nand U6356 (N_6356,N_5526,N_5690);
nor U6357 (N_6357,N_4390,N_5830);
xnor U6358 (N_6358,N_4277,N_4983);
or U6359 (N_6359,N_5277,N_4091);
and U6360 (N_6360,N_4924,N_4517);
and U6361 (N_6361,N_4420,N_5942);
or U6362 (N_6362,N_5392,N_5073);
or U6363 (N_6363,N_5917,N_5015);
or U6364 (N_6364,N_4190,N_4071);
nor U6365 (N_6365,N_4727,N_4852);
or U6366 (N_6366,N_4409,N_5104);
and U6367 (N_6367,N_4261,N_4468);
nor U6368 (N_6368,N_4537,N_4639);
nand U6369 (N_6369,N_5251,N_4593);
or U6370 (N_6370,N_4320,N_4089);
nor U6371 (N_6371,N_4762,N_4193);
and U6372 (N_6372,N_5615,N_5833);
nor U6373 (N_6373,N_4263,N_5415);
or U6374 (N_6374,N_4315,N_5421);
nor U6375 (N_6375,N_5897,N_4480);
or U6376 (N_6376,N_5788,N_5649);
and U6377 (N_6377,N_5567,N_4444);
nand U6378 (N_6378,N_5395,N_5953);
nand U6379 (N_6379,N_4742,N_5433);
or U6380 (N_6380,N_4000,N_4291);
and U6381 (N_6381,N_5748,N_5171);
nor U6382 (N_6382,N_4870,N_5486);
xnor U6383 (N_6383,N_5155,N_5027);
nor U6384 (N_6384,N_4219,N_4775);
nand U6385 (N_6385,N_5635,N_5163);
or U6386 (N_6386,N_4581,N_4970);
xnor U6387 (N_6387,N_4078,N_4767);
xnor U6388 (N_6388,N_4830,N_4575);
or U6389 (N_6389,N_4750,N_5562);
nor U6390 (N_6390,N_4329,N_4552);
nor U6391 (N_6391,N_5714,N_4921);
or U6392 (N_6392,N_5453,N_4496);
and U6393 (N_6393,N_5365,N_4451);
and U6394 (N_6394,N_4515,N_4246);
nand U6395 (N_6395,N_4171,N_4396);
xnor U6396 (N_6396,N_4399,N_4752);
xor U6397 (N_6397,N_4598,N_5205);
xor U6398 (N_6398,N_4901,N_4206);
and U6399 (N_6399,N_5971,N_5848);
nor U6400 (N_6400,N_4848,N_4336);
xnor U6401 (N_6401,N_5282,N_4483);
nor U6402 (N_6402,N_4358,N_4780);
or U6403 (N_6403,N_5972,N_4743);
and U6404 (N_6404,N_5377,N_5665);
xor U6405 (N_6405,N_4275,N_4834);
nand U6406 (N_6406,N_4677,N_5327);
nor U6407 (N_6407,N_4285,N_4695);
nor U6408 (N_6408,N_4866,N_4868);
nand U6409 (N_6409,N_5723,N_4975);
or U6410 (N_6410,N_4448,N_5367);
xor U6411 (N_6411,N_5086,N_5147);
and U6412 (N_6412,N_4751,N_5725);
xnor U6413 (N_6413,N_4492,N_4513);
and U6414 (N_6414,N_5571,N_5356);
nor U6415 (N_6415,N_5125,N_5604);
nand U6416 (N_6416,N_4891,N_4838);
nor U6417 (N_6417,N_4046,N_4841);
or U6418 (N_6418,N_5854,N_5061);
nand U6419 (N_6419,N_4093,N_5733);
nor U6420 (N_6420,N_4653,N_5949);
nand U6421 (N_6421,N_5116,N_4693);
nor U6422 (N_6422,N_4019,N_4844);
nand U6423 (N_6423,N_5466,N_4997);
or U6424 (N_6424,N_5865,N_5681);
or U6425 (N_6425,N_4564,N_4155);
or U6426 (N_6426,N_5549,N_5592);
xnor U6427 (N_6427,N_4954,N_4122);
nor U6428 (N_6428,N_4276,N_5558);
nor U6429 (N_6429,N_4661,N_4505);
nor U6430 (N_6430,N_4958,N_4638);
xor U6431 (N_6431,N_5946,N_5339);
or U6432 (N_6432,N_4539,N_5602);
or U6433 (N_6433,N_4271,N_4332);
xor U6434 (N_6434,N_4562,N_4058);
or U6435 (N_6435,N_5024,N_5374);
nand U6436 (N_6436,N_4342,N_5876);
or U6437 (N_6437,N_5625,N_5136);
and U6438 (N_6438,N_4467,N_5341);
or U6439 (N_6439,N_5348,N_5581);
or U6440 (N_6440,N_5895,N_4528);
and U6441 (N_6441,N_5328,N_4253);
nand U6442 (N_6442,N_4355,N_4686);
nor U6443 (N_6443,N_4906,N_4945);
nand U6444 (N_6444,N_5842,N_4754);
nor U6445 (N_6445,N_4055,N_5058);
and U6446 (N_6446,N_4453,N_4393);
nor U6447 (N_6447,N_5406,N_4938);
nand U6448 (N_6448,N_5789,N_4658);
and U6449 (N_6449,N_5742,N_4064);
nor U6450 (N_6450,N_5797,N_4699);
xor U6451 (N_6451,N_5192,N_4371);
and U6452 (N_6452,N_5671,N_5133);
nor U6453 (N_6453,N_5375,N_4186);
or U6454 (N_6454,N_5983,N_4735);
and U6455 (N_6455,N_5349,N_4450);
xnor U6456 (N_6456,N_4815,N_5631);
or U6457 (N_6457,N_4243,N_5705);
nand U6458 (N_6458,N_4251,N_4755);
nand U6459 (N_6459,N_5936,N_5319);
nor U6460 (N_6460,N_4134,N_4296);
nor U6461 (N_6461,N_5600,N_5785);
xnor U6462 (N_6462,N_4618,N_4230);
nand U6463 (N_6463,N_4597,N_4356);
nor U6464 (N_6464,N_5888,N_4084);
nor U6465 (N_6465,N_5503,N_5270);
xnor U6466 (N_6466,N_4963,N_5203);
nor U6467 (N_6467,N_5213,N_4824);
nand U6468 (N_6468,N_4379,N_5745);
and U6469 (N_6469,N_5941,N_4418);
or U6470 (N_6470,N_5221,N_5332);
nor U6471 (N_6471,N_5245,N_5864);
xor U6472 (N_6472,N_4242,N_5036);
xnor U6473 (N_6473,N_4520,N_5207);
nor U6474 (N_6474,N_4381,N_5080);
and U6475 (N_6475,N_4613,N_5059);
or U6476 (N_6476,N_5845,N_4679);
or U6477 (N_6477,N_5077,N_4606);
and U6478 (N_6478,N_4832,N_4099);
nor U6479 (N_6479,N_5399,N_4779);
nor U6480 (N_6480,N_5031,N_5535);
nand U6481 (N_6481,N_4081,N_5629);
nor U6482 (N_6482,N_5072,N_4907);
nor U6483 (N_6483,N_4541,N_5932);
nand U6484 (N_6484,N_4534,N_4514);
or U6485 (N_6485,N_4057,N_5818);
and U6486 (N_6486,N_4549,N_5300);
nor U6487 (N_6487,N_5057,N_5117);
nor U6488 (N_6488,N_5680,N_5034);
nand U6489 (N_6489,N_5140,N_5677);
or U6490 (N_6490,N_4554,N_5488);
xor U6491 (N_6491,N_5199,N_5633);
and U6492 (N_6492,N_5875,N_5394);
nand U6493 (N_6493,N_4666,N_4154);
and U6494 (N_6494,N_5505,N_4730);
xor U6495 (N_6495,N_5174,N_4650);
or U6496 (N_6496,N_4800,N_4257);
or U6497 (N_6497,N_4053,N_5746);
xor U6498 (N_6498,N_5632,N_5190);
and U6499 (N_6499,N_4309,N_5547);
nor U6500 (N_6500,N_4555,N_4706);
xnor U6501 (N_6501,N_4362,N_4278);
or U6502 (N_6502,N_5905,N_5153);
nor U6503 (N_6503,N_5294,N_5997);
xor U6504 (N_6504,N_4252,N_4937);
or U6505 (N_6505,N_4977,N_5315);
and U6506 (N_6506,N_4522,N_4732);
nor U6507 (N_6507,N_5330,N_4068);
nand U6508 (N_6508,N_4136,N_4006);
nor U6509 (N_6509,N_5860,N_4481);
nor U6510 (N_6510,N_5410,N_4843);
or U6511 (N_6511,N_5607,N_4939);
xnor U6512 (N_6512,N_4435,N_4828);
nand U6513 (N_6513,N_4389,N_4140);
nand U6514 (N_6514,N_5920,N_4391);
and U6515 (N_6515,N_5741,N_5814);
and U6516 (N_6516,N_5551,N_4645);
nor U6517 (N_6517,N_4201,N_5880);
and U6518 (N_6518,N_4231,N_5267);
xor U6519 (N_6519,N_4382,N_5296);
and U6520 (N_6520,N_4675,N_4577);
nand U6521 (N_6521,N_5141,N_5079);
or U6522 (N_6522,N_4341,N_4258);
and U6523 (N_6523,N_4395,N_5546);
xor U6524 (N_6524,N_5342,N_5575);
and U6525 (N_6525,N_4733,N_4065);
xnor U6526 (N_6526,N_4016,N_5777);
or U6527 (N_6527,N_4162,N_4592);
or U6528 (N_6528,N_4183,N_4164);
and U6529 (N_6529,N_4508,N_5775);
xnor U6530 (N_6530,N_4268,N_5208);
nand U6531 (N_6531,N_5576,N_5815);
nor U6532 (N_6532,N_4551,N_4161);
nor U6533 (N_6533,N_4226,N_5618);
and U6534 (N_6534,N_5379,N_5135);
xnor U6535 (N_6535,N_4682,N_5175);
xor U6536 (N_6536,N_4900,N_4432);
xnor U6537 (N_6537,N_5716,N_4521);
nand U6538 (N_6538,N_5757,N_4538);
xor U6539 (N_6539,N_4101,N_5259);
or U6540 (N_6540,N_5204,N_5694);
nor U6541 (N_6541,N_5909,N_4818);
or U6542 (N_6542,N_4457,N_5796);
nand U6543 (N_6543,N_4842,N_4172);
or U6544 (N_6544,N_4138,N_4488);
and U6545 (N_6545,N_5679,N_5256);
and U6546 (N_6546,N_5066,N_4440);
xor U6547 (N_6547,N_4020,N_5362);
or U6548 (N_6548,N_5883,N_5429);
or U6549 (N_6549,N_4927,N_4088);
and U6550 (N_6550,N_5197,N_5986);
and U6551 (N_6551,N_5506,N_5658);
nor U6552 (N_6552,N_5987,N_5962);
nand U6553 (N_6553,N_4596,N_5157);
nor U6554 (N_6554,N_4023,N_4272);
xor U6555 (N_6555,N_4279,N_4310);
nor U6556 (N_6556,N_4090,N_4075);
nand U6557 (N_6557,N_4673,N_4765);
nand U6558 (N_6558,N_5913,N_5193);
nor U6559 (N_6559,N_5802,N_5102);
nand U6560 (N_6560,N_5585,N_5250);
and U6561 (N_6561,N_5313,N_4773);
nand U6562 (N_6562,N_5083,N_5911);
and U6563 (N_6563,N_4609,N_4105);
or U6564 (N_6564,N_5760,N_5984);
and U6565 (N_6565,N_4477,N_5887);
nor U6566 (N_6566,N_4194,N_4990);
xor U6567 (N_6567,N_5947,N_4929);
nand U6568 (N_6568,N_5664,N_4940);
or U6569 (N_6569,N_5901,N_5218);
nand U6570 (N_6570,N_5007,N_4859);
and U6571 (N_6571,N_5594,N_4404);
or U6572 (N_6572,N_5766,N_5424);
nand U6573 (N_6573,N_4031,N_4923);
xor U6574 (N_6574,N_5890,N_5858);
nor U6575 (N_6575,N_4211,N_4791);
or U6576 (N_6576,N_5914,N_4188);
nand U6577 (N_6577,N_5795,N_4525);
nor U6578 (N_6578,N_5022,N_4969);
xnor U6579 (N_6579,N_5427,N_4247);
and U6580 (N_6580,N_5657,N_5634);
nor U6581 (N_6581,N_5563,N_5288);
nor U6582 (N_6582,N_5990,N_4170);
nor U6583 (N_6583,N_4799,N_4512);
nor U6584 (N_6584,N_5461,N_4500);
and U6585 (N_6585,N_5654,N_4061);
nand U6586 (N_6586,N_5196,N_4223);
nand U6587 (N_6587,N_5704,N_4649);
and U6588 (N_6588,N_4856,N_4098);
xor U6589 (N_6589,N_5088,N_5943);
or U6590 (N_6590,N_5035,N_5528);
nand U6591 (N_6591,N_5274,N_5307);
and U6592 (N_6592,N_5803,N_5660);
or U6593 (N_6593,N_5874,N_4303);
and U6594 (N_6594,N_5359,N_5026);
nand U6595 (N_6595,N_5314,N_4096);
nor U6596 (N_6596,N_4957,N_4056);
xnor U6597 (N_6597,N_4671,N_4412);
nand U6598 (N_6598,N_4667,N_4888);
nor U6599 (N_6599,N_4425,N_5676);
and U6600 (N_6600,N_4368,N_4080);
nor U6601 (N_6601,N_5559,N_5265);
xor U6602 (N_6602,N_4062,N_5149);
xor U6603 (N_6603,N_4572,N_4566);
nand U6604 (N_6604,N_4674,N_4300);
or U6605 (N_6605,N_4656,N_4439);
or U6606 (N_6606,N_5085,N_5109);
or U6607 (N_6607,N_4148,N_5127);
xnor U6608 (N_6608,N_4360,N_4405);
nor U6609 (N_6609,N_5060,N_5521);
nand U6610 (N_6610,N_5998,N_4920);
or U6611 (N_6611,N_4793,N_5408);
and U6612 (N_6612,N_5434,N_5812);
nand U6613 (N_6613,N_4713,N_4304);
nand U6614 (N_6614,N_4151,N_5955);
or U6615 (N_6615,N_4898,N_4670);
or U6616 (N_6616,N_4777,N_5656);
nand U6617 (N_6617,N_4010,N_4414);
or U6618 (N_6618,N_4102,N_4228);
nand U6619 (N_6619,N_5701,N_4416);
and U6620 (N_6620,N_4701,N_4616);
or U6621 (N_6621,N_4849,N_4669);
nor U6622 (N_6622,N_5154,N_5201);
nand U6623 (N_6623,N_4208,N_4556);
xnor U6624 (N_6624,N_4111,N_5309);
nor U6625 (N_6625,N_4013,N_5822);
xor U6626 (N_6626,N_4166,N_4996);
nor U6627 (N_6627,N_4587,N_5569);
nand U6628 (N_6628,N_4696,N_4857);
nor U6629 (N_6629,N_5885,N_5819);
nor U6630 (N_6630,N_4130,N_5471);
xor U6631 (N_6631,N_4033,N_4168);
xnor U6632 (N_6632,N_5792,N_4603);
or U6633 (N_6633,N_4802,N_4595);
nand U6634 (N_6634,N_5597,N_5188);
or U6635 (N_6635,N_4157,N_5740);
and U6636 (N_6636,N_5974,N_4608);
nor U6637 (N_6637,N_4372,N_5794);
or U6638 (N_6638,N_4394,N_5809);
or U6639 (N_6639,N_4427,N_4403);
nor U6640 (N_6640,N_4486,N_5908);
and U6641 (N_6641,N_5293,N_4629);
xor U6642 (N_6642,N_4115,N_4165);
xnor U6643 (N_6643,N_4182,N_5939);
xnor U6644 (N_6644,N_4784,N_4107);
nor U6645 (N_6645,N_4839,N_5755);
and U6646 (N_6646,N_5312,N_5383);
nor U6647 (N_6647,N_4224,N_5525);
or U6648 (N_6648,N_5577,N_5431);
xor U6649 (N_6649,N_4256,N_4067);
and U6650 (N_6650,N_5343,N_4647);
xnor U6651 (N_6651,N_4829,N_5534);
nor U6652 (N_6652,N_4222,N_5227);
nand U6653 (N_6653,N_4912,N_4308);
or U6654 (N_6654,N_4401,N_4249);
or U6655 (N_6655,N_4778,N_5906);
and U6656 (N_6656,N_5167,N_5925);
nor U6657 (N_6657,N_5706,N_4043);
nand U6658 (N_6658,N_4652,N_4079);
xnor U6659 (N_6659,N_4156,N_4458);
nor U6660 (N_6660,N_4764,N_4614);
nand U6661 (N_6661,N_5520,N_4734);
nand U6662 (N_6662,N_5231,N_4959);
nand U6663 (N_6663,N_4460,N_4143);
nand U6664 (N_6664,N_4152,N_4991);
nand U6665 (N_6665,N_4264,N_5780);
xnor U6666 (N_6666,N_5065,N_5918);
xnor U6667 (N_6667,N_4908,N_5126);
and U6668 (N_6668,N_4709,N_5460);
or U6669 (N_6669,N_4041,N_4344);
nand U6670 (N_6670,N_5229,N_4049);
nand U6671 (N_6671,N_5165,N_5385);
or U6672 (N_6672,N_4744,N_4324);
xnor U6673 (N_6673,N_4133,N_5062);
or U6674 (N_6674,N_4611,N_5110);
and U6675 (N_6675,N_5560,N_4623);
xor U6676 (N_6676,N_5894,N_5961);
nor U6677 (N_6677,N_5419,N_4992);
nor U6678 (N_6678,N_5436,N_5613);
nand U6679 (N_6679,N_5182,N_4761);
and U6680 (N_6680,N_4684,N_4988);
nor U6681 (N_6681,N_4936,N_5899);
nor U6682 (N_6682,N_5973,N_4579);
nand U6683 (N_6683,N_4305,N_4307);
or U6684 (N_6684,N_4872,N_4419);
or U6685 (N_6685,N_5176,N_5473);
nand U6686 (N_6686,N_5017,N_5092);
xor U6687 (N_6687,N_5695,N_5142);
xnor U6688 (N_6688,N_5770,N_4017);
nor U6689 (N_6689,N_4550,N_5318);
or U6690 (N_6690,N_5184,N_5444);
nor U6691 (N_6691,N_4889,N_5579);
nor U6692 (N_6692,N_5257,N_4139);
or U6693 (N_6693,N_4103,N_5401);
nand U6694 (N_6694,N_4001,N_4349);
and U6695 (N_6695,N_4127,N_4169);
xnor U6696 (N_6696,N_5021,N_4117);
or U6697 (N_6697,N_4180,N_5605);
or U6698 (N_6698,N_4146,N_5452);
nor U6699 (N_6699,N_5516,N_5846);
xor U6700 (N_6700,N_5254,N_5236);
xor U6701 (N_6701,N_4008,N_4254);
or U6702 (N_6702,N_4066,N_5290);
nor U6703 (N_6703,N_4493,N_5769);
nor U6704 (N_6704,N_5855,N_5981);
nor U6705 (N_6705,N_4437,N_4322);
and U6706 (N_6706,N_5590,N_5219);
nor U6707 (N_6707,N_5965,N_5950);
nor U6708 (N_6708,N_5324,N_5396);
nand U6709 (N_6709,N_4094,N_5724);
and U6710 (N_6710,N_5655,N_5614);
nand U6711 (N_6711,N_5335,N_4325);
and U6712 (N_6712,N_5596,N_4925);
nor U6713 (N_6713,N_4524,N_4756);
or U6714 (N_6714,N_5956,N_5485);
nor U6715 (N_6715,N_5347,N_4976);
nand U6716 (N_6716,N_4660,N_5357);
nand U6717 (N_6717,N_5198,N_4578);
xnor U6718 (N_6718,N_4880,N_5608);
nand U6719 (N_6719,N_4112,N_5388);
nand U6720 (N_6720,N_4298,N_5800);
and U6721 (N_6721,N_4119,N_5457);
nand U6722 (N_6722,N_5684,N_4808);
nor U6723 (N_6723,N_4619,N_5698);
xor U6724 (N_6724,N_5390,N_4757);
nor U6725 (N_6725,N_4109,N_4373);
nand U6726 (N_6726,N_4331,N_5497);
and U6727 (N_6727,N_5715,N_5010);
nor U6728 (N_6728,N_5443,N_5853);
nor U6729 (N_6729,N_4063,N_5354);
nand U6730 (N_6730,N_5484,N_5781);
and U6731 (N_6731,N_4625,N_4125);
or U6732 (N_6732,N_4297,N_5306);
nor U6733 (N_6733,N_5214,N_5050);
nor U6734 (N_6734,N_5425,N_4604);
or U6735 (N_6735,N_4359,N_5426);
xor U6736 (N_6736,N_4809,N_5737);
or U6737 (N_6737,N_5502,N_5643);
nor U6738 (N_6738,N_4723,N_5363);
or U6739 (N_6739,N_5253,N_4826);
or U6740 (N_6740,N_4160,N_5263);
nor U6741 (N_6741,N_5759,N_4951);
nand U6742 (N_6742,N_4837,N_4343);
or U6743 (N_6743,N_5004,N_5156);
and U6744 (N_6744,N_5337,N_5122);
nor U6745 (N_6745,N_4783,N_4262);
xnor U6746 (N_6746,N_5179,N_4946);
xor U6747 (N_6747,N_5480,N_4317);
xor U6748 (N_6748,N_5697,N_5699);
nand U6749 (N_6749,N_5487,N_4312);
and U6750 (N_6750,N_5556,N_5416);
nor U6751 (N_6751,N_5580,N_4935);
nand U6752 (N_6752,N_5996,N_4321);
nand U6753 (N_6753,N_4916,N_5382);
and U6754 (N_6754,N_4196,N_4470);
xnor U6755 (N_6755,N_4563,N_5029);
xor U6756 (N_6756,N_5130,N_5915);
and U6757 (N_6757,N_5200,N_4707);
and U6758 (N_6758,N_5586,N_4567);
nand U6759 (N_6759,N_5114,N_4502);
or U6760 (N_6760,N_4831,N_4179);
xor U6761 (N_6761,N_5612,N_5490);
xnor U6762 (N_6762,N_5583,N_4865);
xnor U6763 (N_6763,N_4397,N_4770);
nor U6764 (N_6764,N_5272,N_5637);
and U6765 (N_6765,N_5709,N_5384);
xor U6766 (N_6766,N_4461,N_4311);
nand U6767 (N_6767,N_5049,N_4482);
or U6768 (N_6768,N_4212,N_4452);
and U6769 (N_6769,N_5935,N_4428);
or U6770 (N_6770,N_4741,N_5513);
nand U6771 (N_6771,N_5510,N_4782);
nor U6772 (N_6772,N_4375,N_5323);
xor U6773 (N_6773,N_5281,N_4768);
and U6774 (N_6774,N_4801,N_4886);
nand U6775 (N_6775,N_5467,N_5640);
or U6776 (N_6776,N_5889,N_5405);
nand U6777 (N_6777,N_4299,N_4045);
nand U6778 (N_6778,N_5512,N_5373);
nor U6779 (N_6779,N_5181,N_4620);
nand U6780 (N_6780,N_4690,N_5386);
and U6781 (N_6781,N_5912,N_5233);
and U6782 (N_6782,N_4318,N_4610);
nor U6783 (N_6783,N_5570,N_5496);
or U6784 (N_6784,N_4191,N_5498);
nand U6785 (N_6785,N_5626,N_4973);
nand U6786 (N_6786,N_5477,N_5025);
xnor U6787 (N_6787,N_5609,N_5209);
or U6788 (N_6788,N_5376,N_4786);
xor U6789 (N_6789,N_4612,N_5544);
and U6790 (N_6790,N_5435,N_4511);
and U6791 (N_6791,N_5844,N_5930);
nand U6792 (N_6792,N_4794,N_4267);
nor U6793 (N_6793,N_5787,N_5273);
xnor U6794 (N_6794,N_5292,N_4571);
or U6795 (N_6795,N_4637,N_5369);
xor U6796 (N_6796,N_5094,N_5269);
xnor U6797 (N_6797,N_4407,N_4728);
nor U6798 (N_6798,N_4576,N_4234);
or U6799 (N_6799,N_4039,N_4931);
and U6800 (N_6800,N_4788,N_4600);
nand U6801 (N_6801,N_4860,N_5378);
or U6802 (N_6802,N_5721,N_4198);
nand U6803 (N_6803,N_5850,N_4892);
nand U6804 (N_6804,N_5468,N_4383);
nor U6805 (N_6805,N_4209,N_4987);
nor U6806 (N_6806,N_5978,N_5038);
nor U6807 (N_6807,N_5353,N_5071);
or U6808 (N_6808,N_4999,N_5976);
xor U6809 (N_6809,N_4560,N_5438);
nand U6810 (N_6810,N_4497,N_5744);
nand U6811 (N_6811,N_5067,N_5320);
xnor U6812 (N_6812,N_4965,N_4059);
nor U6813 (N_6813,N_4797,N_4367);
and U6814 (N_6814,N_4430,N_4350);
or U6815 (N_6815,N_5234,N_4890);
nor U6816 (N_6816,N_4584,N_5753);
nor U6817 (N_6817,N_5826,N_5729);
xnor U6818 (N_6818,N_4498,N_5669);
nor U6819 (N_6819,N_5778,N_5492);
nor U6820 (N_6820,N_5689,N_5852);
and U6821 (N_6821,N_4574,N_5098);
nand U6822 (N_6822,N_5210,N_5877);
or U6823 (N_6823,N_4979,N_5500);
and U6824 (N_6824,N_5168,N_4220);
nor U6825 (N_6825,N_5187,N_5884);
xor U6826 (N_6826,N_4417,N_5898);
nand U6827 (N_6827,N_5051,N_5099);
or U6828 (N_6828,N_4123,N_4456);
xnor U6829 (N_6829,N_5816,N_4175);
nor U6830 (N_6830,N_5145,N_4085);
nand U6831 (N_6831,N_4617,N_5249);
or U6832 (N_6832,N_4636,N_4398);
xnor U6833 (N_6833,N_4313,N_4044);
or U6834 (N_6834,N_5807,N_5222);
nor U6835 (N_6835,N_4269,N_4195);
nand U6836 (N_6836,N_4526,N_5336);
and U6837 (N_6837,N_5989,N_5472);
or U6838 (N_6838,N_4863,N_4804);
or U6839 (N_6839,N_5380,N_5302);
nor U6840 (N_6840,N_5666,N_5806);
xnor U6841 (N_6841,N_4028,N_4542);
nor U6842 (N_6842,N_5970,N_4758);
xor U6843 (N_6843,N_4914,N_4510);
and U6844 (N_6844,N_4789,N_5782);
nor U6845 (N_6845,N_5799,N_5371);
xor U6846 (N_6846,N_4173,N_5994);
nor U6847 (N_6847,N_5720,N_4934);
nand U6848 (N_6848,N_4431,N_4487);
and U6849 (N_6849,N_5838,N_5834);
and U6850 (N_6850,N_4601,N_4594);
or U6851 (N_6851,N_5355,N_5166);
or U6852 (N_6852,N_5242,N_4376);
nor U6853 (N_6853,N_4518,N_4002);
nor U6854 (N_6854,N_5151,N_4504);
nor U6855 (N_6855,N_5475,N_4607);
nor U6856 (N_6856,N_4739,N_5866);
nand U6857 (N_6857,N_5459,N_4698);
or U6858 (N_6858,N_5944,N_5557);
xor U6859 (N_6859,N_5651,N_4506);
nand U6860 (N_6860,N_5247,N_5896);
nand U6861 (N_6861,N_4199,N_4676);
and U6862 (N_6862,N_4216,N_4887);
and U6863 (N_6863,N_5966,N_4918);
xnor U6864 (N_6864,N_4930,N_5710);
and U6865 (N_6865,N_5886,N_5078);
and U6866 (N_6866,N_4740,N_4702);
nor U6867 (N_6867,N_4628,N_5591);
or U6868 (N_6868,N_5121,N_4316);
xor U6869 (N_6869,N_5326,N_4110);
nand U6870 (N_6870,N_4032,N_5417);
or U6871 (N_6871,N_4944,N_5240);
xnor U6872 (N_6872,N_5717,N_4455);
or U6873 (N_6873,N_5501,N_5968);
and U6874 (N_6874,N_5752,N_4422);
nand U6875 (N_6875,N_5432,N_4948);
and U6876 (N_6876,N_4875,N_5507);
nand U6877 (N_6877,N_5619,N_5627);
xnor U6878 (N_6878,N_4116,N_5951);
xnor U6879 (N_6879,N_5793,N_4509);
and U6880 (N_6880,N_4725,N_5761);
xnor U6881 (N_6881,N_5504,N_4070);
nor U6882 (N_6882,N_4131,N_4083);
nor U6883 (N_6883,N_4129,N_5646);
nor U6884 (N_6884,N_4781,N_5304);
nor U6885 (N_6885,N_4366,N_4664);
or U6886 (N_6886,N_5479,N_5517);
nand U6887 (N_6887,N_4573,N_5448);
and U6888 (N_6888,N_4237,N_4189);
or U6889 (N_6889,N_4438,N_5389);
xor U6890 (N_6890,N_5995,N_5252);
xor U6891 (N_6891,N_4960,N_5158);
nand U6892 (N_6892,N_5095,N_4124);
xnor U6893 (N_6893,N_4964,N_4651);
xnor U6894 (N_6894,N_5628,N_4215);
xnor U6895 (N_6895,N_5979,N_5641);
or U6896 (N_6896,N_5442,N_4042);
nand U6897 (N_6897,N_5940,N_5093);
and U6898 (N_6898,N_5747,N_5541);
nor U6899 (N_6899,N_4035,N_5574);
xor U6900 (N_6900,N_4466,N_5482);
nor U6901 (N_6901,N_5702,N_5566);
xor U6902 (N_6902,N_4406,N_5248);
nand U6903 (N_6903,N_4433,N_4328);
nand U6904 (N_6904,N_4805,N_5732);
nand U6905 (N_6905,N_4385,N_4989);
nand U6906 (N_6906,N_5111,N_5454);
or U6907 (N_6907,N_4731,N_4747);
nor U6908 (N_6908,N_5285,N_4472);
xnor U6909 (N_6909,N_4149,N_4476);
nand U6910 (N_6910,N_5511,N_5447);
or U6911 (N_6911,N_5246,N_5215);
xor U6912 (N_6912,N_4501,N_5261);
xor U6913 (N_6913,N_5536,N_4494);
nand U6914 (N_6914,N_5331,N_5264);
and U6915 (N_6915,N_4855,N_4490);
nor U6916 (N_6916,N_5582,N_5707);
and U6917 (N_6917,N_4014,N_5280);
or U6918 (N_6918,N_4302,N_4225);
or U6919 (N_6919,N_4640,N_5474);
or U6920 (N_6920,N_4392,N_5470);
nor U6921 (N_6921,N_5005,N_4132);
and U6922 (N_6922,N_5045,N_4836);
xor U6923 (N_6923,N_4869,N_5297);
and U6924 (N_6924,N_5194,N_4745);
nand U6925 (N_6925,N_5783,N_4426);
nand U6926 (N_6926,N_4798,N_4873);
nand U6927 (N_6927,N_5469,N_4445);
nand U6928 (N_6928,N_5691,N_5902);
or U6929 (N_6929,N_5052,N_5805);
nand U6930 (N_6930,N_5738,N_5089);
xnor U6931 (N_6931,N_5084,N_4054);
and U6932 (N_6932,N_5266,N_4266);
and U6933 (N_6933,N_4568,N_5598);
nor U6934 (N_6934,N_5584,N_4210);
nand U6935 (N_6935,N_4114,N_5881);
nand U6936 (N_6936,N_4363,N_4051);
xnor U6937 (N_6937,N_5321,N_4917);
or U6938 (N_6938,N_5124,N_5090);
or U6939 (N_6939,N_4290,N_5703);
or U6940 (N_6940,N_5161,N_5483);
and U6941 (N_6941,N_4259,N_4876);
nand U6942 (N_6942,N_5056,N_5069);
and U6943 (N_6943,N_4854,N_4662);
and U6944 (N_6944,N_4792,N_5352);
nor U6945 (N_6945,N_4475,N_5927);
nand U6946 (N_6946,N_5238,N_4630);
or U6947 (N_6947,N_4011,N_4087);
nand U6948 (N_6948,N_4025,N_5958);
nor U6949 (N_6949,N_4217,N_5397);
nor U6950 (N_6950,N_5538,N_4353);
nor U6951 (N_6951,N_4523,N_4972);
xnor U6952 (N_6952,N_5682,N_4994);
or U6953 (N_6953,N_4441,N_5413);
and U6954 (N_6954,N_4174,N_4229);
nor U6955 (N_6955,N_5295,N_5402);
xor U6956 (N_6956,N_5119,N_5722);
and U6957 (N_6957,N_5711,N_5960);
nor U6958 (N_6958,N_5143,N_4895);
xnor U6959 (N_6959,N_5286,N_5372);
or U6960 (N_6960,N_5622,N_5804);
nand U6961 (N_6961,N_4319,N_5823);
xnor U6962 (N_6962,N_5554,N_4928);
and U6963 (N_6963,N_5963,N_4301);
or U6964 (N_6964,N_5185,N_5593);
nor U6965 (N_6965,N_5687,N_5006);
or U6966 (N_6966,N_5055,N_4819);
nand U6967 (N_6967,N_4167,N_5346);
xor U6968 (N_6968,N_5776,N_5638);
and U6969 (N_6969,N_5977,N_4634);
nor U6970 (N_6970,N_5418,N_4955);
nor U6971 (N_6971,N_4822,N_4052);
nor U6972 (N_6972,N_5561,N_4746);
or U6973 (N_6973,N_5403,N_5159);
and U6974 (N_6974,N_4248,N_4753);
xnor U6975 (N_6975,N_4769,N_4288);
nor U6976 (N_6976,N_5189,N_5762);
and U6977 (N_6977,N_5790,N_5985);
xnor U6978 (N_6978,N_4546,N_5255);
nor U6979 (N_6979,N_4694,N_5728);
and U6980 (N_6980,N_4377,N_4012);
xor U6981 (N_6981,N_4339,N_4034);
nand U6982 (N_6982,N_4289,N_5801);
or U6983 (N_6983,N_5648,N_5652);
nand U6984 (N_6984,N_5553,N_4583);
xnor U6985 (N_6985,N_5101,N_5412);
or U6986 (N_6986,N_5642,N_4821);
or U6987 (N_6987,N_5478,N_4471);
or U6988 (N_6988,N_5767,N_4436);
or U6989 (N_6989,N_5817,N_5217);
xor U6990 (N_6990,N_4434,N_4178);
or U6991 (N_6991,N_5647,N_4274);
or U6992 (N_6992,N_5751,N_5481);
and U6993 (N_6993,N_5064,N_5672);
xnor U6994 (N_6994,N_5624,N_4177);
or U6995 (N_6995,N_4446,N_4949);
or U6996 (N_6996,N_5225,N_4704);
xnor U6997 (N_6997,N_5611,N_5028);
nand U6998 (N_6998,N_5232,N_4411);
nor U6999 (N_6999,N_5843,N_5530);
nand U7000 (N_7000,N_4175,N_4170);
and U7001 (N_7001,N_5792,N_5428);
xor U7002 (N_7002,N_5113,N_5091);
and U7003 (N_7003,N_4586,N_5002);
xnor U7004 (N_7004,N_5167,N_4185);
xnor U7005 (N_7005,N_4994,N_4776);
nand U7006 (N_7006,N_5236,N_5742);
or U7007 (N_7007,N_5051,N_4914);
and U7008 (N_7008,N_5790,N_4140);
and U7009 (N_7009,N_4250,N_5141);
nand U7010 (N_7010,N_4585,N_4358);
xor U7011 (N_7011,N_4673,N_5006);
and U7012 (N_7012,N_5828,N_5569);
xor U7013 (N_7013,N_5744,N_4806);
nor U7014 (N_7014,N_4113,N_4165);
xnor U7015 (N_7015,N_5186,N_4085);
or U7016 (N_7016,N_5632,N_4720);
or U7017 (N_7017,N_4476,N_4791);
xnor U7018 (N_7018,N_5817,N_4349);
nor U7019 (N_7019,N_4214,N_4478);
nor U7020 (N_7020,N_5623,N_5118);
and U7021 (N_7021,N_5358,N_5606);
nand U7022 (N_7022,N_5872,N_4985);
nor U7023 (N_7023,N_4531,N_5465);
xor U7024 (N_7024,N_5431,N_5324);
nor U7025 (N_7025,N_4648,N_5779);
nand U7026 (N_7026,N_5876,N_5804);
or U7027 (N_7027,N_5406,N_5246);
and U7028 (N_7028,N_4643,N_4286);
or U7029 (N_7029,N_5634,N_5612);
nand U7030 (N_7030,N_4891,N_5576);
nor U7031 (N_7031,N_5131,N_4171);
xnor U7032 (N_7032,N_5698,N_4322);
and U7033 (N_7033,N_5534,N_4978);
nor U7034 (N_7034,N_4429,N_5784);
or U7035 (N_7035,N_5696,N_5970);
xor U7036 (N_7036,N_5960,N_4300);
and U7037 (N_7037,N_4894,N_4933);
or U7038 (N_7038,N_5011,N_5893);
nand U7039 (N_7039,N_5105,N_5099);
xnor U7040 (N_7040,N_5580,N_5781);
nor U7041 (N_7041,N_4795,N_5086);
and U7042 (N_7042,N_4528,N_4640);
nand U7043 (N_7043,N_5722,N_5813);
and U7044 (N_7044,N_4909,N_5136);
nor U7045 (N_7045,N_5775,N_4817);
or U7046 (N_7046,N_5849,N_4203);
or U7047 (N_7047,N_5033,N_5343);
xnor U7048 (N_7048,N_5374,N_4983);
or U7049 (N_7049,N_5122,N_4554);
nand U7050 (N_7050,N_4397,N_5193);
nor U7051 (N_7051,N_4468,N_5419);
or U7052 (N_7052,N_4892,N_5466);
or U7053 (N_7053,N_4678,N_5811);
xor U7054 (N_7054,N_4164,N_4980);
nand U7055 (N_7055,N_5442,N_4176);
xnor U7056 (N_7056,N_4712,N_5998);
or U7057 (N_7057,N_4410,N_5646);
xor U7058 (N_7058,N_4453,N_4431);
nor U7059 (N_7059,N_5136,N_4585);
and U7060 (N_7060,N_5724,N_5605);
nand U7061 (N_7061,N_5028,N_4914);
or U7062 (N_7062,N_5122,N_5128);
and U7063 (N_7063,N_5221,N_5087);
nand U7064 (N_7064,N_4426,N_4759);
nand U7065 (N_7065,N_4939,N_5140);
or U7066 (N_7066,N_5353,N_5762);
nor U7067 (N_7067,N_4415,N_4511);
xor U7068 (N_7068,N_4945,N_4902);
nand U7069 (N_7069,N_4710,N_4216);
nor U7070 (N_7070,N_4492,N_4480);
nand U7071 (N_7071,N_4537,N_4471);
xor U7072 (N_7072,N_4649,N_5049);
or U7073 (N_7073,N_4147,N_4370);
xnor U7074 (N_7074,N_4607,N_5473);
and U7075 (N_7075,N_4057,N_4424);
nor U7076 (N_7076,N_5617,N_4389);
nand U7077 (N_7077,N_4757,N_5544);
xor U7078 (N_7078,N_5212,N_5474);
xor U7079 (N_7079,N_4779,N_5093);
and U7080 (N_7080,N_4015,N_4070);
nand U7081 (N_7081,N_5362,N_5926);
or U7082 (N_7082,N_5272,N_4012);
nand U7083 (N_7083,N_5001,N_5954);
or U7084 (N_7084,N_5053,N_5324);
xnor U7085 (N_7085,N_5678,N_4198);
xor U7086 (N_7086,N_4147,N_4928);
xor U7087 (N_7087,N_4974,N_5885);
xnor U7088 (N_7088,N_4421,N_4783);
nand U7089 (N_7089,N_5476,N_5235);
nand U7090 (N_7090,N_4677,N_5258);
or U7091 (N_7091,N_4236,N_5630);
and U7092 (N_7092,N_5354,N_5586);
and U7093 (N_7093,N_4109,N_5137);
xor U7094 (N_7094,N_5926,N_5230);
nand U7095 (N_7095,N_5233,N_4375);
and U7096 (N_7096,N_4476,N_5012);
and U7097 (N_7097,N_4393,N_4354);
and U7098 (N_7098,N_4386,N_4854);
xnor U7099 (N_7099,N_4412,N_4735);
xnor U7100 (N_7100,N_4523,N_5713);
and U7101 (N_7101,N_5335,N_4069);
or U7102 (N_7102,N_4764,N_5923);
and U7103 (N_7103,N_5575,N_4578);
or U7104 (N_7104,N_4133,N_4196);
and U7105 (N_7105,N_5212,N_5719);
xnor U7106 (N_7106,N_5286,N_4617);
nor U7107 (N_7107,N_5105,N_5184);
nand U7108 (N_7108,N_5351,N_5575);
or U7109 (N_7109,N_5418,N_4624);
or U7110 (N_7110,N_4576,N_4821);
xor U7111 (N_7111,N_5199,N_4997);
xor U7112 (N_7112,N_5819,N_4074);
xor U7113 (N_7113,N_5029,N_5975);
xor U7114 (N_7114,N_5684,N_5960);
nor U7115 (N_7115,N_4834,N_5602);
or U7116 (N_7116,N_4000,N_4487);
nand U7117 (N_7117,N_5956,N_5248);
or U7118 (N_7118,N_5778,N_4334);
xor U7119 (N_7119,N_5229,N_4481);
nor U7120 (N_7120,N_5177,N_4368);
xor U7121 (N_7121,N_4964,N_4343);
xor U7122 (N_7122,N_5497,N_5609);
nor U7123 (N_7123,N_5318,N_4059);
and U7124 (N_7124,N_5636,N_4827);
nand U7125 (N_7125,N_5226,N_5700);
or U7126 (N_7126,N_4315,N_4820);
or U7127 (N_7127,N_5631,N_5558);
or U7128 (N_7128,N_4583,N_4330);
and U7129 (N_7129,N_5672,N_4314);
nand U7130 (N_7130,N_5576,N_4024);
and U7131 (N_7131,N_4498,N_5478);
nor U7132 (N_7132,N_5421,N_4557);
nor U7133 (N_7133,N_4628,N_4743);
xor U7134 (N_7134,N_5340,N_5858);
nor U7135 (N_7135,N_4135,N_5313);
nand U7136 (N_7136,N_5507,N_4197);
nand U7137 (N_7137,N_5622,N_4973);
or U7138 (N_7138,N_4974,N_4945);
nor U7139 (N_7139,N_4422,N_5370);
nand U7140 (N_7140,N_5497,N_4286);
nand U7141 (N_7141,N_4567,N_4031);
xor U7142 (N_7142,N_5717,N_4590);
or U7143 (N_7143,N_4913,N_4754);
and U7144 (N_7144,N_5615,N_5465);
xnor U7145 (N_7145,N_4725,N_4664);
nor U7146 (N_7146,N_4300,N_4406);
nor U7147 (N_7147,N_5408,N_4294);
or U7148 (N_7148,N_4464,N_5334);
xnor U7149 (N_7149,N_4814,N_4976);
or U7150 (N_7150,N_5149,N_5727);
nand U7151 (N_7151,N_5741,N_5803);
nor U7152 (N_7152,N_5288,N_4589);
and U7153 (N_7153,N_5456,N_5321);
nor U7154 (N_7154,N_5192,N_4576);
xnor U7155 (N_7155,N_5084,N_4305);
nor U7156 (N_7156,N_5845,N_5865);
xnor U7157 (N_7157,N_5705,N_5490);
and U7158 (N_7158,N_4819,N_4558);
and U7159 (N_7159,N_5367,N_4760);
or U7160 (N_7160,N_4052,N_4645);
xor U7161 (N_7161,N_5985,N_4877);
xor U7162 (N_7162,N_4874,N_4107);
nand U7163 (N_7163,N_5842,N_5437);
nor U7164 (N_7164,N_5471,N_5220);
or U7165 (N_7165,N_4452,N_5857);
and U7166 (N_7166,N_5151,N_4121);
xor U7167 (N_7167,N_4004,N_5895);
and U7168 (N_7168,N_4017,N_5609);
nor U7169 (N_7169,N_5929,N_5968);
xnor U7170 (N_7170,N_4867,N_4435);
xnor U7171 (N_7171,N_5228,N_5332);
or U7172 (N_7172,N_5967,N_5252);
xnor U7173 (N_7173,N_5596,N_4187);
nor U7174 (N_7174,N_5423,N_4183);
and U7175 (N_7175,N_5012,N_4959);
nor U7176 (N_7176,N_5604,N_4633);
nand U7177 (N_7177,N_4733,N_5663);
and U7178 (N_7178,N_5738,N_4963);
or U7179 (N_7179,N_4252,N_4272);
nand U7180 (N_7180,N_4250,N_4273);
and U7181 (N_7181,N_4579,N_4834);
xnor U7182 (N_7182,N_5640,N_4107);
and U7183 (N_7183,N_5055,N_4000);
nor U7184 (N_7184,N_4538,N_4688);
xnor U7185 (N_7185,N_5609,N_4093);
or U7186 (N_7186,N_5281,N_5928);
xor U7187 (N_7187,N_4846,N_4264);
or U7188 (N_7188,N_5972,N_4090);
or U7189 (N_7189,N_4204,N_5729);
and U7190 (N_7190,N_4240,N_4244);
and U7191 (N_7191,N_4394,N_4779);
xor U7192 (N_7192,N_4963,N_4660);
nor U7193 (N_7193,N_4647,N_5457);
or U7194 (N_7194,N_5700,N_5458);
or U7195 (N_7195,N_4537,N_5891);
nand U7196 (N_7196,N_5998,N_5890);
and U7197 (N_7197,N_5756,N_5309);
nand U7198 (N_7198,N_5733,N_4391);
nand U7199 (N_7199,N_4287,N_4330);
nand U7200 (N_7200,N_4056,N_5611);
nand U7201 (N_7201,N_5937,N_5424);
or U7202 (N_7202,N_5332,N_5627);
xor U7203 (N_7203,N_5182,N_5798);
and U7204 (N_7204,N_5972,N_4221);
or U7205 (N_7205,N_5580,N_5395);
nor U7206 (N_7206,N_4169,N_4843);
nand U7207 (N_7207,N_5681,N_5663);
nand U7208 (N_7208,N_4032,N_5702);
xnor U7209 (N_7209,N_4257,N_4691);
and U7210 (N_7210,N_4393,N_5091);
and U7211 (N_7211,N_4696,N_4746);
nor U7212 (N_7212,N_5909,N_4839);
xor U7213 (N_7213,N_5386,N_4765);
xnor U7214 (N_7214,N_4909,N_5706);
and U7215 (N_7215,N_4482,N_4562);
and U7216 (N_7216,N_4317,N_4755);
or U7217 (N_7217,N_4353,N_4547);
nand U7218 (N_7218,N_4152,N_4778);
nor U7219 (N_7219,N_4891,N_5856);
and U7220 (N_7220,N_4414,N_5758);
or U7221 (N_7221,N_5267,N_4463);
or U7222 (N_7222,N_5979,N_5922);
nor U7223 (N_7223,N_5975,N_4049);
and U7224 (N_7224,N_4046,N_4301);
or U7225 (N_7225,N_5831,N_5025);
xor U7226 (N_7226,N_4826,N_4449);
or U7227 (N_7227,N_5791,N_4714);
or U7228 (N_7228,N_5586,N_5717);
nand U7229 (N_7229,N_5459,N_4485);
or U7230 (N_7230,N_4865,N_5683);
or U7231 (N_7231,N_4306,N_4893);
nand U7232 (N_7232,N_4771,N_5761);
and U7233 (N_7233,N_4826,N_4035);
xor U7234 (N_7234,N_5714,N_5700);
and U7235 (N_7235,N_5463,N_4144);
and U7236 (N_7236,N_4281,N_5823);
or U7237 (N_7237,N_5869,N_5048);
or U7238 (N_7238,N_5641,N_4873);
and U7239 (N_7239,N_5956,N_4216);
and U7240 (N_7240,N_4363,N_5345);
nor U7241 (N_7241,N_4299,N_4439);
nor U7242 (N_7242,N_4492,N_5806);
or U7243 (N_7243,N_5433,N_5782);
xor U7244 (N_7244,N_5870,N_5088);
nand U7245 (N_7245,N_4157,N_4109);
nor U7246 (N_7246,N_5980,N_5462);
nor U7247 (N_7247,N_4633,N_4907);
nor U7248 (N_7248,N_4375,N_5150);
and U7249 (N_7249,N_4732,N_4448);
nand U7250 (N_7250,N_5295,N_4314);
nand U7251 (N_7251,N_5003,N_4590);
nand U7252 (N_7252,N_5863,N_4090);
nand U7253 (N_7253,N_5398,N_5419);
and U7254 (N_7254,N_5180,N_5855);
xor U7255 (N_7255,N_4833,N_5099);
or U7256 (N_7256,N_5656,N_4341);
or U7257 (N_7257,N_5181,N_5902);
and U7258 (N_7258,N_5292,N_5711);
xnor U7259 (N_7259,N_5682,N_4397);
xor U7260 (N_7260,N_4992,N_4456);
or U7261 (N_7261,N_5115,N_5934);
and U7262 (N_7262,N_4908,N_4445);
or U7263 (N_7263,N_4541,N_5267);
xnor U7264 (N_7264,N_4505,N_5880);
nand U7265 (N_7265,N_4622,N_5989);
or U7266 (N_7266,N_4464,N_4859);
and U7267 (N_7267,N_4097,N_5009);
nor U7268 (N_7268,N_4020,N_4116);
xnor U7269 (N_7269,N_5175,N_4174);
nor U7270 (N_7270,N_4410,N_4927);
xor U7271 (N_7271,N_5080,N_5231);
and U7272 (N_7272,N_5630,N_4985);
nand U7273 (N_7273,N_4085,N_4955);
nand U7274 (N_7274,N_5613,N_4804);
xnor U7275 (N_7275,N_4072,N_5716);
nor U7276 (N_7276,N_4006,N_5669);
or U7277 (N_7277,N_4317,N_5658);
nor U7278 (N_7278,N_4581,N_5857);
xnor U7279 (N_7279,N_4157,N_4652);
nor U7280 (N_7280,N_4825,N_4592);
nand U7281 (N_7281,N_4043,N_4429);
and U7282 (N_7282,N_4014,N_5785);
nor U7283 (N_7283,N_4362,N_4471);
and U7284 (N_7284,N_5410,N_4595);
and U7285 (N_7285,N_5666,N_4625);
nor U7286 (N_7286,N_4737,N_5327);
nand U7287 (N_7287,N_5411,N_5564);
nor U7288 (N_7288,N_5058,N_5140);
or U7289 (N_7289,N_5427,N_4673);
nand U7290 (N_7290,N_5140,N_5570);
and U7291 (N_7291,N_4477,N_4097);
and U7292 (N_7292,N_4982,N_4370);
xor U7293 (N_7293,N_5876,N_5651);
nor U7294 (N_7294,N_5503,N_5738);
nor U7295 (N_7295,N_4433,N_4850);
nand U7296 (N_7296,N_4345,N_4376);
nand U7297 (N_7297,N_4930,N_4296);
or U7298 (N_7298,N_4075,N_4192);
or U7299 (N_7299,N_5674,N_4672);
nor U7300 (N_7300,N_5024,N_4266);
xnor U7301 (N_7301,N_4036,N_5355);
and U7302 (N_7302,N_4531,N_5036);
nand U7303 (N_7303,N_4955,N_4111);
xor U7304 (N_7304,N_4434,N_5163);
and U7305 (N_7305,N_5378,N_4352);
or U7306 (N_7306,N_4368,N_5258);
nor U7307 (N_7307,N_5490,N_5286);
nand U7308 (N_7308,N_4347,N_5662);
xnor U7309 (N_7309,N_4128,N_4759);
xnor U7310 (N_7310,N_4379,N_5556);
and U7311 (N_7311,N_5019,N_5605);
nand U7312 (N_7312,N_5271,N_4878);
or U7313 (N_7313,N_4470,N_5695);
or U7314 (N_7314,N_4070,N_5452);
nor U7315 (N_7315,N_4636,N_5561);
and U7316 (N_7316,N_4068,N_4601);
xor U7317 (N_7317,N_4968,N_5862);
and U7318 (N_7318,N_4861,N_5671);
or U7319 (N_7319,N_5568,N_4976);
or U7320 (N_7320,N_5488,N_4750);
or U7321 (N_7321,N_5295,N_5114);
or U7322 (N_7322,N_4946,N_5187);
nor U7323 (N_7323,N_5358,N_4986);
xnor U7324 (N_7324,N_5576,N_5337);
or U7325 (N_7325,N_4759,N_4817);
nand U7326 (N_7326,N_5132,N_5830);
or U7327 (N_7327,N_4788,N_5734);
nor U7328 (N_7328,N_5231,N_5813);
and U7329 (N_7329,N_5915,N_4899);
nand U7330 (N_7330,N_5064,N_4760);
and U7331 (N_7331,N_4843,N_4912);
or U7332 (N_7332,N_5882,N_4121);
nand U7333 (N_7333,N_4489,N_5214);
or U7334 (N_7334,N_4965,N_4599);
nor U7335 (N_7335,N_5790,N_4091);
nand U7336 (N_7336,N_4814,N_5230);
or U7337 (N_7337,N_5727,N_4984);
xor U7338 (N_7338,N_4789,N_4621);
xor U7339 (N_7339,N_4078,N_5521);
or U7340 (N_7340,N_4831,N_5185);
xnor U7341 (N_7341,N_5292,N_5137);
xor U7342 (N_7342,N_5409,N_4631);
and U7343 (N_7343,N_4901,N_4084);
xor U7344 (N_7344,N_5301,N_4832);
or U7345 (N_7345,N_5911,N_4550);
or U7346 (N_7346,N_4732,N_5546);
nand U7347 (N_7347,N_4177,N_4131);
or U7348 (N_7348,N_5395,N_5358);
and U7349 (N_7349,N_4709,N_5659);
nor U7350 (N_7350,N_5069,N_5963);
or U7351 (N_7351,N_4795,N_5611);
nand U7352 (N_7352,N_4778,N_4363);
xor U7353 (N_7353,N_4314,N_5010);
nand U7354 (N_7354,N_5413,N_5752);
nor U7355 (N_7355,N_4286,N_4889);
xnor U7356 (N_7356,N_4734,N_4963);
nor U7357 (N_7357,N_4716,N_4007);
nor U7358 (N_7358,N_4460,N_5023);
or U7359 (N_7359,N_5568,N_5454);
nor U7360 (N_7360,N_5002,N_4532);
xor U7361 (N_7361,N_4162,N_4761);
nor U7362 (N_7362,N_4753,N_5227);
nand U7363 (N_7363,N_4453,N_5220);
nand U7364 (N_7364,N_5638,N_5600);
nor U7365 (N_7365,N_5468,N_4657);
or U7366 (N_7366,N_4343,N_5285);
xor U7367 (N_7367,N_4946,N_4920);
or U7368 (N_7368,N_4432,N_5033);
xnor U7369 (N_7369,N_4166,N_4715);
or U7370 (N_7370,N_4409,N_4408);
nor U7371 (N_7371,N_5796,N_5770);
nand U7372 (N_7372,N_4533,N_4404);
or U7373 (N_7373,N_4822,N_4392);
or U7374 (N_7374,N_5800,N_5274);
nor U7375 (N_7375,N_4634,N_4211);
nand U7376 (N_7376,N_5336,N_4967);
nand U7377 (N_7377,N_5173,N_4211);
nor U7378 (N_7378,N_5682,N_5119);
nor U7379 (N_7379,N_5096,N_5126);
nand U7380 (N_7380,N_5389,N_4122);
nand U7381 (N_7381,N_4535,N_4315);
and U7382 (N_7382,N_4791,N_5240);
nand U7383 (N_7383,N_5106,N_5735);
and U7384 (N_7384,N_5817,N_5396);
xor U7385 (N_7385,N_5568,N_4143);
or U7386 (N_7386,N_5463,N_5325);
xnor U7387 (N_7387,N_4227,N_5421);
nor U7388 (N_7388,N_4024,N_5540);
or U7389 (N_7389,N_5511,N_5036);
or U7390 (N_7390,N_5127,N_4895);
nor U7391 (N_7391,N_5141,N_4176);
nor U7392 (N_7392,N_4909,N_4235);
xnor U7393 (N_7393,N_5468,N_4575);
nand U7394 (N_7394,N_5968,N_4629);
nand U7395 (N_7395,N_4954,N_4902);
nand U7396 (N_7396,N_4985,N_5098);
or U7397 (N_7397,N_4922,N_4201);
and U7398 (N_7398,N_4040,N_4338);
and U7399 (N_7399,N_4281,N_4188);
nand U7400 (N_7400,N_4816,N_5425);
or U7401 (N_7401,N_4718,N_5666);
xor U7402 (N_7402,N_5454,N_4357);
xor U7403 (N_7403,N_5083,N_5149);
nand U7404 (N_7404,N_5793,N_4918);
or U7405 (N_7405,N_5153,N_4486);
xnor U7406 (N_7406,N_4523,N_5635);
or U7407 (N_7407,N_5689,N_4735);
nand U7408 (N_7408,N_5624,N_4771);
or U7409 (N_7409,N_4055,N_4574);
nand U7410 (N_7410,N_5370,N_4199);
and U7411 (N_7411,N_4149,N_5471);
or U7412 (N_7412,N_4929,N_4210);
nand U7413 (N_7413,N_4845,N_4388);
xor U7414 (N_7414,N_4745,N_4347);
or U7415 (N_7415,N_4237,N_4793);
or U7416 (N_7416,N_4361,N_4549);
xnor U7417 (N_7417,N_5870,N_4784);
nand U7418 (N_7418,N_5693,N_5364);
or U7419 (N_7419,N_4433,N_5721);
or U7420 (N_7420,N_4169,N_5837);
and U7421 (N_7421,N_5816,N_5387);
xnor U7422 (N_7422,N_5086,N_5979);
nor U7423 (N_7423,N_5478,N_4521);
nor U7424 (N_7424,N_5555,N_5689);
or U7425 (N_7425,N_4611,N_5418);
xor U7426 (N_7426,N_4712,N_5327);
and U7427 (N_7427,N_5999,N_4206);
or U7428 (N_7428,N_5907,N_5167);
and U7429 (N_7429,N_4757,N_5301);
or U7430 (N_7430,N_5604,N_5282);
nand U7431 (N_7431,N_5036,N_4237);
nand U7432 (N_7432,N_5588,N_4878);
and U7433 (N_7433,N_4522,N_5812);
nor U7434 (N_7434,N_4703,N_5597);
and U7435 (N_7435,N_5420,N_4576);
nand U7436 (N_7436,N_5954,N_4394);
xor U7437 (N_7437,N_5021,N_5448);
nand U7438 (N_7438,N_5105,N_4236);
xnor U7439 (N_7439,N_5344,N_4810);
and U7440 (N_7440,N_5886,N_4538);
nor U7441 (N_7441,N_5989,N_5848);
nor U7442 (N_7442,N_4633,N_5119);
and U7443 (N_7443,N_5527,N_4229);
nor U7444 (N_7444,N_4716,N_5557);
and U7445 (N_7445,N_4894,N_4251);
nand U7446 (N_7446,N_4996,N_5523);
nand U7447 (N_7447,N_4490,N_5773);
nand U7448 (N_7448,N_5954,N_5124);
and U7449 (N_7449,N_4016,N_4677);
and U7450 (N_7450,N_4219,N_5608);
and U7451 (N_7451,N_4464,N_5864);
and U7452 (N_7452,N_5178,N_4475);
xor U7453 (N_7453,N_5125,N_4076);
nand U7454 (N_7454,N_5431,N_5831);
nor U7455 (N_7455,N_4675,N_4118);
xnor U7456 (N_7456,N_4626,N_5547);
or U7457 (N_7457,N_4432,N_5504);
xnor U7458 (N_7458,N_4257,N_4011);
xnor U7459 (N_7459,N_5004,N_4440);
nor U7460 (N_7460,N_5211,N_5577);
xor U7461 (N_7461,N_5428,N_5304);
and U7462 (N_7462,N_5332,N_5612);
nor U7463 (N_7463,N_5980,N_5311);
nor U7464 (N_7464,N_5416,N_5839);
xor U7465 (N_7465,N_4226,N_5792);
nand U7466 (N_7466,N_4619,N_4333);
nor U7467 (N_7467,N_5662,N_4708);
nor U7468 (N_7468,N_5069,N_5865);
or U7469 (N_7469,N_5646,N_4803);
nor U7470 (N_7470,N_4827,N_5800);
nor U7471 (N_7471,N_5043,N_4697);
nand U7472 (N_7472,N_4657,N_4487);
xor U7473 (N_7473,N_5261,N_4974);
nand U7474 (N_7474,N_4387,N_5954);
or U7475 (N_7475,N_5193,N_4578);
and U7476 (N_7476,N_4120,N_5388);
and U7477 (N_7477,N_4075,N_5686);
and U7478 (N_7478,N_5674,N_5663);
or U7479 (N_7479,N_5402,N_5898);
or U7480 (N_7480,N_5382,N_5037);
or U7481 (N_7481,N_5561,N_5088);
or U7482 (N_7482,N_5048,N_5692);
or U7483 (N_7483,N_4910,N_4925);
nand U7484 (N_7484,N_5983,N_5395);
nand U7485 (N_7485,N_5785,N_4537);
nand U7486 (N_7486,N_5082,N_4107);
or U7487 (N_7487,N_4059,N_4547);
and U7488 (N_7488,N_5010,N_5470);
and U7489 (N_7489,N_5776,N_5213);
and U7490 (N_7490,N_4611,N_5829);
nand U7491 (N_7491,N_5428,N_4650);
nor U7492 (N_7492,N_5131,N_5310);
nand U7493 (N_7493,N_5717,N_5722);
nand U7494 (N_7494,N_4288,N_5837);
and U7495 (N_7495,N_4043,N_4894);
nor U7496 (N_7496,N_4292,N_5730);
nor U7497 (N_7497,N_5860,N_5169);
nor U7498 (N_7498,N_4816,N_4622);
nand U7499 (N_7499,N_4302,N_4326);
nor U7500 (N_7500,N_4416,N_5658);
or U7501 (N_7501,N_4506,N_5659);
nor U7502 (N_7502,N_5601,N_5733);
or U7503 (N_7503,N_4794,N_5830);
xnor U7504 (N_7504,N_5443,N_5749);
nor U7505 (N_7505,N_5011,N_5976);
or U7506 (N_7506,N_5035,N_5063);
and U7507 (N_7507,N_5650,N_5087);
or U7508 (N_7508,N_4768,N_4544);
nor U7509 (N_7509,N_4316,N_4320);
and U7510 (N_7510,N_4708,N_5688);
nand U7511 (N_7511,N_4664,N_4080);
nor U7512 (N_7512,N_5328,N_5311);
xnor U7513 (N_7513,N_5166,N_5544);
nor U7514 (N_7514,N_5130,N_4277);
and U7515 (N_7515,N_5059,N_4530);
nand U7516 (N_7516,N_5501,N_5866);
nor U7517 (N_7517,N_5862,N_5131);
and U7518 (N_7518,N_5859,N_5168);
or U7519 (N_7519,N_4596,N_5200);
and U7520 (N_7520,N_5723,N_5716);
and U7521 (N_7521,N_4040,N_4256);
xor U7522 (N_7522,N_5262,N_5202);
nand U7523 (N_7523,N_4917,N_5301);
nand U7524 (N_7524,N_5733,N_5336);
xnor U7525 (N_7525,N_4236,N_4887);
nand U7526 (N_7526,N_4921,N_5508);
xnor U7527 (N_7527,N_4094,N_4503);
nand U7528 (N_7528,N_5529,N_5803);
and U7529 (N_7529,N_5653,N_5446);
xor U7530 (N_7530,N_5618,N_5759);
and U7531 (N_7531,N_4818,N_5077);
or U7532 (N_7532,N_5672,N_4594);
or U7533 (N_7533,N_5622,N_4075);
or U7534 (N_7534,N_4622,N_5460);
or U7535 (N_7535,N_5093,N_4022);
and U7536 (N_7536,N_4470,N_5666);
or U7537 (N_7537,N_4197,N_4632);
or U7538 (N_7538,N_5465,N_4739);
or U7539 (N_7539,N_5759,N_5382);
nor U7540 (N_7540,N_4016,N_5055);
xnor U7541 (N_7541,N_4628,N_5678);
xor U7542 (N_7542,N_5602,N_5933);
xnor U7543 (N_7543,N_4010,N_4288);
nor U7544 (N_7544,N_4292,N_5574);
nand U7545 (N_7545,N_5749,N_4954);
or U7546 (N_7546,N_5396,N_4224);
nor U7547 (N_7547,N_4695,N_4043);
and U7548 (N_7548,N_4609,N_5098);
xor U7549 (N_7549,N_5507,N_4146);
nand U7550 (N_7550,N_4095,N_4756);
nor U7551 (N_7551,N_4456,N_5290);
and U7552 (N_7552,N_4202,N_4050);
nand U7553 (N_7553,N_5008,N_4558);
or U7554 (N_7554,N_4387,N_5814);
and U7555 (N_7555,N_4091,N_5679);
and U7556 (N_7556,N_5275,N_4009);
xnor U7557 (N_7557,N_4112,N_4147);
xnor U7558 (N_7558,N_4693,N_4830);
or U7559 (N_7559,N_5116,N_5837);
nand U7560 (N_7560,N_4175,N_5797);
and U7561 (N_7561,N_4113,N_5753);
nand U7562 (N_7562,N_4883,N_4726);
xnor U7563 (N_7563,N_4178,N_5042);
or U7564 (N_7564,N_4902,N_4320);
xnor U7565 (N_7565,N_4640,N_4339);
nand U7566 (N_7566,N_5227,N_4284);
xor U7567 (N_7567,N_5508,N_5777);
or U7568 (N_7568,N_4818,N_4439);
nand U7569 (N_7569,N_5324,N_5953);
and U7570 (N_7570,N_4197,N_5118);
or U7571 (N_7571,N_4944,N_4902);
nand U7572 (N_7572,N_4852,N_5181);
nor U7573 (N_7573,N_5057,N_4275);
nor U7574 (N_7574,N_5947,N_4903);
and U7575 (N_7575,N_5003,N_4811);
nor U7576 (N_7576,N_5350,N_5310);
nand U7577 (N_7577,N_4521,N_4171);
nor U7578 (N_7578,N_5150,N_5125);
nand U7579 (N_7579,N_4720,N_5927);
xnor U7580 (N_7580,N_4220,N_5909);
xnor U7581 (N_7581,N_5779,N_5420);
and U7582 (N_7582,N_4037,N_4364);
and U7583 (N_7583,N_4837,N_5415);
nor U7584 (N_7584,N_5875,N_5599);
xor U7585 (N_7585,N_5022,N_5468);
or U7586 (N_7586,N_4485,N_4761);
nor U7587 (N_7587,N_4679,N_4756);
nand U7588 (N_7588,N_4133,N_4285);
and U7589 (N_7589,N_5899,N_4148);
or U7590 (N_7590,N_5686,N_5436);
or U7591 (N_7591,N_4147,N_5612);
xnor U7592 (N_7592,N_5294,N_5526);
or U7593 (N_7593,N_4662,N_4861);
and U7594 (N_7594,N_4779,N_4531);
nor U7595 (N_7595,N_4851,N_5956);
nor U7596 (N_7596,N_5995,N_5221);
and U7597 (N_7597,N_4907,N_5509);
nor U7598 (N_7598,N_5154,N_5205);
or U7599 (N_7599,N_4868,N_4409);
nand U7600 (N_7600,N_5168,N_4861);
and U7601 (N_7601,N_5881,N_4124);
and U7602 (N_7602,N_4279,N_4172);
nor U7603 (N_7603,N_5791,N_5343);
nand U7604 (N_7604,N_4155,N_5601);
nand U7605 (N_7605,N_4181,N_4807);
or U7606 (N_7606,N_5233,N_5898);
nor U7607 (N_7607,N_5699,N_4582);
and U7608 (N_7608,N_4201,N_4311);
or U7609 (N_7609,N_5059,N_5861);
xnor U7610 (N_7610,N_5998,N_5288);
and U7611 (N_7611,N_5599,N_4223);
nand U7612 (N_7612,N_4096,N_5315);
nand U7613 (N_7613,N_4118,N_4697);
xnor U7614 (N_7614,N_4931,N_4395);
or U7615 (N_7615,N_4860,N_4189);
or U7616 (N_7616,N_5515,N_4512);
nand U7617 (N_7617,N_5902,N_5308);
nand U7618 (N_7618,N_4143,N_4157);
nand U7619 (N_7619,N_5143,N_5825);
and U7620 (N_7620,N_4718,N_4884);
nor U7621 (N_7621,N_5341,N_5537);
nor U7622 (N_7622,N_5250,N_4424);
xnor U7623 (N_7623,N_4821,N_5635);
and U7624 (N_7624,N_5267,N_4514);
nand U7625 (N_7625,N_4006,N_4400);
xnor U7626 (N_7626,N_5198,N_4097);
nand U7627 (N_7627,N_5375,N_5323);
nor U7628 (N_7628,N_4930,N_4676);
and U7629 (N_7629,N_5589,N_4022);
xor U7630 (N_7630,N_5909,N_5170);
and U7631 (N_7631,N_4704,N_5646);
nor U7632 (N_7632,N_5651,N_4262);
nand U7633 (N_7633,N_4555,N_5954);
nor U7634 (N_7634,N_4530,N_5946);
and U7635 (N_7635,N_5420,N_4201);
nor U7636 (N_7636,N_4074,N_4547);
xor U7637 (N_7637,N_4935,N_5780);
or U7638 (N_7638,N_5996,N_4394);
nand U7639 (N_7639,N_5818,N_5145);
xnor U7640 (N_7640,N_5151,N_4265);
and U7641 (N_7641,N_5467,N_5518);
or U7642 (N_7642,N_4552,N_4709);
and U7643 (N_7643,N_5956,N_5402);
xor U7644 (N_7644,N_4910,N_5461);
and U7645 (N_7645,N_4173,N_5412);
xor U7646 (N_7646,N_5075,N_5956);
xnor U7647 (N_7647,N_4144,N_4548);
or U7648 (N_7648,N_4022,N_4665);
and U7649 (N_7649,N_4677,N_4383);
xnor U7650 (N_7650,N_5738,N_4808);
nand U7651 (N_7651,N_5044,N_4158);
and U7652 (N_7652,N_4226,N_5487);
and U7653 (N_7653,N_4039,N_5207);
nand U7654 (N_7654,N_4870,N_5441);
nor U7655 (N_7655,N_4692,N_5500);
and U7656 (N_7656,N_5029,N_5929);
nand U7657 (N_7657,N_4245,N_5940);
xor U7658 (N_7658,N_4927,N_4898);
nor U7659 (N_7659,N_4163,N_5648);
and U7660 (N_7660,N_5128,N_5759);
xor U7661 (N_7661,N_4467,N_5918);
or U7662 (N_7662,N_5321,N_5049);
xnor U7663 (N_7663,N_5408,N_5102);
or U7664 (N_7664,N_5089,N_5997);
and U7665 (N_7665,N_5342,N_4562);
or U7666 (N_7666,N_4940,N_5567);
xor U7667 (N_7667,N_4487,N_5024);
xor U7668 (N_7668,N_4604,N_4421);
nor U7669 (N_7669,N_5604,N_4859);
nor U7670 (N_7670,N_4058,N_5404);
nor U7671 (N_7671,N_5264,N_5880);
or U7672 (N_7672,N_5863,N_5062);
or U7673 (N_7673,N_4531,N_5474);
xnor U7674 (N_7674,N_4816,N_5138);
nor U7675 (N_7675,N_4485,N_5174);
nand U7676 (N_7676,N_5217,N_5507);
xor U7677 (N_7677,N_4284,N_5973);
nand U7678 (N_7678,N_4380,N_5789);
nor U7679 (N_7679,N_4838,N_4875);
nor U7680 (N_7680,N_4287,N_5035);
xnor U7681 (N_7681,N_5413,N_4914);
or U7682 (N_7682,N_5508,N_4689);
nor U7683 (N_7683,N_5044,N_5017);
and U7684 (N_7684,N_5607,N_4471);
or U7685 (N_7685,N_5681,N_4869);
or U7686 (N_7686,N_4201,N_5786);
and U7687 (N_7687,N_4708,N_5811);
and U7688 (N_7688,N_5157,N_5681);
or U7689 (N_7689,N_5546,N_5742);
or U7690 (N_7690,N_5649,N_5185);
nand U7691 (N_7691,N_4680,N_5564);
nor U7692 (N_7692,N_5129,N_4583);
nor U7693 (N_7693,N_4008,N_4795);
or U7694 (N_7694,N_5879,N_4961);
nand U7695 (N_7695,N_5927,N_5253);
or U7696 (N_7696,N_5762,N_5988);
or U7697 (N_7697,N_5311,N_5501);
nand U7698 (N_7698,N_5082,N_5772);
xnor U7699 (N_7699,N_4050,N_4515);
and U7700 (N_7700,N_5643,N_5850);
and U7701 (N_7701,N_4184,N_5627);
nor U7702 (N_7702,N_5857,N_5043);
and U7703 (N_7703,N_4418,N_4396);
or U7704 (N_7704,N_5162,N_4300);
or U7705 (N_7705,N_4122,N_5872);
nor U7706 (N_7706,N_5606,N_5315);
or U7707 (N_7707,N_4005,N_4327);
and U7708 (N_7708,N_4524,N_4294);
and U7709 (N_7709,N_4515,N_4203);
and U7710 (N_7710,N_5892,N_4854);
or U7711 (N_7711,N_5346,N_5609);
nor U7712 (N_7712,N_4206,N_4159);
or U7713 (N_7713,N_4772,N_4088);
xnor U7714 (N_7714,N_5538,N_4828);
xnor U7715 (N_7715,N_4173,N_4614);
xnor U7716 (N_7716,N_5469,N_5353);
xor U7717 (N_7717,N_5171,N_5370);
and U7718 (N_7718,N_4699,N_5091);
and U7719 (N_7719,N_4579,N_5682);
and U7720 (N_7720,N_5621,N_4772);
or U7721 (N_7721,N_5699,N_4074);
nor U7722 (N_7722,N_4124,N_5976);
nor U7723 (N_7723,N_4401,N_5281);
nand U7724 (N_7724,N_4542,N_4552);
or U7725 (N_7725,N_4322,N_5000);
or U7726 (N_7726,N_4097,N_4027);
or U7727 (N_7727,N_4782,N_4384);
and U7728 (N_7728,N_5850,N_4394);
and U7729 (N_7729,N_4985,N_5087);
or U7730 (N_7730,N_5776,N_4026);
nor U7731 (N_7731,N_5032,N_5335);
xnor U7732 (N_7732,N_4522,N_4257);
or U7733 (N_7733,N_4657,N_4125);
and U7734 (N_7734,N_5070,N_5161);
xor U7735 (N_7735,N_5769,N_4734);
xnor U7736 (N_7736,N_4092,N_4825);
and U7737 (N_7737,N_5471,N_5423);
or U7738 (N_7738,N_5821,N_4029);
xor U7739 (N_7739,N_5727,N_5439);
nor U7740 (N_7740,N_4580,N_4923);
nor U7741 (N_7741,N_4773,N_5092);
and U7742 (N_7742,N_5498,N_4761);
or U7743 (N_7743,N_5093,N_5434);
nand U7744 (N_7744,N_4793,N_5295);
nor U7745 (N_7745,N_5749,N_5592);
nor U7746 (N_7746,N_4356,N_4518);
nand U7747 (N_7747,N_5544,N_5528);
nand U7748 (N_7748,N_5717,N_5735);
and U7749 (N_7749,N_5801,N_5289);
and U7750 (N_7750,N_5470,N_5239);
and U7751 (N_7751,N_5215,N_5079);
xnor U7752 (N_7752,N_5439,N_5923);
and U7753 (N_7753,N_5677,N_5136);
and U7754 (N_7754,N_5432,N_5859);
xnor U7755 (N_7755,N_4690,N_4212);
or U7756 (N_7756,N_4981,N_5280);
and U7757 (N_7757,N_5136,N_5822);
xor U7758 (N_7758,N_5494,N_4955);
nor U7759 (N_7759,N_4284,N_4788);
and U7760 (N_7760,N_5356,N_4091);
nor U7761 (N_7761,N_5026,N_4372);
nand U7762 (N_7762,N_4957,N_4399);
or U7763 (N_7763,N_5514,N_5896);
nand U7764 (N_7764,N_4985,N_4937);
and U7765 (N_7765,N_5153,N_5775);
or U7766 (N_7766,N_4932,N_4992);
xor U7767 (N_7767,N_5126,N_4722);
or U7768 (N_7768,N_4984,N_5003);
and U7769 (N_7769,N_4304,N_4990);
and U7770 (N_7770,N_5045,N_5898);
nor U7771 (N_7771,N_5915,N_5585);
or U7772 (N_7772,N_5134,N_5343);
nand U7773 (N_7773,N_5943,N_5676);
xor U7774 (N_7774,N_4021,N_4586);
and U7775 (N_7775,N_4908,N_5107);
or U7776 (N_7776,N_4788,N_5592);
xor U7777 (N_7777,N_4294,N_5098);
xnor U7778 (N_7778,N_5143,N_5543);
xnor U7779 (N_7779,N_5105,N_4605);
and U7780 (N_7780,N_5757,N_4041);
or U7781 (N_7781,N_5019,N_4071);
xnor U7782 (N_7782,N_4959,N_4519);
and U7783 (N_7783,N_5133,N_5027);
nand U7784 (N_7784,N_4076,N_5012);
nand U7785 (N_7785,N_5804,N_5975);
nand U7786 (N_7786,N_4875,N_5992);
xnor U7787 (N_7787,N_4889,N_5537);
nor U7788 (N_7788,N_5860,N_5088);
nor U7789 (N_7789,N_5626,N_4882);
or U7790 (N_7790,N_5673,N_5414);
xnor U7791 (N_7791,N_4595,N_4469);
and U7792 (N_7792,N_5834,N_5873);
nand U7793 (N_7793,N_5827,N_4697);
xor U7794 (N_7794,N_4411,N_4568);
nor U7795 (N_7795,N_5715,N_5683);
nor U7796 (N_7796,N_5928,N_5744);
xor U7797 (N_7797,N_4523,N_4127);
nor U7798 (N_7798,N_4606,N_5456);
xor U7799 (N_7799,N_4212,N_5871);
or U7800 (N_7800,N_4783,N_5550);
and U7801 (N_7801,N_4785,N_5219);
nand U7802 (N_7802,N_4474,N_4486);
xor U7803 (N_7803,N_5350,N_4674);
xnor U7804 (N_7804,N_4649,N_5181);
and U7805 (N_7805,N_4553,N_4537);
nand U7806 (N_7806,N_4515,N_5985);
or U7807 (N_7807,N_4573,N_5926);
or U7808 (N_7808,N_5195,N_5305);
and U7809 (N_7809,N_4981,N_4477);
nand U7810 (N_7810,N_5054,N_5276);
and U7811 (N_7811,N_5546,N_5588);
or U7812 (N_7812,N_4754,N_5092);
and U7813 (N_7813,N_5654,N_5546);
nor U7814 (N_7814,N_4717,N_4346);
xnor U7815 (N_7815,N_4827,N_4069);
nand U7816 (N_7816,N_5827,N_4734);
nor U7817 (N_7817,N_4939,N_4329);
nand U7818 (N_7818,N_5564,N_4383);
nor U7819 (N_7819,N_4467,N_4764);
and U7820 (N_7820,N_4881,N_4444);
and U7821 (N_7821,N_5422,N_5170);
and U7822 (N_7822,N_4442,N_4828);
nor U7823 (N_7823,N_5555,N_4006);
nor U7824 (N_7824,N_4491,N_4425);
nor U7825 (N_7825,N_4937,N_4083);
nand U7826 (N_7826,N_4143,N_5894);
and U7827 (N_7827,N_5291,N_5207);
xnor U7828 (N_7828,N_4890,N_5414);
and U7829 (N_7829,N_5924,N_4829);
nor U7830 (N_7830,N_5010,N_4097);
or U7831 (N_7831,N_5471,N_5259);
or U7832 (N_7832,N_5924,N_5873);
nand U7833 (N_7833,N_5649,N_5329);
or U7834 (N_7834,N_5108,N_5531);
xnor U7835 (N_7835,N_4063,N_5411);
nor U7836 (N_7836,N_4181,N_5824);
or U7837 (N_7837,N_4285,N_4619);
nand U7838 (N_7838,N_4416,N_4309);
xor U7839 (N_7839,N_4267,N_5406);
and U7840 (N_7840,N_4442,N_4290);
or U7841 (N_7841,N_5541,N_4166);
and U7842 (N_7842,N_4788,N_4685);
xor U7843 (N_7843,N_4851,N_5306);
nor U7844 (N_7844,N_5781,N_5378);
and U7845 (N_7845,N_4731,N_4822);
xnor U7846 (N_7846,N_4349,N_4193);
or U7847 (N_7847,N_5299,N_4576);
xor U7848 (N_7848,N_5134,N_4722);
and U7849 (N_7849,N_5846,N_4356);
and U7850 (N_7850,N_5274,N_4672);
or U7851 (N_7851,N_5167,N_5715);
and U7852 (N_7852,N_4058,N_4629);
xor U7853 (N_7853,N_5437,N_5838);
and U7854 (N_7854,N_4454,N_4044);
nand U7855 (N_7855,N_5903,N_5885);
xor U7856 (N_7856,N_4676,N_5187);
and U7857 (N_7857,N_5451,N_5605);
nand U7858 (N_7858,N_5015,N_5467);
and U7859 (N_7859,N_4567,N_4350);
nor U7860 (N_7860,N_5358,N_5378);
or U7861 (N_7861,N_4335,N_5585);
xor U7862 (N_7862,N_4933,N_4549);
nor U7863 (N_7863,N_4117,N_4310);
xnor U7864 (N_7864,N_4379,N_5737);
xnor U7865 (N_7865,N_5823,N_5386);
or U7866 (N_7866,N_4879,N_5477);
or U7867 (N_7867,N_5280,N_5007);
and U7868 (N_7868,N_4693,N_5552);
nand U7869 (N_7869,N_4582,N_4244);
xnor U7870 (N_7870,N_4245,N_4950);
xnor U7871 (N_7871,N_4170,N_5370);
and U7872 (N_7872,N_4677,N_4361);
nor U7873 (N_7873,N_4041,N_5030);
nand U7874 (N_7874,N_5692,N_5635);
xnor U7875 (N_7875,N_5291,N_4535);
nor U7876 (N_7876,N_4601,N_5137);
nand U7877 (N_7877,N_4372,N_4498);
xor U7878 (N_7878,N_4752,N_4760);
or U7879 (N_7879,N_5647,N_5729);
nand U7880 (N_7880,N_4812,N_5864);
nor U7881 (N_7881,N_5889,N_5493);
nor U7882 (N_7882,N_4958,N_5069);
xnor U7883 (N_7883,N_4156,N_4199);
or U7884 (N_7884,N_5541,N_5588);
and U7885 (N_7885,N_5134,N_5671);
nor U7886 (N_7886,N_4886,N_5462);
or U7887 (N_7887,N_5580,N_5629);
or U7888 (N_7888,N_4182,N_5842);
nor U7889 (N_7889,N_5287,N_5175);
xor U7890 (N_7890,N_5943,N_4030);
and U7891 (N_7891,N_5611,N_5977);
and U7892 (N_7892,N_4013,N_5651);
and U7893 (N_7893,N_4276,N_4913);
nor U7894 (N_7894,N_5909,N_4234);
or U7895 (N_7895,N_5701,N_5872);
and U7896 (N_7896,N_5714,N_4838);
and U7897 (N_7897,N_5538,N_5045);
xor U7898 (N_7898,N_4781,N_4290);
and U7899 (N_7899,N_5027,N_4955);
nor U7900 (N_7900,N_5581,N_4056);
xnor U7901 (N_7901,N_4707,N_4569);
nand U7902 (N_7902,N_4956,N_4677);
xor U7903 (N_7903,N_4747,N_5575);
and U7904 (N_7904,N_5451,N_4810);
nor U7905 (N_7905,N_4957,N_5203);
nand U7906 (N_7906,N_5674,N_4081);
and U7907 (N_7907,N_4419,N_5805);
and U7908 (N_7908,N_5715,N_5793);
nand U7909 (N_7909,N_5963,N_4983);
nand U7910 (N_7910,N_4243,N_4075);
xor U7911 (N_7911,N_4894,N_5708);
nor U7912 (N_7912,N_4424,N_4460);
or U7913 (N_7913,N_4070,N_4940);
nor U7914 (N_7914,N_5336,N_4713);
nor U7915 (N_7915,N_4718,N_4668);
nand U7916 (N_7916,N_5358,N_5329);
xor U7917 (N_7917,N_4696,N_5843);
nor U7918 (N_7918,N_4919,N_4793);
and U7919 (N_7919,N_4479,N_4768);
nor U7920 (N_7920,N_4731,N_5832);
xor U7921 (N_7921,N_4311,N_5410);
or U7922 (N_7922,N_5950,N_4824);
xor U7923 (N_7923,N_5931,N_4455);
nand U7924 (N_7924,N_5481,N_5278);
and U7925 (N_7925,N_5309,N_5007);
or U7926 (N_7926,N_5036,N_5189);
xor U7927 (N_7927,N_5456,N_4164);
and U7928 (N_7928,N_4307,N_4208);
and U7929 (N_7929,N_4132,N_5524);
nor U7930 (N_7930,N_4834,N_5698);
xnor U7931 (N_7931,N_4158,N_4557);
nand U7932 (N_7932,N_5327,N_4949);
or U7933 (N_7933,N_5115,N_5569);
or U7934 (N_7934,N_5106,N_5972);
xnor U7935 (N_7935,N_4503,N_5317);
or U7936 (N_7936,N_4750,N_5156);
nor U7937 (N_7937,N_5469,N_4516);
nor U7938 (N_7938,N_5333,N_4015);
nor U7939 (N_7939,N_5329,N_4623);
xnor U7940 (N_7940,N_5850,N_4879);
nor U7941 (N_7941,N_4211,N_4509);
nand U7942 (N_7942,N_5698,N_4760);
xnor U7943 (N_7943,N_5721,N_5919);
or U7944 (N_7944,N_5224,N_4265);
nor U7945 (N_7945,N_4011,N_5120);
nor U7946 (N_7946,N_4723,N_5050);
xnor U7947 (N_7947,N_4795,N_4846);
xor U7948 (N_7948,N_5337,N_5071);
nor U7949 (N_7949,N_5228,N_5222);
or U7950 (N_7950,N_4669,N_5082);
nand U7951 (N_7951,N_4622,N_4480);
and U7952 (N_7952,N_5182,N_4659);
xnor U7953 (N_7953,N_4962,N_5873);
or U7954 (N_7954,N_5324,N_4923);
or U7955 (N_7955,N_4786,N_5489);
nor U7956 (N_7956,N_5553,N_5663);
xor U7957 (N_7957,N_5751,N_4667);
xnor U7958 (N_7958,N_4296,N_5990);
nand U7959 (N_7959,N_4235,N_4990);
nor U7960 (N_7960,N_5990,N_4937);
xnor U7961 (N_7961,N_5361,N_5017);
nand U7962 (N_7962,N_4109,N_4919);
nand U7963 (N_7963,N_4412,N_4660);
and U7964 (N_7964,N_5607,N_5245);
nand U7965 (N_7965,N_5640,N_4637);
and U7966 (N_7966,N_5027,N_4118);
nand U7967 (N_7967,N_5309,N_4816);
nand U7968 (N_7968,N_4045,N_4777);
xor U7969 (N_7969,N_5379,N_4129);
xnor U7970 (N_7970,N_4109,N_4913);
nor U7971 (N_7971,N_5431,N_5529);
and U7972 (N_7972,N_4403,N_5566);
nand U7973 (N_7973,N_5883,N_4095);
and U7974 (N_7974,N_4256,N_4601);
xor U7975 (N_7975,N_4275,N_5868);
nand U7976 (N_7976,N_4487,N_5576);
nand U7977 (N_7977,N_4173,N_4959);
nand U7978 (N_7978,N_5898,N_4160);
or U7979 (N_7979,N_5192,N_5516);
xnor U7980 (N_7980,N_4794,N_4024);
xnor U7981 (N_7981,N_5853,N_5658);
and U7982 (N_7982,N_4038,N_4150);
nand U7983 (N_7983,N_4517,N_5576);
and U7984 (N_7984,N_5146,N_5206);
or U7985 (N_7985,N_4858,N_5993);
nand U7986 (N_7986,N_5684,N_5958);
nand U7987 (N_7987,N_5911,N_4908);
nand U7988 (N_7988,N_5875,N_5201);
xor U7989 (N_7989,N_4874,N_4067);
or U7990 (N_7990,N_4756,N_4712);
nand U7991 (N_7991,N_5079,N_5572);
nor U7992 (N_7992,N_4243,N_5718);
and U7993 (N_7993,N_4626,N_5276);
nand U7994 (N_7994,N_4534,N_4271);
nor U7995 (N_7995,N_4778,N_4397);
nand U7996 (N_7996,N_4353,N_5435);
or U7997 (N_7997,N_4338,N_5116);
nand U7998 (N_7998,N_4995,N_4036);
xnor U7999 (N_7999,N_4319,N_5295);
and U8000 (N_8000,N_6760,N_6036);
nand U8001 (N_8001,N_6836,N_7642);
and U8002 (N_8002,N_6929,N_7127);
or U8003 (N_8003,N_7148,N_6613);
nand U8004 (N_8004,N_6794,N_7549);
and U8005 (N_8005,N_7825,N_6268);
or U8006 (N_8006,N_7136,N_6704);
nor U8007 (N_8007,N_7230,N_6729);
nor U8008 (N_8008,N_7791,N_7391);
and U8009 (N_8009,N_6712,N_6383);
xor U8010 (N_8010,N_6233,N_7122);
or U8011 (N_8011,N_7857,N_7265);
xnor U8012 (N_8012,N_7451,N_7026);
xor U8013 (N_8013,N_6379,N_7793);
or U8014 (N_8014,N_6719,N_7517);
nor U8015 (N_8015,N_7236,N_7606);
and U8016 (N_8016,N_7344,N_7157);
nor U8017 (N_8017,N_7577,N_6968);
xnor U8018 (N_8018,N_6990,N_7775);
and U8019 (N_8019,N_6981,N_7761);
nor U8020 (N_8020,N_7429,N_7990);
xor U8021 (N_8021,N_6937,N_7578);
and U8022 (N_8022,N_6798,N_7333);
and U8023 (N_8023,N_7605,N_6894);
nor U8024 (N_8024,N_6955,N_7471);
xor U8025 (N_8025,N_7010,N_6009);
xnor U8026 (N_8026,N_7315,N_7591);
nand U8027 (N_8027,N_6427,N_6634);
or U8028 (N_8028,N_6530,N_6102);
or U8029 (N_8029,N_7670,N_7497);
or U8030 (N_8030,N_7530,N_7736);
nand U8031 (N_8031,N_7334,N_6272);
nor U8032 (N_8032,N_6576,N_7361);
and U8033 (N_8033,N_6607,N_7755);
and U8034 (N_8034,N_6092,N_7760);
and U8035 (N_8035,N_6595,N_7522);
xnor U8036 (N_8036,N_6288,N_6062);
nor U8037 (N_8037,N_6480,N_7741);
and U8038 (N_8038,N_7737,N_7149);
xor U8039 (N_8039,N_7051,N_7563);
and U8040 (N_8040,N_7012,N_6557);
xnor U8041 (N_8041,N_6289,N_6965);
and U8042 (N_8042,N_7986,N_6699);
nand U8043 (N_8043,N_7652,N_7327);
nor U8044 (N_8044,N_7330,N_7102);
and U8045 (N_8045,N_6481,N_7116);
xnor U8046 (N_8046,N_7616,N_7464);
nand U8047 (N_8047,N_7831,N_6916);
or U8048 (N_8048,N_7194,N_6763);
or U8049 (N_8049,N_7679,N_6204);
nand U8050 (N_8050,N_7492,N_7185);
xor U8051 (N_8051,N_7800,N_6360);
and U8052 (N_8052,N_7463,N_7699);
nor U8053 (N_8053,N_7768,N_7725);
nand U8054 (N_8054,N_6469,N_7233);
nand U8055 (N_8055,N_6920,N_7034);
or U8056 (N_8056,N_7664,N_6168);
and U8057 (N_8057,N_7774,N_6215);
xor U8058 (N_8058,N_7139,N_6787);
or U8059 (N_8059,N_7974,N_7628);
xor U8060 (N_8060,N_7897,N_6389);
nor U8061 (N_8061,N_6082,N_7573);
xor U8062 (N_8062,N_7908,N_7917);
nor U8063 (N_8063,N_6142,N_6212);
or U8064 (N_8064,N_7106,N_6335);
or U8065 (N_8065,N_6552,N_7830);
and U8066 (N_8066,N_6477,N_7469);
xor U8067 (N_8067,N_6733,N_6474);
and U8068 (N_8068,N_7306,N_6216);
or U8069 (N_8069,N_7581,N_6198);
and U8070 (N_8070,N_6554,N_6495);
or U8071 (N_8071,N_6878,N_6718);
xor U8072 (N_8072,N_7502,N_7883);
and U8073 (N_8073,N_7217,N_6635);
or U8074 (N_8074,N_7686,N_6988);
or U8075 (N_8075,N_7702,N_6522);
nand U8076 (N_8076,N_6182,N_7526);
nor U8077 (N_8077,N_7131,N_6121);
nor U8078 (N_8078,N_7576,N_7049);
and U8079 (N_8079,N_6592,N_6668);
nand U8080 (N_8080,N_7602,N_6166);
xor U8081 (N_8081,N_6919,N_7952);
xor U8082 (N_8082,N_7767,N_7704);
and U8083 (N_8083,N_7023,N_6374);
nor U8084 (N_8084,N_6282,N_6447);
and U8085 (N_8085,N_7337,N_7872);
xor U8086 (N_8086,N_7675,N_6912);
xor U8087 (N_8087,N_7635,N_7209);
or U8088 (N_8088,N_7821,N_6609);
xor U8089 (N_8089,N_7382,N_7164);
and U8090 (N_8090,N_6870,N_6663);
xnor U8091 (N_8091,N_6029,N_7972);
nand U8092 (N_8092,N_6783,N_7044);
nand U8093 (N_8093,N_6779,N_7389);
xnor U8094 (N_8094,N_7622,N_7846);
xor U8095 (N_8095,N_7600,N_7251);
and U8096 (N_8096,N_6297,N_7826);
xnor U8097 (N_8097,N_7575,N_7143);
nor U8098 (N_8098,N_7071,N_7880);
and U8099 (N_8099,N_6568,N_6349);
or U8100 (N_8100,N_6569,N_6977);
xnor U8101 (N_8101,N_7811,N_7415);
xnor U8102 (N_8102,N_7910,N_6337);
and U8103 (N_8103,N_6115,N_7873);
nand U8104 (N_8104,N_6502,N_6854);
xor U8105 (N_8105,N_6243,N_7968);
nor U8106 (N_8106,N_7351,N_7216);
xor U8107 (N_8107,N_7716,N_7903);
nand U8108 (N_8108,N_6433,N_7085);
xor U8109 (N_8109,N_6016,N_7850);
and U8110 (N_8110,N_7483,N_7435);
and U8111 (N_8111,N_6695,N_6581);
xnor U8112 (N_8112,N_7640,N_7863);
nand U8113 (N_8113,N_6726,N_7020);
xnor U8114 (N_8114,N_7611,N_6853);
and U8115 (N_8115,N_7944,N_6253);
xnor U8116 (N_8116,N_6312,N_7182);
nor U8117 (N_8117,N_7130,N_7884);
or U8118 (N_8118,N_6037,N_6890);
or U8119 (N_8119,N_6943,N_7378);
and U8120 (N_8120,N_7158,N_7824);
xor U8121 (N_8121,N_7356,N_7015);
nand U8122 (N_8122,N_7173,N_7776);
nor U8123 (N_8123,N_6597,N_6367);
and U8124 (N_8124,N_7866,N_6621);
xnor U8125 (N_8125,N_7519,N_6318);
or U8126 (N_8126,N_7346,N_7156);
or U8127 (N_8127,N_7171,N_6347);
nor U8128 (N_8128,N_7203,N_7060);
or U8129 (N_8129,N_7103,N_6294);
or U8130 (N_8130,N_7543,N_6336);
and U8131 (N_8131,N_6227,N_6651);
nand U8132 (N_8132,N_6299,N_7264);
and U8133 (N_8133,N_7545,N_6584);
and U8134 (N_8134,N_7078,N_6610);
xor U8135 (N_8135,N_6490,N_7927);
nand U8136 (N_8136,N_6966,N_7095);
or U8137 (N_8137,N_7410,N_7646);
or U8138 (N_8138,N_7252,N_7763);
xor U8139 (N_8139,N_6775,N_7003);
and U8140 (N_8140,N_7262,N_7960);
nor U8141 (N_8141,N_6366,N_7542);
or U8142 (N_8142,N_7208,N_7630);
nor U8143 (N_8143,N_7552,N_7401);
or U8144 (N_8144,N_7007,N_7281);
nor U8145 (N_8145,N_6744,N_6542);
xnor U8146 (N_8146,N_7181,N_7461);
xnor U8147 (N_8147,N_6834,N_7744);
or U8148 (N_8148,N_6135,N_6317);
and U8149 (N_8149,N_7282,N_7115);
xnor U8150 (N_8150,N_6230,N_7393);
xor U8151 (N_8151,N_7387,N_6580);
or U8152 (N_8152,N_6618,N_6112);
or U8153 (N_8153,N_7887,N_7810);
xnor U8154 (N_8154,N_6326,N_6371);
and U8155 (N_8155,N_6386,N_6908);
nand U8156 (N_8156,N_6298,N_6202);
or U8157 (N_8157,N_7627,N_6039);
nor U8158 (N_8158,N_6922,N_7144);
or U8159 (N_8159,N_7154,N_6857);
or U8160 (N_8160,N_6874,N_6756);
nand U8161 (N_8161,N_6363,N_6497);
nor U8162 (N_8162,N_6641,N_7677);
or U8163 (N_8163,N_7256,N_7397);
and U8164 (N_8164,N_7042,N_7478);
xnor U8165 (N_8165,N_6440,N_6285);
or U8166 (N_8166,N_7822,N_6707);
nand U8167 (N_8167,N_6746,N_6616);
nand U8168 (N_8168,N_7762,N_7341);
nor U8169 (N_8169,N_6333,N_6703);
and U8170 (N_8170,N_7091,N_7817);
nor U8171 (N_8171,N_7304,N_7260);
or U8172 (N_8172,N_7257,N_6833);
nand U8173 (N_8173,N_6509,N_6883);
xor U8174 (N_8174,N_6117,N_6263);
nor U8175 (N_8175,N_6862,N_6657);
and U8176 (N_8176,N_7503,N_7877);
nor U8177 (N_8177,N_6698,N_6023);
nand U8178 (N_8178,N_6751,N_6287);
and U8179 (N_8179,N_6515,N_6239);
xor U8180 (N_8180,N_7609,N_7384);
nor U8181 (N_8181,N_6560,N_6740);
nor U8182 (N_8182,N_7970,N_6742);
nand U8183 (N_8183,N_7058,N_6021);
or U8184 (N_8184,N_6049,N_7321);
nor U8185 (N_8185,N_6661,N_6627);
and U8186 (N_8186,N_6748,N_6544);
and U8187 (N_8187,N_7374,N_6197);
or U8188 (N_8188,N_6348,N_6320);
and U8189 (N_8189,N_6632,N_6681);
xor U8190 (N_8190,N_7859,N_6653);
or U8191 (N_8191,N_6801,N_6717);
or U8192 (N_8192,N_6210,N_6761);
or U8193 (N_8193,N_7184,N_6310);
nand U8194 (N_8194,N_7816,N_7929);
or U8195 (N_8195,N_7739,N_7275);
nor U8196 (N_8196,N_7660,N_6517);
xor U8197 (N_8197,N_7982,N_7062);
and U8198 (N_8198,N_7566,N_7721);
or U8199 (N_8199,N_6057,N_7661);
nor U8200 (N_8200,N_7047,N_7514);
or U8201 (N_8201,N_6601,N_7644);
xor U8202 (N_8202,N_7889,N_7586);
and U8203 (N_8203,N_6405,N_7898);
or U8204 (N_8204,N_7211,N_6421);
and U8205 (N_8205,N_7249,N_7707);
nor U8206 (N_8206,N_6242,N_6437);
nor U8207 (N_8207,N_6265,N_7740);
or U8208 (N_8208,N_6626,N_6945);
or U8209 (N_8209,N_7009,N_7924);
or U8210 (N_8210,N_6031,N_6940);
xnor U8211 (N_8211,N_6078,N_7786);
or U8212 (N_8212,N_7842,N_7562);
xnor U8213 (N_8213,N_6255,N_7004);
and U8214 (N_8214,N_7326,N_6871);
xor U8215 (N_8215,N_6593,N_6532);
and U8216 (N_8216,N_7806,N_7367);
xor U8217 (N_8217,N_7915,N_6629);
nor U8218 (N_8218,N_6088,N_7777);
nor U8219 (N_8219,N_7297,N_7520);
or U8220 (N_8220,N_6162,N_7293);
nor U8221 (N_8221,N_7146,N_7134);
and U8222 (N_8222,N_7608,N_6460);
nor U8223 (N_8223,N_7765,N_7390);
or U8224 (N_8224,N_6806,N_7662);
nand U8225 (N_8225,N_6973,N_7162);
and U8226 (N_8226,N_7723,N_7967);
nor U8227 (N_8227,N_7727,N_6244);
nand U8228 (N_8228,N_6847,N_7829);
xor U8229 (N_8229,N_7213,N_6054);
xor U8230 (N_8230,N_6611,N_6582);
xnor U8231 (N_8231,N_7681,N_6464);
nand U8232 (N_8232,N_6047,N_6482);
nor U8233 (N_8233,N_7784,N_6248);
nor U8234 (N_8234,N_7920,N_6165);
nand U8235 (N_8235,N_6643,N_6511);
xor U8236 (N_8236,N_6174,N_7813);
xnor U8237 (N_8237,N_7244,N_7518);
nand U8238 (N_8238,N_7750,N_7094);
nand U8239 (N_8239,N_7035,N_7205);
nor U8240 (N_8240,N_7687,N_6391);
and U8241 (N_8241,N_6208,N_6205);
or U8242 (N_8242,N_6426,N_6076);
nand U8243 (N_8243,N_7432,N_7731);
and U8244 (N_8244,N_7779,N_6504);
and U8245 (N_8245,N_6796,N_7076);
and U8246 (N_8246,N_7352,N_6368);
nand U8247 (N_8247,N_6987,N_6789);
or U8248 (N_8248,N_7964,N_7104);
xor U8249 (N_8249,N_7037,N_7837);
nand U8250 (N_8250,N_7939,N_7419);
nor U8251 (N_8251,N_6066,N_7701);
and U8252 (N_8252,N_7521,N_6434);
nor U8253 (N_8253,N_6927,N_6290);
nand U8254 (N_8254,N_6868,N_7882);
xor U8255 (N_8255,N_6415,N_6984);
xor U8256 (N_8256,N_6279,N_7900);
xnor U8257 (N_8257,N_6266,N_7947);
nand U8258 (N_8258,N_7240,N_6065);
xnor U8259 (N_8259,N_6025,N_7796);
nand U8260 (N_8260,N_6491,N_7992);
xnor U8261 (N_8261,N_7220,N_6694);
xnor U8262 (N_8262,N_7331,N_7589);
xnor U8263 (N_8263,N_6455,N_6328);
nor U8264 (N_8264,N_7153,N_7730);
or U8265 (N_8265,N_7500,N_6218);
xor U8266 (N_8266,N_7224,N_7703);
or U8267 (N_8267,N_6808,N_7250);
or U8268 (N_8268,N_7133,N_7090);
nor U8269 (N_8269,N_7467,N_7450);
or U8270 (N_8270,N_6633,N_7676);
or U8271 (N_8271,N_6251,N_6714);
nor U8272 (N_8272,N_6624,N_6046);
and U8273 (N_8273,N_6045,N_6267);
and U8274 (N_8274,N_7803,N_7945);
and U8275 (N_8275,N_7234,N_6380);
nand U8276 (N_8276,N_6416,N_7038);
xnor U8277 (N_8277,N_6083,N_7486);
and U8278 (N_8278,N_7527,N_7089);
nor U8279 (N_8279,N_6068,N_6399);
and U8280 (N_8280,N_7465,N_6193);
and U8281 (N_8281,N_6252,N_7183);
xnor U8282 (N_8282,N_6479,N_7443);
nand U8283 (N_8283,N_7700,N_6483);
or U8284 (N_8284,N_6799,N_6106);
xnor U8285 (N_8285,N_7350,N_6030);
xnor U8286 (N_8286,N_6234,N_7436);
nand U8287 (N_8287,N_7061,N_6180);
nor U8288 (N_8288,N_6369,N_7266);
nand U8289 (N_8289,N_6505,N_7040);
nor U8290 (N_8290,N_6444,N_7501);
nor U8291 (N_8291,N_6586,N_7879);
or U8292 (N_8292,N_6989,N_7749);
nand U8293 (N_8293,N_7312,N_7834);
xnor U8294 (N_8294,N_7787,N_7305);
or U8295 (N_8295,N_6867,N_6113);
nand U8296 (N_8296,N_7229,N_6978);
xnor U8297 (N_8297,N_7655,N_6488);
and U8298 (N_8298,N_7869,N_6196);
nor U8299 (N_8299,N_7358,N_6710);
or U8300 (N_8300,N_7567,N_6144);
xor U8301 (N_8301,N_7174,N_6866);
nand U8302 (N_8302,N_6343,N_7316);
nand U8303 (N_8303,N_6956,N_7400);
and U8304 (N_8304,N_6848,N_6716);
nand U8305 (N_8305,N_6508,N_6075);
and U8306 (N_8306,N_7757,N_6010);
nand U8307 (N_8307,N_6456,N_6201);
xor U8308 (N_8308,N_7011,N_7099);
xnor U8309 (N_8309,N_7215,N_6492);
nand U8310 (N_8310,N_7114,N_7693);
nand U8311 (N_8311,N_6501,N_6750);
or U8312 (N_8312,N_7618,N_7176);
and U8313 (N_8313,N_7325,N_7409);
nor U8314 (N_8314,N_7385,N_6758);
nand U8315 (N_8315,N_6003,N_6468);
and U8316 (N_8316,N_7999,N_6686);
xnor U8317 (N_8317,N_6818,N_7854);
xor U8318 (N_8318,N_6462,N_7766);
and U8319 (N_8319,N_6048,N_6553);
xnor U8320 (N_8320,N_7446,N_7150);
xor U8321 (N_8321,N_6089,N_7491);
or U8322 (N_8322,N_6177,N_7674);
or U8323 (N_8323,N_6425,N_6189);
xnor U8324 (N_8324,N_7783,N_6124);
xor U8325 (N_8325,N_7663,N_6362);
nand U8326 (N_8326,N_7444,N_6013);
nor U8327 (N_8327,N_7938,N_7033);
xnor U8328 (N_8328,N_6953,N_6295);
and U8329 (N_8329,N_7018,N_7287);
and U8330 (N_8330,N_7084,N_7864);
nor U8331 (N_8331,N_6932,N_6804);
nor U8332 (N_8332,N_7805,N_6564);
xnor U8333 (N_8333,N_6947,N_6478);
or U8334 (N_8334,N_6667,N_6388);
nand U8335 (N_8335,N_7484,N_7568);
xor U8336 (N_8336,N_7392,N_7504);
or U8337 (N_8337,N_7665,N_7083);
or U8338 (N_8338,N_6536,N_7347);
nor U8339 (N_8339,N_6178,N_6538);
nor U8340 (N_8340,N_7571,N_7685);
nor U8341 (N_8341,N_6518,N_7141);
xor U8342 (N_8342,N_6005,N_6123);
nor U8343 (N_8343,N_6543,N_7862);
and U8344 (N_8344,N_6837,N_6731);
nor U8345 (N_8345,N_6708,N_6452);
or U8346 (N_8346,N_7402,N_6454);
nand U8347 (N_8347,N_7780,N_7554);
xnor U8348 (N_8348,N_7057,N_6350);
xor U8349 (N_8349,N_7666,N_6158);
and U8350 (N_8350,N_7289,N_6228);
xnor U8351 (N_8351,N_7557,N_6845);
nand U8352 (N_8352,N_7291,N_6514);
nor U8353 (N_8353,N_7838,N_6438);
xor U8354 (N_8354,N_6156,N_7943);
nor U8355 (N_8355,N_6306,N_7770);
and U8356 (N_8356,N_7546,N_6160);
xor U8357 (N_8357,N_6644,N_6291);
nand U8358 (N_8358,N_6428,N_6258);
nand U8359 (N_8359,N_7868,N_6939);
or U8360 (N_8360,N_7511,N_6222);
or U8361 (N_8361,N_7029,N_6110);
xnor U8362 (N_8362,N_7186,N_6126);
nor U8363 (N_8363,N_6418,N_6527);
nor U8364 (N_8364,N_7457,N_6407);
or U8365 (N_8365,N_6942,N_6241);
xor U8366 (N_8366,N_6506,N_7626);
or U8367 (N_8367,N_6771,N_7790);
or U8368 (N_8368,N_6463,N_7911);
nand U8369 (N_8369,N_6614,N_6175);
or U8370 (N_8370,N_6043,N_7189);
xnor U8371 (N_8371,N_6225,N_6958);
and U8372 (N_8372,N_7547,N_7909);
and U8373 (N_8373,N_7081,N_6419);
xor U8374 (N_8374,N_6356,N_6302);
xor U8375 (N_8375,N_7993,N_6286);
and U8376 (N_8376,N_6622,N_7441);
or U8377 (N_8377,N_7753,N_6843);
xnor U8378 (N_8378,N_6963,N_7523);
and U8379 (N_8379,N_7548,N_6476);
xnor U8380 (N_8380,N_6666,N_6090);
and U8381 (N_8381,N_7550,N_6959);
nand U8382 (N_8382,N_6293,N_7764);
nor U8383 (N_8383,N_6727,N_7695);
and U8384 (N_8384,N_6820,N_7930);
nand U8385 (N_8385,N_6807,N_7498);
nand U8386 (N_8386,N_6145,N_7191);
and U8387 (N_8387,N_6019,N_7207);
and U8388 (N_8388,N_7473,N_6974);
and U8389 (N_8389,N_7232,N_7420);
and U8390 (N_8390,N_7241,N_7560);
nand U8391 (N_8391,N_6612,N_7294);
nor U8392 (N_8392,N_6520,N_6675);
xnor U8393 (N_8393,N_6809,N_7319);
nor U8394 (N_8394,N_7769,N_7894);
nor U8395 (N_8395,N_6884,N_7659);
or U8396 (N_8396,N_7980,N_6101);
nor U8397 (N_8397,N_6277,N_6720);
and U8398 (N_8398,N_6948,N_7427);
nand U8399 (N_8399,N_6946,N_7610);
xnor U8400 (N_8400,N_6640,N_7778);
nand U8401 (N_8401,N_6998,N_6986);
and U8402 (N_8402,N_7978,N_6450);
nor U8403 (N_8403,N_7537,N_7603);
xnor U8404 (N_8404,N_6015,N_6994);
nor U8405 (N_8405,N_6556,N_6376);
xnor U8406 (N_8406,N_7735,N_6898);
or U8407 (N_8407,N_6394,N_6417);
or U8408 (N_8408,N_7671,N_6623);
nor U8409 (N_8409,N_6930,N_6143);
xor U8410 (N_8410,N_6097,N_7629);
or U8411 (N_8411,N_7430,N_7407);
and U8412 (N_8412,N_6603,N_6436);
and U8413 (N_8413,N_7533,N_7614);
or U8414 (N_8414,N_6677,N_7353);
xnor U8415 (N_8415,N_6096,N_7905);
xor U8416 (N_8416,N_6402,N_7615);
or U8417 (N_8417,N_6952,N_7445);
xor U8418 (N_8418,N_6431,N_6964);
nor U8419 (N_8419,N_7277,N_7795);
nor U8420 (N_8420,N_7070,N_6207);
nand U8421 (N_8421,N_6654,N_6274);
and U8422 (N_8422,N_7544,N_6551);
nand U8423 (N_8423,N_6683,N_7206);
and U8424 (N_8424,N_6381,N_7273);
or U8425 (N_8425,N_7455,N_7155);
or U8426 (N_8426,N_7957,N_6052);
and U8427 (N_8427,N_7468,N_7950);
nor U8428 (N_8428,N_6697,N_7098);
or U8429 (N_8429,N_7604,N_7195);
or U8430 (N_8430,N_7654,N_6249);
or U8431 (N_8431,N_6264,N_7271);
nand U8432 (N_8432,N_7891,N_6678);
or U8433 (N_8433,N_6035,N_6849);
nor U8434 (N_8434,N_6034,N_6038);
nand U8435 (N_8435,N_7657,N_6770);
nand U8436 (N_8436,N_7798,N_7794);
or U8437 (N_8437,N_7583,N_6192);
nor U8438 (N_8438,N_6445,N_6014);
nor U8439 (N_8439,N_7988,N_7188);
nand U8440 (N_8440,N_6615,N_7893);
nand U8441 (N_8441,N_6103,N_6313);
nand U8442 (N_8442,N_7984,N_7414);
or U8443 (N_8443,N_7395,N_6459);
or U8444 (N_8444,N_7454,N_6133);
or U8445 (N_8445,N_6442,N_6850);
nand U8446 (N_8446,N_6766,N_7585);
nor U8447 (N_8447,N_6276,N_7120);
nand U8448 (N_8448,N_7895,N_6583);
xnor U8449 (N_8449,N_7717,N_7222);
xor U8450 (N_8450,N_6131,N_6390);
xor U8451 (N_8451,N_7074,N_7555);
nand U8452 (N_8452,N_7733,N_6283);
and U8453 (N_8453,N_7138,N_6194);
nor U8454 (N_8454,N_7332,N_7310);
xor U8455 (N_8455,N_7223,N_7607);
nand U8456 (N_8456,N_7386,N_7705);
and U8457 (N_8457,N_7752,N_6100);
and U8458 (N_8458,N_6709,N_7792);
or U8459 (N_8459,N_6221,N_6649);
or U8460 (N_8460,N_6831,N_7204);
and U8461 (N_8461,N_7052,N_6600);
or U8462 (N_8462,N_6879,N_6358);
xor U8463 (N_8463,N_6602,N_6254);
or U8464 (N_8464,N_6385,N_7914);
and U8465 (N_8465,N_6108,N_6599);
and U8466 (N_8466,N_6278,N_6510);
xor U8467 (N_8467,N_7166,N_6687);
nor U8468 (N_8468,N_6410,N_6688);
nor U8469 (N_8469,N_6590,N_6852);
nand U8470 (N_8470,N_7270,N_7132);
or U8471 (N_8471,N_7975,N_7192);
nor U8472 (N_8472,N_6396,N_7480);
nor U8473 (N_8473,N_7449,N_6059);
or U8474 (N_8474,N_6921,N_7918);
nor U8475 (N_8475,N_6087,N_7565);
and U8476 (N_8476,N_6020,N_6665);
and U8477 (N_8477,N_6296,N_7963);
or U8478 (N_8478,N_6420,N_7147);
xor U8479 (N_8479,N_6472,N_6400);
nor U8480 (N_8480,N_7118,N_7933);
or U8481 (N_8481,N_6545,N_6658);
xor U8482 (N_8482,N_7021,N_6475);
or U8483 (N_8483,N_7403,N_7899);
xnor U8484 (N_8484,N_7027,N_7954);
and U8485 (N_8485,N_7802,N_6872);
xnor U8486 (N_8486,N_7376,N_7849);
or U8487 (N_8487,N_6821,N_7499);
xnor U8488 (N_8488,N_6606,N_6992);
or U8489 (N_8489,N_7743,N_6315);
or U8490 (N_8490,N_6967,N_7167);
or U8491 (N_8491,N_6753,N_6997);
or U8492 (N_8492,N_6918,N_7828);
nor U8493 (N_8493,N_6361,N_6637);
and U8494 (N_8494,N_6625,N_7558);
or U8495 (N_8495,N_6487,N_7948);
nor U8496 (N_8496,N_7688,N_6304);
and U8497 (N_8497,N_7474,N_7667);
nand U8498 (N_8498,N_6811,N_7039);
and U8499 (N_8499,N_6069,N_6067);
nor U8500 (N_8500,N_6261,N_6149);
and U8501 (N_8501,N_6713,N_6896);
nor U8502 (N_8502,N_6702,N_7683);
or U8503 (N_8503,N_7845,N_7551);
and U8504 (N_8504,N_7758,N_6881);
xor U8505 (N_8505,N_6764,N_6200);
xnor U8506 (N_8506,N_6167,N_6790);
nand U8507 (N_8507,N_6684,N_7263);
and U8508 (N_8508,N_7177,N_6140);
or U8509 (N_8509,N_6863,N_6245);
nor U8510 (N_8510,N_6095,N_6503);
xnor U8511 (N_8511,N_6188,N_7756);
nor U8512 (N_8512,N_7534,N_6840);
and U8513 (N_8513,N_6851,N_7937);
xor U8514 (N_8514,N_7729,N_7276);
xor U8515 (N_8515,N_7073,N_6646);
nand U8516 (N_8516,N_7482,N_7309);
nor U8517 (N_8517,N_7564,N_6860);
and U8518 (N_8518,N_6519,N_6961);
or U8519 (N_8519,N_6886,N_6949);
xor U8520 (N_8520,N_7338,N_6535);
and U8521 (N_8521,N_7570,N_7109);
xor U8522 (N_8522,N_6555,N_6319);
nor U8523 (N_8523,N_7710,N_6938);
or U8524 (N_8524,N_6835,N_7272);
nand U8525 (N_8525,N_6673,N_7801);
nand U8526 (N_8526,N_7231,N_7137);
or U8527 (N_8527,N_6706,N_7372);
and U8528 (N_8528,N_7279,N_7125);
xnor U8529 (N_8529,N_7528,N_6524);
nand U8530 (N_8530,N_6042,N_7019);
nor U8531 (N_8531,N_6864,N_6563);
and U8532 (N_8532,N_6004,N_7298);
nand U8533 (N_8533,N_6589,N_6724);
nor U8534 (N_8534,N_7080,N_7966);
nor U8535 (N_8535,N_6181,N_6220);
or U8536 (N_8536,N_6786,N_7307);
nor U8537 (N_8537,N_6715,N_7690);
and U8538 (N_8538,N_7969,N_7151);
xor U8539 (N_8539,N_7935,N_7175);
or U8540 (N_8540,N_7008,N_7101);
nand U8541 (N_8541,N_6723,N_7302);
nand U8542 (N_8542,N_6271,N_6122);
nand U8543 (N_8543,N_6734,N_6539);
xor U8544 (N_8544,N_6690,N_6301);
nor U8545 (N_8545,N_6755,N_7274);
or U8546 (N_8546,N_7673,N_6936);
and U8547 (N_8547,N_6824,N_7906);
nor U8548 (N_8548,N_7582,N_7301);
or U8549 (N_8549,N_7043,N_7433);
nor U8550 (N_8550,N_7363,N_7199);
and U8551 (N_8551,N_7013,N_7732);
xnor U8552 (N_8552,N_6594,N_7054);
nor U8553 (N_8553,N_6050,N_6950);
or U8554 (N_8554,N_6179,N_7242);
or U8555 (N_8555,N_6061,N_7470);
xor U8556 (N_8556,N_7595,N_6570);
nand U8557 (N_8557,N_6591,N_7934);
nor U8558 (N_8558,N_6473,N_6888);
xnor U8559 (N_8559,N_7371,N_7283);
or U8560 (N_8560,N_7985,N_7005);
or U8561 (N_8561,N_7902,N_6769);
nand U8562 (N_8562,N_6772,N_7092);
xor U8563 (N_8563,N_6063,N_7682);
and U8564 (N_8564,N_7643,N_7324);
or U8565 (N_8565,N_7152,N_7773);
xor U8566 (N_8566,N_6211,N_6044);
or U8567 (N_8567,N_6325,N_6485);
xnor U8568 (N_8568,N_7738,N_6040);
nand U8569 (N_8569,N_6983,N_7759);
xor U8570 (N_8570,N_7921,N_6493);
or U8571 (N_8571,N_6905,N_7226);
and U8572 (N_8572,N_7587,N_7785);
and U8573 (N_8573,N_7812,N_7841);
or U8574 (N_8574,N_7525,N_6074);
xnor U8575 (N_8575,N_6105,N_6841);
or U8576 (N_8576,N_6002,N_6001);
nor U8577 (N_8577,N_7031,N_6334);
xnor U8578 (N_8578,N_7653,N_7979);
or U8579 (N_8579,N_7329,N_6338);
xnor U8580 (N_8580,N_6669,N_6674);
xor U8581 (N_8581,N_6907,N_7079);
nor U8582 (N_8582,N_7179,N_7065);
nand U8583 (N_8583,N_7269,N_7580);
nor U8584 (N_8584,N_7941,N_7965);
nor U8585 (N_8585,N_6164,N_6127);
or U8586 (N_8586,N_7995,N_7028);
and U8587 (N_8587,N_7314,N_7366);
nand U8588 (N_8588,N_6012,N_7159);
or U8589 (N_8589,N_7932,N_7645);
nand U8590 (N_8590,N_7772,N_6280);
or U8591 (N_8591,N_7442,N_6534);
or U8592 (N_8592,N_7067,N_6671);
xor U8593 (N_8593,N_7823,N_6055);
xor U8594 (N_8594,N_6214,N_7505);
nand U8595 (N_8595,N_6257,N_7976);
and U8596 (N_8596,N_7197,N_6909);
nor U8597 (N_8597,N_6782,N_6639);
nand U8598 (N_8598,N_7926,N_6757);
and U8599 (N_8599,N_6439,N_6846);
nor U8600 (N_8600,N_6153,N_7870);
nand U8601 (N_8601,N_6403,N_7145);
xnor U8602 (N_8602,N_6813,N_6951);
nor U8603 (N_8603,N_6507,N_6759);
and U8604 (N_8604,N_6136,N_7355);
nand U8605 (N_8605,N_7459,N_7201);
and U8606 (N_8606,N_7068,N_7658);
xnor U8607 (N_8607,N_6575,N_6270);
or U8608 (N_8608,N_6784,N_6887);
xor U8609 (N_8609,N_7292,N_6027);
or U8610 (N_8610,N_6924,N_6979);
nor U8611 (N_8611,N_6281,N_7165);
and U8612 (N_8612,N_6893,N_6605);
and U8613 (N_8613,N_7405,N_7875);
or U8614 (N_8614,N_6081,N_7408);
nor U8615 (N_8615,N_7851,N_7448);
xor U8616 (N_8616,N_6026,N_7135);
nand U8617 (N_8617,N_7977,N_6899);
nand U8618 (N_8618,N_7267,N_7804);
nand U8619 (N_8619,N_6780,N_7025);
and U8620 (N_8620,N_6917,N_6330);
and U8621 (N_8621,N_7340,N_7063);
xor U8622 (N_8622,N_7107,N_7190);
or U8623 (N_8623,N_7633,N_7286);
and U8624 (N_8624,N_7170,N_6696);
and U8625 (N_8625,N_7048,N_6976);
or U8626 (N_8626,N_7513,N_7874);
and U8627 (N_8627,N_7839,N_7623);
nand U8628 (N_8628,N_6224,N_6231);
or U8629 (N_8629,N_6926,N_6754);
and U8630 (N_8630,N_6645,N_7261);
xor U8631 (N_8631,N_7259,N_6762);
and U8632 (N_8632,N_7055,N_7989);
nand U8633 (N_8633,N_7524,N_6559);
or U8634 (N_8634,N_7412,N_7247);
nand U8635 (N_8635,N_7509,N_6980);
nor U8636 (N_8636,N_7650,N_7858);
nand U8637 (N_8637,N_6148,N_7856);
nor U8638 (N_8638,N_6397,N_7540);
or U8639 (N_8639,N_6869,N_6341);
nand U8640 (N_8640,N_7904,N_7246);
nand U8641 (N_8641,N_7064,N_7187);
xnor U8642 (N_8642,N_7434,N_7477);
and U8643 (N_8643,N_6838,N_7097);
or U8644 (N_8644,N_7239,N_7913);
xnor U8645 (N_8645,N_6232,N_7620);
nor U8646 (N_8646,N_6284,N_7510);
nand U8647 (N_8647,N_6596,N_6387);
xnor U8648 (N_8648,N_6457,N_7431);
and U8649 (N_8649,N_6414,N_7452);
xnor U8650 (N_8650,N_7364,N_6537);
and U8651 (N_8651,N_7077,N_7840);
nor U8652 (N_8652,N_6091,N_6512);
or U8653 (N_8653,N_7647,N_7559);
xnor U8654 (N_8654,N_6941,N_7592);
xnor U8655 (N_8655,N_7819,N_6154);
nand U8656 (N_8656,N_6996,N_6778);
and U8657 (N_8657,N_7715,N_6747);
and U8658 (N_8658,N_7508,N_7308);
nor U8659 (N_8659,N_7886,N_6650);
and U8660 (N_8660,N_7598,N_7493);
nand U8661 (N_8661,N_6017,N_6152);
and U8662 (N_8662,N_6359,N_7956);
xnor U8663 (N_8663,N_6785,N_6238);
nand U8664 (N_8664,N_7072,N_6107);
nor U8665 (N_8665,N_6705,N_6453);
and U8666 (N_8666,N_6486,N_6546);
nor U8667 (N_8667,N_7258,N_7348);
or U8668 (N_8668,N_6229,N_6209);
or U8669 (N_8669,N_7722,N_6139);
or U8670 (N_8670,N_6931,N_6372);
and U8671 (N_8671,N_7489,N_7439);
xnor U8672 (N_8672,N_7649,N_7680);
xor U8673 (N_8673,N_7128,N_6256);
or U8674 (N_8674,N_6412,N_7601);
xor U8675 (N_8675,N_6913,N_6119);
nor U8676 (N_8676,N_6300,N_7121);
xnor U8677 (N_8677,N_7782,N_7714);
xnor U8678 (N_8678,N_6985,N_7593);
nand U8679 (N_8679,N_7745,N_7219);
nand U8680 (N_8680,N_6885,N_7368);
and U8681 (N_8681,N_7867,N_7971);
nand U8682 (N_8682,N_6470,N_6411);
nor U8683 (N_8683,N_6353,N_7169);
and U8684 (N_8684,N_7030,N_6880);
nand U8685 (N_8685,N_7360,N_6316);
nand U8686 (N_8686,N_7100,N_7789);
and U8687 (N_8687,N_7200,N_7142);
and U8688 (N_8688,N_6170,N_6911);
nand U8689 (N_8689,N_7692,N_7050);
nand U8690 (N_8690,N_6173,N_7637);
nor U8691 (N_8691,N_7268,N_6079);
and U8692 (N_8692,N_6865,N_6814);
and U8693 (N_8693,N_7996,N_6803);
nor U8694 (N_8694,N_7617,N_6752);
xnor U8695 (N_8695,N_6157,N_7691);
nor U8696 (N_8696,N_7836,N_6749);
nand U8697 (N_8697,N_6382,N_6873);
nor U8698 (N_8698,N_7290,N_7599);
and U8699 (N_8699,N_7108,N_6080);
xnor U8700 (N_8700,N_6226,N_7288);
nor U8701 (N_8701,N_7456,N_7619);
nand U8702 (N_8702,N_6236,N_7425);
or U8703 (N_8703,N_6307,N_6448);
xor U8704 (N_8704,N_7113,N_6672);
nand U8705 (N_8705,N_6466,N_6184);
xor U8706 (N_8706,N_7852,N_7383);
nor U8707 (N_8707,N_6118,N_6000);
and U8708 (N_8708,N_7724,N_6562);
nand U8709 (N_8709,N_7284,N_7373);
nand U8710 (N_8710,N_6736,N_6577);
nand U8711 (N_8711,N_6791,N_6906);
nor U8712 (N_8712,N_6829,N_7485);
nand U8713 (N_8713,N_7962,N_7853);
nand U8714 (N_8714,N_7888,N_7214);
and U8715 (N_8715,N_6598,N_6648);
xor U8716 (N_8716,N_6680,N_7313);
and U8717 (N_8717,N_7404,N_6033);
xnor U8718 (N_8718,N_6077,N_6138);
nor U8719 (N_8719,N_7014,N_7163);
nor U8720 (N_8720,N_6999,N_6073);
xor U8721 (N_8721,N_6354,N_7706);
nor U8722 (N_8722,N_6768,N_6084);
xor U8723 (N_8723,N_6822,N_7336);
nor U8724 (N_8724,N_7597,N_7002);
or U8725 (N_8725,N_6743,N_6859);
or U8726 (N_8726,N_7539,N_7998);
or U8727 (N_8727,N_7032,N_7951);
and U8728 (N_8728,N_6109,N_7369);
and U8729 (N_8729,N_7253,N_7949);
nor U8730 (N_8730,N_7983,N_7000);
or U8731 (N_8731,N_6721,N_6314);
nor U8732 (N_8732,N_6732,N_7438);
nor U8733 (N_8733,N_7088,N_7847);
and U8734 (N_8734,N_7579,N_7896);
nor U8735 (N_8735,N_7399,N_6086);
xnor U8736 (N_8736,N_6891,N_6132);
nand U8737 (N_8737,N_6842,N_7168);
and U8738 (N_8738,N_6636,N_7631);
xor U8739 (N_8739,N_6370,N_7720);
and U8740 (N_8740,N_7516,N_7561);
or U8741 (N_8741,N_6430,N_7160);
xnor U8742 (N_8742,N_7621,N_7912);
nor U8743 (N_8743,N_6006,N_7734);
and U8744 (N_8744,N_7590,N_6876);
nand U8745 (N_8745,N_6111,N_6561);
nand U8746 (N_8746,N_7458,N_6900);
nand U8747 (N_8747,N_7299,N_6954);
nor U8748 (N_8748,N_7238,N_7045);
and U8749 (N_8749,N_6812,N_7447);
nand U8750 (N_8750,N_7129,N_7180);
or U8751 (N_8751,N_7418,N_6604);
nand U8752 (N_8752,N_6659,N_6855);
and U8753 (N_8753,N_7123,N_6461);
nand U8754 (N_8754,N_7713,N_6567);
nor U8755 (N_8755,N_6378,N_6484);
nand U8756 (N_8756,N_6159,N_6064);
nand U8757 (N_8757,N_7082,N_7919);
and U8758 (N_8758,N_7781,N_6155);
nor U8759 (N_8759,N_6915,N_6085);
and U8760 (N_8760,N_7953,N_6793);
xnor U8761 (N_8761,N_6056,N_6129);
nor U8762 (N_8762,N_6311,N_7335);
and U8763 (N_8763,N_7475,N_7928);
xor U8764 (N_8764,N_6032,N_6500);
and U8765 (N_8765,N_7462,N_7117);
and U8766 (N_8766,N_7507,N_6655);
or U8767 (N_8767,N_7428,N_6620);
or U8768 (N_8768,N_6513,N_6691);
xor U8769 (N_8769,N_7285,N_6332);
or U8770 (N_8770,N_6523,N_6161);
nand U8771 (N_8771,N_7844,N_7843);
nand U8772 (N_8772,N_6443,N_6275);
nor U8773 (N_8773,N_6219,N_7440);
or U8774 (N_8774,N_7708,N_7380);
or U8775 (N_8775,N_7678,N_6856);
and U8776 (N_8776,N_6777,N_7668);
nand U8777 (N_8777,N_7379,N_6738);
xor U8778 (N_8778,N_7394,N_7512);
nand U8779 (N_8779,N_6128,N_7634);
or U8780 (N_8780,N_6321,N_7172);
or U8781 (N_8781,N_6269,N_6467);
nand U8782 (N_8782,N_6739,N_6125);
xor U8783 (N_8783,N_7728,N_6094);
and U8784 (N_8784,N_6099,N_6323);
or U8785 (N_8785,N_7916,N_7535);
nor U8786 (N_8786,N_6765,N_7890);
and U8787 (N_8787,N_7398,N_7417);
and U8788 (N_8788,N_7411,N_6817);
or U8789 (N_8789,N_7066,N_6449);
nor U8790 (N_8790,N_6262,N_7001);
xnor U8791 (N_8791,N_7788,N_7771);
or U8792 (N_8792,N_7709,N_6700);
or U8793 (N_8793,N_7624,N_7712);
xnor U8794 (N_8794,N_7124,N_6471);
nor U8795 (N_8795,N_7105,N_7472);
and U8796 (N_8796,N_6191,N_7377);
nand U8797 (N_8797,N_7754,N_7632);
or U8798 (N_8798,N_7541,N_7365);
xnor U8799 (N_8799,N_6692,N_7718);
xor U8800 (N_8800,N_6451,N_6889);
and U8801 (N_8801,N_6810,N_6795);
xor U8802 (N_8802,N_7227,N_6957);
and U8803 (N_8803,N_7481,N_6364);
and U8804 (N_8804,N_7556,N_6676);
or U8805 (N_8805,N_7041,N_7907);
nand U8806 (N_8806,N_7696,N_7613);
nand U8807 (N_8807,N_7255,N_7479);
nand U8808 (N_8808,N_7698,N_6340);
xnor U8809 (N_8809,N_7087,N_7112);
or U8810 (N_8810,N_7490,N_6187);
and U8811 (N_8811,N_6877,N_7476);
and U8812 (N_8812,N_7370,N_7046);
and U8813 (N_8813,N_6566,N_7574);
nor U8814 (N_8814,N_6800,N_6022);
or U8815 (N_8815,N_7006,N_6186);
or U8816 (N_8816,N_6693,N_6458);
xnor U8817 (N_8817,N_6875,N_6767);
nand U8818 (N_8818,N_7726,N_6788);
nand U8819 (N_8819,N_6670,N_6151);
or U8820 (N_8820,N_6934,N_7311);
xnor U8821 (N_8821,N_7648,N_6465);
and U8822 (N_8822,N_7876,N_6446);
nor U8823 (N_8823,N_7245,N_6585);
nor U8824 (N_8824,N_7317,N_6730);
and U8825 (N_8825,N_6176,N_7495);
and U8826 (N_8826,N_6571,N_7396);
nand U8827 (N_8827,N_6826,N_6346);
or U8828 (N_8828,N_6413,N_6774);
and U8829 (N_8829,N_7538,N_6260);
or U8830 (N_8830,N_6339,N_6685);
nand U8831 (N_8831,N_6529,N_6617);
and U8832 (N_8832,N_6970,N_7955);
or U8833 (N_8833,N_7056,N_6689);
nand U8834 (N_8834,N_7320,N_7212);
nand U8835 (N_8835,N_6933,N_6060);
nand U8836 (N_8836,N_7178,N_6104);
xnor U8837 (N_8837,N_6944,N_6324);
xnor U8838 (N_8838,N_6816,N_6185);
and U8839 (N_8839,N_6574,N_6628);
and U8840 (N_8840,N_6398,N_6409);
xnor U8841 (N_8841,N_6432,N_6342);
and U8842 (N_8842,N_6935,N_7987);
and U8843 (N_8843,N_6839,N_7636);
or U8844 (N_8844,N_6496,N_6579);
nor U8845 (N_8845,N_7639,N_7861);
or U8846 (N_8846,N_7198,N_6550);
xor U8847 (N_8847,N_7746,N_6327);
nor U8848 (N_8848,N_6541,N_7111);
nand U8849 (N_8849,N_6711,N_6352);
and U8850 (N_8850,N_7466,N_7202);
and U8851 (N_8851,N_6141,N_7295);
nand U8852 (N_8852,N_7697,N_7237);
and U8853 (N_8853,N_7413,N_7093);
nand U8854 (N_8854,N_6982,N_7053);
nor U8855 (N_8855,N_6011,N_7300);
and U8856 (N_8856,N_6823,N_7669);
nor U8857 (N_8857,N_7747,N_7488);
or U8858 (N_8858,N_7672,N_7748);
xnor U8859 (N_8859,N_6116,N_6815);
or U8860 (N_8860,N_6053,N_6051);
nand U8861 (N_8861,N_7359,N_7807);
nor U8862 (N_8862,N_6422,N_6024);
xnor U8863 (N_8863,N_7799,N_6169);
xor U8864 (N_8864,N_6638,N_7453);
xor U8865 (N_8865,N_7024,N_7881);
and U8866 (N_8866,N_6147,N_6521);
and U8867 (N_8867,N_7638,N_7096);
nor U8868 (N_8868,N_6773,N_6832);
and U8869 (N_8869,N_7641,N_7381);
nand U8870 (N_8870,N_6547,N_7625);
nor U8871 (N_8871,N_6384,N_6533);
nor U8872 (N_8872,N_6203,N_6424);
and U8873 (N_8873,N_6401,N_7572);
nor U8874 (N_8874,N_6345,N_6375);
xnor U8875 (N_8875,N_6355,N_6489);
xnor U8876 (N_8876,N_6357,N_7196);
and U8877 (N_8877,N_6028,N_7711);
and U8878 (N_8878,N_6494,N_7689);
nor U8879 (N_8879,N_7961,N_6199);
nand U8880 (N_8880,N_7349,N_7925);
xnor U8881 (N_8881,N_6163,N_7210);
nor U8882 (N_8882,N_7280,N_6558);
nand U8883 (N_8883,N_6827,N_6792);
xnor U8884 (N_8884,N_6656,N_7494);
and U8885 (N_8885,N_7588,N_6901);
nor U8886 (N_8886,N_6525,N_6171);
or U8887 (N_8887,N_6093,N_7126);
or U8888 (N_8888,N_6516,N_6728);
nor U8889 (N_8889,N_6351,N_6292);
nor U8890 (N_8890,N_7931,N_7892);
xor U8891 (N_8891,N_6041,N_7742);
or U8892 (N_8892,N_7422,N_7940);
and U8893 (N_8893,N_7322,N_7901);
nor U8894 (N_8894,N_6797,N_6897);
xor U8895 (N_8895,N_7296,N_6630);
and U8896 (N_8896,N_7835,N_7529);
and U8897 (N_8897,N_7254,N_6805);
and U8898 (N_8898,N_7860,N_7569);
nand U8899 (N_8899,N_6395,N_6737);
or U8900 (N_8900,N_6975,N_7553);
or U8901 (N_8901,N_7339,N_6903);
nand U8902 (N_8902,N_6882,N_6273);
nand U8903 (N_8903,N_7820,N_7228);
and U8904 (N_8904,N_6701,N_7248);
nand U8905 (N_8905,N_6392,N_6682);
and U8906 (N_8906,N_6741,N_6962);
nor U8907 (N_8907,N_6608,N_7651);
and U8908 (N_8908,N_7075,N_6098);
xor U8909 (N_8909,N_6365,N_7885);
nand U8910 (N_8910,N_7416,N_6008);
or U8911 (N_8911,N_6531,N_6830);
or U8912 (N_8912,N_7532,N_7584);
and U8913 (N_8913,N_6373,N_7069);
or U8914 (N_8914,N_7460,N_6745);
nand U8915 (N_8915,N_6660,N_7140);
and U8916 (N_8916,N_7036,N_7751);
xnor U8917 (N_8917,N_7437,N_6240);
or U8918 (N_8918,N_7656,N_6928);
nor U8919 (N_8919,N_6435,N_6250);
xnor U8920 (N_8920,N_7426,N_6344);
nand U8921 (N_8921,N_7161,N_7303);
or U8922 (N_8922,N_6664,N_6247);
xor U8923 (N_8923,N_6309,N_6120);
xnor U8924 (N_8924,N_6825,N_7424);
and U8925 (N_8925,N_7594,N_7221);
nand U8926 (N_8926,N_7942,N_7694);
nand U8927 (N_8927,N_6329,N_6423);
or U8928 (N_8928,N_6619,N_6910);
or U8929 (N_8929,N_7959,N_6776);
xor U8930 (N_8930,N_6861,N_6925);
and U8931 (N_8931,N_7328,N_7375);
xor U8932 (N_8932,N_6662,N_7362);
nand U8933 (N_8933,N_7423,N_6572);
nand U8934 (N_8934,N_7981,N_6303);
xnor U8935 (N_8935,N_7421,N_6018);
nor U8936 (N_8936,N_6923,N_6071);
nor U8937 (N_8937,N_6058,N_6499);
nor U8938 (N_8938,N_6072,N_7923);
nor U8939 (N_8939,N_6828,N_7016);
or U8940 (N_8940,N_7318,N_7973);
nor U8941 (N_8941,N_6429,N_6969);
xor U8942 (N_8942,N_7991,N_6995);
or U8943 (N_8943,N_7017,N_7818);
xnor U8944 (N_8944,N_7832,N_7865);
xor U8945 (N_8945,N_6130,N_6528);
xor U8946 (N_8946,N_7059,N_7343);
and U8947 (N_8947,N_6548,N_6993);
xor U8948 (N_8948,N_6725,N_6393);
nor U8949 (N_8949,N_7684,N_6526);
nor U8950 (N_8950,N_7225,N_6137);
xnor U8951 (N_8951,N_7855,N_6781);
xnor U8952 (N_8952,N_6331,N_7596);
or U8953 (N_8953,N_7278,N_6246);
xor U8954 (N_8954,N_6213,N_7506);
nand U8955 (N_8955,N_6652,N_7342);
nor U8956 (N_8956,N_7809,N_6972);
and U8957 (N_8957,N_7218,N_6587);
nor U8958 (N_8958,N_6007,N_6183);
or U8959 (N_8959,N_7323,N_6206);
and U8960 (N_8960,N_6858,N_7994);
or U8961 (N_8961,N_6895,N_7946);
or U8962 (N_8962,N_6195,N_6588);
nand U8963 (N_8963,N_6070,N_6991);
xor U8964 (N_8964,N_7827,N_6914);
xor U8965 (N_8965,N_6441,N_6114);
and U8966 (N_8966,N_7815,N_7958);
or U8967 (N_8967,N_7345,N_7536);
nor U8968 (N_8968,N_6631,N_7354);
xnor U8969 (N_8969,N_7814,N_7406);
xnor U8970 (N_8970,N_7871,N_6844);
nor U8971 (N_8971,N_7797,N_6642);
and U8972 (N_8972,N_6573,N_7515);
nand U8973 (N_8973,N_6578,N_7022);
and U8974 (N_8974,N_7086,N_6735);
and U8975 (N_8975,N_6647,N_7487);
or U8976 (N_8976,N_7936,N_7193);
and U8977 (N_8977,N_7833,N_7119);
nor U8978 (N_8978,N_6150,N_6404);
xnor U8979 (N_8979,N_6406,N_6217);
xnor U8980 (N_8980,N_7878,N_6722);
nor U8981 (N_8981,N_7110,N_6549);
xor U8982 (N_8982,N_6819,N_7496);
xor U8983 (N_8983,N_7388,N_7243);
nand U8984 (N_8984,N_7922,N_6904);
xor U8985 (N_8985,N_6322,N_7848);
or U8986 (N_8986,N_6223,N_7719);
nand U8987 (N_8987,N_6408,N_6377);
nor U8988 (N_8988,N_6540,N_6237);
nand U8989 (N_8989,N_7808,N_6146);
nand U8990 (N_8990,N_7357,N_6902);
and U8991 (N_8991,N_6802,N_7235);
xor U8992 (N_8992,N_7531,N_6259);
nor U8993 (N_8993,N_6190,N_6679);
nand U8994 (N_8994,N_6134,N_6565);
xor U8995 (N_8995,N_6892,N_7612);
nand U8996 (N_8996,N_6305,N_6960);
or U8997 (N_8997,N_6308,N_7997);
and U8998 (N_8998,N_6235,N_6971);
or U8999 (N_8999,N_6172,N_6498);
nor U9000 (N_9000,N_7297,N_7580);
and U9001 (N_9001,N_6729,N_7950);
nand U9002 (N_9002,N_6576,N_7534);
or U9003 (N_9003,N_6209,N_6902);
or U9004 (N_9004,N_6439,N_6641);
nor U9005 (N_9005,N_7736,N_7411);
nor U9006 (N_9006,N_7908,N_6489);
xor U9007 (N_9007,N_7392,N_6105);
xor U9008 (N_9008,N_7166,N_7160);
or U9009 (N_9009,N_7309,N_7753);
xnor U9010 (N_9010,N_7387,N_7886);
xor U9011 (N_9011,N_6657,N_6683);
and U9012 (N_9012,N_6538,N_7975);
or U9013 (N_9013,N_7609,N_7591);
nor U9014 (N_9014,N_7140,N_6127);
or U9015 (N_9015,N_7394,N_6620);
nand U9016 (N_9016,N_7247,N_7629);
xor U9017 (N_9017,N_7588,N_7906);
and U9018 (N_9018,N_6132,N_7731);
or U9019 (N_9019,N_6092,N_6100);
nand U9020 (N_9020,N_7011,N_7567);
xnor U9021 (N_9021,N_6699,N_6601);
and U9022 (N_9022,N_7338,N_6512);
xor U9023 (N_9023,N_6849,N_7182);
or U9024 (N_9024,N_7446,N_7995);
and U9025 (N_9025,N_7219,N_6499);
nor U9026 (N_9026,N_7881,N_7338);
and U9027 (N_9027,N_7641,N_6308);
or U9028 (N_9028,N_6028,N_6960);
or U9029 (N_9029,N_7764,N_7129);
and U9030 (N_9030,N_6518,N_7122);
and U9031 (N_9031,N_6094,N_7223);
nor U9032 (N_9032,N_7680,N_6244);
and U9033 (N_9033,N_7114,N_7858);
and U9034 (N_9034,N_6850,N_7080);
nand U9035 (N_9035,N_7298,N_7449);
xnor U9036 (N_9036,N_6002,N_6562);
or U9037 (N_9037,N_7923,N_6580);
nor U9038 (N_9038,N_6529,N_6777);
nor U9039 (N_9039,N_6841,N_6067);
xnor U9040 (N_9040,N_6557,N_7192);
or U9041 (N_9041,N_7144,N_7881);
xnor U9042 (N_9042,N_6326,N_6393);
xor U9043 (N_9043,N_7390,N_7586);
xor U9044 (N_9044,N_7473,N_6613);
or U9045 (N_9045,N_7483,N_6731);
or U9046 (N_9046,N_7984,N_6231);
nor U9047 (N_9047,N_7030,N_6371);
nand U9048 (N_9048,N_6032,N_7725);
nand U9049 (N_9049,N_6971,N_7540);
xnor U9050 (N_9050,N_6271,N_6959);
or U9051 (N_9051,N_7195,N_6761);
nand U9052 (N_9052,N_7023,N_6711);
xnor U9053 (N_9053,N_6986,N_7948);
xnor U9054 (N_9054,N_6442,N_6589);
or U9055 (N_9055,N_6657,N_6236);
or U9056 (N_9056,N_7222,N_7227);
xnor U9057 (N_9057,N_6246,N_7169);
and U9058 (N_9058,N_7994,N_7710);
nor U9059 (N_9059,N_6777,N_7418);
or U9060 (N_9060,N_6637,N_7069);
or U9061 (N_9061,N_6595,N_6318);
or U9062 (N_9062,N_7728,N_7357);
nor U9063 (N_9063,N_7131,N_7840);
and U9064 (N_9064,N_6424,N_6505);
nand U9065 (N_9065,N_6229,N_7224);
nand U9066 (N_9066,N_6809,N_7957);
or U9067 (N_9067,N_6292,N_6435);
xor U9068 (N_9068,N_6022,N_6942);
and U9069 (N_9069,N_6069,N_7736);
nand U9070 (N_9070,N_6638,N_7734);
or U9071 (N_9071,N_6610,N_7505);
xor U9072 (N_9072,N_7337,N_6317);
nand U9073 (N_9073,N_6440,N_7840);
xnor U9074 (N_9074,N_6028,N_6651);
xor U9075 (N_9075,N_6335,N_7864);
nor U9076 (N_9076,N_7838,N_6504);
and U9077 (N_9077,N_7445,N_7398);
and U9078 (N_9078,N_7876,N_6486);
nor U9079 (N_9079,N_7590,N_7578);
and U9080 (N_9080,N_6118,N_6473);
or U9081 (N_9081,N_6854,N_6362);
nor U9082 (N_9082,N_7980,N_6026);
nand U9083 (N_9083,N_7431,N_7902);
nand U9084 (N_9084,N_7441,N_6107);
nand U9085 (N_9085,N_7281,N_7012);
or U9086 (N_9086,N_7376,N_7490);
nor U9087 (N_9087,N_7605,N_6651);
xor U9088 (N_9088,N_7898,N_7734);
or U9089 (N_9089,N_6624,N_7237);
nand U9090 (N_9090,N_6683,N_6589);
and U9091 (N_9091,N_6868,N_7346);
nand U9092 (N_9092,N_7949,N_6870);
nand U9093 (N_9093,N_6419,N_6495);
xor U9094 (N_9094,N_7043,N_6791);
or U9095 (N_9095,N_7410,N_7118);
nand U9096 (N_9096,N_7727,N_6584);
nand U9097 (N_9097,N_6496,N_7668);
or U9098 (N_9098,N_6802,N_6204);
or U9099 (N_9099,N_6169,N_7822);
xor U9100 (N_9100,N_6688,N_6925);
nor U9101 (N_9101,N_6014,N_6337);
nor U9102 (N_9102,N_6858,N_7067);
or U9103 (N_9103,N_6057,N_6456);
or U9104 (N_9104,N_6798,N_6193);
or U9105 (N_9105,N_7695,N_7910);
or U9106 (N_9106,N_6951,N_7944);
nor U9107 (N_9107,N_6668,N_7691);
nand U9108 (N_9108,N_7436,N_6400);
or U9109 (N_9109,N_7420,N_7939);
and U9110 (N_9110,N_6195,N_6682);
and U9111 (N_9111,N_6961,N_6228);
and U9112 (N_9112,N_7698,N_6702);
nor U9113 (N_9113,N_6698,N_7007);
and U9114 (N_9114,N_6405,N_7804);
or U9115 (N_9115,N_6631,N_7604);
nor U9116 (N_9116,N_7583,N_6549);
or U9117 (N_9117,N_7138,N_7699);
xor U9118 (N_9118,N_6668,N_7475);
nand U9119 (N_9119,N_6073,N_6838);
nand U9120 (N_9120,N_7086,N_6484);
or U9121 (N_9121,N_6152,N_7839);
and U9122 (N_9122,N_7002,N_6285);
xor U9123 (N_9123,N_6438,N_7496);
nor U9124 (N_9124,N_6818,N_6056);
nand U9125 (N_9125,N_6776,N_7774);
nor U9126 (N_9126,N_6828,N_7254);
nand U9127 (N_9127,N_6267,N_7808);
or U9128 (N_9128,N_6913,N_7032);
nor U9129 (N_9129,N_7549,N_6179);
xor U9130 (N_9130,N_6006,N_6532);
xnor U9131 (N_9131,N_7991,N_7089);
nand U9132 (N_9132,N_6972,N_6559);
or U9133 (N_9133,N_7870,N_7250);
nor U9134 (N_9134,N_6382,N_6257);
xor U9135 (N_9135,N_7967,N_7364);
and U9136 (N_9136,N_7341,N_7268);
xor U9137 (N_9137,N_6554,N_7627);
and U9138 (N_9138,N_7874,N_6612);
nor U9139 (N_9139,N_6053,N_6533);
nand U9140 (N_9140,N_6984,N_7129);
and U9141 (N_9141,N_6509,N_7032);
xnor U9142 (N_9142,N_7392,N_7137);
xnor U9143 (N_9143,N_6418,N_7623);
xor U9144 (N_9144,N_7316,N_6467);
nor U9145 (N_9145,N_7984,N_7004);
nor U9146 (N_9146,N_6450,N_6597);
or U9147 (N_9147,N_7735,N_6559);
and U9148 (N_9148,N_6736,N_7030);
nor U9149 (N_9149,N_6358,N_6434);
xnor U9150 (N_9150,N_6725,N_7739);
xor U9151 (N_9151,N_7166,N_6947);
nand U9152 (N_9152,N_7826,N_6300);
xnor U9153 (N_9153,N_6352,N_6655);
xnor U9154 (N_9154,N_6022,N_7497);
xor U9155 (N_9155,N_6475,N_6960);
and U9156 (N_9156,N_7781,N_7668);
xor U9157 (N_9157,N_6952,N_7672);
xor U9158 (N_9158,N_7105,N_6861);
nor U9159 (N_9159,N_7370,N_7640);
nor U9160 (N_9160,N_6688,N_6231);
or U9161 (N_9161,N_7964,N_6027);
nand U9162 (N_9162,N_6083,N_7891);
and U9163 (N_9163,N_6042,N_6326);
or U9164 (N_9164,N_6657,N_6595);
nand U9165 (N_9165,N_6713,N_6393);
nand U9166 (N_9166,N_6728,N_7364);
or U9167 (N_9167,N_6130,N_6924);
xor U9168 (N_9168,N_7863,N_7397);
or U9169 (N_9169,N_6762,N_6312);
nor U9170 (N_9170,N_6683,N_6613);
or U9171 (N_9171,N_6376,N_7810);
xnor U9172 (N_9172,N_6074,N_6695);
xnor U9173 (N_9173,N_7590,N_6031);
nor U9174 (N_9174,N_6982,N_6523);
and U9175 (N_9175,N_7748,N_7914);
nor U9176 (N_9176,N_6603,N_6403);
or U9177 (N_9177,N_6206,N_6432);
nand U9178 (N_9178,N_7737,N_7215);
and U9179 (N_9179,N_6193,N_7722);
and U9180 (N_9180,N_6841,N_6818);
nand U9181 (N_9181,N_6638,N_7465);
xnor U9182 (N_9182,N_7640,N_7494);
xor U9183 (N_9183,N_7451,N_6442);
and U9184 (N_9184,N_7409,N_6162);
nor U9185 (N_9185,N_7661,N_6917);
or U9186 (N_9186,N_6599,N_7932);
and U9187 (N_9187,N_6979,N_7266);
xor U9188 (N_9188,N_6647,N_6181);
or U9189 (N_9189,N_7509,N_7429);
nor U9190 (N_9190,N_7302,N_6613);
nor U9191 (N_9191,N_7857,N_7903);
or U9192 (N_9192,N_6662,N_6435);
or U9193 (N_9193,N_7729,N_6158);
or U9194 (N_9194,N_6523,N_7081);
nand U9195 (N_9195,N_6562,N_7497);
nand U9196 (N_9196,N_6476,N_6259);
nor U9197 (N_9197,N_6091,N_6195);
xor U9198 (N_9198,N_6007,N_7008);
or U9199 (N_9199,N_7707,N_7753);
nor U9200 (N_9200,N_7339,N_6055);
or U9201 (N_9201,N_6204,N_6681);
nor U9202 (N_9202,N_6234,N_6374);
nand U9203 (N_9203,N_7702,N_6301);
xnor U9204 (N_9204,N_7995,N_6370);
or U9205 (N_9205,N_6504,N_7537);
and U9206 (N_9206,N_7987,N_6049);
and U9207 (N_9207,N_6574,N_6375);
nor U9208 (N_9208,N_7942,N_6553);
nand U9209 (N_9209,N_7776,N_7652);
or U9210 (N_9210,N_7784,N_6388);
or U9211 (N_9211,N_7721,N_6057);
nor U9212 (N_9212,N_6580,N_7460);
or U9213 (N_9213,N_6857,N_7656);
nand U9214 (N_9214,N_6852,N_6983);
or U9215 (N_9215,N_6706,N_7455);
and U9216 (N_9216,N_6095,N_6167);
or U9217 (N_9217,N_6705,N_6133);
and U9218 (N_9218,N_6020,N_7631);
nand U9219 (N_9219,N_6402,N_6114);
nand U9220 (N_9220,N_7507,N_7282);
and U9221 (N_9221,N_6213,N_6227);
and U9222 (N_9222,N_6282,N_6707);
xor U9223 (N_9223,N_6191,N_6835);
nor U9224 (N_9224,N_7351,N_7425);
xor U9225 (N_9225,N_7345,N_6186);
or U9226 (N_9226,N_7942,N_6932);
or U9227 (N_9227,N_7451,N_6936);
nor U9228 (N_9228,N_6413,N_6602);
nor U9229 (N_9229,N_6295,N_6061);
and U9230 (N_9230,N_7959,N_6586);
nor U9231 (N_9231,N_7664,N_7009);
nand U9232 (N_9232,N_7414,N_6679);
nand U9233 (N_9233,N_6294,N_7512);
or U9234 (N_9234,N_6883,N_6920);
and U9235 (N_9235,N_6368,N_6681);
and U9236 (N_9236,N_7457,N_7815);
and U9237 (N_9237,N_6875,N_7602);
nand U9238 (N_9238,N_7017,N_7492);
nand U9239 (N_9239,N_6017,N_7423);
nor U9240 (N_9240,N_6855,N_6839);
nor U9241 (N_9241,N_6001,N_6115);
nand U9242 (N_9242,N_7926,N_6615);
nand U9243 (N_9243,N_6062,N_6823);
and U9244 (N_9244,N_6269,N_7916);
nand U9245 (N_9245,N_7614,N_6799);
nor U9246 (N_9246,N_6734,N_7864);
nand U9247 (N_9247,N_7069,N_6523);
or U9248 (N_9248,N_6138,N_6549);
nor U9249 (N_9249,N_7009,N_7461);
or U9250 (N_9250,N_6047,N_6950);
nor U9251 (N_9251,N_7332,N_6234);
nor U9252 (N_9252,N_7871,N_6797);
xnor U9253 (N_9253,N_6471,N_6915);
xnor U9254 (N_9254,N_7369,N_6758);
and U9255 (N_9255,N_7370,N_7921);
nor U9256 (N_9256,N_6310,N_7231);
nand U9257 (N_9257,N_6456,N_7081);
or U9258 (N_9258,N_6508,N_6266);
or U9259 (N_9259,N_7461,N_6323);
xor U9260 (N_9260,N_6717,N_7293);
nand U9261 (N_9261,N_6050,N_6446);
nor U9262 (N_9262,N_7376,N_7600);
xor U9263 (N_9263,N_6975,N_6596);
nand U9264 (N_9264,N_7758,N_7288);
nor U9265 (N_9265,N_7213,N_6076);
nor U9266 (N_9266,N_7706,N_7154);
nor U9267 (N_9267,N_7973,N_7321);
xor U9268 (N_9268,N_7698,N_7704);
nor U9269 (N_9269,N_6286,N_6008);
or U9270 (N_9270,N_7874,N_6111);
nand U9271 (N_9271,N_6455,N_6864);
nor U9272 (N_9272,N_6800,N_6955);
nor U9273 (N_9273,N_7786,N_6931);
nand U9274 (N_9274,N_7982,N_7433);
and U9275 (N_9275,N_7090,N_6830);
xor U9276 (N_9276,N_7615,N_7143);
and U9277 (N_9277,N_7251,N_6982);
or U9278 (N_9278,N_7940,N_7192);
or U9279 (N_9279,N_6027,N_7064);
or U9280 (N_9280,N_6336,N_6590);
nand U9281 (N_9281,N_7647,N_6044);
and U9282 (N_9282,N_7574,N_6339);
xnor U9283 (N_9283,N_7452,N_7408);
xor U9284 (N_9284,N_6995,N_6113);
nand U9285 (N_9285,N_7903,N_6110);
nor U9286 (N_9286,N_6657,N_6134);
nor U9287 (N_9287,N_6119,N_7388);
nor U9288 (N_9288,N_6553,N_6624);
or U9289 (N_9289,N_7435,N_6633);
nor U9290 (N_9290,N_6907,N_6303);
and U9291 (N_9291,N_7981,N_6702);
xor U9292 (N_9292,N_7901,N_6523);
and U9293 (N_9293,N_6854,N_6327);
and U9294 (N_9294,N_6224,N_6751);
nor U9295 (N_9295,N_6868,N_7803);
nand U9296 (N_9296,N_6921,N_7544);
nand U9297 (N_9297,N_6919,N_7667);
nor U9298 (N_9298,N_6827,N_6154);
nand U9299 (N_9299,N_6382,N_6877);
nor U9300 (N_9300,N_6194,N_7484);
nor U9301 (N_9301,N_6916,N_7981);
xor U9302 (N_9302,N_7035,N_7631);
nor U9303 (N_9303,N_7260,N_7652);
or U9304 (N_9304,N_6805,N_7700);
or U9305 (N_9305,N_7909,N_7293);
xor U9306 (N_9306,N_6858,N_6662);
xor U9307 (N_9307,N_6790,N_7370);
or U9308 (N_9308,N_6223,N_7818);
or U9309 (N_9309,N_7992,N_7379);
nor U9310 (N_9310,N_6344,N_7927);
or U9311 (N_9311,N_7033,N_7981);
or U9312 (N_9312,N_6580,N_7391);
xnor U9313 (N_9313,N_6295,N_7179);
nor U9314 (N_9314,N_7077,N_7731);
xnor U9315 (N_9315,N_7610,N_7909);
nand U9316 (N_9316,N_6875,N_7964);
and U9317 (N_9317,N_6134,N_6647);
nand U9318 (N_9318,N_6336,N_6486);
or U9319 (N_9319,N_7864,N_6550);
and U9320 (N_9320,N_6425,N_6129);
and U9321 (N_9321,N_6119,N_7469);
xnor U9322 (N_9322,N_6828,N_7709);
nand U9323 (N_9323,N_7936,N_7654);
or U9324 (N_9324,N_6282,N_6891);
nand U9325 (N_9325,N_6219,N_6604);
nor U9326 (N_9326,N_6644,N_6524);
nand U9327 (N_9327,N_7801,N_6066);
nor U9328 (N_9328,N_7950,N_7230);
or U9329 (N_9329,N_7341,N_6723);
nor U9330 (N_9330,N_6525,N_7806);
nor U9331 (N_9331,N_6779,N_6628);
or U9332 (N_9332,N_6893,N_6465);
nand U9333 (N_9333,N_7318,N_6612);
nand U9334 (N_9334,N_6102,N_7077);
and U9335 (N_9335,N_6476,N_6014);
or U9336 (N_9336,N_6973,N_6241);
xor U9337 (N_9337,N_6312,N_6166);
and U9338 (N_9338,N_7133,N_6994);
or U9339 (N_9339,N_6567,N_7263);
nand U9340 (N_9340,N_6456,N_6737);
nor U9341 (N_9341,N_6824,N_7305);
nor U9342 (N_9342,N_7001,N_7913);
or U9343 (N_9343,N_7516,N_7898);
and U9344 (N_9344,N_7662,N_7067);
or U9345 (N_9345,N_7941,N_6191);
nor U9346 (N_9346,N_6198,N_7026);
nor U9347 (N_9347,N_7398,N_7270);
and U9348 (N_9348,N_6902,N_6601);
nor U9349 (N_9349,N_7064,N_7245);
or U9350 (N_9350,N_6668,N_7596);
or U9351 (N_9351,N_6122,N_7472);
or U9352 (N_9352,N_7232,N_6944);
nor U9353 (N_9353,N_7088,N_6913);
or U9354 (N_9354,N_6544,N_6476);
or U9355 (N_9355,N_7198,N_7041);
and U9356 (N_9356,N_6000,N_7904);
nand U9357 (N_9357,N_7204,N_6827);
nand U9358 (N_9358,N_7373,N_7902);
xor U9359 (N_9359,N_7604,N_7289);
nand U9360 (N_9360,N_7007,N_6727);
and U9361 (N_9361,N_7681,N_7904);
nand U9362 (N_9362,N_7221,N_6797);
and U9363 (N_9363,N_7879,N_6897);
xnor U9364 (N_9364,N_6622,N_6883);
nor U9365 (N_9365,N_7572,N_6723);
and U9366 (N_9366,N_6303,N_6007);
xor U9367 (N_9367,N_7283,N_6106);
or U9368 (N_9368,N_7847,N_7654);
nand U9369 (N_9369,N_7282,N_7878);
nand U9370 (N_9370,N_6807,N_7631);
xor U9371 (N_9371,N_7788,N_6857);
nand U9372 (N_9372,N_6262,N_6764);
or U9373 (N_9373,N_6214,N_6428);
nor U9374 (N_9374,N_7444,N_7180);
nor U9375 (N_9375,N_6331,N_6569);
and U9376 (N_9376,N_7770,N_6158);
or U9377 (N_9377,N_6263,N_6518);
xnor U9378 (N_9378,N_6489,N_7242);
xor U9379 (N_9379,N_6707,N_7847);
xnor U9380 (N_9380,N_6120,N_7272);
and U9381 (N_9381,N_7013,N_6816);
nand U9382 (N_9382,N_7753,N_7775);
or U9383 (N_9383,N_6674,N_7361);
and U9384 (N_9384,N_6207,N_6719);
nor U9385 (N_9385,N_6698,N_6658);
and U9386 (N_9386,N_7950,N_6233);
and U9387 (N_9387,N_7896,N_7446);
nor U9388 (N_9388,N_7440,N_6698);
or U9389 (N_9389,N_6210,N_6750);
nand U9390 (N_9390,N_6059,N_7134);
nor U9391 (N_9391,N_6837,N_7195);
or U9392 (N_9392,N_7134,N_7679);
and U9393 (N_9393,N_6118,N_7883);
or U9394 (N_9394,N_6653,N_7758);
or U9395 (N_9395,N_6811,N_7176);
or U9396 (N_9396,N_7093,N_6914);
or U9397 (N_9397,N_7669,N_6343);
xnor U9398 (N_9398,N_7396,N_7938);
xor U9399 (N_9399,N_6508,N_7159);
or U9400 (N_9400,N_7873,N_7159);
or U9401 (N_9401,N_7999,N_6719);
xnor U9402 (N_9402,N_7910,N_7195);
or U9403 (N_9403,N_6967,N_7045);
nand U9404 (N_9404,N_6020,N_6851);
xor U9405 (N_9405,N_7467,N_7724);
nor U9406 (N_9406,N_6379,N_7001);
xnor U9407 (N_9407,N_7542,N_7823);
nand U9408 (N_9408,N_7565,N_6627);
or U9409 (N_9409,N_6989,N_6846);
nor U9410 (N_9410,N_7329,N_7351);
or U9411 (N_9411,N_7615,N_7639);
nor U9412 (N_9412,N_6293,N_6728);
or U9413 (N_9413,N_7546,N_7926);
or U9414 (N_9414,N_7705,N_7559);
or U9415 (N_9415,N_6893,N_6067);
nand U9416 (N_9416,N_6577,N_7105);
or U9417 (N_9417,N_6570,N_6972);
or U9418 (N_9418,N_7797,N_7054);
and U9419 (N_9419,N_6681,N_6400);
xor U9420 (N_9420,N_6527,N_6005);
nand U9421 (N_9421,N_7496,N_6102);
and U9422 (N_9422,N_6582,N_6281);
and U9423 (N_9423,N_7508,N_7783);
nor U9424 (N_9424,N_6110,N_7109);
and U9425 (N_9425,N_7447,N_7282);
nand U9426 (N_9426,N_7316,N_7241);
and U9427 (N_9427,N_6070,N_6949);
xnor U9428 (N_9428,N_7395,N_6896);
xor U9429 (N_9429,N_7108,N_7580);
nor U9430 (N_9430,N_7195,N_7639);
xor U9431 (N_9431,N_7579,N_6052);
or U9432 (N_9432,N_6718,N_7711);
nor U9433 (N_9433,N_6998,N_7921);
nand U9434 (N_9434,N_6160,N_7699);
nand U9435 (N_9435,N_6212,N_7620);
and U9436 (N_9436,N_7288,N_6770);
xnor U9437 (N_9437,N_7236,N_7597);
and U9438 (N_9438,N_6286,N_7037);
and U9439 (N_9439,N_6316,N_7682);
nand U9440 (N_9440,N_6918,N_6790);
nand U9441 (N_9441,N_6116,N_7364);
nor U9442 (N_9442,N_6173,N_6862);
xor U9443 (N_9443,N_6233,N_7391);
or U9444 (N_9444,N_7124,N_7431);
and U9445 (N_9445,N_7134,N_6457);
xnor U9446 (N_9446,N_7631,N_7180);
or U9447 (N_9447,N_6037,N_6749);
nor U9448 (N_9448,N_7627,N_6868);
nor U9449 (N_9449,N_6117,N_6169);
and U9450 (N_9450,N_6132,N_6402);
xnor U9451 (N_9451,N_6977,N_7546);
or U9452 (N_9452,N_6977,N_6004);
or U9453 (N_9453,N_7231,N_7009);
or U9454 (N_9454,N_6500,N_7283);
xnor U9455 (N_9455,N_6881,N_7220);
or U9456 (N_9456,N_7616,N_6326);
nor U9457 (N_9457,N_6642,N_6915);
nand U9458 (N_9458,N_6975,N_6010);
and U9459 (N_9459,N_6029,N_6527);
xor U9460 (N_9460,N_6236,N_6588);
xnor U9461 (N_9461,N_7128,N_7413);
and U9462 (N_9462,N_6980,N_6810);
xor U9463 (N_9463,N_7003,N_6845);
and U9464 (N_9464,N_6947,N_7541);
or U9465 (N_9465,N_6739,N_6006);
or U9466 (N_9466,N_6377,N_6850);
xnor U9467 (N_9467,N_7080,N_6361);
nand U9468 (N_9468,N_7312,N_6627);
or U9469 (N_9469,N_6484,N_6980);
and U9470 (N_9470,N_7316,N_7084);
or U9471 (N_9471,N_7245,N_6804);
nor U9472 (N_9472,N_7718,N_7032);
xor U9473 (N_9473,N_7138,N_6705);
and U9474 (N_9474,N_7842,N_7092);
and U9475 (N_9475,N_6245,N_7033);
or U9476 (N_9476,N_6798,N_6176);
xnor U9477 (N_9477,N_7264,N_6782);
and U9478 (N_9478,N_6321,N_7804);
nand U9479 (N_9479,N_6362,N_6451);
xor U9480 (N_9480,N_6757,N_7026);
and U9481 (N_9481,N_6899,N_6644);
or U9482 (N_9482,N_6043,N_7928);
nand U9483 (N_9483,N_7529,N_6549);
and U9484 (N_9484,N_6138,N_7482);
xor U9485 (N_9485,N_7663,N_6505);
nand U9486 (N_9486,N_7472,N_6882);
and U9487 (N_9487,N_6121,N_7602);
or U9488 (N_9488,N_7524,N_6299);
and U9489 (N_9489,N_7293,N_7083);
xnor U9490 (N_9490,N_7210,N_6647);
or U9491 (N_9491,N_6241,N_6144);
nand U9492 (N_9492,N_6640,N_7745);
nand U9493 (N_9493,N_6098,N_6504);
nand U9494 (N_9494,N_7228,N_6750);
and U9495 (N_9495,N_7865,N_6320);
nand U9496 (N_9496,N_6146,N_7493);
nor U9497 (N_9497,N_6544,N_6533);
nor U9498 (N_9498,N_7738,N_6135);
nor U9499 (N_9499,N_7066,N_7528);
or U9500 (N_9500,N_7557,N_6508);
xnor U9501 (N_9501,N_6243,N_7655);
nand U9502 (N_9502,N_7699,N_7397);
nor U9503 (N_9503,N_6011,N_6635);
nor U9504 (N_9504,N_6875,N_7835);
nand U9505 (N_9505,N_6176,N_7576);
nor U9506 (N_9506,N_7258,N_6191);
or U9507 (N_9507,N_6345,N_6148);
nand U9508 (N_9508,N_6402,N_6621);
nor U9509 (N_9509,N_6116,N_7587);
xnor U9510 (N_9510,N_6163,N_6178);
nand U9511 (N_9511,N_7508,N_7018);
or U9512 (N_9512,N_6244,N_7424);
or U9513 (N_9513,N_6272,N_6156);
xnor U9514 (N_9514,N_7918,N_7258);
xnor U9515 (N_9515,N_6175,N_6489);
nor U9516 (N_9516,N_7271,N_7901);
or U9517 (N_9517,N_6367,N_6771);
nand U9518 (N_9518,N_7317,N_7032);
nand U9519 (N_9519,N_7714,N_7883);
nand U9520 (N_9520,N_6905,N_7571);
and U9521 (N_9521,N_6975,N_6738);
xor U9522 (N_9522,N_7664,N_6273);
nand U9523 (N_9523,N_6883,N_7820);
and U9524 (N_9524,N_6203,N_7473);
nor U9525 (N_9525,N_6306,N_7420);
and U9526 (N_9526,N_6324,N_7033);
or U9527 (N_9527,N_6224,N_7827);
nor U9528 (N_9528,N_7865,N_6941);
and U9529 (N_9529,N_7500,N_6392);
and U9530 (N_9530,N_6875,N_7853);
nand U9531 (N_9531,N_6886,N_6522);
and U9532 (N_9532,N_6294,N_7651);
and U9533 (N_9533,N_6616,N_6906);
nand U9534 (N_9534,N_6728,N_6125);
and U9535 (N_9535,N_6007,N_6163);
or U9536 (N_9536,N_7370,N_7721);
and U9537 (N_9537,N_6134,N_7112);
nor U9538 (N_9538,N_7036,N_6130);
nand U9539 (N_9539,N_7447,N_7561);
or U9540 (N_9540,N_6262,N_6968);
nand U9541 (N_9541,N_7843,N_7772);
nand U9542 (N_9542,N_6826,N_6629);
or U9543 (N_9543,N_7661,N_7060);
and U9544 (N_9544,N_6619,N_7854);
nand U9545 (N_9545,N_6705,N_7198);
and U9546 (N_9546,N_6302,N_7099);
or U9547 (N_9547,N_6541,N_6368);
xor U9548 (N_9548,N_7360,N_6566);
nand U9549 (N_9549,N_6037,N_6508);
nor U9550 (N_9550,N_7596,N_7191);
nand U9551 (N_9551,N_6606,N_7685);
nand U9552 (N_9552,N_7363,N_6605);
xor U9553 (N_9553,N_7819,N_6802);
xor U9554 (N_9554,N_7086,N_7683);
nand U9555 (N_9555,N_7693,N_6978);
and U9556 (N_9556,N_6386,N_7275);
nor U9557 (N_9557,N_6083,N_7387);
xor U9558 (N_9558,N_7394,N_7071);
nand U9559 (N_9559,N_7903,N_7386);
or U9560 (N_9560,N_6070,N_7004);
nor U9561 (N_9561,N_6009,N_7359);
xnor U9562 (N_9562,N_7838,N_7650);
nor U9563 (N_9563,N_7453,N_6160);
nand U9564 (N_9564,N_6913,N_7867);
nand U9565 (N_9565,N_6797,N_7918);
nor U9566 (N_9566,N_7539,N_6734);
nand U9567 (N_9567,N_7109,N_6686);
xor U9568 (N_9568,N_7546,N_7472);
nor U9569 (N_9569,N_7053,N_6469);
and U9570 (N_9570,N_7863,N_6160);
xnor U9571 (N_9571,N_7390,N_6544);
nor U9572 (N_9572,N_7094,N_7872);
nand U9573 (N_9573,N_6065,N_6606);
and U9574 (N_9574,N_6879,N_6661);
nand U9575 (N_9575,N_6458,N_7148);
xnor U9576 (N_9576,N_6644,N_6240);
and U9577 (N_9577,N_6927,N_7398);
or U9578 (N_9578,N_7097,N_6844);
nor U9579 (N_9579,N_6273,N_7446);
and U9580 (N_9580,N_7217,N_6403);
nor U9581 (N_9581,N_7456,N_7729);
xor U9582 (N_9582,N_6722,N_6658);
xnor U9583 (N_9583,N_7022,N_7893);
nor U9584 (N_9584,N_6160,N_7844);
nor U9585 (N_9585,N_6967,N_7704);
or U9586 (N_9586,N_6082,N_7717);
xnor U9587 (N_9587,N_7297,N_7681);
nand U9588 (N_9588,N_7594,N_7962);
nor U9589 (N_9589,N_6566,N_7636);
nand U9590 (N_9590,N_6671,N_7882);
or U9591 (N_9591,N_6899,N_6036);
and U9592 (N_9592,N_7477,N_7336);
xor U9593 (N_9593,N_7355,N_7789);
nor U9594 (N_9594,N_6195,N_7278);
and U9595 (N_9595,N_7376,N_7007);
nand U9596 (N_9596,N_6965,N_6077);
or U9597 (N_9597,N_6264,N_7822);
xnor U9598 (N_9598,N_6738,N_7075);
xor U9599 (N_9599,N_6757,N_6205);
and U9600 (N_9600,N_6897,N_7950);
nand U9601 (N_9601,N_6191,N_6787);
and U9602 (N_9602,N_7056,N_7443);
nand U9603 (N_9603,N_6119,N_7803);
xnor U9604 (N_9604,N_6492,N_7622);
and U9605 (N_9605,N_6623,N_7591);
nand U9606 (N_9606,N_7487,N_7689);
xnor U9607 (N_9607,N_6812,N_7137);
and U9608 (N_9608,N_7568,N_6804);
nor U9609 (N_9609,N_6658,N_7637);
or U9610 (N_9610,N_6459,N_6887);
nor U9611 (N_9611,N_6102,N_6271);
xnor U9612 (N_9612,N_6211,N_6196);
xor U9613 (N_9613,N_6495,N_7076);
and U9614 (N_9614,N_6290,N_6775);
nor U9615 (N_9615,N_6206,N_6227);
or U9616 (N_9616,N_6606,N_6594);
nand U9617 (N_9617,N_7355,N_7890);
or U9618 (N_9618,N_7271,N_6335);
nand U9619 (N_9619,N_7701,N_7040);
xnor U9620 (N_9620,N_7821,N_7557);
xor U9621 (N_9621,N_7471,N_7436);
nand U9622 (N_9622,N_7352,N_6046);
and U9623 (N_9623,N_7165,N_6703);
and U9624 (N_9624,N_7481,N_7880);
nand U9625 (N_9625,N_7014,N_7715);
nor U9626 (N_9626,N_6815,N_6288);
xnor U9627 (N_9627,N_7199,N_7212);
nand U9628 (N_9628,N_7683,N_6709);
xnor U9629 (N_9629,N_7218,N_6576);
nor U9630 (N_9630,N_6065,N_6059);
nand U9631 (N_9631,N_6330,N_7555);
and U9632 (N_9632,N_7987,N_7301);
nand U9633 (N_9633,N_7376,N_7927);
or U9634 (N_9634,N_6363,N_6294);
nor U9635 (N_9635,N_6714,N_7436);
and U9636 (N_9636,N_6516,N_6671);
nand U9637 (N_9637,N_6955,N_7528);
and U9638 (N_9638,N_7938,N_7315);
or U9639 (N_9639,N_7961,N_6435);
and U9640 (N_9640,N_6606,N_6344);
nand U9641 (N_9641,N_7814,N_6825);
or U9642 (N_9642,N_7853,N_6168);
xnor U9643 (N_9643,N_6208,N_6726);
nor U9644 (N_9644,N_7768,N_7171);
xnor U9645 (N_9645,N_7889,N_7575);
xnor U9646 (N_9646,N_7832,N_7014);
xor U9647 (N_9647,N_7304,N_6170);
or U9648 (N_9648,N_6242,N_7540);
xor U9649 (N_9649,N_7704,N_7778);
and U9650 (N_9650,N_7105,N_7381);
xor U9651 (N_9651,N_6054,N_7991);
nor U9652 (N_9652,N_7705,N_6380);
xor U9653 (N_9653,N_6064,N_6184);
and U9654 (N_9654,N_7370,N_7758);
nor U9655 (N_9655,N_6833,N_7334);
or U9656 (N_9656,N_7247,N_7035);
xnor U9657 (N_9657,N_6795,N_7318);
nor U9658 (N_9658,N_6692,N_6879);
nor U9659 (N_9659,N_7613,N_6852);
and U9660 (N_9660,N_6354,N_6839);
xor U9661 (N_9661,N_6095,N_6826);
xor U9662 (N_9662,N_6028,N_6268);
or U9663 (N_9663,N_6463,N_7147);
xnor U9664 (N_9664,N_6215,N_6700);
xnor U9665 (N_9665,N_7473,N_7016);
and U9666 (N_9666,N_7280,N_6918);
or U9667 (N_9667,N_7828,N_6114);
nor U9668 (N_9668,N_7087,N_7031);
xor U9669 (N_9669,N_6119,N_7105);
or U9670 (N_9670,N_6825,N_6948);
or U9671 (N_9671,N_7940,N_6997);
xor U9672 (N_9672,N_7287,N_7366);
nor U9673 (N_9673,N_7972,N_7800);
nand U9674 (N_9674,N_7858,N_6269);
nor U9675 (N_9675,N_6773,N_6573);
nand U9676 (N_9676,N_7568,N_6355);
xnor U9677 (N_9677,N_7632,N_6107);
nand U9678 (N_9678,N_7587,N_6105);
or U9679 (N_9679,N_6185,N_7689);
or U9680 (N_9680,N_6659,N_7903);
nand U9681 (N_9681,N_7958,N_6370);
nor U9682 (N_9682,N_7866,N_6536);
xor U9683 (N_9683,N_6796,N_6985);
and U9684 (N_9684,N_7028,N_6130);
or U9685 (N_9685,N_7409,N_7104);
or U9686 (N_9686,N_7847,N_6158);
and U9687 (N_9687,N_6278,N_6091);
xor U9688 (N_9688,N_7818,N_7158);
nor U9689 (N_9689,N_7390,N_6603);
and U9690 (N_9690,N_6796,N_7260);
xor U9691 (N_9691,N_7026,N_6833);
or U9692 (N_9692,N_6117,N_7479);
and U9693 (N_9693,N_7015,N_6075);
nor U9694 (N_9694,N_6995,N_6798);
nor U9695 (N_9695,N_6346,N_6733);
nor U9696 (N_9696,N_7137,N_7075);
and U9697 (N_9697,N_6488,N_6423);
and U9698 (N_9698,N_7241,N_6181);
xnor U9699 (N_9699,N_6424,N_7510);
xor U9700 (N_9700,N_6905,N_7270);
nand U9701 (N_9701,N_7220,N_7295);
or U9702 (N_9702,N_7614,N_7764);
nand U9703 (N_9703,N_6139,N_6768);
nor U9704 (N_9704,N_6079,N_6379);
xor U9705 (N_9705,N_6635,N_6525);
or U9706 (N_9706,N_6750,N_7763);
nor U9707 (N_9707,N_6972,N_6923);
nor U9708 (N_9708,N_6004,N_6044);
xor U9709 (N_9709,N_7751,N_7775);
nand U9710 (N_9710,N_7175,N_6541);
nand U9711 (N_9711,N_6509,N_7247);
or U9712 (N_9712,N_6672,N_6676);
nand U9713 (N_9713,N_7622,N_7221);
and U9714 (N_9714,N_6199,N_7494);
nor U9715 (N_9715,N_7693,N_7156);
xnor U9716 (N_9716,N_7292,N_6761);
and U9717 (N_9717,N_6654,N_6194);
and U9718 (N_9718,N_7018,N_6826);
nand U9719 (N_9719,N_7275,N_6701);
nor U9720 (N_9720,N_6704,N_6941);
and U9721 (N_9721,N_6586,N_6360);
xnor U9722 (N_9722,N_7808,N_7227);
or U9723 (N_9723,N_6353,N_7721);
nor U9724 (N_9724,N_7834,N_6587);
nand U9725 (N_9725,N_7139,N_7152);
or U9726 (N_9726,N_6895,N_7559);
and U9727 (N_9727,N_6081,N_6611);
or U9728 (N_9728,N_6880,N_7381);
or U9729 (N_9729,N_6137,N_7652);
xnor U9730 (N_9730,N_6920,N_6848);
or U9731 (N_9731,N_7342,N_7866);
and U9732 (N_9732,N_7117,N_7860);
nand U9733 (N_9733,N_7233,N_7573);
or U9734 (N_9734,N_7921,N_6791);
nand U9735 (N_9735,N_7335,N_7126);
and U9736 (N_9736,N_6122,N_7025);
nand U9737 (N_9737,N_6645,N_6641);
xnor U9738 (N_9738,N_6890,N_6641);
xor U9739 (N_9739,N_7923,N_6811);
and U9740 (N_9740,N_6905,N_6098);
xnor U9741 (N_9741,N_6020,N_7108);
nand U9742 (N_9742,N_7216,N_7563);
xnor U9743 (N_9743,N_6801,N_7940);
nor U9744 (N_9744,N_6372,N_6309);
or U9745 (N_9745,N_7814,N_6557);
and U9746 (N_9746,N_6118,N_6751);
nand U9747 (N_9747,N_7613,N_6976);
or U9748 (N_9748,N_6406,N_6005);
xnor U9749 (N_9749,N_6066,N_7099);
and U9750 (N_9750,N_6244,N_6024);
nand U9751 (N_9751,N_7063,N_6964);
nand U9752 (N_9752,N_6473,N_7575);
xor U9753 (N_9753,N_7539,N_6286);
xor U9754 (N_9754,N_6050,N_6131);
or U9755 (N_9755,N_6640,N_7994);
xnor U9756 (N_9756,N_6611,N_6105);
and U9757 (N_9757,N_6701,N_7930);
xor U9758 (N_9758,N_6700,N_7984);
and U9759 (N_9759,N_6411,N_7320);
and U9760 (N_9760,N_7428,N_6120);
nor U9761 (N_9761,N_7959,N_6372);
xor U9762 (N_9762,N_7273,N_6834);
nand U9763 (N_9763,N_7922,N_7987);
xnor U9764 (N_9764,N_7571,N_6645);
nand U9765 (N_9765,N_6732,N_6553);
and U9766 (N_9766,N_6746,N_7186);
xnor U9767 (N_9767,N_6177,N_7728);
or U9768 (N_9768,N_6956,N_6202);
or U9769 (N_9769,N_7725,N_6846);
and U9770 (N_9770,N_6374,N_7793);
nor U9771 (N_9771,N_6417,N_7342);
or U9772 (N_9772,N_7275,N_7373);
and U9773 (N_9773,N_6964,N_6985);
nand U9774 (N_9774,N_7526,N_6782);
xor U9775 (N_9775,N_6497,N_7995);
or U9776 (N_9776,N_6045,N_6893);
or U9777 (N_9777,N_6704,N_6054);
nor U9778 (N_9778,N_6591,N_7939);
and U9779 (N_9779,N_6639,N_7231);
xor U9780 (N_9780,N_7714,N_6167);
and U9781 (N_9781,N_6447,N_6509);
nor U9782 (N_9782,N_7706,N_7760);
nor U9783 (N_9783,N_7737,N_6128);
xor U9784 (N_9784,N_6472,N_7174);
or U9785 (N_9785,N_6466,N_7206);
xor U9786 (N_9786,N_7560,N_6344);
and U9787 (N_9787,N_7342,N_7489);
nand U9788 (N_9788,N_6821,N_7324);
or U9789 (N_9789,N_7086,N_7503);
nand U9790 (N_9790,N_6597,N_7519);
nand U9791 (N_9791,N_6743,N_7492);
nand U9792 (N_9792,N_6808,N_6930);
xor U9793 (N_9793,N_6619,N_7615);
nor U9794 (N_9794,N_7824,N_7902);
and U9795 (N_9795,N_7625,N_7956);
nand U9796 (N_9796,N_6452,N_6242);
and U9797 (N_9797,N_7370,N_6484);
nand U9798 (N_9798,N_7179,N_6810);
and U9799 (N_9799,N_6819,N_7272);
xnor U9800 (N_9800,N_6345,N_7117);
xnor U9801 (N_9801,N_6683,N_6696);
nor U9802 (N_9802,N_6994,N_7386);
or U9803 (N_9803,N_6685,N_6717);
nor U9804 (N_9804,N_6156,N_7703);
and U9805 (N_9805,N_7266,N_7856);
or U9806 (N_9806,N_6828,N_7917);
xor U9807 (N_9807,N_6185,N_7699);
xor U9808 (N_9808,N_6236,N_7699);
nor U9809 (N_9809,N_6614,N_6759);
nand U9810 (N_9810,N_7982,N_6502);
xor U9811 (N_9811,N_6291,N_6423);
or U9812 (N_9812,N_7377,N_6578);
nand U9813 (N_9813,N_6595,N_7091);
and U9814 (N_9814,N_6823,N_6248);
nand U9815 (N_9815,N_6686,N_7502);
nand U9816 (N_9816,N_7043,N_6462);
and U9817 (N_9817,N_7614,N_6435);
or U9818 (N_9818,N_6751,N_7559);
and U9819 (N_9819,N_7232,N_6618);
or U9820 (N_9820,N_7153,N_6477);
nor U9821 (N_9821,N_6951,N_6544);
xnor U9822 (N_9822,N_7452,N_7035);
and U9823 (N_9823,N_7337,N_6703);
nand U9824 (N_9824,N_6468,N_7126);
and U9825 (N_9825,N_6263,N_6553);
or U9826 (N_9826,N_6944,N_6818);
nand U9827 (N_9827,N_6966,N_7181);
nor U9828 (N_9828,N_6555,N_7610);
or U9829 (N_9829,N_6080,N_7349);
nor U9830 (N_9830,N_6148,N_6042);
or U9831 (N_9831,N_6117,N_7251);
xnor U9832 (N_9832,N_7632,N_7338);
xnor U9833 (N_9833,N_7413,N_6875);
or U9834 (N_9834,N_7773,N_7873);
xnor U9835 (N_9835,N_6126,N_6197);
nor U9836 (N_9836,N_6761,N_6822);
nor U9837 (N_9837,N_7854,N_6505);
nor U9838 (N_9838,N_6663,N_6295);
nor U9839 (N_9839,N_7718,N_6434);
nand U9840 (N_9840,N_7322,N_7885);
and U9841 (N_9841,N_7284,N_6887);
xnor U9842 (N_9842,N_6279,N_6302);
and U9843 (N_9843,N_7733,N_6489);
nand U9844 (N_9844,N_7498,N_7157);
nor U9845 (N_9845,N_7837,N_7647);
xnor U9846 (N_9846,N_6740,N_6698);
nand U9847 (N_9847,N_7369,N_7606);
nand U9848 (N_9848,N_7029,N_6583);
and U9849 (N_9849,N_6400,N_6427);
and U9850 (N_9850,N_6226,N_6213);
xnor U9851 (N_9851,N_6039,N_7063);
nand U9852 (N_9852,N_6998,N_7385);
nand U9853 (N_9853,N_6330,N_7077);
xor U9854 (N_9854,N_7223,N_7055);
or U9855 (N_9855,N_7340,N_7440);
or U9856 (N_9856,N_6562,N_6894);
and U9857 (N_9857,N_6134,N_6463);
and U9858 (N_9858,N_6916,N_6149);
and U9859 (N_9859,N_7245,N_6285);
nand U9860 (N_9860,N_7540,N_7754);
nor U9861 (N_9861,N_7049,N_6000);
nand U9862 (N_9862,N_7658,N_6198);
and U9863 (N_9863,N_6669,N_6863);
nor U9864 (N_9864,N_7384,N_7295);
xnor U9865 (N_9865,N_6878,N_6217);
nand U9866 (N_9866,N_6214,N_6141);
nand U9867 (N_9867,N_6455,N_6764);
nand U9868 (N_9868,N_6128,N_7458);
or U9869 (N_9869,N_6141,N_7951);
and U9870 (N_9870,N_7912,N_6441);
or U9871 (N_9871,N_7325,N_6980);
xor U9872 (N_9872,N_6868,N_7030);
and U9873 (N_9873,N_7013,N_7110);
xnor U9874 (N_9874,N_6976,N_6446);
or U9875 (N_9875,N_6072,N_7859);
or U9876 (N_9876,N_6938,N_6292);
nor U9877 (N_9877,N_7677,N_7676);
xor U9878 (N_9878,N_7789,N_7898);
xnor U9879 (N_9879,N_6782,N_7339);
nor U9880 (N_9880,N_6140,N_6728);
or U9881 (N_9881,N_7114,N_6242);
nor U9882 (N_9882,N_6330,N_7453);
nand U9883 (N_9883,N_7805,N_7976);
and U9884 (N_9884,N_7931,N_7312);
nand U9885 (N_9885,N_6009,N_6157);
xnor U9886 (N_9886,N_7532,N_6249);
nor U9887 (N_9887,N_6145,N_7881);
nand U9888 (N_9888,N_6838,N_7426);
or U9889 (N_9889,N_7200,N_7492);
nor U9890 (N_9890,N_7088,N_6318);
nor U9891 (N_9891,N_6947,N_6756);
xnor U9892 (N_9892,N_6973,N_7850);
and U9893 (N_9893,N_6733,N_7068);
nand U9894 (N_9894,N_7108,N_7616);
or U9895 (N_9895,N_6459,N_6650);
xor U9896 (N_9896,N_6994,N_6864);
xor U9897 (N_9897,N_7390,N_6574);
or U9898 (N_9898,N_7008,N_6705);
and U9899 (N_9899,N_7744,N_7639);
nor U9900 (N_9900,N_7303,N_7774);
nand U9901 (N_9901,N_7866,N_6308);
xor U9902 (N_9902,N_6540,N_7589);
and U9903 (N_9903,N_7714,N_6737);
nor U9904 (N_9904,N_6832,N_7802);
and U9905 (N_9905,N_6625,N_7247);
nand U9906 (N_9906,N_6998,N_6092);
or U9907 (N_9907,N_6365,N_6998);
xnor U9908 (N_9908,N_6749,N_6532);
nor U9909 (N_9909,N_6630,N_7692);
nand U9910 (N_9910,N_6206,N_7955);
and U9911 (N_9911,N_6804,N_6103);
nor U9912 (N_9912,N_6144,N_6518);
nand U9913 (N_9913,N_6715,N_6912);
xnor U9914 (N_9914,N_7713,N_6849);
nor U9915 (N_9915,N_7745,N_7177);
nand U9916 (N_9916,N_6370,N_7767);
xnor U9917 (N_9917,N_7987,N_6184);
nor U9918 (N_9918,N_6335,N_6652);
or U9919 (N_9919,N_7631,N_6386);
and U9920 (N_9920,N_7145,N_7835);
nor U9921 (N_9921,N_7542,N_7251);
and U9922 (N_9922,N_6400,N_7975);
and U9923 (N_9923,N_6527,N_6453);
nand U9924 (N_9924,N_6801,N_6706);
or U9925 (N_9925,N_6395,N_6154);
nor U9926 (N_9926,N_7243,N_6906);
xor U9927 (N_9927,N_6516,N_6452);
nor U9928 (N_9928,N_7620,N_6380);
and U9929 (N_9929,N_7604,N_6240);
or U9930 (N_9930,N_6840,N_6040);
xnor U9931 (N_9931,N_6311,N_6557);
or U9932 (N_9932,N_7241,N_7631);
or U9933 (N_9933,N_6987,N_7062);
nand U9934 (N_9934,N_6443,N_6317);
nor U9935 (N_9935,N_6985,N_6704);
and U9936 (N_9936,N_6262,N_6851);
nand U9937 (N_9937,N_7180,N_7422);
nand U9938 (N_9938,N_6978,N_7225);
xnor U9939 (N_9939,N_7304,N_6993);
and U9940 (N_9940,N_7540,N_7820);
nor U9941 (N_9941,N_7547,N_6058);
xnor U9942 (N_9942,N_6264,N_6426);
xor U9943 (N_9943,N_6899,N_7766);
nor U9944 (N_9944,N_7972,N_7321);
nand U9945 (N_9945,N_7471,N_7124);
or U9946 (N_9946,N_7247,N_6791);
nor U9947 (N_9947,N_7871,N_6998);
or U9948 (N_9948,N_7174,N_7653);
nor U9949 (N_9949,N_7268,N_7432);
nor U9950 (N_9950,N_7985,N_6933);
nand U9951 (N_9951,N_6195,N_7525);
or U9952 (N_9952,N_6769,N_7141);
and U9953 (N_9953,N_6843,N_6512);
nor U9954 (N_9954,N_6165,N_7993);
and U9955 (N_9955,N_6665,N_7545);
nor U9956 (N_9956,N_6408,N_6265);
nand U9957 (N_9957,N_7192,N_6890);
and U9958 (N_9958,N_7192,N_7022);
nor U9959 (N_9959,N_7886,N_7144);
xnor U9960 (N_9960,N_7529,N_6086);
nor U9961 (N_9961,N_6130,N_6722);
or U9962 (N_9962,N_7427,N_6625);
or U9963 (N_9963,N_6768,N_7549);
and U9964 (N_9964,N_7732,N_6647);
nand U9965 (N_9965,N_6876,N_6088);
xnor U9966 (N_9966,N_7571,N_6274);
nand U9967 (N_9967,N_6932,N_6613);
nor U9968 (N_9968,N_6970,N_7745);
or U9969 (N_9969,N_7616,N_7564);
and U9970 (N_9970,N_6748,N_6143);
nand U9971 (N_9971,N_7778,N_7886);
nor U9972 (N_9972,N_7470,N_7511);
and U9973 (N_9973,N_7794,N_6160);
xor U9974 (N_9974,N_6375,N_6881);
or U9975 (N_9975,N_6203,N_7535);
or U9976 (N_9976,N_6689,N_6472);
or U9977 (N_9977,N_6721,N_6051);
or U9978 (N_9978,N_6552,N_6188);
nor U9979 (N_9979,N_7379,N_7060);
nor U9980 (N_9980,N_7062,N_7939);
and U9981 (N_9981,N_6893,N_7773);
and U9982 (N_9982,N_6268,N_6115);
nor U9983 (N_9983,N_7129,N_6908);
or U9984 (N_9984,N_7967,N_6681);
nor U9985 (N_9985,N_7684,N_7159);
nand U9986 (N_9986,N_7466,N_7469);
nor U9987 (N_9987,N_6210,N_7790);
xor U9988 (N_9988,N_7330,N_7056);
nor U9989 (N_9989,N_7772,N_7527);
nand U9990 (N_9990,N_7189,N_7614);
xnor U9991 (N_9991,N_6460,N_6800);
or U9992 (N_9992,N_6451,N_7855);
and U9993 (N_9993,N_7999,N_6221);
xor U9994 (N_9994,N_6199,N_6348);
xnor U9995 (N_9995,N_7613,N_7849);
nor U9996 (N_9996,N_6795,N_7616);
or U9997 (N_9997,N_7953,N_6691);
nor U9998 (N_9998,N_7741,N_6195);
nor U9999 (N_9999,N_7842,N_7324);
nand UO_0 (O_0,N_8465,N_8260);
nand UO_1 (O_1,N_8309,N_9424);
and UO_2 (O_2,N_8963,N_8106);
nand UO_3 (O_3,N_9375,N_9290);
or UO_4 (O_4,N_9719,N_8801);
and UO_5 (O_5,N_9260,N_8211);
xnor UO_6 (O_6,N_9744,N_9156);
nor UO_7 (O_7,N_9953,N_8476);
nand UO_8 (O_8,N_8618,N_8179);
and UO_9 (O_9,N_9635,N_8520);
xnor UO_10 (O_10,N_9237,N_9247);
nand UO_11 (O_11,N_9298,N_8331);
nor UO_12 (O_12,N_8605,N_9798);
nor UO_13 (O_13,N_9334,N_9741);
or UO_14 (O_14,N_8158,N_9687);
xor UO_15 (O_15,N_8032,N_8300);
and UO_16 (O_16,N_9745,N_8351);
nand UO_17 (O_17,N_9531,N_9326);
nor UO_18 (O_18,N_9792,N_9048);
or UO_19 (O_19,N_9561,N_8288);
nor UO_20 (O_20,N_8339,N_8171);
and UO_21 (O_21,N_9128,N_9279);
nand UO_22 (O_22,N_8431,N_8494);
or UO_23 (O_23,N_8362,N_8663);
or UO_24 (O_24,N_9732,N_8048);
nor UO_25 (O_25,N_9336,N_8312);
nand UO_26 (O_26,N_8680,N_9416);
nor UO_27 (O_27,N_9180,N_8940);
xor UO_28 (O_28,N_8974,N_8917);
or UO_29 (O_29,N_8567,N_8482);
or UO_30 (O_30,N_8378,N_8376);
nor UO_31 (O_31,N_9082,N_9870);
xnor UO_32 (O_32,N_9008,N_8207);
xor UO_33 (O_33,N_9500,N_8898);
nor UO_34 (O_34,N_8695,N_8070);
nand UO_35 (O_35,N_9620,N_9931);
xor UO_36 (O_36,N_9928,N_8538);
and UO_37 (O_37,N_9236,N_9311);
nand UO_38 (O_38,N_9878,N_8959);
or UO_39 (O_39,N_9027,N_9625);
and UO_40 (O_40,N_9495,N_9589);
nor UO_41 (O_41,N_9426,N_9694);
xnor UO_42 (O_42,N_8140,N_8793);
or UO_43 (O_43,N_9276,N_9886);
xor UO_44 (O_44,N_8706,N_9302);
or UO_45 (O_45,N_9513,N_8560);
nand UO_46 (O_46,N_8303,N_9806);
nand UO_47 (O_47,N_8758,N_9618);
nand UO_48 (O_48,N_8224,N_8647);
and UO_49 (O_49,N_8009,N_9482);
xnor UO_50 (O_50,N_9207,N_8664);
or UO_51 (O_51,N_8841,N_9445);
xnor UO_52 (O_52,N_8532,N_9571);
nor UO_53 (O_53,N_8585,N_9564);
xnor UO_54 (O_54,N_8789,N_9491);
or UO_55 (O_55,N_8530,N_9056);
nand UO_56 (O_56,N_8537,N_9164);
nor UO_57 (O_57,N_9391,N_8846);
and UO_58 (O_58,N_9986,N_8993);
nor UO_59 (O_59,N_8285,N_8772);
and UO_60 (O_60,N_8679,N_9652);
nor UO_61 (O_61,N_8548,N_9304);
nand UO_62 (O_62,N_9592,N_9348);
nand UO_63 (O_63,N_8791,N_9922);
nor UO_64 (O_64,N_9095,N_8095);
or UO_65 (O_65,N_8135,N_8019);
or UO_66 (O_66,N_8874,N_9990);
and UO_67 (O_67,N_9672,N_8341);
xnor UO_68 (O_68,N_9114,N_8077);
xnor UO_69 (O_69,N_8924,N_8512);
nor UO_70 (O_70,N_8083,N_8643);
and UO_71 (O_71,N_8030,N_9425);
nor UO_72 (O_72,N_9154,N_9457);
nand UO_73 (O_73,N_9765,N_8258);
nor UO_74 (O_74,N_9427,N_8667);
nor UO_75 (O_75,N_9955,N_9402);
nor UO_76 (O_76,N_8594,N_8380);
nand UO_77 (O_77,N_9357,N_8366);
or UO_78 (O_78,N_8901,N_9176);
and UO_79 (O_79,N_8755,N_8635);
or UO_80 (O_80,N_9573,N_8481);
and UO_81 (O_81,N_9373,N_8435);
nor UO_82 (O_82,N_8098,N_8005);
nor UO_83 (O_83,N_8557,N_8725);
xor UO_84 (O_84,N_9430,N_8167);
nor UO_85 (O_85,N_9684,N_8323);
nor UO_86 (O_86,N_9774,N_9847);
and UO_87 (O_87,N_8017,N_9674);
xnor UO_88 (O_88,N_9204,N_9789);
nor UO_89 (O_89,N_8790,N_9935);
or UO_90 (O_90,N_9645,N_9855);
nor UO_91 (O_91,N_9602,N_9601);
xor UO_92 (O_92,N_9567,N_9401);
nor UO_93 (O_93,N_8838,N_8797);
or UO_94 (O_94,N_8177,N_9605);
xnor UO_95 (O_95,N_8774,N_9079);
and UO_96 (O_96,N_8081,N_9775);
and UO_97 (O_97,N_9845,N_8469);
xor UO_98 (O_98,N_9581,N_9702);
nor UO_99 (O_99,N_8650,N_9210);
nand UO_100 (O_100,N_9570,N_8393);
xnor UO_101 (O_101,N_9244,N_8641);
xnor UO_102 (O_102,N_8632,N_9211);
nand UO_103 (O_103,N_8737,N_9381);
nand UO_104 (O_104,N_8620,N_8525);
xnor UO_105 (O_105,N_9643,N_9671);
and UO_106 (O_106,N_9194,N_8496);
nor UO_107 (O_107,N_9469,N_9165);
nor UO_108 (O_108,N_8299,N_8052);
nand UO_109 (O_109,N_9738,N_8832);
nand UO_110 (O_110,N_8584,N_8455);
nand UO_111 (O_111,N_8028,N_9594);
xor UO_112 (O_112,N_9320,N_9012);
and UO_113 (O_113,N_8085,N_9834);
nor UO_114 (O_114,N_9523,N_8876);
nand UO_115 (O_115,N_9026,N_8619);
nor UO_116 (O_116,N_9436,N_9807);
or UO_117 (O_117,N_8792,N_8571);
and UO_118 (O_118,N_9428,N_8405);
and UO_119 (O_119,N_8382,N_9413);
nor UO_120 (O_120,N_9393,N_8069);
xor UO_121 (O_121,N_9225,N_8346);
xnor UO_122 (O_122,N_8960,N_9317);
and UO_123 (O_123,N_8334,N_8989);
nand UO_124 (O_124,N_9239,N_8973);
or UO_125 (O_125,N_9733,N_9188);
xnor UO_126 (O_126,N_9748,N_9031);
and UO_127 (O_127,N_9212,N_9910);
nor UO_128 (O_128,N_8250,N_9947);
nor UO_129 (O_129,N_8996,N_9734);
and UO_130 (O_130,N_9174,N_9119);
or UO_131 (O_131,N_8319,N_9690);
nand UO_132 (O_132,N_8436,N_9499);
nor UO_133 (O_133,N_8698,N_9576);
nand UO_134 (O_134,N_9527,N_8452);
xnor UO_135 (O_135,N_9150,N_8416);
nand UO_136 (O_136,N_9988,N_8534);
or UO_137 (O_137,N_9053,N_9697);
nand UO_138 (O_138,N_9784,N_8675);
or UO_139 (O_139,N_8872,N_8753);
and UO_140 (O_140,N_9562,N_8951);
nor UO_141 (O_141,N_9462,N_8297);
nand UO_142 (O_142,N_8308,N_8626);
and UO_143 (O_143,N_8131,N_8552);
or UO_144 (O_144,N_9369,N_8591);
nor UO_145 (O_145,N_8249,N_8922);
and UO_146 (O_146,N_9431,N_8780);
nand UO_147 (O_147,N_8875,N_8350);
nand UO_148 (O_148,N_8153,N_9812);
xnor UO_149 (O_149,N_9315,N_9217);
or UO_150 (O_150,N_9778,N_8598);
and UO_151 (O_151,N_8910,N_9704);
or UO_152 (O_152,N_8451,N_9017);
and UO_153 (O_153,N_9899,N_8742);
nor UO_154 (O_154,N_8592,N_9448);
and UO_155 (O_155,N_8627,N_8155);
nor UO_156 (O_156,N_8479,N_8168);
and UO_157 (O_157,N_9088,N_9216);
or UO_158 (O_158,N_9429,N_8244);
nor UO_159 (O_159,N_8890,N_8246);
nand UO_160 (O_160,N_9084,N_8292);
or UO_161 (O_161,N_9337,N_9591);
nor UO_162 (O_162,N_8317,N_9264);
and UO_163 (O_163,N_9065,N_9747);
xnor UO_164 (O_164,N_8007,N_9032);
nand UO_165 (O_165,N_9912,N_9272);
and UO_166 (O_166,N_9406,N_8716);
xnor UO_167 (O_167,N_9545,N_9742);
xor UO_168 (O_168,N_8337,N_8550);
and UO_169 (O_169,N_8196,N_8603);
xor UO_170 (O_170,N_8900,N_9900);
nor UO_171 (O_171,N_9363,N_9170);
nor UO_172 (O_172,N_9725,N_9287);
xor UO_173 (O_173,N_9916,N_9408);
xor UO_174 (O_174,N_9177,N_9667);
and UO_175 (O_175,N_8929,N_8835);
nand UO_176 (O_176,N_8545,N_9437);
nor UO_177 (O_177,N_9965,N_9465);
or UO_178 (O_178,N_8105,N_8180);
or UO_179 (O_179,N_9354,N_9121);
xor UO_180 (O_180,N_9658,N_9246);
xor UO_181 (O_181,N_8785,N_8713);
nand UO_182 (O_182,N_8779,N_8810);
and UO_183 (O_183,N_9587,N_8109);
or UO_184 (O_184,N_8216,N_9875);
or UO_185 (O_185,N_8390,N_9766);
nor UO_186 (O_186,N_9650,N_8414);
nand UO_187 (O_187,N_9323,N_9321);
nand UO_188 (O_188,N_9187,N_8665);
xnor UO_189 (O_189,N_8885,N_9838);
or UO_190 (O_190,N_8076,N_9286);
nand UO_191 (O_191,N_9941,N_9699);
nor UO_192 (O_192,N_9484,N_9062);
xnor UO_193 (O_193,N_8824,N_9535);
nand UO_194 (O_194,N_9863,N_9023);
xnor UO_195 (O_195,N_9479,N_9314);
nand UO_196 (O_196,N_9559,N_9473);
nand UO_197 (O_197,N_8068,N_8651);
nor UO_198 (O_198,N_8072,N_9481);
xnor UO_199 (O_199,N_8638,N_8247);
or UO_200 (O_200,N_9558,N_8873);
and UO_201 (O_201,N_8046,N_9809);
nor UO_202 (O_202,N_9035,N_9967);
xor UO_203 (O_203,N_8808,N_9383);
nor UO_204 (O_204,N_9782,N_9621);
nor UO_205 (O_205,N_8287,N_8492);
nand UO_206 (O_206,N_9994,N_9140);
xnor UO_207 (O_207,N_8542,N_8255);
nor UO_208 (O_208,N_9772,N_8554);
xnor UO_209 (O_209,N_9464,N_8031);
and UO_210 (O_210,N_9821,N_9917);
and UO_211 (O_211,N_9388,N_9395);
nor UO_212 (O_212,N_9692,N_9467);
and UO_213 (O_213,N_8986,N_8368);
nand UO_214 (O_214,N_9322,N_8558);
nand UO_215 (O_215,N_9136,N_9492);
and UO_216 (O_216,N_8189,N_9629);
nor UO_217 (O_217,N_9546,N_8187);
nor UO_218 (O_218,N_9390,N_9030);
nand UO_219 (O_219,N_8448,N_9028);
nor UO_220 (O_220,N_8373,N_9083);
xnor UO_221 (O_221,N_8485,N_8021);
nor UO_222 (O_222,N_9593,N_9989);
nand UO_223 (O_223,N_8833,N_9544);
and UO_224 (O_224,N_9743,N_9574);
and UO_225 (O_225,N_9312,N_9343);
xor UO_226 (O_226,N_8461,N_9832);
nand UO_227 (O_227,N_8689,N_8787);
and UO_228 (O_228,N_8209,N_8112);
xor UO_229 (O_229,N_8355,N_9072);
nor UO_230 (O_230,N_9112,N_9793);
or UO_231 (O_231,N_8977,N_9346);
or UO_232 (O_232,N_8907,N_9355);
xnor UO_233 (O_233,N_8181,N_8256);
nor UO_234 (O_234,N_9708,N_9046);
xnor UO_235 (O_235,N_9496,N_9514);
nand UO_236 (O_236,N_8904,N_8369);
or UO_237 (O_237,N_8082,N_8043);
nand UO_238 (O_238,N_9737,N_9915);
nand UO_239 (O_239,N_8434,N_9685);
nand UO_240 (O_240,N_8586,N_9932);
nand UO_241 (O_241,N_9344,N_8002);
xor UO_242 (O_242,N_9435,N_8061);
nand UO_243 (O_243,N_8908,N_8652);
nand UO_244 (O_244,N_9754,N_8212);
nor UO_245 (O_245,N_9963,N_8734);
or UO_246 (O_246,N_8051,N_9584);
nand UO_247 (O_247,N_8539,N_9485);
xnor UO_248 (O_248,N_8225,N_9328);
xor UO_249 (O_249,N_9161,N_8912);
xor UO_250 (O_250,N_9192,N_9933);
and UO_251 (O_251,N_9862,N_8536);
and UO_252 (O_252,N_9813,N_9257);
xnor UO_253 (O_253,N_8463,N_8524);
or UO_254 (O_254,N_8543,N_9971);
xor UO_255 (O_255,N_8360,N_8844);
or UO_256 (O_256,N_8422,N_8157);
nor UO_257 (O_257,N_9477,N_9403);
xnor UO_258 (O_258,N_9706,N_9679);
or UO_259 (O_259,N_9631,N_9441);
xor UO_260 (O_260,N_9162,N_9528);
and UO_261 (O_261,N_8279,N_8273);
or UO_262 (O_262,N_8175,N_9104);
and UO_263 (O_263,N_8549,N_8709);
nand UO_264 (O_264,N_9726,N_8577);
or UO_265 (O_265,N_9245,N_8745);
or UO_266 (O_266,N_9221,N_9010);
nand UO_267 (O_267,N_8636,N_9157);
or UO_268 (O_268,N_8869,N_9506);
and UO_269 (O_269,N_8442,N_9033);
and UO_270 (O_270,N_9099,N_9818);
nor UO_271 (O_271,N_8354,N_8814);
nand UO_272 (O_272,N_8796,N_8428);
or UO_273 (O_273,N_9583,N_8163);
nor UO_274 (O_274,N_8719,N_9773);
and UO_275 (O_275,N_9653,N_9108);
nand UO_276 (O_276,N_8639,N_8381);
xnor UO_277 (O_277,N_8278,N_8722);
nand UO_278 (O_278,N_9327,N_9872);
nand UO_279 (O_279,N_9608,N_9801);
nand UO_280 (O_280,N_9868,N_8164);
xnor UO_281 (O_281,N_8941,N_9181);
nand UO_282 (O_282,N_8768,N_9888);
xnor UO_283 (O_283,N_8637,N_8377);
nand UO_284 (O_284,N_8795,N_8860);
or UO_285 (O_285,N_9525,N_9103);
and UO_286 (O_286,N_9020,N_9768);
nor UO_287 (O_287,N_8113,N_9616);
and UO_288 (O_288,N_8305,N_9648);
and UO_289 (O_289,N_8692,N_9294);
or UO_290 (O_290,N_9848,N_9764);
and UO_291 (O_291,N_9399,N_8065);
or UO_292 (O_292,N_9330,N_9249);
nor UO_293 (O_293,N_8822,N_9577);
nor UO_294 (O_294,N_9689,N_9052);
nor UO_295 (O_295,N_9045,N_8899);
or UO_296 (O_296,N_8235,N_9665);
nand UO_297 (O_297,N_8983,N_8561);
xor UO_298 (O_298,N_8602,N_8282);
xor UO_299 (O_299,N_9384,N_9533);
xnor UO_300 (O_300,N_9242,N_8483);
nor UO_301 (O_301,N_8347,N_9149);
nand UO_302 (O_302,N_9278,N_8818);
nor UO_303 (O_303,N_9755,N_9041);
xor UO_304 (O_304,N_8114,N_9777);
or UO_305 (O_305,N_9534,N_8424);
xor UO_306 (O_306,N_8480,N_8261);
xor UO_307 (O_307,N_8867,N_8671);
nor UO_308 (O_308,N_8587,N_8437);
nand UO_309 (O_309,N_9034,N_9815);
and UO_310 (O_310,N_9106,N_8272);
and UO_311 (O_311,N_9632,N_8848);
nor UO_312 (O_312,N_8013,N_8966);
xnor UO_313 (O_313,N_9289,N_8553);
or UO_314 (O_314,N_9021,N_9305);
nand UO_315 (O_315,N_9865,N_8868);
nor UO_316 (O_316,N_8429,N_8462);
or UO_317 (O_317,N_8402,N_9869);
xor UO_318 (O_318,N_8029,N_9705);
nor UO_319 (O_319,N_9978,N_9120);
and UO_320 (O_320,N_8457,N_9229);
nor UO_321 (O_321,N_9368,N_9579);
xnor UO_322 (O_322,N_8947,N_8329);
nand UO_323 (O_323,N_8311,N_8470);
nor UO_324 (O_324,N_8840,N_8967);
nand UO_325 (O_325,N_8981,N_8863);
nand UO_326 (O_326,N_8693,N_9440);
nor UO_327 (O_327,N_8805,N_8034);
or UO_328 (O_328,N_8396,N_8385);
or UO_329 (O_329,N_9316,N_8746);
and UO_330 (O_330,N_8950,N_8439);
nor UO_331 (O_331,N_9728,N_9780);
nor UO_332 (O_332,N_9508,N_9148);
nor UO_333 (O_333,N_8562,N_9400);
xnor UO_334 (O_334,N_9735,N_8806);
nor UO_335 (O_335,N_9449,N_8925);
nor UO_336 (O_336,N_8606,N_8233);
xor UO_337 (O_337,N_8729,N_9285);
or UO_338 (O_338,N_8609,N_9200);
xnor UO_339 (O_339,N_8870,N_8128);
xor UO_340 (O_340,N_9439,N_9940);
nor UO_341 (O_341,N_8582,N_8836);
xor UO_342 (O_342,N_9904,N_8526);
or UO_343 (O_343,N_9359,N_8964);
nor UO_344 (O_344,N_9243,N_9392);
nor UO_345 (O_345,N_8799,N_8893);
and UO_346 (O_346,N_8302,N_8741);
xor UO_347 (O_347,N_9998,N_8356);
and UO_348 (O_348,N_9520,N_9678);
nand UO_349 (O_349,N_8714,N_9398);
nor UO_350 (O_350,N_8767,N_8064);
and UO_351 (O_351,N_8686,N_8306);
nand UO_352 (O_352,N_8395,N_9668);
nand UO_353 (O_353,N_8324,N_9526);
or UO_354 (O_354,N_8134,N_9474);
and UO_355 (O_355,N_9421,N_9167);
nor UO_356 (O_356,N_9790,N_8828);
xor UO_357 (O_357,N_8294,N_9881);
nor UO_358 (O_358,N_8430,N_8475);
and UO_359 (O_359,N_9946,N_8712);
nor UO_360 (O_360,N_9649,N_9580);
nand UO_361 (O_361,N_9929,N_8523);
nor UO_362 (O_362,N_8044,N_9490);
xnor UO_363 (O_363,N_8364,N_8559);
and UO_364 (O_364,N_9342,N_8597);
nand UO_365 (O_365,N_9914,N_9516);
or UO_366 (O_366,N_9475,N_8332);
xor UO_367 (O_367,N_8055,N_8459);
nor UO_368 (O_368,N_9255,N_9044);
nor UO_369 (O_369,N_8842,N_8958);
nor UO_370 (O_370,N_9447,N_8121);
and UO_371 (O_371,N_8788,N_8668);
xnor UO_372 (O_372,N_9604,N_8419);
xor UO_373 (O_373,N_9151,N_9854);
nand UO_374 (O_374,N_8677,N_9228);
xor UO_375 (O_375,N_9038,N_8147);
nand UO_376 (O_376,N_8268,N_8401);
or UO_377 (O_377,N_9884,N_8037);
nor UO_378 (O_378,N_9213,N_8054);
or UO_379 (O_379,N_8718,N_9468);
nand UO_380 (O_380,N_8493,N_9394);
or UO_381 (O_381,N_9152,N_8415);
or UO_382 (O_382,N_8253,N_8945);
nand UO_383 (O_383,N_8145,N_9991);
nand UO_384 (O_384,N_9205,N_9879);
or UO_385 (O_385,N_9051,N_8197);
xor UO_386 (O_386,N_8176,N_8160);
and UO_387 (O_387,N_8408,N_8264);
nor UO_388 (O_388,N_9091,N_9892);
nor UO_389 (O_389,N_9351,N_9866);
nand UO_390 (O_390,N_9329,N_9105);
xnor UO_391 (O_391,N_8896,N_9804);
nor UO_392 (O_392,N_8757,N_9663);
xnor UO_393 (O_393,N_9776,N_9727);
or UO_394 (O_394,N_8497,N_9675);
nand UO_395 (O_395,N_9111,N_8218);
nor UO_396 (O_396,N_9131,N_8291);
or UO_397 (O_397,N_8612,N_8949);
nand UO_398 (O_398,N_9976,N_9611);
xnor UO_399 (O_399,N_8450,N_8194);
or UO_400 (O_400,N_9543,N_8972);
and UO_401 (O_401,N_9758,N_9182);
nor UO_402 (O_402,N_9999,N_9539);
xnor UO_403 (O_403,N_9144,N_9197);
and UO_404 (O_404,N_8773,N_8691);
nand UO_405 (O_405,N_9666,N_8809);
and UO_406 (O_406,N_8999,N_8556);
nor UO_407 (O_407,N_9158,N_8702);
and UO_408 (O_408,N_8533,N_8555);
or UO_409 (O_409,N_9352,N_9831);
or UO_410 (O_410,N_9123,N_9387);
or UO_411 (O_411,N_9443,N_8624);
or UO_412 (O_412,N_8607,N_8012);
nand UO_413 (O_413,N_9063,N_8736);
nor UO_414 (O_414,N_8855,N_9833);
nand UO_415 (O_415,N_8340,N_9937);
or UO_416 (O_416,N_9254,N_8733);
nand UO_417 (O_417,N_8454,N_9610);
xnor UO_418 (O_418,N_8708,N_9896);
nand UO_419 (O_419,N_8472,N_8622);
or UO_420 (O_420,N_8777,N_8230);
xnor UO_421 (O_421,N_8979,N_8975);
xor UO_422 (O_422,N_8953,N_8723);
nor UO_423 (O_423,N_9830,N_8214);
xor UO_424 (O_424,N_8120,N_8094);
and UO_425 (O_425,N_8815,N_8418);
xor UO_426 (O_426,N_8041,N_9299);
xnor UO_427 (O_427,N_8634,N_8521);
and UO_428 (O_428,N_9214,N_8886);
or UO_429 (O_429,N_9227,N_8367);
and UO_430 (O_430,N_9488,N_9655);
xnor UO_431 (O_431,N_8456,N_8962);
and UO_432 (O_432,N_9893,N_8406);
nand UO_433 (O_433,N_8397,N_8883);
nand UO_434 (O_434,N_8409,N_8984);
nand UO_435 (O_435,N_9498,N_9731);
xor UO_436 (O_436,N_8769,N_9980);
xor UO_437 (O_437,N_9709,N_8915);
nand UO_438 (O_438,N_9951,N_9767);
nor UO_439 (O_439,N_8357,N_9036);
or UO_440 (O_440,N_9934,N_9301);
and UO_441 (O_441,N_9964,N_9258);
and UO_442 (O_442,N_8572,N_9199);
xnor UO_443 (O_443,N_8750,N_8099);
nor UO_444 (O_444,N_9614,N_8948);
or UO_445 (O_445,N_9005,N_9538);
or UO_446 (O_446,N_8786,N_8124);
xnor UO_447 (O_447,N_9340,N_8060);
or UO_448 (O_448,N_9628,N_9198);
and UO_449 (O_449,N_8998,N_9944);
nand UO_450 (O_450,N_8073,N_8670);
nor UO_451 (O_451,N_9799,N_9186);
and UO_452 (O_452,N_9647,N_8823);
and UO_453 (O_453,N_9811,N_8227);
nand UO_454 (O_454,N_9313,N_8241);
or UO_455 (O_455,N_8871,N_9511);
nand UO_456 (O_456,N_8980,N_8003);
and UO_457 (O_457,N_9905,N_9960);
or UO_458 (O_458,N_9000,N_8473);
or UO_459 (O_459,N_9771,N_8086);
and UO_460 (O_460,N_9493,N_9850);
nand UO_461 (O_461,N_9948,N_9563);
nand UO_462 (O_462,N_8731,N_8392);
nand UO_463 (O_463,N_9503,N_8453);
and UO_464 (O_464,N_9347,N_8939);
nand UO_465 (O_465,N_8839,N_8115);
or UO_466 (O_466,N_9828,N_8930);
and UO_467 (O_467,N_8441,N_8122);
or UO_468 (O_468,N_9478,N_8327);
nand UO_469 (O_469,N_8229,N_9296);
nand UO_470 (O_470,N_8277,N_8970);
and UO_471 (O_471,N_9407,N_9876);
nand UO_472 (O_472,N_9683,N_9795);
or UO_473 (O_473,N_9471,N_9757);
or UO_474 (O_474,N_9080,N_8477);
and UO_475 (O_475,N_9992,N_8499);
nand UO_476 (O_476,N_8386,N_9117);
xnor UO_477 (O_477,N_9231,N_9711);
or UO_478 (O_478,N_8100,N_9550);
nor UO_479 (O_479,N_8906,N_8820);
and UO_480 (O_480,N_9997,N_9308);
and UO_481 (O_481,N_9092,N_8889);
and UO_482 (O_482,N_9006,N_8759);
xnor UO_483 (O_483,N_9522,N_8541);
and UO_484 (O_484,N_9494,N_8172);
nand UO_485 (O_485,N_9410,N_8661);
nor UO_486 (O_486,N_9566,N_9716);
and UO_487 (O_487,N_8240,N_8894);
and UO_488 (O_488,N_8022,N_9714);
nand UO_489 (O_489,N_8266,N_8365);
nor UO_490 (O_490,N_9267,N_8236);
xnor UO_491 (O_491,N_8053,N_8564);
xor UO_492 (O_492,N_9590,N_9295);
xor UO_493 (O_493,N_8267,N_9456);
nand UO_494 (O_494,N_9979,N_9097);
or UO_495 (O_495,N_9661,N_9222);
nor UO_496 (O_496,N_9450,N_9163);
and UO_497 (O_497,N_8760,N_8678);
and UO_498 (O_498,N_9024,N_8976);
nand UO_499 (O_499,N_9486,N_9853);
nand UO_500 (O_500,N_8566,N_9926);
nand UO_501 (O_501,N_9560,N_9843);
and UO_502 (O_502,N_8659,N_8704);
nand UO_503 (O_503,N_8961,N_9047);
and UO_504 (O_504,N_9921,N_8756);
nor UO_505 (O_505,N_8006,N_9098);
nor UO_506 (O_506,N_8690,N_8024);
and UO_507 (O_507,N_8501,N_9861);
and UO_508 (O_508,N_8248,N_9568);
xor UO_509 (O_509,N_8588,N_9004);
and UO_510 (O_510,N_8466,N_8590);
or UO_511 (O_511,N_9142,N_9309);
or UO_512 (O_512,N_9756,N_8352);
and UO_513 (O_513,N_9851,N_9202);
or UO_514 (O_514,N_9993,N_9913);
nand UO_515 (O_515,N_8909,N_8563);
nand UO_516 (O_516,N_8518,N_9633);
and UO_517 (O_517,N_8383,N_9670);
nand UO_518 (O_518,N_8800,N_9969);
nand UO_519 (O_519,N_9127,N_8701);
nand UO_520 (O_520,N_9483,N_9081);
nand UO_521 (O_521,N_8994,N_9397);
or UO_522 (O_522,N_8201,N_8184);
xnor UO_523 (O_523,N_8110,N_8169);
and UO_524 (O_524,N_9586,N_9133);
and UO_525 (O_525,N_8583,N_9089);
nand UO_526 (O_526,N_8781,N_8857);
nand UO_527 (O_527,N_9537,N_9054);
or UO_528 (O_528,N_9248,N_9957);
nand UO_529 (O_529,N_9292,N_8919);
and UO_530 (O_530,N_8239,N_8969);
xnor UO_531 (O_531,N_8092,N_8174);
nand UO_532 (O_532,N_9691,N_9377);
or UO_533 (O_533,N_8579,N_8881);
nand UO_534 (O_534,N_8880,N_9906);
and UO_535 (O_535,N_8517,N_9066);
xnor UO_536 (O_536,N_8642,N_9235);
xnor UO_537 (O_537,N_9209,N_9595);
nand UO_538 (O_538,N_9224,N_8954);
nor UO_539 (O_539,N_9507,N_9920);
xnor UO_540 (O_540,N_8293,N_9693);
xor UO_541 (O_541,N_9356,N_8097);
nand UO_542 (O_542,N_9109,N_9497);
xor UO_543 (O_543,N_8794,N_8730);
or UO_544 (O_544,N_9753,N_9319);
and UO_545 (O_545,N_8765,N_8672);
nand UO_546 (O_546,N_9442,N_8243);
nor UO_547 (O_547,N_9680,N_9603);
or UO_548 (O_548,N_9064,N_9835);
nor UO_549 (O_549,N_8088,N_9578);
nor UO_550 (O_550,N_9250,N_9240);
nor UO_551 (O_551,N_9263,N_9293);
and UO_552 (O_552,N_8026,N_9972);
nor UO_553 (O_553,N_8202,N_8039);
or UO_554 (O_554,N_8226,N_8952);
and UO_555 (O_555,N_8371,N_8004);
nor UO_556 (O_556,N_9037,N_9409);
xor UO_557 (O_557,N_9588,N_9599);
and UO_558 (O_558,N_8738,N_9009);
or UO_559 (O_559,N_9644,N_8301);
nand UO_560 (O_560,N_8569,N_9761);
or UO_561 (O_561,N_8198,N_9268);
and UO_562 (O_562,N_8059,N_9619);
and UO_563 (O_563,N_8850,N_8208);
nor UO_564 (O_564,N_8399,N_8444);
nor UO_565 (O_565,N_9480,N_8505);
nor UO_566 (O_566,N_8613,N_8771);
xor UO_567 (O_567,N_8223,N_9637);
and UO_568 (O_568,N_8807,N_9110);
nor UO_569 (O_569,N_9077,N_9512);
nand UO_570 (O_570,N_8803,N_8071);
xnor UO_571 (O_571,N_8804,N_8220);
xnor UO_572 (O_572,N_8995,N_8487);
or UO_573 (O_573,N_9085,N_8335);
nand UO_574 (O_574,N_9043,N_9961);
nand UO_575 (O_575,N_8655,N_8042);
and UO_576 (O_576,N_9219,N_9007);
and UO_577 (O_577,N_9039,N_8152);
nand UO_578 (O_578,N_8856,N_8067);
and UO_579 (O_579,N_8133,N_8298);
or UO_580 (O_580,N_9987,N_8204);
nor UO_581 (O_581,N_8262,N_8000);
and UO_582 (O_582,N_8551,N_8215);
xnor UO_583 (O_583,N_8107,N_8942);
xor UO_584 (O_584,N_9265,N_8957);
and UO_585 (O_585,N_8968,N_8640);
nand UO_586 (O_586,N_8228,N_8978);
or UO_587 (O_587,N_8502,N_8269);
nor UO_588 (O_588,N_9371,N_8117);
nand UO_589 (O_589,N_9078,N_9455);
and UO_590 (O_590,N_9836,N_8063);
nor UO_591 (O_591,N_8685,N_9885);
xor UO_592 (O_592,N_8049,N_9291);
and UO_593 (O_593,N_8864,N_8433);
xnor UO_594 (O_594,N_9367,N_8816);
nand UO_595 (O_595,N_9277,N_8798);
nand UO_596 (O_596,N_8727,N_8190);
nor UO_597 (O_597,N_8657,N_8232);
and UO_598 (O_598,N_8827,N_8575);
and UO_599 (O_599,N_8096,N_9382);
nand UO_600 (O_600,N_9458,N_8884);
or UO_601 (O_601,N_9206,N_8862);
and UO_602 (O_602,N_9651,N_9918);
or UO_603 (O_603,N_9686,N_9779);
xor UO_604 (O_604,N_9662,N_9378);
and UO_605 (O_605,N_9332,N_9118);
nor UO_606 (O_606,N_8763,N_9215);
nor UO_607 (O_607,N_8861,N_8656);
nor UO_608 (O_608,N_8735,N_9871);
nand UO_609 (O_609,N_8132,N_9349);
and UO_610 (O_610,N_8035,N_9617);
and UO_611 (O_611,N_9890,N_9810);
nand UO_612 (O_612,N_9420,N_9360);
nand UO_613 (O_613,N_9489,N_9977);
xnor UO_614 (O_614,N_9808,N_9094);
nand UO_615 (O_615,N_9130,N_8178);
nor UO_616 (O_616,N_8581,N_8688);
or UO_617 (O_617,N_8407,N_8126);
nor UO_618 (O_618,N_9001,N_9827);
nand UO_619 (O_619,N_9132,N_8118);
xnor UO_620 (O_620,N_8304,N_8159);
nor UO_621 (O_621,N_8394,N_9069);
nand UO_622 (O_622,N_8933,N_9852);
and UO_623 (O_623,N_8747,N_8372);
nand UO_624 (O_624,N_9597,N_8956);
nand UO_625 (O_625,N_9470,N_9746);
and UO_626 (O_626,N_8057,N_9003);
nor UO_627 (O_627,N_8217,N_8784);
nor UO_628 (O_628,N_9639,N_8016);
xor UO_629 (O_629,N_8621,N_8330);
xnor UO_630 (O_630,N_9417,N_9984);
nor UO_631 (O_631,N_9762,N_9274);
and UO_632 (O_632,N_8314,N_8283);
and UO_633 (O_633,N_9770,N_8715);
nand UO_634 (O_634,N_9016,N_9466);
or UO_635 (O_635,N_9476,N_9883);
and UO_636 (O_636,N_9688,N_8263);
and UO_637 (O_637,N_9724,N_9284);
xor UO_638 (O_638,N_9814,N_8404);
and UO_639 (O_639,N_8751,N_9556);
xor UO_640 (O_640,N_9936,N_9251);
or UO_641 (O_641,N_9752,N_8851);
xor UO_642 (O_642,N_8125,N_9434);
and UO_643 (O_643,N_9310,N_9681);
nand UO_644 (O_644,N_8749,N_8510);
nand UO_645 (O_645,N_9093,N_8971);
or UO_646 (O_646,N_9138,N_8812);
xnor UO_647 (O_647,N_8726,N_8275);
or UO_648 (O_648,N_8008,N_8913);
nor UO_649 (O_649,N_8859,N_9822);
xnor UO_650 (O_650,N_9877,N_8252);
nand UO_651 (O_651,N_9849,N_9252);
or UO_652 (O_652,N_8257,N_8744);
xnor UO_653 (O_653,N_8762,N_9682);
nor UO_654 (O_654,N_9502,N_8412);
or UO_655 (O_655,N_9509,N_9540);
xor UO_656 (O_656,N_8601,N_8509);
and UO_657 (O_657,N_8102,N_8423);
nor UO_658 (O_658,N_9943,N_9196);
xnor UO_659 (O_659,N_8123,N_8687);
and UO_660 (O_660,N_8015,N_8858);
xnor UO_661 (O_661,N_8484,N_8905);
xor UO_662 (O_662,N_8144,N_8375);
nand UO_663 (O_663,N_9551,N_8615);
and UO_664 (O_664,N_9606,N_9839);
and UO_665 (O_665,N_9677,N_8349);
nor UO_666 (O_666,N_8500,N_9911);
or UO_667 (O_667,N_9259,N_8440);
nand UO_668 (O_668,N_8724,N_8669);
nand UO_669 (O_669,N_8150,N_8464);
or UO_670 (O_670,N_8928,N_8238);
xor UO_671 (O_671,N_9014,N_9414);
xnor UO_672 (O_672,N_9086,N_8119);
or UO_673 (O_673,N_9803,N_9460);
xnor UO_674 (O_674,N_9365,N_9624);
xnor UO_675 (O_675,N_8315,N_9751);
and UO_676 (O_676,N_8997,N_8920);
xor UO_677 (O_677,N_9938,N_8717);
nand UO_678 (O_678,N_9145,N_9923);
nand UO_679 (O_679,N_9897,N_8937);
nor UO_680 (O_680,N_8449,N_8916);
nor UO_681 (O_681,N_9759,N_9903);
or UO_682 (O_682,N_9572,N_8358);
and UO_683 (O_683,N_9233,N_9100);
nand UO_684 (O_684,N_8221,N_9124);
nor UO_685 (O_685,N_9379,N_8237);
nor UO_686 (O_686,N_9656,N_8540);
nor UO_687 (O_687,N_8420,N_9710);
nor UO_688 (O_688,N_9134,N_9950);
and UO_689 (O_689,N_9880,N_9404);
or UO_690 (O_690,N_8234,N_8991);
xor UO_691 (O_691,N_9195,N_8443);
nand UO_692 (O_692,N_8091,N_9664);
xor UO_693 (O_693,N_9739,N_8565);
or UO_694 (O_694,N_8333,N_8137);
and UO_695 (O_695,N_8516,N_9241);
and UO_696 (O_696,N_8775,N_8438);
and UO_697 (O_697,N_9113,N_9824);
xnor UO_698 (O_698,N_9841,N_8388);
or UO_699 (O_699,N_9331,N_9018);
or UO_700 (O_700,N_9864,N_9894);
xnor UO_701 (O_701,N_9137,N_9022);
nand UO_702 (O_702,N_8633,N_8284);
xnor UO_703 (O_703,N_9411,N_8752);
nand UO_704 (O_704,N_9575,N_8281);
nand UO_705 (O_705,N_8183,N_8782);
nand UO_706 (O_706,N_8192,N_8020);
or UO_707 (O_707,N_9116,N_8398);
and UO_708 (O_708,N_8531,N_9362);
xnor UO_709 (O_709,N_9541,N_9419);
xnor UO_710 (O_710,N_8050,N_9557);
and UO_711 (O_711,N_9873,N_9676);
nor UO_712 (O_712,N_8432,N_9908);
or UO_713 (O_713,N_8242,N_9669);
xnor UO_714 (O_714,N_8825,N_9825);
nand UO_715 (O_715,N_9721,N_9060);
xnor UO_716 (O_716,N_8474,N_9630);
nand UO_717 (O_717,N_8813,N_9125);
and UO_718 (O_718,N_9820,N_8625);
nand UO_719 (O_719,N_8826,N_8935);
nor UO_720 (O_720,N_9927,N_8421);
or UO_721 (O_721,N_8089,N_8700);
and UO_722 (O_722,N_9423,N_9919);
or UO_723 (O_723,N_9548,N_9909);
and UO_724 (O_724,N_9203,N_8811);
or UO_725 (O_725,N_9472,N_8985);
nor UO_726 (O_726,N_8568,N_8699);
and UO_727 (O_727,N_9444,N_9015);
nand UO_728 (O_728,N_8931,N_8721);
and UO_729 (O_729,N_8188,N_9366);
or UO_730 (O_730,N_9983,N_8265);
xnor UO_731 (O_731,N_9517,N_8478);
and UO_732 (O_732,N_9433,N_9335);
xor UO_733 (O_733,N_9549,N_8515);
and UO_734 (O_734,N_9612,N_8654);
nor UO_735 (O_735,N_9800,N_9942);
xnor UO_736 (O_736,N_8946,N_9569);
and UO_737 (O_737,N_9902,N_8720);
nand UO_738 (O_738,N_9640,N_8673);
xor UO_739 (O_739,N_8630,N_9280);
or UO_740 (O_740,N_9703,N_9952);
or UO_741 (O_741,N_8578,N_9788);
nor UO_742 (O_742,N_9386,N_8280);
nand UO_743 (O_743,N_8644,N_8982);
xnor UO_744 (O_744,N_9717,N_9191);
or UO_745 (O_745,N_9025,N_8684);
xnor UO_746 (O_746,N_8343,N_9925);
or UO_747 (O_747,N_8819,N_9019);
xnor UO_748 (O_748,N_8142,N_9271);
nor UO_749 (O_749,N_8326,N_9646);
xor UO_750 (O_750,N_8154,N_8271);
xor UO_751 (O_751,N_9505,N_9954);
or UO_752 (O_752,N_8703,N_8467);
xor UO_753 (O_753,N_9168,N_8023);
and UO_754 (O_754,N_8066,N_9817);
or UO_755 (O_755,N_9882,N_9266);
and UO_756 (O_756,N_8471,N_8748);
nand UO_757 (O_757,N_8544,N_8093);
nor UO_758 (O_758,N_9826,N_9554);
nor UO_759 (O_759,N_8514,N_9510);
nand UO_760 (O_760,N_9996,N_9325);
nand UO_761 (O_761,N_8705,N_8576);
nand UO_762 (O_762,N_9609,N_9707);
xor UO_763 (O_763,N_9627,N_8136);
xnor UO_764 (O_764,N_8027,N_9057);
nor UO_765 (O_765,N_8193,N_8921);
or UO_766 (O_766,N_9238,N_9958);
xnor UO_767 (O_767,N_9829,N_8513);
xor UO_768 (O_768,N_8010,N_9418);
nand UO_769 (O_769,N_9122,N_9422);
and UO_770 (O_770,N_9061,N_9729);
or UO_771 (O_771,N_8766,N_8829);
or UO_772 (O_772,N_8116,N_9201);
xor UO_773 (O_773,N_9553,N_8200);
and UO_774 (O_774,N_8310,N_8033);
or UO_775 (O_775,N_8927,N_8080);
xor UO_776 (O_776,N_9867,N_8038);
nand UO_777 (O_777,N_9155,N_8830);
xnor UO_778 (O_778,N_8146,N_8486);
or UO_779 (O_779,N_8739,N_8251);
xor UO_780 (O_780,N_9185,N_8646);
and UO_781 (O_781,N_8345,N_8210);
xnor UO_782 (O_782,N_9461,N_8645);
and UO_783 (O_783,N_9701,N_9802);
nor UO_784 (O_784,N_8990,N_9338);
and UO_785 (O_785,N_8849,N_9857);
nor UO_786 (O_786,N_9547,N_9598);
nand UO_787 (O_787,N_9532,N_8186);
nor UO_788 (O_788,N_8413,N_8161);
nor UO_789 (O_789,N_9129,N_9273);
or UO_790 (O_790,N_8213,N_9324);
nand UO_791 (O_791,N_9405,N_9791);
and UO_792 (O_792,N_8546,N_8918);
nor UO_793 (O_793,N_8595,N_9380);
nor UO_794 (O_794,N_8058,N_9641);
nand UO_795 (O_795,N_9518,N_8458);
nand UO_796 (O_796,N_9234,N_8955);
xor UO_797 (O_797,N_9654,N_8325);
nand UO_798 (O_798,N_9115,N_8079);
xnor UO_799 (O_799,N_8062,N_8488);
xor UO_800 (O_800,N_8570,N_9613);
or UO_801 (O_801,N_8084,N_8610);
or UO_802 (O_802,N_9956,N_8108);
xnor UO_803 (O_803,N_8934,N_8837);
or UO_804 (O_804,N_8025,N_9147);
or UO_805 (O_805,N_8865,N_9076);
nand UO_806 (O_806,N_9846,N_9153);
nor UO_807 (O_807,N_9797,N_8519);
and UO_808 (O_808,N_9179,N_9183);
xnor UO_809 (O_809,N_8206,N_8783);
nor UO_810 (O_810,N_9102,N_8231);
nor UO_811 (O_811,N_9805,N_8754);
nand UO_812 (O_812,N_8321,N_9438);
xnor UO_813 (O_813,N_9524,N_8666);
and UO_814 (O_814,N_9190,N_8491);
and UO_815 (O_815,N_8845,N_8182);
nand UO_816 (O_816,N_9529,N_9223);
and UO_817 (O_817,N_9530,N_9565);
and UO_818 (O_818,N_8389,N_9785);
nor UO_819 (O_819,N_8600,N_9521);
and UO_820 (O_820,N_9842,N_8817);
and UO_821 (O_821,N_9962,N_8648);
and UO_822 (O_822,N_8173,N_8529);
and UO_823 (O_823,N_9370,N_9341);
nor UO_824 (O_824,N_8987,N_8361);
and UO_825 (O_825,N_8130,N_8988);
or UO_826 (O_826,N_8014,N_8040);
and UO_827 (O_827,N_8599,N_9740);
xor UO_828 (O_828,N_8318,N_8141);
nand UO_829 (O_829,N_8507,N_8162);
nor UO_830 (O_830,N_9353,N_8580);
or UO_831 (O_831,N_9819,N_8447);
nand UO_832 (O_832,N_9722,N_9139);
and UO_833 (O_833,N_8342,N_9749);
nand UO_834 (O_834,N_9275,N_8629);
xor UO_835 (O_835,N_9975,N_8087);
and UO_836 (O_836,N_9160,N_9715);
nor UO_837 (O_837,N_8902,N_8460);
nor UO_838 (O_838,N_9253,N_9073);
nor UO_839 (O_839,N_8374,N_8338);
or UO_840 (O_840,N_9141,N_9013);
nand UO_841 (O_841,N_9159,N_8847);
xor UO_842 (O_842,N_8888,N_8129);
and UO_843 (O_843,N_8764,N_8504);
or UO_844 (O_844,N_9226,N_9859);
and UO_845 (O_845,N_9372,N_9781);
nor UO_846 (O_846,N_9501,N_8320);
and UO_847 (O_847,N_8854,N_8891);
and UO_848 (O_848,N_9966,N_8892);
xor UO_849 (O_849,N_9463,N_8426);
nor UO_850 (O_850,N_8574,N_8138);
or UO_851 (O_851,N_8696,N_8148);
xnor UO_852 (O_852,N_9898,N_9985);
xor UO_853 (O_853,N_8274,N_8370);
xnor UO_854 (O_854,N_9459,N_8653);
and UO_855 (O_855,N_9718,N_9364);
or UO_856 (O_856,N_9659,N_8943);
nand UO_857 (O_857,N_8743,N_9055);
and UO_858 (O_858,N_8307,N_9700);
nor UO_859 (O_859,N_9698,N_8259);
or UO_860 (O_860,N_8853,N_9582);
or UO_861 (O_861,N_8821,N_9696);
xor UO_862 (O_862,N_9011,N_9769);
xor UO_863 (O_863,N_9358,N_8878);
or UO_864 (O_864,N_9657,N_9736);
nor UO_865 (O_865,N_8270,N_9446);
and UO_866 (O_866,N_9070,N_8384);
nand UO_867 (O_867,N_9172,N_8143);
and UO_868 (O_868,N_9634,N_8489);
and UO_869 (O_869,N_8631,N_8879);
nand UO_870 (O_870,N_8660,N_9058);
and UO_871 (O_871,N_8882,N_9712);
nor UO_872 (O_872,N_8589,N_8427);
or UO_873 (O_873,N_9837,N_8662);
nand UO_874 (O_874,N_9981,N_8468);
nor UO_875 (O_875,N_8649,N_8276);
nor UO_876 (O_876,N_9723,N_8834);
and UO_877 (O_877,N_8728,N_8018);
and UO_878 (O_878,N_8965,N_9973);
nor UO_879 (O_879,N_8710,N_8936);
nand UO_880 (O_880,N_8001,N_9303);
or UO_881 (O_881,N_9763,N_9075);
and UO_882 (O_882,N_9096,N_9389);
and UO_883 (O_883,N_8914,N_8203);
and UO_884 (O_884,N_9361,N_9071);
and UO_885 (O_885,N_8403,N_9306);
or UO_886 (O_886,N_9874,N_9002);
and UO_887 (O_887,N_9945,N_8674);
nand UO_888 (O_888,N_9783,N_8111);
xor UO_889 (O_889,N_9184,N_9067);
nand UO_890 (O_890,N_9042,N_8011);
nor UO_891 (O_891,N_8611,N_8151);
and UO_892 (O_892,N_8877,N_8313);
nand UO_893 (O_893,N_8078,N_9504);
and UO_894 (O_894,N_8170,N_8547);
and UO_895 (O_895,N_8036,N_9282);
or UO_896 (O_896,N_8614,N_9891);
or UO_897 (O_897,N_8363,N_8411);
xor UO_898 (O_898,N_8391,N_8191);
nand UO_899 (O_899,N_8296,N_9949);
and UO_900 (O_900,N_8944,N_8417);
nor UO_901 (O_901,N_8498,N_8379);
nand UO_902 (O_902,N_8535,N_9126);
nand UO_903 (O_903,N_8490,N_9262);
nand UO_904 (O_904,N_8682,N_9297);
and UO_905 (O_905,N_9786,N_9907);
nor UO_906 (O_906,N_8056,N_8295);
nor UO_907 (O_907,N_9760,N_9796);
nand UO_908 (O_908,N_8604,N_9300);
nand UO_909 (O_909,N_8628,N_9895);
and UO_910 (O_910,N_9536,N_9615);
or UO_911 (O_911,N_8425,N_8761);
xor UO_912 (O_912,N_8495,N_8344);
nand UO_913 (O_913,N_9995,N_9143);
xor UO_914 (O_914,N_9901,N_8286);
or UO_915 (O_915,N_9339,N_8697);
nand UO_916 (O_916,N_8732,N_9823);
and UO_917 (O_917,N_9816,N_9415);
and UO_918 (O_918,N_9787,N_9166);
nand UO_919 (O_919,N_9959,N_9939);
nor UO_920 (O_920,N_9270,N_8503);
xnor UO_921 (O_921,N_8075,N_8289);
and UO_922 (O_922,N_8623,N_9432);
nor UO_923 (O_923,N_8831,N_8676);
nor UO_924 (O_924,N_8149,N_9452);
xor UO_925 (O_925,N_9695,N_9230);
nor UO_926 (O_926,N_8895,N_8254);
xor UO_927 (O_927,N_8694,N_9515);
nand UO_928 (O_928,N_9345,N_9269);
or UO_929 (O_929,N_8387,N_9135);
and UO_930 (O_930,N_9585,N_9374);
and UO_931 (O_931,N_9029,N_9626);
nand UO_932 (O_932,N_9090,N_8681);
xor UO_933 (O_933,N_9068,N_8047);
nand UO_934 (O_934,N_9281,N_9175);
and UO_935 (O_935,N_9860,N_9542);
nor UO_936 (O_936,N_9636,N_9552);
nand UO_937 (O_937,N_8127,N_8527);
xor UO_938 (O_938,N_9974,N_8205);
nor UO_939 (O_939,N_8090,N_9318);
xnor UO_940 (O_940,N_8897,N_9107);
and UO_941 (O_941,N_8165,N_9519);
xor UO_942 (O_942,N_9189,N_9887);
nor UO_943 (O_943,N_8336,N_8446);
or UO_944 (O_944,N_9794,N_9256);
and UO_945 (O_945,N_8522,N_8353);
nor UO_946 (O_946,N_8707,N_9261);
and UO_947 (O_947,N_9220,N_9396);
and UO_948 (O_948,N_9607,N_8528);
or UO_949 (O_949,N_8852,N_9858);
and UO_950 (O_950,N_8322,N_8776);
nand UO_951 (O_951,N_9307,N_9844);
and UO_952 (O_952,N_9059,N_8511);
xor UO_953 (O_953,N_8616,N_9453);
nor UO_954 (O_954,N_8683,N_9660);
nor UO_955 (O_955,N_9555,N_9074);
nor UO_956 (O_956,N_8992,N_8185);
nor UO_957 (O_957,N_8923,N_8290);
or UO_958 (O_958,N_9173,N_8222);
or UO_959 (O_959,N_9600,N_8926);
xnor UO_960 (O_960,N_8778,N_9333);
nor UO_961 (O_961,N_9673,N_8101);
xnor UO_962 (O_962,N_9622,N_9968);
nor UO_963 (O_963,N_8348,N_8400);
or UO_964 (O_964,N_9178,N_8506);
xor UO_965 (O_965,N_8617,N_8608);
nand UO_966 (O_966,N_8445,N_8596);
nor UO_967 (O_967,N_8887,N_9171);
or UO_968 (O_968,N_8245,N_9049);
nor UO_969 (O_969,N_9288,N_9487);
xnor UO_970 (O_970,N_9924,N_8932);
xnor UO_971 (O_971,N_8359,N_9642);
and UO_972 (O_972,N_9208,N_9376);
or UO_973 (O_973,N_8316,N_9623);
nor UO_974 (O_974,N_9730,N_9218);
nor UO_975 (O_975,N_8219,N_8328);
and UO_976 (O_976,N_9454,N_9856);
and UO_977 (O_977,N_9101,N_9193);
and UO_978 (O_978,N_9087,N_8843);
xnor UO_979 (O_979,N_8770,N_8410);
and UO_980 (O_980,N_8866,N_8802);
or UO_981 (O_981,N_9889,N_9930);
and UO_982 (O_982,N_8195,N_9982);
nand UO_983 (O_983,N_8199,N_9040);
xnor UO_984 (O_984,N_9232,N_8911);
nor UO_985 (O_985,N_8593,N_8740);
xnor UO_986 (O_986,N_8166,N_9750);
nor UO_987 (O_987,N_9638,N_8658);
nor UO_988 (O_988,N_8903,N_9412);
and UO_989 (O_989,N_8573,N_9169);
nor UO_990 (O_990,N_8103,N_9720);
or UO_991 (O_991,N_8139,N_9146);
nor UO_992 (O_992,N_9385,N_9840);
and UO_993 (O_993,N_8104,N_9713);
or UO_994 (O_994,N_9596,N_9451);
nor UO_995 (O_995,N_9970,N_8045);
xnor UO_996 (O_996,N_9350,N_9050);
and UO_997 (O_997,N_8074,N_8711);
nand UO_998 (O_998,N_8508,N_9283);
xnor UO_999 (O_999,N_8938,N_8156);
nor UO_1000 (O_1000,N_8498,N_8660);
and UO_1001 (O_1001,N_8700,N_8971);
nand UO_1002 (O_1002,N_9502,N_8815);
xor UO_1003 (O_1003,N_8351,N_8635);
and UO_1004 (O_1004,N_9649,N_8507);
nand UO_1005 (O_1005,N_8690,N_9140);
nor UO_1006 (O_1006,N_8235,N_8681);
or UO_1007 (O_1007,N_9698,N_8066);
xnor UO_1008 (O_1008,N_9951,N_8732);
and UO_1009 (O_1009,N_9294,N_9627);
or UO_1010 (O_1010,N_9244,N_8453);
and UO_1011 (O_1011,N_9387,N_9361);
nor UO_1012 (O_1012,N_9271,N_9728);
or UO_1013 (O_1013,N_8858,N_9129);
nand UO_1014 (O_1014,N_9015,N_9673);
nor UO_1015 (O_1015,N_8243,N_8525);
and UO_1016 (O_1016,N_9201,N_8998);
xnor UO_1017 (O_1017,N_9290,N_8739);
and UO_1018 (O_1018,N_9514,N_8100);
or UO_1019 (O_1019,N_9640,N_9079);
and UO_1020 (O_1020,N_9090,N_8169);
nor UO_1021 (O_1021,N_9914,N_8915);
nor UO_1022 (O_1022,N_8597,N_8311);
and UO_1023 (O_1023,N_8529,N_9730);
nor UO_1024 (O_1024,N_9592,N_8992);
xor UO_1025 (O_1025,N_9182,N_9320);
nor UO_1026 (O_1026,N_8361,N_9057);
or UO_1027 (O_1027,N_8236,N_8856);
xor UO_1028 (O_1028,N_8223,N_8449);
and UO_1029 (O_1029,N_8373,N_9171);
nor UO_1030 (O_1030,N_8950,N_8334);
or UO_1031 (O_1031,N_9022,N_9953);
nand UO_1032 (O_1032,N_9822,N_9904);
nand UO_1033 (O_1033,N_9271,N_8760);
nor UO_1034 (O_1034,N_9960,N_9411);
nor UO_1035 (O_1035,N_9667,N_8842);
and UO_1036 (O_1036,N_9747,N_8892);
xnor UO_1037 (O_1037,N_8132,N_8922);
and UO_1038 (O_1038,N_8472,N_9093);
nand UO_1039 (O_1039,N_9332,N_8678);
and UO_1040 (O_1040,N_8214,N_9723);
and UO_1041 (O_1041,N_8109,N_8613);
or UO_1042 (O_1042,N_9466,N_8001);
and UO_1043 (O_1043,N_9245,N_8094);
nor UO_1044 (O_1044,N_8094,N_8086);
and UO_1045 (O_1045,N_9135,N_9558);
and UO_1046 (O_1046,N_8900,N_9125);
nand UO_1047 (O_1047,N_8636,N_9741);
xor UO_1048 (O_1048,N_9766,N_9987);
or UO_1049 (O_1049,N_8787,N_9162);
and UO_1050 (O_1050,N_9151,N_9399);
nor UO_1051 (O_1051,N_8826,N_9334);
nor UO_1052 (O_1052,N_9428,N_8843);
nor UO_1053 (O_1053,N_8930,N_8709);
xnor UO_1054 (O_1054,N_8567,N_9483);
xor UO_1055 (O_1055,N_9929,N_9522);
xnor UO_1056 (O_1056,N_8349,N_9462);
nand UO_1057 (O_1057,N_9821,N_8640);
xnor UO_1058 (O_1058,N_8747,N_8687);
or UO_1059 (O_1059,N_9487,N_8303);
nor UO_1060 (O_1060,N_8988,N_9913);
nor UO_1061 (O_1061,N_9310,N_9242);
nor UO_1062 (O_1062,N_9810,N_9134);
nor UO_1063 (O_1063,N_8946,N_8320);
nand UO_1064 (O_1064,N_8948,N_9536);
nor UO_1065 (O_1065,N_8610,N_9393);
xnor UO_1066 (O_1066,N_9117,N_8645);
xor UO_1067 (O_1067,N_9698,N_8129);
xnor UO_1068 (O_1068,N_8981,N_8709);
nand UO_1069 (O_1069,N_8177,N_8363);
nor UO_1070 (O_1070,N_8856,N_9151);
or UO_1071 (O_1071,N_8159,N_9328);
nand UO_1072 (O_1072,N_8968,N_8090);
or UO_1073 (O_1073,N_9982,N_9943);
nor UO_1074 (O_1074,N_8065,N_9484);
nor UO_1075 (O_1075,N_9037,N_8490);
xor UO_1076 (O_1076,N_8541,N_8993);
xnor UO_1077 (O_1077,N_8770,N_8182);
nor UO_1078 (O_1078,N_9832,N_8084);
or UO_1079 (O_1079,N_9060,N_9001);
xnor UO_1080 (O_1080,N_8836,N_9179);
nand UO_1081 (O_1081,N_8175,N_8064);
or UO_1082 (O_1082,N_8595,N_8889);
nor UO_1083 (O_1083,N_9792,N_9213);
or UO_1084 (O_1084,N_9197,N_9036);
xnor UO_1085 (O_1085,N_9077,N_9603);
and UO_1086 (O_1086,N_9401,N_9458);
nor UO_1087 (O_1087,N_8387,N_9394);
xnor UO_1088 (O_1088,N_9843,N_8010);
nor UO_1089 (O_1089,N_9315,N_9029);
nor UO_1090 (O_1090,N_8070,N_8014);
xor UO_1091 (O_1091,N_9236,N_8435);
and UO_1092 (O_1092,N_8168,N_9986);
and UO_1093 (O_1093,N_9232,N_9574);
xnor UO_1094 (O_1094,N_8087,N_9306);
nand UO_1095 (O_1095,N_9131,N_9630);
nor UO_1096 (O_1096,N_9202,N_9288);
nand UO_1097 (O_1097,N_9393,N_8403);
and UO_1098 (O_1098,N_9767,N_8831);
xor UO_1099 (O_1099,N_9413,N_9996);
nand UO_1100 (O_1100,N_8025,N_8476);
nand UO_1101 (O_1101,N_9029,N_8258);
or UO_1102 (O_1102,N_8766,N_8792);
nor UO_1103 (O_1103,N_8980,N_8506);
and UO_1104 (O_1104,N_9747,N_8850);
and UO_1105 (O_1105,N_8058,N_8696);
nor UO_1106 (O_1106,N_9565,N_9597);
nand UO_1107 (O_1107,N_8570,N_8967);
nor UO_1108 (O_1108,N_9561,N_9276);
nand UO_1109 (O_1109,N_9343,N_9029);
nor UO_1110 (O_1110,N_8087,N_8296);
nand UO_1111 (O_1111,N_8376,N_8038);
nor UO_1112 (O_1112,N_9350,N_9581);
nor UO_1113 (O_1113,N_8445,N_9829);
xnor UO_1114 (O_1114,N_9651,N_9357);
nor UO_1115 (O_1115,N_8041,N_8570);
xor UO_1116 (O_1116,N_8323,N_8583);
and UO_1117 (O_1117,N_9772,N_9200);
nor UO_1118 (O_1118,N_9664,N_9994);
xnor UO_1119 (O_1119,N_8625,N_9398);
nand UO_1120 (O_1120,N_8070,N_8954);
xor UO_1121 (O_1121,N_9188,N_9590);
and UO_1122 (O_1122,N_9970,N_8768);
xnor UO_1123 (O_1123,N_9175,N_9142);
nand UO_1124 (O_1124,N_9018,N_9886);
or UO_1125 (O_1125,N_9253,N_9854);
nand UO_1126 (O_1126,N_9437,N_9568);
nand UO_1127 (O_1127,N_9399,N_9020);
xor UO_1128 (O_1128,N_8891,N_9796);
nor UO_1129 (O_1129,N_8872,N_9633);
nor UO_1130 (O_1130,N_9551,N_9176);
or UO_1131 (O_1131,N_9281,N_8112);
nand UO_1132 (O_1132,N_8883,N_9053);
and UO_1133 (O_1133,N_9970,N_9865);
nand UO_1134 (O_1134,N_8282,N_9468);
xor UO_1135 (O_1135,N_9312,N_8473);
nor UO_1136 (O_1136,N_8154,N_9260);
nor UO_1137 (O_1137,N_9420,N_8529);
xor UO_1138 (O_1138,N_9209,N_8653);
or UO_1139 (O_1139,N_9511,N_9305);
nor UO_1140 (O_1140,N_9112,N_8670);
and UO_1141 (O_1141,N_9223,N_9788);
xor UO_1142 (O_1142,N_8467,N_9446);
xnor UO_1143 (O_1143,N_9379,N_8535);
or UO_1144 (O_1144,N_8855,N_8877);
or UO_1145 (O_1145,N_8335,N_8929);
nand UO_1146 (O_1146,N_9219,N_8575);
nand UO_1147 (O_1147,N_8805,N_8788);
or UO_1148 (O_1148,N_8307,N_8716);
nand UO_1149 (O_1149,N_9647,N_9151);
xnor UO_1150 (O_1150,N_8456,N_8159);
xnor UO_1151 (O_1151,N_9875,N_8932);
and UO_1152 (O_1152,N_8328,N_8390);
and UO_1153 (O_1153,N_8632,N_8225);
and UO_1154 (O_1154,N_9655,N_9815);
nand UO_1155 (O_1155,N_8241,N_8515);
xnor UO_1156 (O_1156,N_9709,N_8506);
nor UO_1157 (O_1157,N_9218,N_9032);
nor UO_1158 (O_1158,N_9381,N_8869);
or UO_1159 (O_1159,N_8867,N_9059);
xor UO_1160 (O_1160,N_8563,N_8614);
nor UO_1161 (O_1161,N_9799,N_8320);
nor UO_1162 (O_1162,N_8439,N_9154);
xnor UO_1163 (O_1163,N_9561,N_9793);
or UO_1164 (O_1164,N_9500,N_9598);
nor UO_1165 (O_1165,N_9839,N_9085);
nor UO_1166 (O_1166,N_9139,N_8780);
xor UO_1167 (O_1167,N_8224,N_9794);
or UO_1168 (O_1168,N_8378,N_9857);
and UO_1169 (O_1169,N_9447,N_9439);
xnor UO_1170 (O_1170,N_8805,N_8419);
nor UO_1171 (O_1171,N_8842,N_9257);
nor UO_1172 (O_1172,N_9179,N_8588);
nor UO_1173 (O_1173,N_8240,N_9583);
xor UO_1174 (O_1174,N_9129,N_9171);
nand UO_1175 (O_1175,N_8733,N_8238);
nor UO_1176 (O_1176,N_9909,N_9632);
nor UO_1177 (O_1177,N_8952,N_9673);
nor UO_1178 (O_1178,N_8263,N_8504);
nand UO_1179 (O_1179,N_9883,N_8252);
nand UO_1180 (O_1180,N_8274,N_9333);
nor UO_1181 (O_1181,N_8680,N_9332);
and UO_1182 (O_1182,N_9577,N_9824);
nand UO_1183 (O_1183,N_9828,N_8818);
nand UO_1184 (O_1184,N_8962,N_9794);
and UO_1185 (O_1185,N_9959,N_8654);
nand UO_1186 (O_1186,N_9765,N_9678);
or UO_1187 (O_1187,N_8173,N_9181);
nand UO_1188 (O_1188,N_9971,N_8505);
or UO_1189 (O_1189,N_9277,N_8440);
nor UO_1190 (O_1190,N_8378,N_8052);
nand UO_1191 (O_1191,N_9711,N_8393);
nor UO_1192 (O_1192,N_8392,N_8136);
and UO_1193 (O_1193,N_9029,N_9859);
xnor UO_1194 (O_1194,N_9930,N_8396);
xor UO_1195 (O_1195,N_8952,N_8783);
nand UO_1196 (O_1196,N_8950,N_8532);
xnor UO_1197 (O_1197,N_9479,N_8156);
or UO_1198 (O_1198,N_9840,N_8292);
nor UO_1199 (O_1199,N_9086,N_8106);
or UO_1200 (O_1200,N_8986,N_8831);
nor UO_1201 (O_1201,N_8241,N_8901);
or UO_1202 (O_1202,N_9497,N_9785);
and UO_1203 (O_1203,N_9236,N_8784);
and UO_1204 (O_1204,N_9018,N_9474);
nor UO_1205 (O_1205,N_8638,N_9672);
or UO_1206 (O_1206,N_8952,N_8154);
nand UO_1207 (O_1207,N_9568,N_9547);
xor UO_1208 (O_1208,N_9061,N_8431);
nor UO_1209 (O_1209,N_9954,N_9481);
or UO_1210 (O_1210,N_8581,N_9415);
nor UO_1211 (O_1211,N_9468,N_9654);
and UO_1212 (O_1212,N_8735,N_8669);
and UO_1213 (O_1213,N_8002,N_9002);
or UO_1214 (O_1214,N_8904,N_8374);
and UO_1215 (O_1215,N_9018,N_9896);
or UO_1216 (O_1216,N_8884,N_8967);
nor UO_1217 (O_1217,N_8583,N_8742);
nor UO_1218 (O_1218,N_9604,N_8858);
or UO_1219 (O_1219,N_8701,N_9254);
xor UO_1220 (O_1220,N_8354,N_9218);
or UO_1221 (O_1221,N_9411,N_8450);
nand UO_1222 (O_1222,N_8087,N_9284);
and UO_1223 (O_1223,N_8126,N_9959);
and UO_1224 (O_1224,N_8430,N_9466);
and UO_1225 (O_1225,N_8682,N_8164);
and UO_1226 (O_1226,N_9037,N_8872);
nand UO_1227 (O_1227,N_9174,N_9415);
nand UO_1228 (O_1228,N_9079,N_9462);
and UO_1229 (O_1229,N_8818,N_8075);
xor UO_1230 (O_1230,N_8059,N_8613);
and UO_1231 (O_1231,N_8434,N_8957);
and UO_1232 (O_1232,N_8667,N_8769);
nor UO_1233 (O_1233,N_8532,N_9179);
nand UO_1234 (O_1234,N_8868,N_8781);
nor UO_1235 (O_1235,N_8373,N_9978);
and UO_1236 (O_1236,N_8957,N_8107);
or UO_1237 (O_1237,N_8796,N_9359);
nand UO_1238 (O_1238,N_8207,N_9193);
or UO_1239 (O_1239,N_9621,N_9510);
or UO_1240 (O_1240,N_9562,N_8306);
and UO_1241 (O_1241,N_9408,N_9563);
nand UO_1242 (O_1242,N_8879,N_8567);
or UO_1243 (O_1243,N_9087,N_9146);
or UO_1244 (O_1244,N_9110,N_9698);
nor UO_1245 (O_1245,N_8838,N_9242);
or UO_1246 (O_1246,N_8460,N_8659);
nor UO_1247 (O_1247,N_9114,N_9344);
xnor UO_1248 (O_1248,N_9538,N_8007);
nor UO_1249 (O_1249,N_8771,N_9107);
xnor UO_1250 (O_1250,N_8269,N_8673);
nand UO_1251 (O_1251,N_8093,N_9309);
nand UO_1252 (O_1252,N_8181,N_9247);
nor UO_1253 (O_1253,N_9176,N_8388);
xnor UO_1254 (O_1254,N_9339,N_9223);
and UO_1255 (O_1255,N_8426,N_8943);
nand UO_1256 (O_1256,N_8336,N_9609);
nand UO_1257 (O_1257,N_8019,N_8780);
and UO_1258 (O_1258,N_9745,N_9826);
nor UO_1259 (O_1259,N_8057,N_9071);
or UO_1260 (O_1260,N_8668,N_9557);
xnor UO_1261 (O_1261,N_9558,N_8889);
or UO_1262 (O_1262,N_9878,N_8684);
nor UO_1263 (O_1263,N_9524,N_9038);
nand UO_1264 (O_1264,N_8937,N_9292);
xor UO_1265 (O_1265,N_8165,N_9614);
nand UO_1266 (O_1266,N_9956,N_9281);
xnor UO_1267 (O_1267,N_9511,N_8833);
or UO_1268 (O_1268,N_9313,N_9897);
xnor UO_1269 (O_1269,N_9589,N_8283);
nor UO_1270 (O_1270,N_8001,N_9357);
nand UO_1271 (O_1271,N_9734,N_8998);
and UO_1272 (O_1272,N_8952,N_9685);
nor UO_1273 (O_1273,N_9972,N_8046);
or UO_1274 (O_1274,N_9112,N_8838);
nor UO_1275 (O_1275,N_9287,N_9954);
nand UO_1276 (O_1276,N_9965,N_9258);
xnor UO_1277 (O_1277,N_8868,N_9059);
nor UO_1278 (O_1278,N_8851,N_8247);
and UO_1279 (O_1279,N_8405,N_9092);
or UO_1280 (O_1280,N_9180,N_9010);
and UO_1281 (O_1281,N_8906,N_8945);
xor UO_1282 (O_1282,N_8895,N_9397);
nor UO_1283 (O_1283,N_8874,N_8037);
nor UO_1284 (O_1284,N_8725,N_9416);
or UO_1285 (O_1285,N_9013,N_9825);
and UO_1286 (O_1286,N_8272,N_9173);
and UO_1287 (O_1287,N_9786,N_9113);
nand UO_1288 (O_1288,N_9122,N_9686);
or UO_1289 (O_1289,N_8674,N_8647);
xnor UO_1290 (O_1290,N_9531,N_9375);
or UO_1291 (O_1291,N_8661,N_9635);
or UO_1292 (O_1292,N_9790,N_8277);
nor UO_1293 (O_1293,N_8484,N_9646);
nor UO_1294 (O_1294,N_8660,N_9316);
xor UO_1295 (O_1295,N_8064,N_9395);
xor UO_1296 (O_1296,N_9413,N_8702);
or UO_1297 (O_1297,N_9404,N_9542);
and UO_1298 (O_1298,N_9681,N_9415);
or UO_1299 (O_1299,N_8386,N_9479);
nand UO_1300 (O_1300,N_8199,N_9227);
xnor UO_1301 (O_1301,N_9878,N_8671);
or UO_1302 (O_1302,N_8139,N_9067);
nor UO_1303 (O_1303,N_9211,N_9874);
and UO_1304 (O_1304,N_9277,N_8158);
nor UO_1305 (O_1305,N_9000,N_9693);
nor UO_1306 (O_1306,N_8729,N_8438);
and UO_1307 (O_1307,N_9050,N_8547);
nand UO_1308 (O_1308,N_9320,N_8764);
nor UO_1309 (O_1309,N_9637,N_9868);
nand UO_1310 (O_1310,N_8158,N_9869);
and UO_1311 (O_1311,N_9811,N_8361);
or UO_1312 (O_1312,N_8871,N_9707);
xor UO_1313 (O_1313,N_9007,N_9864);
nor UO_1314 (O_1314,N_8511,N_8964);
nor UO_1315 (O_1315,N_9877,N_8661);
and UO_1316 (O_1316,N_8642,N_9327);
or UO_1317 (O_1317,N_8424,N_9304);
or UO_1318 (O_1318,N_8715,N_8205);
and UO_1319 (O_1319,N_8356,N_8239);
xor UO_1320 (O_1320,N_8779,N_8117);
xnor UO_1321 (O_1321,N_8024,N_8537);
nor UO_1322 (O_1322,N_8265,N_8256);
nand UO_1323 (O_1323,N_9207,N_8124);
or UO_1324 (O_1324,N_8246,N_8916);
nand UO_1325 (O_1325,N_8882,N_9455);
nand UO_1326 (O_1326,N_9723,N_8308);
nand UO_1327 (O_1327,N_8192,N_8472);
nand UO_1328 (O_1328,N_9236,N_9075);
or UO_1329 (O_1329,N_9962,N_8883);
nand UO_1330 (O_1330,N_9726,N_8712);
or UO_1331 (O_1331,N_8255,N_8038);
xor UO_1332 (O_1332,N_9983,N_9196);
nor UO_1333 (O_1333,N_8468,N_8878);
xor UO_1334 (O_1334,N_9382,N_8464);
or UO_1335 (O_1335,N_9677,N_9848);
xnor UO_1336 (O_1336,N_8969,N_9531);
nor UO_1337 (O_1337,N_8064,N_9801);
nand UO_1338 (O_1338,N_8839,N_8252);
and UO_1339 (O_1339,N_9706,N_8211);
nor UO_1340 (O_1340,N_8151,N_8912);
xor UO_1341 (O_1341,N_8840,N_9859);
and UO_1342 (O_1342,N_9196,N_8086);
nor UO_1343 (O_1343,N_8241,N_8345);
nor UO_1344 (O_1344,N_9044,N_8333);
nor UO_1345 (O_1345,N_9179,N_8899);
nand UO_1346 (O_1346,N_9239,N_9279);
xor UO_1347 (O_1347,N_8694,N_8481);
nand UO_1348 (O_1348,N_9229,N_9569);
nand UO_1349 (O_1349,N_8510,N_9675);
or UO_1350 (O_1350,N_9430,N_9532);
nand UO_1351 (O_1351,N_9925,N_8690);
and UO_1352 (O_1352,N_9217,N_8790);
or UO_1353 (O_1353,N_8891,N_9109);
and UO_1354 (O_1354,N_8968,N_9815);
and UO_1355 (O_1355,N_8926,N_9932);
and UO_1356 (O_1356,N_9355,N_8573);
nand UO_1357 (O_1357,N_8487,N_9292);
nor UO_1358 (O_1358,N_8133,N_9820);
xnor UO_1359 (O_1359,N_8195,N_8349);
and UO_1360 (O_1360,N_9064,N_9480);
and UO_1361 (O_1361,N_8110,N_9981);
nand UO_1362 (O_1362,N_8066,N_8179);
nor UO_1363 (O_1363,N_8645,N_8927);
and UO_1364 (O_1364,N_9262,N_9100);
xnor UO_1365 (O_1365,N_8500,N_8058);
nand UO_1366 (O_1366,N_8643,N_9323);
and UO_1367 (O_1367,N_9137,N_8304);
nor UO_1368 (O_1368,N_8260,N_8387);
nand UO_1369 (O_1369,N_8237,N_9910);
nor UO_1370 (O_1370,N_9525,N_8962);
and UO_1371 (O_1371,N_9592,N_9756);
nor UO_1372 (O_1372,N_8800,N_8958);
nand UO_1373 (O_1373,N_9413,N_9388);
and UO_1374 (O_1374,N_8321,N_9138);
and UO_1375 (O_1375,N_8016,N_8796);
xor UO_1376 (O_1376,N_8602,N_8634);
nor UO_1377 (O_1377,N_9866,N_8263);
nand UO_1378 (O_1378,N_8596,N_8826);
or UO_1379 (O_1379,N_8057,N_9941);
or UO_1380 (O_1380,N_9896,N_9932);
xor UO_1381 (O_1381,N_8399,N_9558);
and UO_1382 (O_1382,N_9347,N_8036);
xnor UO_1383 (O_1383,N_9339,N_9462);
xor UO_1384 (O_1384,N_9060,N_8380);
or UO_1385 (O_1385,N_9414,N_8803);
and UO_1386 (O_1386,N_8196,N_9441);
or UO_1387 (O_1387,N_9446,N_8224);
xnor UO_1388 (O_1388,N_8381,N_8994);
nor UO_1389 (O_1389,N_9880,N_9199);
nand UO_1390 (O_1390,N_8048,N_8642);
and UO_1391 (O_1391,N_9115,N_8590);
and UO_1392 (O_1392,N_8738,N_8637);
xnor UO_1393 (O_1393,N_8919,N_8675);
nor UO_1394 (O_1394,N_9631,N_9270);
and UO_1395 (O_1395,N_9036,N_8585);
xor UO_1396 (O_1396,N_9140,N_9699);
nor UO_1397 (O_1397,N_8457,N_8831);
xnor UO_1398 (O_1398,N_8637,N_9024);
nand UO_1399 (O_1399,N_9428,N_8724);
xnor UO_1400 (O_1400,N_9004,N_9781);
nand UO_1401 (O_1401,N_8883,N_8703);
and UO_1402 (O_1402,N_8928,N_9963);
nand UO_1403 (O_1403,N_9095,N_9955);
or UO_1404 (O_1404,N_9084,N_9664);
nor UO_1405 (O_1405,N_9063,N_8443);
nor UO_1406 (O_1406,N_9357,N_9142);
nor UO_1407 (O_1407,N_9083,N_8156);
and UO_1408 (O_1408,N_8634,N_9278);
and UO_1409 (O_1409,N_8369,N_8747);
nor UO_1410 (O_1410,N_9835,N_9148);
or UO_1411 (O_1411,N_8719,N_9994);
nand UO_1412 (O_1412,N_8293,N_8053);
nand UO_1413 (O_1413,N_9679,N_9903);
nand UO_1414 (O_1414,N_8557,N_8241);
nor UO_1415 (O_1415,N_9450,N_8754);
nor UO_1416 (O_1416,N_8208,N_9311);
or UO_1417 (O_1417,N_9194,N_9679);
nor UO_1418 (O_1418,N_8221,N_9641);
nor UO_1419 (O_1419,N_8789,N_8016);
or UO_1420 (O_1420,N_8182,N_9194);
and UO_1421 (O_1421,N_8967,N_8864);
and UO_1422 (O_1422,N_8970,N_9780);
or UO_1423 (O_1423,N_8229,N_9099);
or UO_1424 (O_1424,N_9020,N_9889);
and UO_1425 (O_1425,N_8521,N_9771);
nor UO_1426 (O_1426,N_8963,N_8452);
nor UO_1427 (O_1427,N_8794,N_9979);
and UO_1428 (O_1428,N_9680,N_8937);
and UO_1429 (O_1429,N_8341,N_9567);
and UO_1430 (O_1430,N_8296,N_8340);
nor UO_1431 (O_1431,N_9293,N_8842);
xnor UO_1432 (O_1432,N_9695,N_9551);
nand UO_1433 (O_1433,N_9916,N_8043);
nor UO_1434 (O_1434,N_9316,N_9627);
or UO_1435 (O_1435,N_9426,N_9844);
nor UO_1436 (O_1436,N_8239,N_9919);
and UO_1437 (O_1437,N_9637,N_9951);
xnor UO_1438 (O_1438,N_9887,N_8484);
or UO_1439 (O_1439,N_9015,N_8729);
and UO_1440 (O_1440,N_8943,N_9780);
xor UO_1441 (O_1441,N_8275,N_8835);
nand UO_1442 (O_1442,N_9892,N_8567);
xnor UO_1443 (O_1443,N_9685,N_8970);
nand UO_1444 (O_1444,N_8106,N_9178);
nor UO_1445 (O_1445,N_8521,N_9629);
nor UO_1446 (O_1446,N_8236,N_8177);
and UO_1447 (O_1447,N_8080,N_9682);
or UO_1448 (O_1448,N_9416,N_9993);
nor UO_1449 (O_1449,N_8397,N_8045);
nor UO_1450 (O_1450,N_9790,N_9273);
xor UO_1451 (O_1451,N_8136,N_8040);
and UO_1452 (O_1452,N_9759,N_9074);
nand UO_1453 (O_1453,N_8453,N_8510);
nand UO_1454 (O_1454,N_8013,N_9704);
xor UO_1455 (O_1455,N_8926,N_8151);
xnor UO_1456 (O_1456,N_9164,N_9174);
and UO_1457 (O_1457,N_8091,N_9058);
nand UO_1458 (O_1458,N_8512,N_8015);
xnor UO_1459 (O_1459,N_9728,N_8065);
and UO_1460 (O_1460,N_8881,N_9484);
xnor UO_1461 (O_1461,N_9384,N_8205);
or UO_1462 (O_1462,N_9063,N_8540);
and UO_1463 (O_1463,N_9429,N_8572);
nor UO_1464 (O_1464,N_8122,N_8474);
and UO_1465 (O_1465,N_9428,N_8010);
or UO_1466 (O_1466,N_8420,N_9784);
or UO_1467 (O_1467,N_9411,N_8073);
or UO_1468 (O_1468,N_9428,N_8796);
nor UO_1469 (O_1469,N_8658,N_8597);
or UO_1470 (O_1470,N_8527,N_8864);
xnor UO_1471 (O_1471,N_8579,N_9178);
nor UO_1472 (O_1472,N_9706,N_8720);
xor UO_1473 (O_1473,N_9368,N_9492);
and UO_1474 (O_1474,N_8553,N_9295);
nor UO_1475 (O_1475,N_8671,N_8512);
nand UO_1476 (O_1476,N_9012,N_9382);
nand UO_1477 (O_1477,N_9150,N_9009);
nor UO_1478 (O_1478,N_9697,N_9155);
nand UO_1479 (O_1479,N_9832,N_9528);
nor UO_1480 (O_1480,N_9771,N_9511);
xor UO_1481 (O_1481,N_8720,N_9707);
xor UO_1482 (O_1482,N_9332,N_9874);
nand UO_1483 (O_1483,N_8326,N_9267);
nor UO_1484 (O_1484,N_9459,N_9881);
xnor UO_1485 (O_1485,N_8654,N_8505);
nor UO_1486 (O_1486,N_8583,N_8189);
xnor UO_1487 (O_1487,N_8326,N_8710);
nor UO_1488 (O_1488,N_9710,N_9920);
or UO_1489 (O_1489,N_8355,N_9099);
or UO_1490 (O_1490,N_8809,N_8989);
and UO_1491 (O_1491,N_8949,N_9511);
and UO_1492 (O_1492,N_8577,N_8127);
and UO_1493 (O_1493,N_9028,N_9367);
nor UO_1494 (O_1494,N_9650,N_8924);
xnor UO_1495 (O_1495,N_8588,N_9225);
nand UO_1496 (O_1496,N_8932,N_9608);
or UO_1497 (O_1497,N_8188,N_9465);
nor UO_1498 (O_1498,N_9206,N_9444);
nand UO_1499 (O_1499,N_8397,N_9690);
endmodule