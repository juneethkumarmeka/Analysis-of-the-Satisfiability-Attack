module basic_2000_20000_2500_40_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
or U0 (N_0,In_173,In_1961);
and U1 (N_1,In_831,In_851);
nand U2 (N_2,In_704,In_361);
xor U3 (N_3,In_339,In_1846);
nor U4 (N_4,In_1051,In_325);
nand U5 (N_5,In_1000,In_781);
or U6 (N_6,In_121,In_1399);
and U7 (N_7,In_433,In_242);
nor U8 (N_8,In_1512,In_64);
and U9 (N_9,In_749,In_837);
xnor U10 (N_10,In_1873,In_1105);
or U11 (N_11,In_1246,In_532);
xor U12 (N_12,In_149,In_683);
nor U13 (N_13,In_1902,In_356);
nand U14 (N_14,In_1714,In_1521);
xor U15 (N_15,In_559,In_510);
or U16 (N_16,In_1911,In_35);
nand U17 (N_17,In_1260,In_1491);
nand U18 (N_18,In_1631,In_595);
nor U19 (N_19,In_529,In_1710);
or U20 (N_20,In_99,In_1914);
or U21 (N_21,In_1906,In_4);
nor U22 (N_22,In_798,In_1212);
nand U23 (N_23,In_1062,In_1186);
nand U24 (N_24,In_232,In_377);
or U25 (N_25,In_1639,In_809);
xnor U26 (N_26,In_946,In_1275);
and U27 (N_27,In_353,In_179);
or U28 (N_28,In_626,In_1336);
nand U29 (N_29,In_1032,In_1099);
nand U30 (N_30,In_625,In_1865);
xnor U31 (N_31,In_1938,In_1030);
nor U32 (N_32,In_509,In_1249);
xor U33 (N_33,In_883,In_1872);
nand U34 (N_34,In_1479,In_1781);
nor U35 (N_35,In_1495,In_1580);
nand U36 (N_36,In_528,In_1951);
or U37 (N_37,In_981,In_867);
nand U38 (N_38,In_240,In_1169);
nor U39 (N_39,In_622,In_460);
nand U40 (N_40,In_941,In_1712);
nor U41 (N_41,In_1632,In_372);
nor U42 (N_42,In_222,In_296);
nor U43 (N_43,In_553,In_824);
xnor U44 (N_44,In_18,In_14);
or U45 (N_45,In_1451,In_212);
or U46 (N_46,In_1385,In_1531);
nor U47 (N_47,In_318,In_645);
or U48 (N_48,In_1729,In_1070);
and U49 (N_49,In_1998,In_37);
nand U50 (N_50,In_1538,In_1356);
or U51 (N_51,In_217,In_1615);
nor U52 (N_52,In_32,In_1421);
and U53 (N_53,In_1994,In_856);
nor U54 (N_54,In_635,In_1822);
nor U55 (N_55,In_524,In_264);
or U56 (N_56,In_1764,In_863);
xnor U57 (N_57,In_1463,In_1835);
and U58 (N_58,In_963,In_247);
and U59 (N_59,In_151,In_1840);
nand U60 (N_60,In_1403,In_210);
or U61 (N_61,In_333,In_1361);
nor U62 (N_62,In_711,In_55);
nor U63 (N_63,In_1815,In_1262);
xor U64 (N_64,In_571,In_381);
nor U65 (N_65,In_921,In_833);
or U66 (N_66,In_1346,In_1226);
and U67 (N_67,In_1210,In_1572);
or U68 (N_68,In_1554,In_1090);
nor U69 (N_69,In_1378,In_125);
nor U70 (N_70,In_458,In_1966);
nor U71 (N_71,In_1027,In_1599);
nor U72 (N_72,In_650,In_709);
nor U73 (N_73,In_1601,In_1214);
nand U74 (N_74,In_535,In_74);
nand U75 (N_75,In_623,In_1585);
or U76 (N_76,In_1168,In_1029);
nor U77 (N_77,In_314,In_829);
xor U78 (N_78,In_1808,In_580);
and U79 (N_79,In_1019,In_1871);
nor U80 (N_80,In_1583,In_873);
and U81 (N_81,In_1597,In_299);
xnor U82 (N_82,In_141,In_1221);
or U83 (N_83,In_1696,In_67);
xnor U84 (N_84,In_669,In_805);
and U85 (N_85,In_1081,In_640);
nand U86 (N_86,In_736,In_281);
or U87 (N_87,In_375,In_1579);
nor U88 (N_88,In_1775,In_1141);
nor U89 (N_89,In_665,In_1444);
xnor U90 (N_90,In_1928,In_194);
xnor U91 (N_91,In_551,In_1636);
nor U92 (N_92,In_329,In_1217);
and U93 (N_93,In_861,In_1205);
or U94 (N_94,In_391,In_1134);
or U95 (N_95,In_1676,In_1702);
or U96 (N_96,In_1423,In_60);
nor U97 (N_97,In_1153,In_814);
xor U98 (N_98,In_359,In_1500);
nor U99 (N_99,In_262,In_1983);
nand U100 (N_100,In_1135,In_1145);
and U101 (N_101,In_957,In_1115);
and U102 (N_102,In_1637,In_839);
or U103 (N_103,In_1279,In_1629);
or U104 (N_104,In_701,In_846);
and U105 (N_105,In_1420,In_762);
and U106 (N_106,In_1080,In_686);
or U107 (N_107,In_1836,In_163);
nand U108 (N_108,In_900,In_1082);
or U109 (N_109,In_287,In_1110);
and U110 (N_110,In_7,In_989);
nand U111 (N_111,In_1063,In_1722);
and U112 (N_112,In_922,In_1433);
and U113 (N_113,In_664,In_358);
xor U114 (N_114,In_1369,In_894);
nand U115 (N_115,In_1357,In_319);
nor U116 (N_116,In_305,In_1190);
xnor U117 (N_117,In_105,In_1593);
nor U118 (N_118,In_82,In_1119);
nor U119 (N_119,In_1731,In_673);
xnor U120 (N_120,In_211,In_1726);
or U121 (N_121,In_1026,In_1044);
and U122 (N_122,In_1040,In_1819);
and U123 (N_123,In_1703,In_504);
or U124 (N_124,In_769,In_279);
nand U125 (N_125,In_459,In_26);
or U126 (N_126,In_864,In_1046);
or U127 (N_127,In_1486,In_542);
xnor U128 (N_128,In_1351,In_1277);
or U129 (N_129,In_1203,In_1142);
xor U130 (N_130,In_1511,In_388);
or U131 (N_131,In_778,In_412);
or U132 (N_132,In_1238,In_271);
nor U133 (N_133,In_1170,In_1409);
xor U134 (N_134,In_298,In_1688);
or U135 (N_135,In_307,In_1912);
nand U136 (N_136,In_935,In_140);
or U137 (N_137,In_1236,In_1100);
and U138 (N_138,In_582,In_658);
xor U139 (N_139,In_1418,In_402);
and U140 (N_140,In_1364,In_1290);
and U141 (N_141,In_954,In_820);
and U142 (N_142,In_849,In_1899);
nor U143 (N_143,In_1448,In_1770);
or U144 (N_144,In_923,In_390);
or U145 (N_145,In_316,In_1680);
nand U146 (N_146,In_322,In_1942);
xnor U147 (N_147,In_1685,In_38);
nor U148 (N_148,In_1452,In_1758);
xor U149 (N_149,In_850,In_1033);
and U150 (N_150,In_251,In_1829);
nand U151 (N_151,In_676,In_1723);
nor U152 (N_152,In_291,In_1969);
and U153 (N_153,In_1450,In_1489);
or U154 (N_154,In_70,In_1031);
or U155 (N_155,In_1691,In_206);
nand U156 (N_156,In_1541,In_899);
or U157 (N_157,In_742,In_1889);
xnor U158 (N_158,In_1661,In_1167);
nor U159 (N_159,In_106,In_1592);
nand U160 (N_160,In_1627,In_1497);
nand U161 (N_161,In_1155,In_477);
and U162 (N_162,In_1015,In_832);
xor U163 (N_163,In_59,In_526);
nor U164 (N_164,In_1827,In_1474);
or U165 (N_165,In_245,In_810);
nand U166 (N_166,In_1784,In_784);
nand U167 (N_167,In_735,In_1122);
and U168 (N_168,In_1093,In_1657);
xnor U169 (N_169,In_1642,In_1774);
xnor U170 (N_170,In_872,In_1769);
or U171 (N_171,In_1481,In_920);
xnor U172 (N_172,In_1013,In_1708);
or U173 (N_173,In_200,In_780);
nor U174 (N_174,In_1201,In_540);
nand U175 (N_175,In_1483,In_1844);
and U176 (N_176,In_1406,In_789);
nor U177 (N_177,In_1305,In_636);
nand U178 (N_178,In_1633,In_1164);
xnor U179 (N_179,In_490,In_266);
or U180 (N_180,In_1957,In_1493);
nor U181 (N_181,In_1747,In_1704);
and U182 (N_182,In_1665,In_227);
nor U183 (N_183,In_1821,In_684);
and U184 (N_184,In_51,In_974);
and U185 (N_185,In_1268,In_878);
and U186 (N_186,In_572,In_1525);
and U187 (N_187,In_1446,In_848);
nand U188 (N_188,In_909,In_1069);
and U189 (N_189,In_594,In_1291);
xor U190 (N_190,In_143,In_1598);
xor U191 (N_191,In_1294,In_773);
or U192 (N_192,In_1408,In_1494);
xnor U193 (N_193,In_1659,In_1831);
and U194 (N_194,In_632,In_303);
nand U195 (N_195,In_85,In_139);
nor U196 (N_196,In_465,In_403);
or U197 (N_197,In_1499,In_277);
nand U198 (N_198,In_1057,In_515);
nand U199 (N_199,In_866,In_159);
and U200 (N_200,In_992,In_1092);
or U201 (N_201,In_1139,In_567);
and U202 (N_202,In_357,In_328);
nand U203 (N_203,In_569,In_570);
nand U204 (N_204,In_1751,In_1877);
and U205 (N_205,In_1207,In_603);
or U206 (N_206,In_1910,In_876);
and U207 (N_207,In_1503,In_836);
and U208 (N_208,In_343,In_1079);
nor U209 (N_209,In_1459,In_426);
xnor U210 (N_210,In_1458,In_463);
or U211 (N_211,In_1753,In_215);
or U212 (N_212,In_525,In_450);
nand U213 (N_213,In_1851,In_1725);
nand U214 (N_214,In_1152,In_892);
nand U215 (N_215,In_112,In_1533);
nor U216 (N_216,In_696,In_1068);
nand U217 (N_217,In_1881,In_50);
and U218 (N_218,In_156,In_1507);
or U219 (N_219,In_39,In_1131);
or U220 (N_220,In_1048,In_681);
or U221 (N_221,In_1176,In_1876);
nand U222 (N_222,In_1237,In_714);
nand U223 (N_223,In_1367,In_1358);
or U224 (N_224,In_1454,In_1682);
nand U225 (N_225,In_561,In_1549);
or U226 (N_226,In_1109,In_1485);
and U227 (N_227,In_1387,In_1341);
and U228 (N_228,In_611,In_313);
nor U229 (N_229,In_1677,In_1327);
or U230 (N_230,In_1529,In_233);
or U231 (N_231,In_998,In_425);
nor U232 (N_232,In_1300,In_693);
or U233 (N_233,In_823,In_1324);
and U234 (N_234,In_1978,In_1316);
nor U235 (N_235,In_1394,In_1028);
nor U236 (N_236,In_902,In_1380);
nand U237 (N_237,In_782,In_468);
nor U238 (N_238,In_1513,In_1247);
nor U239 (N_239,In_1923,In_1133);
xnor U240 (N_240,In_1687,In_950);
or U241 (N_241,In_1544,In_624);
and U242 (N_242,In_83,In_1552);
nor U243 (N_243,In_396,In_1165);
or U244 (N_244,In_285,In_1196);
xor U245 (N_245,In_104,In_1841);
xor U246 (N_246,In_560,In_1445);
or U247 (N_247,In_1065,In_1039);
xor U248 (N_248,In_1239,In_880);
xnor U249 (N_249,In_1299,In_1256);
and U250 (N_250,In_483,In_167);
nand U251 (N_251,In_1776,In_407);
or U252 (N_252,In_1075,In_89);
nor U253 (N_253,In_1606,In_534);
and U254 (N_254,In_1641,In_1879);
nor U255 (N_255,In_1405,In_578);
xnor U256 (N_256,In_444,In_968);
and U257 (N_257,In_1012,In_725);
and U258 (N_258,In_1900,In_746);
xor U259 (N_259,In_1177,In_142);
nor U260 (N_260,In_705,In_68);
and U261 (N_261,In_1522,In_565);
xnor U262 (N_262,In_991,In_48);
or U263 (N_263,In_96,In_928);
nand U264 (N_264,In_618,In_72);
nand U265 (N_265,In_807,In_218);
and U266 (N_266,In_1882,In_445);
nand U267 (N_267,In_269,In_203);
and U268 (N_268,In_420,In_480);
or U269 (N_269,In_1506,In_790);
nand U270 (N_270,In_1449,In_230);
nand U271 (N_271,In_721,In_654);
nand U272 (N_272,In_597,In_964);
xor U273 (N_273,In_1197,In_1958);
nand U274 (N_274,In_1679,In_1698);
xor U275 (N_275,In_710,In_1767);
xor U276 (N_276,In_1947,In_1401);
xnor U277 (N_277,In_1990,In_918);
nor U278 (N_278,In_691,In_1948);
xor U279 (N_279,In_180,In_349);
and U280 (N_280,In_1298,In_1359);
or U281 (N_281,In_1077,In_546);
nor U282 (N_282,In_1895,In_474);
xnor U283 (N_283,In_984,In_648);
and U284 (N_284,In_213,In_1820);
xor U285 (N_285,In_1681,In_1718);
xnor U286 (N_286,In_910,In_983);
and U287 (N_287,In_517,In_1407);
nor U288 (N_288,In_1860,In_838);
nor U289 (N_289,In_548,In_178);
xor U290 (N_290,In_1897,In_1339);
xnor U291 (N_291,In_1055,In_394);
or U292 (N_292,In_817,In_1997);
and U293 (N_293,In_17,In_129);
xnor U294 (N_294,In_614,In_589);
xor U295 (N_295,In_1830,In_1292);
and U296 (N_296,In_926,In_1008);
and U297 (N_297,In_531,In_1794);
and U298 (N_298,In_677,In_1622);
xor U299 (N_299,In_209,In_1996);
nand U300 (N_300,In_1453,In_429);
nand U301 (N_301,In_796,In_638);
nand U302 (N_302,In_1783,In_834);
or U303 (N_303,In_421,In_293);
or U304 (N_304,In_1002,In_1137);
or U305 (N_305,In_988,In_1575);
nor U306 (N_306,In_47,In_442);
and U307 (N_307,In_398,In_1746);
or U308 (N_308,In_1397,In_722);
and U309 (N_309,In_341,In_224);
xnor U310 (N_310,In_270,In_825);
xnor U311 (N_311,In_428,In_1813);
nand U312 (N_312,In_1654,In_12);
and U313 (N_313,In_155,In_1861);
or U314 (N_314,In_172,In_1664);
nand U315 (N_315,In_1315,In_13);
nor U316 (N_316,In_803,In_20);
nor U317 (N_317,In_42,In_1390);
and U318 (N_318,In_586,In_1950);
or U319 (N_319,In_1847,In_552);
or U320 (N_320,In_1288,In_799);
nand U321 (N_321,In_1832,In_793);
or U322 (N_322,In_389,In_868);
or U323 (N_323,In_1293,In_418);
nand U324 (N_324,In_727,In_310);
nor U325 (N_325,In_1054,In_280);
nand U326 (N_326,In_258,In_438);
nor U327 (N_327,In_1591,In_1590);
xnor U328 (N_328,In_1853,In_1671);
xnor U329 (N_329,In_1559,In_932);
nor U330 (N_330,In_122,In_1270);
nor U331 (N_331,In_1608,In_1733);
and U332 (N_332,In_730,In_81);
and U333 (N_333,In_901,In_1834);
nor U334 (N_334,In_1867,In_1626);
or U335 (N_335,In_166,In_808);
xor U336 (N_336,In_1353,In_397);
xnor U337 (N_337,In_996,In_1376);
xnor U338 (N_338,In_1414,In_446);
and U339 (N_339,In_724,In_1120);
xor U340 (N_340,In_1982,In_1945);
nor U341 (N_341,In_27,In_1245);
nand U342 (N_342,In_1673,In_1624);
nand U343 (N_343,In_133,In_462);
or U344 (N_344,In_1655,In_1297);
xor U345 (N_345,In_449,In_812);
and U346 (N_346,In_1595,In_1760);
nand U347 (N_347,In_308,In_95);
nor U348 (N_348,In_1925,In_130);
nand U349 (N_349,In_1344,In_347);
or U350 (N_350,In_666,In_327);
nand U351 (N_351,In_248,In_1265);
and U352 (N_352,In_1618,In_365);
nor U353 (N_353,In_1964,In_1104);
xnor U354 (N_354,In_404,In_417);
and U355 (N_355,In_1755,In_1548);
xor U356 (N_356,In_273,In_1041);
nand U357 (N_357,In_1918,In_40);
and U358 (N_358,In_62,In_1962);
and U359 (N_359,In_1287,In_489);
nor U360 (N_360,In_1927,In_1250);
xor U361 (N_361,In_1586,In_1993);
xor U362 (N_362,In_275,In_1514);
and U363 (N_363,In_1014,In_1219);
and U364 (N_364,In_1926,In_1697);
xor U365 (N_365,In_1372,In_862);
nand U366 (N_366,In_1007,In_813);
and U367 (N_367,In_1974,In_661);
or U368 (N_368,In_1335,In_936);
nand U369 (N_369,In_21,In_1222);
or U370 (N_370,In_1604,In_2);
xnor U371 (N_371,In_1866,In_660);
or U372 (N_372,In_620,In_877);
or U373 (N_373,In_1773,In_193);
nor U374 (N_374,In_1371,In_1232);
xor U375 (N_375,In_119,In_1443);
or U376 (N_376,In_1916,In_409);
nand U377 (N_377,In_84,In_228);
nand U378 (N_378,In_1535,In_708);
nand U379 (N_379,In_961,In_953);
nand U380 (N_380,In_1193,In_342);
xor U381 (N_381,In_126,In_678);
nor U382 (N_382,In_1643,In_858);
or U383 (N_383,In_1052,In_15);
xnor U384 (N_384,In_1343,In_1528);
and U385 (N_385,In_1934,In_56);
or U386 (N_386,In_905,In_1402);
and U387 (N_387,In_731,In_1436);
and U388 (N_388,In_717,In_786);
nand U389 (N_389,In_687,In_1884);
nand U390 (N_390,In_43,In_1505);
or U391 (N_391,In_304,In_1763);
nor U392 (N_392,In_1307,In_1715);
or U393 (N_393,In_1553,In_496);
nor U394 (N_394,In_758,In_630);
or U395 (N_395,In_1482,In_1523);
and U396 (N_396,In_1537,In_1323);
xor U397 (N_397,In_600,In_1972);
and U398 (N_398,In_370,In_405);
or U399 (N_399,In_754,In_103);
nor U400 (N_400,In_1352,In_36);
and U401 (N_401,In_410,In_1765);
nand U402 (N_402,In_1584,In_1053);
nor U403 (N_403,In_1243,In_1875);
and U404 (N_404,In_893,In_1709);
nand U405 (N_405,In_1384,In_874);
nand U406 (N_406,In_1816,In_744);
or U407 (N_407,In_484,In_469);
nand U408 (N_408,In_1652,In_1778);
nor U409 (N_409,In_1242,In_610);
nor U410 (N_410,In_760,In_117);
and U411 (N_411,In_1825,In_1106);
and U412 (N_412,In_290,In_338);
nor U413 (N_413,In_712,In_1588);
or U414 (N_414,In_1071,In_134);
nand U415 (N_415,In_1824,In_827);
or U416 (N_416,In_1883,In_1864);
nor U417 (N_417,In_30,In_1797);
xnor U418 (N_418,In_1125,In_1749);
xor U419 (N_419,In_234,In_1333);
nand U420 (N_420,In_334,In_1550);
or U421 (N_421,In_1609,In_355);
or U422 (N_422,In_1563,In_612);
or U423 (N_423,In_1915,In_1308);
or U424 (N_424,In_1060,In_1587);
nand U425 (N_425,In_1843,In_975);
nor U426 (N_426,In_498,In_1917);
xnor U427 (N_427,In_386,In_642);
or U428 (N_428,In_1461,In_1020);
nor U429 (N_429,In_1484,In_306);
nand U430 (N_430,In_860,In_383);
nand U431 (N_431,In_1258,In_886);
nand U432 (N_432,In_1752,In_958);
or U433 (N_433,In_1151,In_549);
xor U434 (N_434,In_1374,In_127);
and U435 (N_435,In_547,In_1231);
or U436 (N_436,In_649,In_564);
xnor U437 (N_437,In_401,In_1570);
and U438 (N_438,In_1094,In_544);
xor U439 (N_439,In_1025,In_205);
nand U440 (N_440,In_651,In_1762);
nor U441 (N_441,In_1744,In_1230);
nor U442 (N_442,In_584,In_1569);
nand U443 (N_443,In_763,In_1206);
nand U444 (N_444,In_414,In_256);
nor U445 (N_445,In_392,In_1811);
or U446 (N_446,In_1227,In_702);
nand U447 (N_447,In_1189,In_168);
or U448 (N_448,In_853,In_1072);
nand U449 (N_449,In_73,In_1546);
nand U450 (N_450,In_706,In_1276);
nand U451 (N_451,In_1112,In_186);
or U452 (N_452,In_1248,In_1561);
nand U453 (N_453,In_1382,In_1943);
nor U454 (N_454,In_1838,In_1415);
or U455 (N_455,In_447,In_146);
or U456 (N_456,In_777,In_236);
and U457 (N_457,In_573,In_440);
and U458 (N_458,In_1603,In_945);
or U459 (N_459,In_1140,In_1036);
or U460 (N_460,In_656,In_1362);
or U461 (N_461,In_1839,In_183);
nor U462 (N_462,In_801,In_1411);
nor U463 (N_463,In_1022,In_221);
and U464 (N_464,In_728,In_1909);
or U465 (N_465,In_639,In_1891);
nand U466 (N_466,In_362,In_1880);
xnor U467 (N_467,In_1617,In_1267);
nor U468 (N_468,In_1208,In_1024);
and U469 (N_469,In_1194,In_1863);
or U470 (N_470,In_1127,In_993);
nand U471 (N_471,In_225,In_393);
nand U472 (N_472,In_865,In_400);
xor U473 (N_473,In_967,In_972);
and U474 (N_474,In_896,In_175);
nand U475 (N_475,In_1396,In_602);
and U476 (N_476,In_1158,In_160);
nor U477 (N_477,In_145,In_123);
xnor U478 (N_478,In_1973,In_157);
and U479 (N_479,In_1318,In_330);
or U480 (N_480,In_1628,In_1332);
and U481 (N_481,In_1992,In_574);
nor U482 (N_482,In_238,In_520);
nand U483 (N_483,In_1178,In_1520);
and U484 (N_484,In_629,In_0);
or U485 (N_485,In_657,In_1234);
or U486 (N_486,In_1355,In_1791);
nand U487 (N_487,In_767,In_765);
or U488 (N_488,In_302,In_432);
and U489 (N_489,In_1707,In_1724);
nand U490 (N_490,In_680,In_757);
nor U491 (N_491,In_1391,In_1817);
nor U492 (N_492,In_1301,In_550);
nor U493 (N_493,In_1607,In_1255);
and U494 (N_494,In_5,In_1058);
or U495 (N_495,In_252,In_1929);
nand U496 (N_496,In_847,In_1809);
nor U497 (N_497,In_1430,In_1551);
or U498 (N_498,In_1672,In_1796);
or U499 (N_499,In_497,In_1101);
nor U500 (N_500,In_952,N_187);
xor U501 (N_501,In_933,N_314);
and U502 (N_502,N_123,In_1903);
xnor U503 (N_503,In_57,In_1955);
nand U504 (N_504,N_474,In_1904);
nor U505 (N_505,N_368,In_1042);
xnor U506 (N_506,In_276,N_181);
and U507 (N_507,In_406,N_433);
xnor U508 (N_508,N_155,N_1);
nor U509 (N_509,N_416,N_292);
xor U510 (N_510,In_1228,N_197);
xor U511 (N_511,N_403,N_279);
xnor U512 (N_512,In_1547,In_1793);
or U513 (N_513,N_193,In_616);
or U514 (N_514,N_378,N_216);
or U515 (N_515,In_1492,N_44);
xor U516 (N_516,N_158,In_1274);
xor U517 (N_517,In_1623,In_1229);
xor U518 (N_518,In_633,In_815);
nand U519 (N_519,N_432,In_885);
nor U520 (N_520,In_1759,In_162);
or U521 (N_521,N_497,In_1524);
or U522 (N_522,N_390,In_86);
or U523 (N_523,N_365,In_1473);
nor U524 (N_524,In_1566,In_1804);
nor U525 (N_525,In_1991,In_455);
and U526 (N_526,N_159,N_265);
and U527 (N_527,In_1913,N_95);
nor U528 (N_528,In_713,N_436);
nand U529 (N_529,N_163,In_1542);
nand U530 (N_530,In_1183,In_1630);
nand U531 (N_531,In_607,In_1768);
nand U532 (N_532,In_23,In_1750);
and U533 (N_533,In_1157,In_1419);
nor U534 (N_534,In_109,In_755);
or U535 (N_535,In_1066,In_268);
xnor U536 (N_536,N_325,N_201);
xnor U537 (N_537,In_1388,In_472);
nand U538 (N_538,In_1434,N_286);
xnor U539 (N_539,In_1577,In_503);
xnor U540 (N_540,In_1347,N_361);
xor U541 (N_541,In_818,In_1526);
or U542 (N_542,In_58,N_302);
nor U543 (N_543,In_1644,N_277);
xor U544 (N_544,N_349,N_412);
nor U545 (N_545,N_83,N_437);
xor U546 (N_546,In_539,In_617);
and U547 (N_547,In_1216,In_1837);
or U548 (N_548,In_364,N_414);
nand U549 (N_549,In_1565,N_241);
nand U550 (N_550,In_1108,N_63);
nor U551 (N_551,In_1517,In_1322);
nand U552 (N_552,In_1662,In_189);
and U553 (N_553,In_473,N_285);
or U554 (N_554,In_898,In_1215);
xnor U555 (N_555,In_1331,In_1313);
and U556 (N_556,N_162,In_24);
or U557 (N_557,N_221,In_1211);
xnor U558 (N_558,In_1967,In_1146);
nor U559 (N_559,N_269,In_1711);
nand U560 (N_560,In_776,N_25);
nor U561 (N_561,In_802,In_11);
nand U562 (N_562,N_199,In_1304);
nor U563 (N_563,In_897,N_256);
nor U564 (N_564,In_995,In_1354);
and U565 (N_565,N_202,In_697);
xor U566 (N_566,In_246,In_906);
and U567 (N_567,In_887,N_282);
xor U568 (N_568,In_1050,N_106);
and U569 (N_569,In_1124,In_185);
or U570 (N_570,N_224,In_1848);
or U571 (N_571,In_1375,N_463);
nor U572 (N_572,In_239,N_103);
and U573 (N_573,In_312,In_219);
nand U574 (N_574,In_502,N_270);
nor U575 (N_575,In_1818,In_634);
and U576 (N_576,N_179,In_828);
or U577 (N_577,In_326,In_387);
and U578 (N_578,In_135,In_1931);
nor U579 (N_579,In_747,N_172);
nand U580 (N_580,In_1690,N_262);
and U581 (N_581,N_406,In_108);
or U582 (N_582,In_1619,In_323);
and U583 (N_583,N_0,In_1545);
and U584 (N_584,N_465,In_659);
xor U585 (N_585,N_117,In_367);
nand U586 (N_586,N_453,In_184);
or U587 (N_587,In_137,In_1172);
xor U588 (N_588,N_105,In_1496);
xnor U589 (N_589,N_94,In_1191);
xnor U590 (N_590,N_315,In_1435);
nor U591 (N_591,N_442,In_250);
and U592 (N_592,In_260,N_109);
and U593 (N_593,N_407,In_519);
nor U594 (N_594,In_1325,In_487);
and U595 (N_595,In_694,In_715);
and U596 (N_596,N_88,N_276);
nor U597 (N_597,N_230,In_631);
and U598 (N_598,In_1428,In_1386);
nand U599 (N_599,N_419,In_1460);
or U600 (N_600,In_408,N_130);
or U601 (N_601,In_1422,In_1198);
nor U602 (N_602,In_1001,N_231);
or U603 (N_603,In_1612,N_29);
nand U604 (N_604,In_368,In_740);
or U605 (N_605,N_59,In_615);
or U606 (N_606,N_410,In_1845);
or U607 (N_607,In_1807,In_1648);
nand U608 (N_608,N_214,In_1264);
and U609 (N_609,In_152,N_13);
nor U610 (N_610,In_237,N_86);
nor U611 (N_611,In_33,N_447);
and U612 (N_612,N_188,In_336);
nor U613 (N_613,In_1225,In_1660);
nor U614 (N_614,N_135,N_430);
nand U615 (N_615,In_1432,In_692);
nand U616 (N_616,N_423,In_590);
and U617 (N_617,In_1302,In_456);
or U618 (N_618,N_184,N_72);
nand U619 (N_619,N_249,In_120);
xnor U620 (N_620,In_943,In_541);
xor U621 (N_621,N_62,In_320);
nand U622 (N_622,In_170,In_1314);
or U623 (N_623,In_682,In_344);
nor U624 (N_624,In_1534,In_679);
and U625 (N_625,N_321,In_1995);
and U626 (N_626,In_1653,N_154);
nor U627 (N_627,In_1498,In_1850);
and U628 (N_628,In_1894,N_69);
and U629 (N_629,In_1252,In_411);
nor U630 (N_630,In_911,In_1465);
or U631 (N_631,In_576,In_1317);
and U632 (N_632,In_1381,In_951);
and U633 (N_633,In_1266,N_283);
xnor U634 (N_634,In_53,In_1706);
xnor U635 (N_635,In_348,In_628);
nor U636 (N_636,In_745,In_1719);
nand U637 (N_637,N_186,In_966);
xor U638 (N_638,In_192,In_1976);
xor U639 (N_639,N_486,In_939);
xor U640 (N_640,N_76,In_66);
nor U641 (N_641,In_395,In_1209);
or U642 (N_642,In_819,In_598);
and U643 (N_643,In_985,In_1107);
nor U644 (N_644,In_948,N_26);
nor U645 (N_645,In_1855,In_28);
nand U646 (N_646,In_1087,N_48);
nor U647 (N_647,N_347,In_259);
nand U648 (N_648,In_1571,N_431);
or U649 (N_649,N_426,N_32);
and U650 (N_650,In_672,N_64);
nor U651 (N_651,In_1693,N_30);
xor U652 (N_652,In_1568,In_1023);
and U653 (N_653,In_415,In_521);
nand U654 (N_654,In_340,In_366);
nor U655 (N_655,In_999,In_556);
nor U656 (N_656,N_299,In_1102);
and U657 (N_657,N_458,In_774);
nand U658 (N_658,In_1321,In_543);
and U659 (N_659,N_492,In_695);
or U660 (N_660,In_1946,In_804);
xor U661 (N_661,N_456,In_195);
or U662 (N_662,In_566,In_1181);
and U663 (N_663,N_127,In_1431);
nand U664 (N_664,N_384,In_1999);
xnor U665 (N_665,N_359,In_102);
nor U666 (N_666,N_438,N_476);
or U667 (N_667,In_1932,In_331);
nand U668 (N_668,In_1812,N_268);
nand U669 (N_669,N_174,N_6);
or U670 (N_670,N_455,N_56);
or U671 (N_671,In_337,In_1471);
nor U672 (N_672,In_1003,In_1798);
nand U673 (N_673,In_1780,In_508);
and U674 (N_674,In_591,N_39);
nand U675 (N_675,N_337,In_1788);
xnor U676 (N_676,N_137,N_223);
and U677 (N_677,N_290,N_446);
and U678 (N_678,In_144,In_977);
and U679 (N_679,N_40,N_79);
xnor U680 (N_680,In_1620,In_741);
nand U681 (N_681,In_132,In_1732);
nor U682 (N_682,N_136,N_2);
and U683 (N_683,N_257,In_267);
xnor U684 (N_684,In_1779,In_1095);
nand U685 (N_685,N_121,N_112);
nor U686 (N_686,In_1869,N_493);
xor U687 (N_687,In_148,N_18);
nand U688 (N_688,N_78,N_24);
and U689 (N_689,In_98,In_1424);
xor U690 (N_690,N_251,In_1666);
nand U691 (N_691,N_254,In_1038);
nand U692 (N_692,N_93,In_1392);
and U693 (N_693,In_399,In_538);
xor U694 (N_694,In_879,In_1161);
and U695 (N_695,In_978,In_1173);
or U696 (N_696,In_1188,In_315);
nor U697 (N_697,In_970,In_855);
and U698 (N_698,In_1096,In_174);
or U699 (N_699,In_1663,In_435);
xor U700 (N_700,In_1166,In_1083);
or U701 (N_701,In_1117,In_147);
or U702 (N_702,N_483,In_500);
xor U703 (N_703,In_1536,In_522);
nand U704 (N_704,In_113,In_1147);
or U705 (N_705,In_1278,N_461);
xnor U706 (N_706,N_331,N_9);
nand U707 (N_707,In_1220,In_461);
and U708 (N_708,In_720,N_170);
nand U709 (N_709,In_822,In_1656);
nor U710 (N_710,In_707,N_20);
and U711 (N_711,In_716,N_351);
nand U712 (N_712,N_381,N_300);
or U713 (N_713,In_1555,In_1213);
nand U714 (N_714,N_97,N_487);
nor U715 (N_715,In_1074,N_387);
and U716 (N_716,N_28,In_1649);
xnor U717 (N_717,In_1389,In_791);
nor U718 (N_718,In_1005,In_1447);
xor U719 (N_719,In_1366,N_148);
nor U720 (N_720,In_1043,In_1814);
and U721 (N_721,N_211,In_380);
nand U722 (N_722,In_1162,In_1736);
nor U723 (N_723,N_494,In_1941);
nand U724 (N_724,N_98,N_77);
or U725 (N_725,In_568,In_1988);
or U726 (N_726,In_1892,In_1516);
and U727 (N_727,N_180,N_491);
nor U728 (N_728,In_606,In_1795);
nand U729 (N_729,In_138,In_424);
nor U730 (N_730,In_479,In_1097);
or U731 (N_731,N_468,In_1898);
xor U732 (N_732,In_374,In_903);
or U733 (N_733,In_826,N_449);
nand U734 (N_734,N_120,In_309);
or U735 (N_735,In_843,In_1734);
xnor U736 (N_736,In_1741,In_947);
xnor U737 (N_737,In_1118,In_1187);
and U738 (N_738,In_930,In_737);
nand U739 (N_739,In_482,In_1921);
or U740 (N_740,In_587,In_1692);
nand U741 (N_741,In_609,In_588);
xnor U742 (N_742,N_244,N_488);
and U743 (N_743,N_341,N_259);
xnor U744 (N_744,In_283,N_370);
and U745 (N_745,In_783,In_1613);
or U746 (N_746,N_176,N_369);
nand U747 (N_747,In_1800,N_288);
nand U748 (N_748,In_1295,In_1310);
or U749 (N_749,N_37,In_1088);
xnor U750 (N_750,In_1061,In_1530);
or U751 (N_751,In_772,In_949);
and U752 (N_752,In_1338,N_165);
nand U753 (N_753,In_1981,In_698);
nand U754 (N_754,N_82,N_247);
nand U755 (N_755,N_222,N_336);
or U756 (N_756,In_376,In_1416);
or U757 (N_757,In_1413,In_976);
nor U758 (N_758,N_375,In_1509);
nand U759 (N_759,In_1700,In_507);
and U760 (N_760,In_1567,In_1772);
xnor U761 (N_761,N_305,In_1689);
and U762 (N_762,N_206,In_555);
and U763 (N_763,In_384,In_1787);
or U764 (N_764,In_49,In_1686);
xnor U765 (N_765,N_427,N_102);
xor U766 (N_766,In_1398,In_1576);
nor U767 (N_767,In_1478,In_76);
or U768 (N_768,In_1034,In_216);
and U769 (N_769,In_1240,In_527);
nand U770 (N_770,N_298,N_490);
xor U771 (N_771,N_232,In_1261);
nor U772 (N_772,N_475,N_245);
nor U773 (N_773,N_353,In_1907);
or U774 (N_774,In_1457,N_317);
xnor U775 (N_775,In_1244,In_88);
nor U776 (N_776,In_1330,In_1605);
and U777 (N_777,N_100,N_472);
or U778 (N_778,N_91,In_1939);
nand U779 (N_779,N_363,In_31);
nor U780 (N_780,In_1743,N_141);
xnor U781 (N_781,In_1091,N_168);
nor U782 (N_782,In_1823,N_405);
and U783 (N_783,In_1470,In_1614);
and U784 (N_784,In_345,In_292);
nor U785 (N_785,N_225,In_931);
or U786 (N_786,In_107,N_12);
or U787 (N_787,In_243,In_1944);
and U788 (N_788,N_45,In_423);
or U789 (N_789,N_132,In_1987);
xor U790 (N_790,In_1937,In_1658);
nand U791 (N_791,In_1379,In_1647);
nor U792 (N_792,In_1429,In_1121);
and U793 (N_793,In_1084,N_228);
nand U794 (N_794,N_477,In_379);
and U795 (N_795,In_907,In_1011);
xnor U796 (N_796,In_1806,In_1581);
nor U797 (N_797,N_281,N_448);
nor U798 (N_798,In_1144,N_227);
or U799 (N_799,In_1959,In_1532);
nand U800 (N_800,In_1365,N_85);
or U801 (N_801,N_128,In_478);
and U802 (N_802,In_1721,In_1059);
xor U803 (N_803,In_1241,N_460);
or U804 (N_804,In_1574,In_1184);
and U805 (N_805,In_969,In_282);
and U806 (N_806,In_464,In_452);
xor U807 (N_807,In_69,N_415);
and U808 (N_808,In_208,In_1350);
nor U809 (N_809,In_914,In_1984);
and U810 (N_810,In_1968,N_203);
or U811 (N_811,In_668,In_1468);
and U812 (N_812,In_1952,In_1638);
or U813 (N_813,In_845,In_794);
or U814 (N_814,In_637,N_200);
or U815 (N_815,In_1195,In_1740);
and U816 (N_816,N_334,In_752);
nand U817 (N_817,In_1490,In_1833);
xnor U818 (N_818,N_420,In_732);
or U819 (N_819,N_489,In_1803);
or U820 (N_820,In_1936,In_1006);
or U821 (N_821,In_1777,In_821);
nand U822 (N_822,N_146,N_185);
nor U823 (N_823,In_1634,In_1056);
nor U824 (N_824,In_1977,In_1801);
nor U825 (N_825,In_1859,In_766);
and U826 (N_826,In_1701,In_231);
xor U827 (N_827,N_96,In_965);
nor U828 (N_828,In_1395,In_191);
xnor U829 (N_829,In_627,N_480);
or U830 (N_830,In_434,In_1235);
xor U831 (N_831,In_785,N_47);
nand U832 (N_832,In_1905,N_379);
xor U833 (N_833,In_1442,In_371);
or U834 (N_834,In_1103,In_1930);
nor U835 (N_835,In_937,In_263);
or U836 (N_836,In_1456,In_1469);
and U837 (N_837,In_685,N_328);
xor U838 (N_838,N_167,In_214);
or U839 (N_839,N_152,In_3);
xor U840 (N_840,In_1404,In_471);
or U841 (N_841,In_190,In_1621);
xor U842 (N_842,N_71,N_333);
nor U843 (N_843,In_1828,In_1989);
and U844 (N_844,In_223,In_1271);
nor U845 (N_845,N_380,In_1694);
or U846 (N_846,N_342,In_647);
nor U847 (N_847,In_816,In_8);
and U848 (N_848,N_266,In_641);
nor U849 (N_849,In_1480,In_1098);
xnor U850 (N_850,N_464,N_473);
xor U851 (N_851,In_908,In_1334);
or U852 (N_852,N_166,In_244);
nor U853 (N_853,In_675,In_249);
nor U854 (N_854,In_1136,N_445);
nor U855 (N_855,N_233,In_1582);
or U856 (N_856,N_417,In_1284);
nand U857 (N_857,N_373,In_1893);
nand U858 (N_858,In_857,In_101);
and U859 (N_859,N_443,In_311);
nor U860 (N_860,In_1886,In_378);
xnor U861 (N_861,N_87,In_1748);
xnor U862 (N_862,In_605,N_226);
or U863 (N_863,N_338,In_1086);
nor U864 (N_864,In_751,In_593);
nor U865 (N_865,In_363,N_451);
or U866 (N_866,N_175,In_1602);
xor U867 (N_867,In_274,N_422);
xnor U868 (N_868,In_1667,N_21);
or U869 (N_869,N_183,In_439);
nor U870 (N_870,In_895,N_42);
nand U871 (N_871,N_316,In_257);
and U872 (N_872,N_73,N_50);
nand U873 (N_873,N_291,In_457);
and U874 (N_874,In_1427,In_1640);
nand U875 (N_875,In_443,N_385);
xor U876 (N_876,In_1018,In_554);
nor U877 (N_877,N_323,In_917);
or U878 (N_878,In_1437,In_1611);
nor U879 (N_879,In_1852,N_70);
xor U880 (N_880,In_1960,In_199);
nor U881 (N_881,In_46,N_177);
nor U882 (N_882,In_201,In_1171);
and U883 (N_883,In_1610,In_1263);
xnor U884 (N_884,In_1218,In_1280);
nor U885 (N_885,N_74,N_394);
nand U886 (N_886,N_343,In_100);
or U887 (N_887,In_9,N_33);
and U888 (N_888,In_750,In_1971);
nor U889 (N_889,In_493,In_619);
nor U890 (N_890,In_1792,In_1878);
and U891 (N_891,N_114,In_321);
xor U892 (N_892,In_1138,N_296);
nand U893 (N_893,In_700,In_1560);
and U894 (N_894,N_229,In_1017);
nor U895 (N_895,In_1940,N_287);
xor U896 (N_896,N_209,In_198);
xnor U897 (N_897,N_267,In_997);
xnor U898 (N_898,In_770,In_1377);
nor U899 (N_899,In_25,In_1204);
nor U900 (N_900,In_512,N_408);
xor U901 (N_901,In_944,In_779);
xor U902 (N_902,In_253,N_189);
or U903 (N_903,In_416,N_22);
nor U904 (N_904,In_1870,In_499);
and U905 (N_905,In_1130,N_212);
xor U906 (N_906,N_428,In_431);
and U907 (N_907,In_1510,N_462);
xnor U908 (N_908,In_131,In_1);
and U909 (N_909,In_1259,In_1695);
nor U910 (N_910,N_104,In_1283);
nor U911 (N_911,In_994,N_435);
or U912 (N_912,In_1174,In_1123);
nor U913 (N_913,In_1674,N_19);
and U914 (N_914,In_176,N_34);
nor U915 (N_915,In_913,N_150);
nand U916 (N_916,In_115,In_674);
or U917 (N_917,In_385,N_450);
xnor U918 (N_918,In_1802,In_354);
xor U919 (N_919,In_1975,In_93);
or U920 (N_920,In_187,In_491);
nor U921 (N_921,N_5,N_307);
xor U922 (N_922,In_1175,In_422);
xnor U923 (N_923,N_344,In_792);
nor U924 (N_924,N_145,In_1742);
and U925 (N_925,In_1766,N_110);
nor U926 (N_926,In_165,N_354);
nand U927 (N_927,In_536,N_116);
nand U928 (N_928,N_466,N_54);
and U929 (N_929,N_3,In_1924);
xor U930 (N_930,N_391,N_90);
xnor U931 (N_931,N_434,In_1004);
nor U932 (N_932,In_255,In_1578);
nand U933 (N_933,In_844,In_1273);
or U934 (N_934,In_466,In_1342);
nand U935 (N_935,In_884,N_8);
nor U936 (N_936,In_841,N_322);
xnor U937 (N_937,In_1919,In_915);
nor U938 (N_938,N_10,In_1185);
xnor U939 (N_939,In_317,In_1440);
nand U940 (N_940,In_1009,In_1426);
xor U941 (N_941,N_250,In_1757);
xor U942 (N_942,N_35,N_80);
xnor U943 (N_943,In_1067,In_533);
xor U944 (N_944,In_982,N_301);
xor U945 (N_945,In_261,In_662);
and U946 (N_946,In_1085,In_419);
xnor U947 (N_947,In_973,In_1963);
nor U948 (N_948,In_1842,In_492);
nor U949 (N_949,N_15,In_1129);
or U950 (N_950,N_356,In_1558);
nand U951 (N_951,In_1646,N_255);
or U952 (N_952,N_111,In_1908);
nand U953 (N_953,In_1699,In_1306);
or U954 (N_954,N_217,In_52);
or U955 (N_955,N_164,In_663);
xnor U956 (N_956,N_204,In_601);
and U957 (N_957,In_352,N_131);
nor U958 (N_958,N_382,N_320);
and U959 (N_959,In_1200,N_237);
nor U960 (N_960,In_871,In_690);
nor U961 (N_961,In_518,In_1651);
or U962 (N_962,N_210,In_859);
or U963 (N_963,N_439,N_101);
nand U964 (N_964,N_308,N_485);
nor U965 (N_965,N_107,N_471);
and U966 (N_966,In_229,In_1573);
nor U967 (N_967,In_1073,N_459);
and U968 (N_968,In_182,In_1790);
nand U969 (N_969,In_599,In_775);
xnor U970 (N_970,In_427,In_118);
xnor U971 (N_971,N_404,N_306);
nor U972 (N_972,In_1199,In_1363);
nor U973 (N_973,In_1717,N_236);
and U974 (N_974,N_478,In_738);
or U975 (N_975,In_1683,In_1635);
or U976 (N_976,In_764,In_1467);
or U977 (N_977,In_265,In_756);
nand U978 (N_978,In_940,In_78);
or U979 (N_979,N_327,N_386);
nor U980 (N_980,In_1410,N_27);
or U981 (N_981,In_373,In_1488);
xor U982 (N_982,In_869,In_1761);
and U983 (N_983,In_621,In_1557);
nand U984 (N_984,In_16,N_389);
nor U985 (N_985,N_339,In_888);
nor U986 (N_986,In_689,In_557);
nand U987 (N_987,N_470,In_1956);
nor U988 (N_988,In_1849,In_451);
or U989 (N_989,N_424,In_79);
nand U990 (N_990,N_151,In_45);
nor U991 (N_991,N_271,N_348);
and U992 (N_992,In_644,In_718);
or U993 (N_993,In_54,N_293);
or U994 (N_994,In_1735,In_1282);
xnor U995 (N_995,N_261,In_1160);
nor U996 (N_996,In_161,In_1281);
xor U997 (N_997,N_144,In_181);
or U998 (N_998,N_149,In_1862);
or U999 (N_999,In_97,In_1986);
or U1000 (N_1000,In_514,N_584);
and U1001 (N_1001,N_982,In_286);
xor U1002 (N_1002,N_806,N_526);
xnor U1003 (N_1003,In_1462,N_215);
or U1004 (N_1004,N_469,In_297);
nor U1005 (N_1005,N_207,In_643);
nand U1006 (N_1006,N_845,In_987);
nand U1007 (N_1007,N_565,N_196);
or U1008 (N_1008,In_1035,In_1285);
nand U1009 (N_1009,N_401,N_49);
xnor U1010 (N_1010,N_651,N_509);
or U1011 (N_1011,In_77,In_1156);
nor U1012 (N_1012,N_799,In_1349);
nand U1013 (N_1013,In_278,In_369);
xor U1014 (N_1014,In_577,In_585);
nand U1015 (N_1015,N_891,N_392);
xnor U1016 (N_1016,N_671,N_730);
nor U1017 (N_1017,In_1738,N_914);
nand U1018 (N_1018,In_830,N_731);
xor U1019 (N_1019,N_376,In_34);
xnor U1020 (N_1020,In_959,N_388);
xnor U1021 (N_1021,In_1675,In_486);
nor U1022 (N_1022,In_116,In_1857);
or U1023 (N_1023,In_1887,N_623);
xor U1024 (N_1024,N_527,N_878);
or U1025 (N_1025,N_968,N_360);
nor U1026 (N_1026,N_643,N_821);
xor U1027 (N_1027,N_318,N_996);
and U1028 (N_1028,In_870,N_624);
xnor U1029 (N_1029,N_816,N_479);
and U1030 (N_1030,In_1527,In_1425);
nor U1031 (N_1031,In_800,N_846);
nand U1032 (N_1032,N_798,N_734);
and U1033 (N_1033,N_701,N_581);
and U1034 (N_1034,In_1589,N_899);
and U1035 (N_1035,N_708,N_252);
nand U1036 (N_1036,N_830,In_1179);
nand U1037 (N_1037,In_90,N_289);
nand U1038 (N_1038,N_733,N_658);
nand U1039 (N_1039,N_970,In_1312);
nor U1040 (N_1040,In_1466,N_983);
xnor U1041 (N_1041,N_594,N_628);
nand U1042 (N_1042,N_995,In_335);
or U1043 (N_1043,In_912,In_288);
or U1044 (N_1044,N_858,N_129);
or U1045 (N_1045,In_1045,N_761);
nand U1046 (N_1046,N_807,N_310);
or U1047 (N_1047,N_740,In_1475);
or U1048 (N_1048,N_38,N_790);
and U1049 (N_1049,N_894,N_500);
nand U1050 (N_1050,N_794,N_140);
xor U1051 (N_1051,N_429,N_814);
or U1052 (N_1052,N_263,N_568);
and U1053 (N_1053,In_1985,In_1340);
xnor U1054 (N_1054,In_475,In_739);
and U1055 (N_1055,N_864,N_124);
xnor U1056 (N_1056,N_685,N_602);
and U1057 (N_1057,In_1337,In_505);
or U1058 (N_1058,N_910,N_529);
nand U1059 (N_1059,In_1786,In_1251);
and U1060 (N_1060,N_553,N_654);
and U1061 (N_1061,N_742,N_564);
xnor U1062 (N_1062,N_715,In_842);
nor U1063 (N_1063,In_788,N_803);
xnor U1064 (N_1064,N_604,In_840);
nor U1065 (N_1065,N_888,N_340);
and U1066 (N_1066,N_192,N_767);
and U1067 (N_1067,N_980,N_889);
nor U1068 (N_1068,N_661,N_551);
or U1069 (N_1069,N_897,N_853);
xnor U1070 (N_1070,In_1616,In_124);
and U1071 (N_1071,N_134,N_912);
and U1072 (N_1072,N_519,N_366);
nand U1073 (N_1073,N_36,N_514);
or U1074 (N_1074,In_1233,N_242);
and U1075 (N_1075,N_750,N_484);
and U1076 (N_1076,N_670,N_902);
nand U1077 (N_1077,N_738,N_776);
and U1078 (N_1078,N_856,In_891);
and U1079 (N_1079,N_863,N_590);
nand U1080 (N_1080,In_1296,N_900);
nand U1081 (N_1081,N_950,In_1805);
nor U1082 (N_1082,In_1289,In_1720);
and U1083 (N_1083,N_402,N_608);
and U1084 (N_1084,N_178,In_177);
and U1085 (N_1085,In_927,In_1254);
nor U1086 (N_1086,N_92,In_136);
or U1087 (N_1087,In_272,N_14);
and U1088 (N_1088,In_10,N_842);
or U1089 (N_1089,In_1116,In_1154);
or U1090 (N_1090,In_1678,In_220);
and U1091 (N_1091,In_1464,In_1668);
or U1092 (N_1092,N_7,N_707);
xor U1093 (N_1093,N_425,N_552);
and U1094 (N_1094,N_663,N_660);
and U1095 (N_1095,N_358,N_108);
and U1096 (N_1096,N_859,N_672);
xnor U1097 (N_1097,N_711,N_974);
and U1098 (N_1098,N_571,N_765);
nand U1099 (N_1099,In_1890,N_678);
nand U1100 (N_1100,In_934,In_87);
and U1101 (N_1101,In_1920,N_544);
and U1102 (N_1102,N_913,N_617);
nand U1103 (N_1103,In_413,N_138);
and U1104 (N_1104,N_892,N_525);
nand U1105 (N_1105,N_771,N_238);
nor U1106 (N_1106,In_646,N_284);
nor U1107 (N_1107,N_953,N_947);
nor U1108 (N_1108,In_294,N_825);
xnor U1109 (N_1109,N_925,In_1922);
and U1110 (N_1110,In_1782,In_1730);
and U1111 (N_1111,N_992,N_119);
nor U1112 (N_1112,In_324,N_850);
xnor U1113 (N_1113,N_760,N_55);
xnor U1114 (N_1114,N_810,In_1713);
and U1115 (N_1115,In_1441,N_702);
nand U1116 (N_1116,In_153,N_791);
and U1117 (N_1117,N_726,N_880);
or U1118 (N_1118,N_865,N_668);
xnor U1119 (N_1119,In_986,In_1645);
and U1120 (N_1120,In_734,In_506);
and U1121 (N_1121,N_729,N_578);
xor U1122 (N_1122,N_681,In_289);
xnor U1123 (N_1123,In_1360,In_1888);
nor U1124 (N_1124,In_579,In_1487);
or U1125 (N_1125,N_627,In_971);
xnor U1126 (N_1126,In_1901,N_699);
nand U1127 (N_1127,N_887,N_639);
and U1128 (N_1128,N_592,N_793);
or U1129 (N_1129,N_649,N_686);
nand U1130 (N_1130,N_714,N_507);
nor U1131 (N_1131,N_557,N_540);
and U1132 (N_1132,In_44,N_274);
or U1133 (N_1133,N_31,N_647);
nor U1134 (N_1134,N_800,N_600);
xnor U1135 (N_1135,N_796,N_802);
nor U1136 (N_1136,N_543,N_614);
or U1137 (N_1137,N_481,In_164);
nand U1138 (N_1138,N_205,In_806);
and U1139 (N_1139,N_754,In_1540);
xnor U1140 (N_1140,N_777,N_60);
and U1141 (N_1141,N_875,In_1383);
nand U1142 (N_1142,N_737,In_962);
and U1143 (N_1143,N_508,N_667);
nand U1144 (N_1144,In_575,N_998);
and U1145 (N_1145,N_952,N_549);
and U1146 (N_1146,N_143,N_563);
and U1147 (N_1147,In_1163,In_1113);
nor U1148 (N_1148,N_147,N_759);
nor U1149 (N_1149,N_23,In_1064);
nand U1150 (N_1150,N_693,N_393);
xnor U1151 (N_1151,N_809,N_916);
nand U1152 (N_1152,In_795,In_382);
nand U1153 (N_1153,N_890,N_662);
nand U1154 (N_1154,N_683,N_975);
and U1155 (N_1155,N_606,N_930);
or U1156 (N_1156,N_911,N_57);
or U1157 (N_1157,In_653,N_275);
nand U1158 (N_1158,N_752,N_16);
xor U1159 (N_1159,In_1979,In_743);
nor U1160 (N_1160,In_481,In_19);
nor U1161 (N_1161,N_997,N_940);
nor U1162 (N_1162,In_753,N_655);
xnor U1163 (N_1163,In_441,N_503);
and U1164 (N_1164,In_470,N_467);
nor U1165 (N_1165,N_510,In_1180);
xor U1166 (N_1166,N_374,N_786);
xor U1167 (N_1167,In_63,In_1539);
xor U1168 (N_1168,N_235,N_694);
and U1169 (N_1169,In_608,In_797);
xor U1170 (N_1170,In_1329,N_725);
nand U1171 (N_1171,N_781,N_631);
nor U1172 (N_1172,N_775,In_748);
or U1173 (N_1173,N_780,N_522);
and U1174 (N_1174,N_539,In_1477);
and U1175 (N_1175,In_1319,N_966);
or U1176 (N_1176,In_254,N_576);
nor U1177 (N_1177,N_772,N_986);
or U1178 (N_1178,In_604,In_65);
or U1179 (N_1179,In_1705,In_202);
nand U1180 (N_1180,In_1594,N_560);
nor U1181 (N_1181,N_852,N_482);
and U1182 (N_1182,N_808,In_1128);
nand U1183 (N_1183,N_987,N_763);
nand U1184 (N_1184,N_440,In_530);
and U1185 (N_1185,N_43,N_511);
and U1186 (N_1186,N_587,In_516);
nor U1187 (N_1187,N_931,N_618);
and U1188 (N_1188,N_877,N_616);
and U1189 (N_1189,In_980,N_812);
and U1190 (N_1190,In_1954,N_51);
or U1191 (N_1191,N_787,In_6);
and U1192 (N_1192,In_128,In_1754);
xor U1193 (N_1193,N_615,N_535);
xnor U1194 (N_1194,N_951,In_904);
xnor U1195 (N_1195,In_1980,In_1159);
xor U1196 (N_1196,N_973,N_411);
or U1197 (N_1197,In_1223,N_53);
or U1198 (N_1198,In_1149,In_1393);
and U1199 (N_1199,N_961,N_258);
nor U1200 (N_1200,N_941,N_335);
nand U1201 (N_1201,N_886,N_629);
nor U1202 (N_1202,In_1515,N_397);
xor U1203 (N_1203,N_501,N_719);
and U1204 (N_1204,In_158,N_194);
nor U1205 (N_1205,N_332,N_294);
and U1206 (N_1206,N_330,In_1650);
nand U1207 (N_1207,N_400,N_957);
or U1208 (N_1208,In_1269,N_612);
nor U1209 (N_1209,N_67,N_885);
nor U1210 (N_1210,In_925,N_743);
nand U1211 (N_1211,In_1078,In_1368);
xor U1212 (N_1212,N_674,In_882);
nand U1213 (N_1213,N_948,In_811);
nand U1214 (N_1214,N_160,In_1739);
nor U1215 (N_1215,N_990,N_634);
xnor U1216 (N_1216,N_921,N_901);
xnor U1217 (N_1217,In_1501,In_351);
nand U1218 (N_1218,N_868,N_829);
or U1219 (N_1219,N_234,N_831);
xor U1220 (N_1220,N_984,In_1727);
nand U1221 (N_1221,N_240,N_679);
nand U1222 (N_1222,In_1874,N_190);
or U1223 (N_1223,In_1455,N_580);
or U1224 (N_1224,N_766,N_933);
or U1225 (N_1225,In_1669,In_1508);
nor U1226 (N_1226,N_862,N_171);
nor U1227 (N_1227,N_89,N_324);
or U1228 (N_1228,N_591,N_918);
nor U1229 (N_1229,In_1328,In_733);
nand U1230 (N_1230,In_852,N_773);
and U1231 (N_1231,N_346,N_195);
and U1232 (N_1232,N_917,In_1785);
or U1233 (N_1233,N_770,N_303);
nand U1234 (N_1234,N_985,N_836);
and U1235 (N_1235,N_688,In_688);
xor U1236 (N_1236,N_680,N_609);
xor U1237 (N_1237,In_759,N_611);
nor U1238 (N_1238,N_309,N_502);
and U1239 (N_1239,In_61,N_895);
nor U1240 (N_1240,N_642,In_154);
or U1241 (N_1241,N_669,In_448);
nor U1242 (N_1242,In_1150,In_1858);
nor U1243 (N_1243,N_855,In_1286);
nor U1244 (N_1244,In_875,N_304);
xor U1245 (N_1245,In_1826,N_574);
nor U1246 (N_1246,N_905,N_589);
or U1247 (N_1247,N_843,In_110);
xnor U1248 (N_1248,In_71,N_837);
nand U1249 (N_1249,N_955,N_133);
and U1250 (N_1250,N_659,N_444);
and U1251 (N_1251,N_156,N_757);
xnor U1252 (N_1252,N_954,In_1670);
nand U1253 (N_1253,N_677,N_198);
xnor U1254 (N_1254,In_430,N_566);
or U1255 (N_1255,N_546,N_656);
and U1256 (N_1256,N_520,In_92);
and U1257 (N_1257,In_1309,In_723);
nor U1258 (N_1258,In_436,N_869);
and U1259 (N_1259,N_827,N_61);
xnor U1260 (N_1260,N_645,In_1600);
nor U1261 (N_1261,N_876,In_1896);
nor U1262 (N_1262,N_620,N_820);
xor U1263 (N_1263,In_1412,In_523);
and U1264 (N_1264,N_313,N_118);
and U1265 (N_1265,N_739,In_890);
xnor U1266 (N_1266,N_125,In_1810);
xor U1267 (N_1267,In_1562,N_577);
or U1268 (N_1268,N_906,In_1143);
and U1269 (N_1269,N_441,N_908);
nand U1270 (N_1270,N_929,N_619);
nor U1271 (N_1271,N_972,In_1953);
nand U1272 (N_1272,N_942,N_939);
nor U1273 (N_1273,In_729,N_849);
or U1274 (N_1274,N_934,In_924);
nand U1275 (N_1275,N_872,N_977);
xnor U1276 (N_1276,N_847,N_278);
nor U1277 (N_1277,In_91,N_801);
xor U1278 (N_1278,N_521,N_126);
xor U1279 (N_1279,In_485,N_260);
nand U1280 (N_1280,In_1132,N_979);
nor U1281 (N_1281,N_638,In_197);
and U1282 (N_1282,N_532,N_367);
xnor U1283 (N_1283,N_633,N_747);
and U1284 (N_1284,N_547,N_524);
nor U1285 (N_1285,In_1192,N_182);
or U1286 (N_1286,N_833,In_938);
or U1287 (N_1287,N_873,N_635);
nor U1288 (N_1288,In_1417,In_1556);
nand U1289 (N_1289,N_652,In_1021);
and U1290 (N_1290,In_1111,N_828);
and U1291 (N_1291,In_1868,N_946);
or U1292 (N_1292,In_955,N_676);
and U1293 (N_1293,In_596,N_561);
nand U1294 (N_1294,N_545,N_352);
nor U1295 (N_1295,N_851,N_567);
nor U1296 (N_1296,N_622,In_1684);
xnor U1297 (N_1297,N_811,N_835);
or U1298 (N_1298,In_671,N_665);
nor U1299 (N_1299,N_399,In_1126);
and U1300 (N_1300,N_994,In_787);
or U1301 (N_1301,N_826,In_1518);
nor U1302 (N_1302,In_226,N_768);
nor U1303 (N_1303,In_1047,N_924);
xor U1304 (N_1304,In_300,N_848);
and U1305 (N_1305,N_632,In_592);
nand U1306 (N_1306,N_840,N_689);
and U1307 (N_1307,N_345,N_626);
xnor U1308 (N_1308,N_822,N_838);
xor U1309 (N_1309,In_360,In_188);
and U1310 (N_1310,N_644,N_697);
nand U1311 (N_1311,N_797,N_813);
xnor U1312 (N_1312,In_979,N_99);
and U1313 (N_1313,N_542,N_548);
and U1314 (N_1314,N_745,In_1272);
nor U1315 (N_1315,In_1182,In_1049);
nand U1316 (N_1316,N_161,N_784);
or U1317 (N_1317,N_700,N_898);
or U1318 (N_1318,N_506,N_558);
xnor U1319 (N_1319,N_640,N_646);
and U1320 (N_1320,In_1224,N_783);
nand U1321 (N_1321,N_653,N_932);
nor U1322 (N_1322,In_1716,N_844);
xor U1323 (N_1323,N_753,N_637);
and U1324 (N_1324,N_993,N_46);
and U1325 (N_1325,N_976,In_467);
xor U1326 (N_1326,N_841,In_1076);
or U1327 (N_1327,N_295,N_220);
and U1328 (N_1328,N_555,In_171);
xor U1329 (N_1329,In_545,N_153);
nand U1330 (N_1330,N_272,N_744);
nand U1331 (N_1331,In_1037,N_538);
nand U1332 (N_1332,In_1504,In_1756);
xnor U1333 (N_1333,N_706,In_1148);
nand U1334 (N_1334,N_936,N_496);
xnor U1335 (N_1335,N_692,In_284);
nor U1336 (N_1336,N_297,N_579);
xor U1337 (N_1337,N_66,N_874);
and U1338 (N_1338,N_818,N_636);
and U1339 (N_1339,N_113,In_495);
nand U1340 (N_1340,N_588,In_1949);
nand U1341 (N_1341,N_157,N_684);
or U1342 (N_1342,N_421,N_937);
xnor U1343 (N_1343,N_788,In_1854);
xnor U1344 (N_1344,N_965,In_1320);
nand U1345 (N_1345,N_867,In_1564);
or U1346 (N_1346,In_1519,N_949);
nor U1347 (N_1347,N_712,N_748);
xor U1348 (N_1348,N_173,N_530);
nor U1349 (N_1349,In_768,In_513);
or U1350 (N_1350,N_774,N_65);
or U1351 (N_1351,N_716,N_962);
nand U1352 (N_1352,In_114,N_562);
or U1353 (N_1353,N_749,In_346);
nand U1354 (N_1354,N_860,N_703);
nand U1355 (N_1355,N_769,N_690);
nor U1356 (N_1356,N_350,N_915);
nor U1357 (N_1357,In_1737,N_516);
nor U1358 (N_1358,In_511,N_723);
xor U1359 (N_1359,In_703,N_246);
xor U1360 (N_1360,In_1970,N_371);
xnor U1361 (N_1361,N_751,In_1771);
nor U1362 (N_1362,N_960,N_253);
nor U1363 (N_1363,N_989,In_1202);
xor U1364 (N_1364,N_695,N_832);
xnor U1365 (N_1365,In_1856,N_68);
nor U1366 (N_1366,In_761,N_536);
or U1367 (N_1367,In_667,N_139);
xnor U1368 (N_1368,N_713,N_518);
nand U1369 (N_1369,In_494,In_80);
and U1370 (N_1370,In_1345,In_1326);
nand U1371 (N_1371,In_476,N_935);
or U1372 (N_1372,N_903,N_789);
nor U1373 (N_1373,In_652,N_718);
xnor U1374 (N_1374,N_583,N_641);
xnor U1375 (N_1375,N_248,N_815);
or U1376 (N_1376,N_115,N_541);
and U1377 (N_1377,N_597,N_958);
nor U1378 (N_1378,N_978,In_295);
nor U1379 (N_1379,N_728,N_732);
nor U1380 (N_1380,N_504,N_585);
or U1381 (N_1381,N_861,N_409);
xor U1382 (N_1382,N_927,N_537);
nor U1383 (N_1383,N_218,In_1502);
xor U1384 (N_1384,In_111,In_670);
and U1385 (N_1385,N_573,N_329);
nand U1386 (N_1386,In_1476,In_1114);
or U1387 (N_1387,N_517,N_817);
xor U1388 (N_1388,N_778,N_630);
nand U1389 (N_1389,N_896,N_991);
nor U1390 (N_1390,In_1935,N_664);
and U1391 (N_1391,N_792,N_52);
nor U1392 (N_1392,In_1728,In_350);
or U1393 (N_1393,In_1789,N_735);
nand U1394 (N_1394,N_764,In_196);
nand U1395 (N_1395,N_762,N_724);
or U1396 (N_1396,N_823,N_857);
xor U1397 (N_1397,In_558,N_355);
or U1398 (N_1398,In_75,In_929);
nand U1399 (N_1399,N_523,N_923);
xor U1400 (N_1400,In_583,In_1543);
nor U1401 (N_1401,N_657,N_696);
and U1402 (N_1402,In_699,N_741);
nor U1403 (N_1403,N_264,In_916);
nor U1404 (N_1404,N_944,N_311);
nand U1405 (N_1405,In_562,N_919);
nand U1406 (N_1406,N_687,In_1016);
xor U1407 (N_1407,N_512,N_999);
and U1408 (N_1408,N_4,N_717);
and U1409 (N_1409,N_605,In_581);
nand U1410 (N_1410,N_613,N_610);
or U1411 (N_1411,In_1400,N_208);
or U1412 (N_1412,N_554,N_673);
nand U1413 (N_1413,N_582,In_454);
nor U1414 (N_1414,In_1253,N_413);
and U1415 (N_1415,N_499,In_655);
xnor U1416 (N_1416,N_756,N_383);
or U1417 (N_1417,In_235,N_41);
or U1418 (N_1418,In_1439,N_904);
nand U1419 (N_1419,N_17,N_569);
and U1420 (N_1420,N_58,N_705);
nand U1421 (N_1421,N_357,In_919);
or U1422 (N_1422,N_586,N_398);
nor U1423 (N_1423,N_785,N_11);
and U1424 (N_1424,N_312,N_319);
nand U1425 (N_1425,N_377,N_534);
xor U1426 (N_1426,In_854,N_395);
and U1427 (N_1427,In_1965,In_488);
nand U1428 (N_1428,N_326,N_710);
nand U1429 (N_1429,N_926,In_41);
nand U1430 (N_1430,N_691,N_593);
nor U1431 (N_1431,N_531,N_559);
nand U1432 (N_1432,N_866,N_452);
or U1433 (N_1433,N_219,N_570);
xnor U1434 (N_1434,N_839,In_1010);
nand U1435 (N_1435,N_595,N_556);
nand U1436 (N_1436,N_909,In_1885);
nand U1437 (N_1437,In_881,N_505);
or U1438 (N_1438,N_495,N_603);
nor U1439 (N_1439,In_1438,In_1596);
nor U1440 (N_1440,N_81,In_204);
or U1441 (N_1441,N_364,N_273);
or U1442 (N_1442,In_501,N_596);
and U1443 (N_1443,N_533,N_804);
nand U1444 (N_1444,N_213,In_169);
nor U1445 (N_1445,N_920,N_122);
nor U1446 (N_1446,N_698,N_882);
and U1447 (N_1447,N_675,In_301);
nor U1448 (N_1448,N_883,N_945);
nand U1449 (N_1449,N_755,In_1089);
nor U1450 (N_1450,N_142,N_498);
or U1451 (N_1451,In_22,In_563);
nand U1452 (N_1452,In_150,N_746);
or U1453 (N_1453,N_721,N_879);
or U1454 (N_1454,In_613,In_437);
nor U1455 (N_1455,In_889,In_241);
nor U1456 (N_1456,N_824,N_956);
nor U1457 (N_1457,N_709,In_942);
and U1458 (N_1458,N_938,N_601);
nor U1459 (N_1459,N_834,N_457);
or U1460 (N_1460,N_599,N_870);
nand U1461 (N_1461,N_575,In_835);
or U1462 (N_1462,N_191,N_805);
or U1463 (N_1463,N_598,In_719);
nor U1464 (N_1464,In_1625,In_1370);
nor U1465 (N_1465,N_648,N_928);
nand U1466 (N_1466,In_1257,N_819);
nor U1467 (N_1467,In_332,N_943);
and U1468 (N_1468,In_771,N_550);
or U1469 (N_1469,N_650,N_682);
xnor U1470 (N_1470,N_969,N_981);
or U1471 (N_1471,N_736,N_963);
or U1472 (N_1472,N_572,N_372);
nand U1473 (N_1473,N_75,N_795);
nor U1474 (N_1474,In_1472,In_956);
nand U1475 (N_1475,In_94,N_971);
nor U1476 (N_1476,In_1745,In_1799);
nor U1477 (N_1477,In_1373,N_854);
nand U1478 (N_1478,N_881,N_418);
xnor U1479 (N_1479,In_960,N_362);
and U1480 (N_1480,N_779,N_727);
xor U1481 (N_1481,N_396,N_515);
nand U1482 (N_1482,N_893,In_453);
xor U1483 (N_1483,In_29,N_84);
and U1484 (N_1484,In_207,N_621);
or U1485 (N_1485,N_169,N_871);
nor U1486 (N_1486,In_537,In_990);
nand U1487 (N_1487,N_528,N_607);
or U1488 (N_1488,N_967,N_625);
nor U1489 (N_1489,N_988,In_1933);
nand U1490 (N_1490,N_666,In_726);
or U1491 (N_1491,N_243,N_513);
or U1492 (N_1492,N_704,N_959);
xnor U1493 (N_1493,In_1348,N_280);
nand U1494 (N_1494,In_1303,In_1311);
nand U1495 (N_1495,N_884,N_454);
xor U1496 (N_1496,N_922,N_722);
or U1497 (N_1497,N_782,N_720);
or U1498 (N_1498,N_758,N_239);
nand U1499 (N_1499,N_964,N_907);
and U1500 (N_1500,N_1389,N_1392);
nor U1501 (N_1501,N_1085,N_1019);
nor U1502 (N_1502,N_1204,N_1018);
and U1503 (N_1503,N_1480,N_1440);
and U1504 (N_1504,N_1125,N_1215);
or U1505 (N_1505,N_1162,N_1293);
xor U1506 (N_1506,N_1088,N_1044);
nor U1507 (N_1507,N_1498,N_1350);
nor U1508 (N_1508,N_1374,N_1443);
or U1509 (N_1509,N_1174,N_1250);
and U1510 (N_1510,N_1153,N_1321);
and U1511 (N_1511,N_1145,N_1304);
and U1512 (N_1512,N_1324,N_1188);
nor U1513 (N_1513,N_1436,N_1104);
or U1514 (N_1514,N_1242,N_1186);
xor U1515 (N_1515,N_1181,N_1405);
and U1516 (N_1516,N_1397,N_1446);
xor U1517 (N_1517,N_1227,N_1451);
or U1518 (N_1518,N_1468,N_1168);
and U1519 (N_1519,N_1122,N_1233);
or U1520 (N_1520,N_1001,N_1452);
nor U1521 (N_1521,N_1177,N_1040);
xor U1522 (N_1522,N_1158,N_1076);
nand U1523 (N_1523,N_1302,N_1267);
nand U1524 (N_1524,N_1455,N_1245);
and U1525 (N_1525,N_1244,N_1315);
and U1526 (N_1526,N_1165,N_1354);
and U1527 (N_1527,N_1313,N_1131);
nor U1528 (N_1528,N_1022,N_1118);
nor U1529 (N_1529,N_1264,N_1341);
xor U1530 (N_1530,N_1332,N_1035);
nor U1531 (N_1531,N_1295,N_1139);
xor U1532 (N_1532,N_1248,N_1175);
or U1533 (N_1533,N_1370,N_1442);
and U1534 (N_1534,N_1281,N_1167);
nand U1535 (N_1535,N_1147,N_1499);
xor U1536 (N_1536,N_1318,N_1329);
or U1537 (N_1537,N_1172,N_1219);
nor U1538 (N_1538,N_1235,N_1218);
nor U1539 (N_1539,N_1489,N_1146);
nor U1540 (N_1540,N_1340,N_1102);
xnor U1541 (N_1541,N_1071,N_1484);
or U1542 (N_1542,N_1209,N_1087);
nor U1543 (N_1543,N_1409,N_1257);
and U1544 (N_1544,N_1021,N_1299);
xnor U1545 (N_1545,N_1179,N_1323);
xor U1546 (N_1546,N_1116,N_1277);
and U1547 (N_1547,N_1482,N_1107);
and U1548 (N_1548,N_1461,N_1450);
nand U1549 (N_1549,N_1178,N_1020);
xor U1550 (N_1550,N_1060,N_1337);
nand U1551 (N_1551,N_1239,N_1260);
or U1552 (N_1552,N_1183,N_1191);
or U1553 (N_1553,N_1055,N_1207);
nand U1554 (N_1554,N_1421,N_1403);
or U1555 (N_1555,N_1258,N_1189);
xnor U1556 (N_1556,N_1073,N_1200);
nor U1557 (N_1557,N_1095,N_1325);
or U1558 (N_1558,N_1126,N_1028);
nor U1559 (N_1559,N_1120,N_1353);
xor U1560 (N_1560,N_1345,N_1265);
nor U1561 (N_1561,N_1399,N_1445);
nor U1562 (N_1562,N_1271,N_1469);
nand U1563 (N_1563,N_1124,N_1173);
xnor U1564 (N_1564,N_1142,N_1495);
nor U1565 (N_1565,N_1148,N_1472);
nor U1566 (N_1566,N_1128,N_1268);
and U1567 (N_1567,N_1100,N_1041);
nor U1568 (N_1568,N_1097,N_1077);
xor U1569 (N_1569,N_1135,N_1311);
or U1570 (N_1570,N_1049,N_1263);
and U1571 (N_1571,N_1494,N_1180);
and U1572 (N_1572,N_1479,N_1216);
xnor U1573 (N_1573,N_1474,N_1448);
nand U1574 (N_1574,N_1230,N_1276);
nand U1575 (N_1575,N_1052,N_1256);
or U1576 (N_1576,N_1253,N_1042);
or U1577 (N_1577,N_1224,N_1033);
xnor U1578 (N_1578,N_1388,N_1410);
nor U1579 (N_1579,N_1365,N_1220);
or U1580 (N_1580,N_1029,N_1487);
xor U1581 (N_1581,N_1282,N_1110);
nor U1582 (N_1582,N_1053,N_1015);
nor U1583 (N_1583,N_1284,N_1008);
nand U1584 (N_1584,N_1333,N_1016);
or U1585 (N_1585,N_1261,N_1301);
or U1586 (N_1586,N_1202,N_1026);
nor U1587 (N_1587,N_1433,N_1477);
xor U1588 (N_1588,N_1025,N_1082);
and U1589 (N_1589,N_1288,N_1113);
and U1590 (N_1590,N_1138,N_1185);
and U1591 (N_1591,N_1289,N_1381);
nand U1592 (N_1592,N_1369,N_1080);
or U1593 (N_1593,N_1270,N_1030);
and U1594 (N_1594,N_1223,N_1309);
nor U1595 (N_1595,N_1123,N_1098);
or U1596 (N_1596,N_1195,N_1283);
and U1597 (N_1597,N_1368,N_1361);
nor U1598 (N_1598,N_1214,N_1149);
xnor U1599 (N_1599,N_1419,N_1251);
nor U1600 (N_1600,N_1032,N_1217);
xnor U1601 (N_1601,N_1470,N_1467);
and U1602 (N_1602,N_1243,N_1286);
nand U1603 (N_1603,N_1091,N_1473);
or U1604 (N_1604,N_1320,N_1431);
and U1605 (N_1605,N_1000,N_1294);
nor U1606 (N_1606,N_1017,N_1092);
and U1607 (N_1607,N_1130,N_1013);
nand U1608 (N_1608,N_1434,N_1127);
nand U1609 (N_1609,N_1377,N_1305);
or U1610 (N_1610,N_1447,N_1206);
nor U1611 (N_1611,N_1319,N_1047);
xnor U1612 (N_1612,N_1366,N_1093);
nand U1613 (N_1613,N_1231,N_1057);
nor U1614 (N_1614,N_1466,N_1335);
xnor U1615 (N_1615,N_1342,N_1292);
xnor U1616 (N_1616,N_1290,N_1086);
or U1617 (N_1617,N_1221,N_1068);
and U1618 (N_1618,N_1108,N_1266);
nand U1619 (N_1619,N_1492,N_1111);
and U1620 (N_1620,N_1063,N_1156);
and U1621 (N_1621,N_1312,N_1141);
nand U1622 (N_1622,N_1378,N_1164);
xor U1623 (N_1623,N_1346,N_1004);
nor U1624 (N_1624,N_1238,N_1084);
and U1625 (N_1625,N_1255,N_1423);
nand U1626 (N_1626,N_1427,N_1072);
and U1627 (N_1627,N_1367,N_1054);
or U1628 (N_1628,N_1454,N_1420);
or U1629 (N_1629,N_1391,N_1273);
nand U1630 (N_1630,N_1394,N_1196);
nor U1631 (N_1631,N_1363,N_1306);
xnor U1632 (N_1632,N_1330,N_1297);
or U1633 (N_1633,N_1339,N_1056);
or U1634 (N_1634,N_1232,N_1134);
xor U1635 (N_1635,N_1190,N_1356);
or U1636 (N_1636,N_1184,N_1364);
nor U1637 (N_1637,N_1061,N_1051);
and U1638 (N_1638,N_1280,N_1274);
and U1639 (N_1639,N_1036,N_1048);
and U1640 (N_1640,N_1416,N_1449);
xor U1641 (N_1641,N_1117,N_1338);
or U1642 (N_1642,N_1331,N_1067);
nor U1643 (N_1643,N_1010,N_1432);
xor U1644 (N_1644,N_1062,N_1143);
and U1645 (N_1645,N_1096,N_1430);
xor U1646 (N_1646,N_1279,N_1199);
and U1647 (N_1647,N_1422,N_1114);
nand U1648 (N_1648,N_1163,N_1376);
nand U1649 (N_1649,N_1411,N_1005);
xnor U1650 (N_1650,N_1132,N_1458);
or U1651 (N_1651,N_1438,N_1246);
or U1652 (N_1652,N_1404,N_1212);
nor U1653 (N_1653,N_1193,N_1497);
nand U1654 (N_1654,N_1027,N_1327);
xnor U1655 (N_1655,N_1089,N_1460);
and U1656 (N_1656,N_1129,N_1322);
or U1657 (N_1657,N_1441,N_1252);
nor U1658 (N_1658,N_1398,N_1314);
or U1659 (N_1659,N_1343,N_1038);
nor U1660 (N_1660,N_1444,N_1334);
and U1661 (N_1661,N_1382,N_1486);
xnor U1662 (N_1662,N_1155,N_1307);
xor U1663 (N_1663,N_1247,N_1201);
or U1664 (N_1664,N_1426,N_1357);
nand U1665 (N_1665,N_1464,N_1094);
nor U1666 (N_1666,N_1328,N_1002);
and U1667 (N_1667,N_1105,N_1166);
xor U1668 (N_1668,N_1349,N_1228);
and U1669 (N_1669,N_1176,N_1278);
nand U1670 (N_1670,N_1160,N_1310);
nand U1671 (N_1671,N_1425,N_1344);
nor U1672 (N_1672,N_1006,N_1259);
and U1673 (N_1673,N_1285,N_1065);
or U1674 (N_1674,N_1079,N_1300);
or U1675 (N_1675,N_1187,N_1362);
nand U1676 (N_1676,N_1192,N_1046);
nor U1677 (N_1677,N_1024,N_1208);
or U1678 (N_1678,N_1254,N_1115);
or U1679 (N_1679,N_1222,N_1308);
xor U1680 (N_1680,N_1157,N_1483);
and U1681 (N_1681,N_1194,N_1395);
nand U1682 (N_1682,N_1103,N_1347);
or U1683 (N_1683,N_1112,N_1078);
nor U1684 (N_1684,N_1456,N_1303);
or U1685 (N_1685,N_1379,N_1476);
nor U1686 (N_1686,N_1037,N_1203);
nand U1687 (N_1687,N_1069,N_1406);
nand U1688 (N_1688,N_1490,N_1383);
xor U1689 (N_1689,N_1213,N_1465);
xor U1690 (N_1690,N_1023,N_1262);
nand U1691 (N_1691,N_1150,N_1225);
nor U1692 (N_1692,N_1066,N_1402);
xnor U1693 (N_1693,N_1237,N_1478);
and U1694 (N_1694,N_1491,N_1390);
xor U1695 (N_1695,N_1407,N_1418);
nand U1696 (N_1696,N_1317,N_1413);
xor U1697 (N_1697,N_1151,N_1011);
and U1698 (N_1698,N_1401,N_1336);
or U1699 (N_1699,N_1144,N_1488);
nor U1700 (N_1700,N_1372,N_1083);
or U1701 (N_1701,N_1481,N_1373);
nor U1702 (N_1702,N_1385,N_1159);
and U1703 (N_1703,N_1169,N_1296);
nor U1704 (N_1704,N_1170,N_1275);
or U1705 (N_1705,N_1463,N_1236);
nand U1706 (N_1706,N_1355,N_1211);
nor U1707 (N_1707,N_1133,N_1090);
or U1708 (N_1708,N_1012,N_1358);
or U1709 (N_1709,N_1198,N_1070);
xnor U1710 (N_1710,N_1428,N_1171);
nand U1711 (N_1711,N_1140,N_1074);
xnor U1712 (N_1712,N_1197,N_1471);
and U1713 (N_1713,N_1439,N_1415);
xnor U1714 (N_1714,N_1050,N_1387);
and U1715 (N_1715,N_1059,N_1291);
and U1716 (N_1716,N_1384,N_1351);
xnor U1717 (N_1717,N_1316,N_1371);
xor U1718 (N_1718,N_1412,N_1453);
nor U1719 (N_1719,N_1380,N_1475);
and U1720 (N_1720,N_1400,N_1099);
nand U1721 (N_1721,N_1081,N_1437);
xnor U1722 (N_1722,N_1003,N_1154);
nor U1723 (N_1723,N_1229,N_1386);
or U1724 (N_1724,N_1424,N_1287);
xnor U1725 (N_1725,N_1014,N_1429);
nand U1726 (N_1726,N_1462,N_1043);
xor U1727 (N_1727,N_1106,N_1457);
xor U1728 (N_1728,N_1496,N_1161);
nor U1729 (N_1729,N_1396,N_1241);
and U1730 (N_1730,N_1326,N_1352);
or U1731 (N_1731,N_1064,N_1348);
and U1732 (N_1732,N_1182,N_1408);
nand U1733 (N_1733,N_1459,N_1058);
nand U1734 (N_1734,N_1360,N_1210);
or U1735 (N_1735,N_1435,N_1031);
or U1736 (N_1736,N_1101,N_1485);
nand U1737 (N_1737,N_1137,N_1359);
nand U1738 (N_1738,N_1119,N_1375);
nand U1739 (N_1739,N_1075,N_1226);
or U1740 (N_1740,N_1034,N_1007);
and U1741 (N_1741,N_1249,N_1121);
xor U1742 (N_1742,N_1136,N_1240);
nand U1743 (N_1743,N_1109,N_1272);
xor U1744 (N_1744,N_1493,N_1039);
nand U1745 (N_1745,N_1393,N_1152);
and U1746 (N_1746,N_1298,N_1205);
or U1747 (N_1747,N_1045,N_1009);
and U1748 (N_1748,N_1234,N_1269);
and U1749 (N_1749,N_1417,N_1414);
nand U1750 (N_1750,N_1054,N_1162);
nor U1751 (N_1751,N_1322,N_1154);
xnor U1752 (N_1752,N_1423,N_1230);
xnor U1753 (N_1753,N_1283,N_1243);
and U1754 (N_1754,N_1405,N_1408);
nor U1755 (N_1755,N_1005,N_1457);
nor U1756 (N_1756,N_1140,N_1075);
xnor U1757 (N_1757,N_1180,N_1055);
and U1758 (N_1758,N_1447,N_1209);
xor U1759 (N_1759,N_1092,N_1282);
or U1760 (N_1760,N_1253,N_1475);
nand U1761 (N_1761,N_1278,N_1293);
xnor U1762 (N_1762,N_1471,N_1495);
and U1763 (N_1763,N_1478,N_1118);
xor U1764 (N_1764,N_1053,N_1115);
nor U1765 (N_1765,N_1031,N_1317);
nand U1766 (N_1766,N_1263,N_1103);
nand U1767 (N_1767,N_1307,N_1234);
nor U1768 (N_1768,N_1165,N_1175);
and U1769 (N_1769,N_1426,N_1079);
and U1770 (N_1770,N_1218,N_1219);
and U1771 (N_1771,N_1276,N_1266);
xor U1772 (N_1772,N_1476,N_1086);
nand U1773 (N_1773,N_1202,N_1168);
nor U1774 (N_1774,N_1343,N_1188);
nor U1775 (N_1775,N_1278,N_1160);
nor U1776 (N_1776,N_1381,N_1343);
or U1777 (N_1777,N_1375,N_1462);
or U1778 (N_1778,N_1148,N_1055);
nor U1779 (N_1779,N_1451,N_1180);
xor U1780 (N_1780,N_1149,N_1406);
nand U1781 (N_1781,N_1337,N_1227);
nand U1782 (N_1782,N_1272,N_1152);
nand U1783 (N_1783,N_1056,N_1477);
and U1784 (N_1784,N_1265,N_1475);
or U1785 (N_1785,N_1110,N_1093);
nor U1786 (N_1786,N_1449,N_1400);
and U1787 (N_1787,N_1488,N_1264);
nand U1788 (N_1788,N_1066,N_1046);
xnor U1789 (N_1789,N_1480,N_1299);
nor U1790 (N_1790,N_1002,N_1003);
and U1791 (N_1791,N_1081,N_1131);
nand U1792 (N_1792,N_1467,N_1256);
nand U1793 (N_1793,N_1363,N_1376);
or U1794 (N_1794,N_1411,N_1262);
xor U1795 (N_1795,N_1212,N_1250);
nor U1796 (N_1796,N_1315,N_1259);
nor U1797 (N_1797,N_1448,N_1006);
and U1798 (N_1798,N_1079,N_1061);
nand U1799 (N_1799,N_1240,N_1073);
nand U1800 (N_1800,N_1450,N_1160);
or U1801 (N_1801,N_1114,N_1247);
or U1802 (N_1802,N_1328,N_1475);
or U1803 (N_1803,N_1378,N_1196);
nand U1804 (N_1804,N_1430,N_1007);
or U1805 (N_1805,N_1013,N_1351);
xor U1806 (N_1806,N_1171,N_1241);
xor U1807 (N_1807,N_1143,N_1427);
xnor U1808 (N_1808,N_1435,N_1227);
nand U1809 (N_1809,N_1311,N_1369);
or U1810 (N_1810,N_1037,N_1440);
and U1811 (N_1811,N_1061,N_1109);
nand U1812 (N_1812,N_1407,N_1240);
and U1813 (N_1813,N_1141,N_1351);
nand U1814 (N_1814,N_1229,N_1282);
nand U1815 (N_1815,N_1058,N_1143);
or U1816 (N_1816,N_1259,N_1138);
nand U1817 (N_1817,N_1180,N_1489);
nand U1818 (N_1818,N_1319,N_1406);
and U1819 (N_1819,N_1228,N_1475);
nand U1820 (N_1820,N_1416,N_1133);
or U1821 (N_1821,N_1371,N_1086);
xor U1822 (N_1822,N_1255,N_1000);
or U1823 (N_1823,N_1106,N_1072);
or U1824 (N_1824,N_1289,N_1117);
xnor U1825 (N_1825,N_1305,N_1005);
nand U1826 (N_1826,N_1324,N_1190);
and U1827 (N_1827,N_1020,N_1203);
or U1828 (N_1828,N_1245,N_1287);
xor U1829 (N_1829,N_1227,N_1143);
or U1830 (N_1830,N_1116,N_1402);
nand U1831 (N_1831,N_1034,N_1137);
xnor U1832 (N_1832,N_1262,N_1113);
nand U1833 (N_1833,N_1017,N_1206);
or U1834 (N_1834,N_1410,N_1114);
or U1835 (N_1835,N_1090,N_1299);
xor U1836 (N_1836,N_1202,N_1086);
and U1837 (N_1837,N_1007,N_1111);
and U1838 (N_1838,N_1248,N_1108);
and U1839 (N_1839,N_1292,N_1059);
nand U1840 (N_1840,N_1236,N_1437);
nand U1841 (N_1841,N_1352,N_1181);
xor U1842 (N_1842,N_1155,N_1347);
nand U1843 (N_1843,N_1155,N_1270);
and U1844 (N_1844,N_1037,N_1421);
or U1845 (N_1845,N_1449,N_1079);
and U1846 (N_1846,N_1346,N_1353);
xnor U1847 (N_1847,N_1199,N_1232);
xor U1848 (N_1848,N_1298,N_1344);
nor U1849 (N_1849,N_1336,N_1363);
nand U1850 (N_1850,N_1067,N_1049);
xor U1851 (N_1851,N_1238,N_1487);
nor U1852 (N_1852,N_1170,N_1146);
nor U1853 (N_1853,N_1420,N_1026);
nor U1854 (N_1854,N_1474,N_1153);
nor U1855 (N_1855,N_1073,N_1376);
nand U1856 (N_1856,N_1239,N_1006);
or U1857 (N_1857,N_1371,N_1156);
and U1858 (N_1858,N_1191,N_1228);
and U1859 (N_1859,N_1304,N_1326);
or U1860 (N_1860,N_1164,N_1402);
nand U1861 (N_1861,N_1157,N_1000);
and U1862 (N_1862,N_1304,N_1467);
nor U1863 (N_1863,N_1398,N_1279);
or U1864 (N_1864,N_1030,N_1455);
nor U1865 (N_1865,N_1340,N_1219);
nand U1866 (N_1866,N_1220,N_1063);
nor U1867 (N_1867,N_1145,N_1096);
and U1868 (N_1868,N_1260,N_1300);
nand U1869 (N_1869,N_1172,N_1414);
and U1870 (N_1870,N_1456,N_1477);
nand U1871 (N_1871,N_1325,N_1352);
and U1872 (N_1872,N_1286,N_1355);
xor U1873 (N_1873,N_1246,N_1443);
or U1874 (N_1874,N_1333,N_1403);
nand U1875 (N_1875,N_1363,N_1299);
or U1876 (N_1876,N_1378,N_1423);
and U1877 (N_1877,N_1173,N_1170);
nor U1878 (N_1878,N_1013,N_1024);
or U1879 (N_1879,N_1212,N_1353);
nand U1880 (N_1880,N_1040,N_1118);
or U1881 (N_1881,N_1020,N_1257);
and U1882 (N_1882,N_1185,N_1476);
xnor U1883 (N_1883,N_1209,N_1354);
xor U1884 (N_1884,N_1359,N_1432);
nand U1885 (N_1885,N_1492,N_1138);
nand U1886 (N_1886,N_1262,N_1263);
nand U1887 (N_1887,N_1297,N_1140);
xor U1888 (N_1888,N_1070,N_1433);
nand U1889 (N_1889,N_1171,N_1377);
xnor U1890 (N_1890,N_1218,N_1475);
and U1891 (N_1891,N_1184,N_1233);
nand U1892 (N_1892,N_1466,N_1099);
or U1893 (N_1893,N_1368,N_1229);
nand U1894 (N_1894,N_1057,N_1380);
or U1895 (N_1895,N_1460,N_1133);
nand U1896 (N_1896,N_1397,N_1089);
nor U1897 (N_1897,N_1165,N_1281);
nor U1898 (N_1898,N_1370,N_1105);
nand U1899 (N_1899,N_1320,N_1048);
and U1900 (N_1900,N_1102,N_1237);
nor U1901 (N_1901,N_1301,N_1245);
xnor U1902 (N_1902,N_1402,N_1443);
or U1903 (N_1903,N_1312,N_1188);
nand U1904 (N_1904,N_1066,N_1310);
and U1905 (N_1905,N_1439,N_1175);
and U1906 (N_1906,N_1007,N_1380);
nand U1907 (N_1907,N_1115,N_1021);
and U1908 (N_1908,N_1000,N_1093);
or U1909 (N_1909,N_1214,N_1244);
xor U1910 (N_1910,N_1011,N_1040);
nand U1911 (N_1911,N_1207,N_1303);
and U1912 (N_1912,N_1436,N_1028);
and U1913 (N_1913,N_1342,N_1412);
nand U1914 (N_1914,N_1479,N_1178);
xnor U1915 (N_1915,N_1377,N_1442);
nand U1916 (N_1916,N_1226,N_1142);
xor U1917 (N_1917,N_1131,N_1488);
and U1918 (N_1918,N_1381,N_1011);
or U1919 (N_1919,N_1137,N_1205);
xor U1920 (N_1920,N_1197,N_1108);
or U1921 (N_1921,N_1215,N_1415);
xnor U1922 (N_1922,N_1126,N_1056);
nand U1923 (N_1923,N_1123,N_1117);
xor U1924 (N_1924,N_1311,N_1235);
or U1925 (N_1925,N_1020,N_1126);
xnor U1926 (N_1926,N_1217,N_1099);
nor U1927 (N_1927,N_1124,N_1427);
nand U1928 (N_1928,N_1270,N_1202);
or U1929 (N_1929,N_1339,N_1114);
and U1930 (N_1930,N_1314,N_1251);
nand U1931 (N_1931,N_1435,N_1135);
nor U1932 (N_1932,N_1070,N_1394);
xnor U1933 (N_1933,N_1308,N_1012);
xnor U1934 (N_1934,N_1022,N_1264);
nand U1935 (N_1935,N_1025,N_1294);
xnor U1936 (N_1936,N_1439,N_1239);
and U1937 (N_1937,N_1329,N_1247);
xnor U1938 (N_1938,N_1185,N_1093);
and U1939 (N_1939,N_1073,N_1268);
and U1940 (N_1940,N_1314,N_1305);
nand U1941 (N_1941,N_1313,N_1024);
nor U1942 (N_1942,N_1417,N_1307);
or U1943 (N_1943,N_1389,N_1368);
and U1944 (N_1944,N_1284,N_1454);
nand U1945 (N_1945,N_1446,N_1048);
nand U1946 (N_1946,N_1408,N_1092);
or U1947 (N_1947,N_1147,N_1423);
or U1948 (N_1948,N_1187,N_1337);
nand U1949 (N_1949,N_1147,N_1183);
and U1950 (N_1950,N_1093,N_1022);
nor U1951 (N_1951,N_1281,N_1060);
nand U1952 (N_1952,N_1001,N_1188);
nand U1953 (N_1953,N_1448,N_1307);
nor U1954 (N_1954,N_1474,N_1271);
nor U1955 (N_1955,N_1384,N_1275);
or U1956 (N_1956,N_1039,N_1263);
and U1957 (N_1957,N_1401,N_1024);
nand U1958 (N_1958,N_1434,N_1404);
or U1959 (N_1959,N_1364,N_1469);
and U1960 (N_1960,N_1043,N_1132);
or U1961 (N_1961,N_1493,N_1343);
nand U1962 (N_1962,N_1340,N_1058);
xnor U1963 (N_1963,N_1390,N_1060);
xnor U1964 (N_1964,N_1328,N_1218);
xor U1965 (N_1965,N_1104,N_1318);
and U1966 (N_1966,N_1224,N_1163);
xnor U1967 (N_1967,N_1325,N_1302);
nand U1968 (N_1968,N_1149,N_1365);
nor U1969 (N_1969,N_1402,N_1386);
or U1970 (N_1970,N_1264,N_1069);
or U1971 (N_1971,N_1146,N_1169);
or U1972 (N_1972,N_1213,N_1222);
nor U1973 (N_1973,N_1081,N_1165);
xnor U1974 (N_1974,N_1419,N_1142);
xnor U1975 (N_1975,N_1167,N_1295);
xor U1976 (N_1976,N_1033,N_1090);
and U1977 (N_1977,N_1226,N_1094);
or U1978 (N_1978,N_1276,N_1140);
and U1979 (N_1979,N_1172,N_1215);
xor U1980 (N_1980,N_1490,N_1331);
nor U1981 (N_1981,N_1380,N_1458);
or U1982 (N_1982,N_1423,N_1270);
nor U1983 (N_1983,N_1141,N_1290);
xnor U1984 (N_1984,N_1326,N_1462);
and U1985 (N_1985,N_1069,N_1423);
nand U1986 (N_1986,N_1494,N_1470);
or U1987 (N_1987,N_1109,N_1326);
nand U1988 (N_1988,N_1338,N_1407);
and U1989 (N_1989,N_1488,N_1249);
xor U1990 (N_1990,N_1197,N_1481);
or U1991 (N_1991,N_1476,N_1031);
xor U1992 (N_1992,N_1428,N_1039);
xnor U1993 (N_1993,N_1089,N_1469);
nor U1994 (N_1994,N_1191,N_1141);
nand U1995 (N_1995,N_1341,N_1342);
nand U1996 (N_1996,N_1269,N_1296);
xnor U1997 (N_1997,N_1098,N_1497);
nor U1998 (N_1998,N_1285,N_1461);
nand U1999 (N_1999,N_1340,N_1033);
nand U2000 (N_2000,N_1584,N_1719);
xor U2001 (N_2001,N_1580,N_1586);
xnor U2002 (N_2002,N_1601,N_1571);
or U2003 (N_2003,N_1998,N_1517);
nand U2004 (N_2004,N_1962,N_1864);
or U2005 (N_2005,N_1841,N_1741);
and U2006 (N_2006,N_1913,N_1717);
xnor U2007 (N_2007,N_1805,N_1617);
xor U2008 (N_2008,N_1981,N_1982);
or U2009 (N_2009,N_1831,N_1605);
and U2010 (N_2010,N_1797,N_1651);
xnor U2011 (N_2011,N_1904,N_1914);
nand U2012 (N_2012,N_1699,N_1549);
and U2013 (N_2013,N_1630,N_1877);
nor U2014 (N_2014,N_1681,N_1589);
xnor U2015 (N_2015,N_1692,N_1602);
or U2016 (N_2016,N_1876,N_1745);
nor U2017 (N_2017,N_1955,N_1504);
xor U2018 (N_2018,N_1939,N_1560);
xor U2019 (N_2019,N_1989,N_1514);
nor U2020 (N_2020,N_1579,N_1842);
nor U2021 (N_2021,N_1974,N_1680);
nor U2022 (N_2022,N_1661,N_1813);
nor U2023 (N_2023,N_1619,N_1623);
or U2024 (N_2024,N_1853,N_1624);
nand U2025 (N_2025,N_1888,N_1952);
and U2026 (N_2026,N_1666,N_1505);
nand U2027 (N_2027,N_1771,N_1844);
xor U2028 (N_2028,N_1554,N_1764);
nand U2029 (N_2029,N_1610,N_1582);
and U2030 (N_2030,N_1795,N_1802);
xnor U2031 (N_2031,N_1973,N_1621);
xnor U2032 (N_2032,N_1678,N_1837);
xnor U2033 (N_2033,N_1523,N_1575);
and U2034 (N_2034,N_1570,N_1603);
or U2035 (N_2035,N_1927,N_1716);
and U2036 (N_2036,N_1783,N_1595);
or U2037 (N_2037,N_1714,N_1519);
xnor U2038 (N_2038,N_1984,N_1881);
nor U2039 (N_2039,N_1943,N_1917);
nand U2040 (N_2040,N_1880,N_1569);
or U2041 (N_2041,N_1901,N_1926);
xor U2042 (N_2042,N_1632,N_1938);
nor U2043 (N_2043,N_1810,N_1676);
or U2044 (N_2044,N_1960,N_1792);
nor U2045 (N_2045,N_1700,N_1767);
xor U2046 (N_2046,N_1949,N_1520);
and U2047 (N_2047,N_1965,N_1856);
xnor U2048 (N_2048,N_1903,N_1704);
or U2049 (N_2049,N_1996,N_1874);
nor U2050 (N_2050,N_1636,N_1667);
xnor U2051 (N_2051,N_1510,N_1501);
and U2052 (N_2052,N_1766,N_1834);
xnor U2053 (N_2053,N_1657,N_1663);
xor U2054 (N_2054,N_1525,N_1776);
nor U2055 (N_2055,N_1832,N_1542);
nand U2056 (N_2056,N_1866,N_1635);
nor U2057 (N_2057,N_1838,N_1941);
nor U2058 (N_2058,N_1591,N_1654);
nor U2059 (N_2059,N_1997,N_1550);
or U2060 (N_2060,N_1670,N_1684);
xnor U2061 (N_2061,N_1909,N_1506);
and U2062 (N_2062,N_1851,N_1801);
xor U2063 (N_2063,N_1945,N_1685);
or U2064 (N_2064,N_1855,N_1983);
nor U2065 (N_2065,N_1556,N_1746);
or U2066 (N_2066,N_1759,N_1961);
and U2067 (N_2067,N_1883,N_1648);
nor U2068 (N_2068,N_1780,N_1902);
nand U2069 (N_2069,N_1691,N_1843);
or U2070 (N_2070,N_1588,N_1777);
and U2071 (N_2071,N_1991,N_1976);
nand U2072 (N_2072,N_1957,N_1507);
nand U2073 (N_2073,N_1731,N_1791);
nor U2074 (N_2074,N_1835,N_1786);
xor U2075 (N_2075,N_1628,N_1944);
or U2076 (N_2076,N_1540,N_1977);
or U2077 (N_2077,N_1869,N_1641);
and U2078 (N_2078,N_1953,N_1748);
xnor U2079 (N_2079,N_1994,N_1808);
xnor U2080 (N_2080,N_1912,N_1733);
or U2081 (N_2081,N_1990,N_1705);
xor U2082 (N_2082,N_1544,N_1915);
xor U2083 (N_2083,N_1793,N_1756);
nand U2084 (N_2084,N_1847,N_1749);
nand U2085 (N_2085,N_1911,N_1701);
nand U2086 (N_2086,N_1633,N_1583);
xor U2087 (N_2087,N_1593,N_1599);
and U2088 (N_2088,N_1658,N_1708);
nor U2089 (N_2089,N_1898,N_1942);
xor U2090 (N_2090,N_1634,N_1590);
and U2091 (N_2091,N_1643,N_1723);
xor U2092 (N_2092,N_1796,N_1536);
xnor U2093 (N_2093,N_1566,N_1627);
nor U2094 (N_2094,N_1607,N_1739);
xor U2095 (N_2095,N_1891,N_1581);
and U2096 (N_2096,N_1649,N_1932);
nor U2097 (N_2097,N_1778,N_1873);
and U2098 (N_2098,N_1528,N_1823);
or U2099 (N_2099,N_1713,N_1916);
xnor U2100 (N_2100,N_1697,N_1794);
xnor U2101 (N_2101,N_1897,N_1726);
xnor U2102 (N_2102,N_1850,N_1600);
nor U2103 (N_2103,N_1702,N_1948);
nand U2104 (N_2104,N_1553,N_1679);
or U2105 (N_2105,N_1720,N_1650);
xnor U2106 (N_2106,N_1598,N_1668);
or U2107 (N_2107,N_1821,N_1735);
and U2108 (N_2108,N_1809,N_1555);
or U2109 (N_2109,N_1951,N_1769);
and U2110 (N_2110,N_1924,N_1980);
xnor U2111 (N_2111,N_1761,N_1545);
nor U2112 (N_2112,N_1559,N_1928);
nand U2113 (N_2113,N_1563,N_1518);
or U2114 (N_2114,N_1644,N_1524);
and U2115 (N_2115,N_1640,N_1816);
xnor U2116 (N_2116,N_1988,N_1686);
nor U2117 (N_2117,N_1740,N_1787);
nand U2118 (N_2118,N_1611,N_1537);
nor U2119 (N_2119,N_1752,N_1655);
and U2120 (N_2120,N_1721,N_1529);
xor U2121 (N_2121,N_1712,N_1845);
nor U2122 (N_2122,N_1872,N_1867);
and U2123 (N_2123,N_1933,N_1878);
or U2124 (N_2124,N_1516,N_1659);
and U2125 (N_2125,N_1959,N_1889);
nand U2126 (N_2126,N_1722,N_1750);
nor U2127 (N_2127,N_1711,N_1937);
or U2128 (N_2128,N_1899,N_1615);
nor U2129 (N_2129,N_1687,N_1754);
nor U2130 (N_2130,N_1620,N_1671);
nor U2131 (N_2131,N_1882,N_1987);
nor U2132 (N_2132,N_1758,N_1859);
or U2133 (N_2133,N_1660,N_1995);
nand U2134 (N_2134,N_1585,N_1568);
nor U2135 (N_2135,N_1870,N_1531);
nor U2136 (N_2136,N_1830,N_1541);
and U2137 (N_2137,N_1703,N_1829);
nand U2138 (N_2138,N_1806,N_1594);
nand U2139 (N_2139,N_1696,N_1609);
nor U2140 (N_2140,N_1652,N_1637);
xnor U2141 (N_2141,N_1653,N_1508);
nand U2142 (N_2142,N_1751,N_1828);
xnor U2143 (N_2143,N_1817,N_1790);
or U2144 (N_2144,N_1858,N_1757);
nor U2145 (N_2145,N_1535,N_1857);
xor U2146 (N_2146,N_1985,N_1500);
and U2147 (N_2147,N_1646,N_1782);
nand U2148 (N_2148,N_1895,N_1683);
nor U2149 (N_2149,N_1728,N_1825);
and U2150 (N_2150,N_1564,N_1532);
nor U2151 (N_2151,N_1718,N_1682);
nor U2152 (N_2152,N_1577,N_1673);
and U2153 (N_2153,N_1732,N_1999);
nor U2154 (N_2154,N_1592,N_1613);
or U2155 (N_2155,N_1789,N_1972);
nand U2156 (N_2156,N_1645,N_1747);
nor U2157 (N_2157,N_1921,N_1688);
and U2158 (N_2158,N_1526,N_1647);
or U2159 (N_2159,N_1715,N_1730);
nand U2160 (N_2160,N_1954,N_1665);
nor U2161 (N_2161,N_1967,N_1618);
nor U2162 (N_2162,N_1975,N_1811);
nor U2163 (N_2163,N_1934,N_1743);
or U2164 (N_2164,N_1694,N_1992);
nand U2165 (N_2165,N_1890,N_1521);
or U2166 (N_2166,N_1963,N_1784);
and U2167 (N_2167,N_1935,N_1744);
nor U2168 (N_2168,N_1539,N_1677);
nand U2169 (N_2169,N_1894,N_1587);
nand U2170 (N_2170,N_1753,N_1738);
or U2171 (N_2171,N_1511,N_1885);
nand U2172 (N_2172,N_1538,N_1737);
nand U2173 (N_2173,N_1596,N_1547);
and U2174 (N_2174,N_1512,N_1574);
nand U2175 (N_2175,N_1727,N_1772);
xor U2176 (N_2176,N_1840,N_1839);
or U2177 (N_2177,N_1923,N_1551);
xnor U2178 (N_2178,N_1781,N_1736);
nand U2179 (N_2179,N_1966,N_1562);
xor U2180 (N_2180,N_1706,N_1768);
and U2181 (N_2181,N_1827,N_1978);
or U2182 (N_2182,N_1868,N_1662);
nor U2183 (N_2183,N_1631,N_1760);
xnor U2184 (N_2184,N_1573,N_1725);
and U2185 (N_2185,N_1971,N_1950);
nand U2186 (N_2186,N_1558,N_1892);
nand U2187 (N_2187,N_1622,N_1956);
and U2188 (N_2188,N_1690,N_1875);
or U2189 (N_2189,N_1509,N_1884);
nor U2190 (N_2190,N_1871,N_1552);
xnor U2191 (N_2191,N_1773,N_1695);
xnor U2192 (N_2192,N_1762,N_1968);
and U2193 (N_2193,N_1572,N_1807);
or U2194 (N_2194,N_1906,N_1815);
or U2195 (N_2195,N_1612,N_1625);
nand U2196 (N_2196,N_1861,N_1887);
nand U2197 (N_2197,N_1742,N_1833);
xor U2198 (N_2198,N_1724,N_1546);
or U2199 (N_2199,N_1534,N_1788);
nand U2200 (N_2200,N_1849,N_1765);
xnor U2201 (N_2201,N_1922,N_1799);
or U2202 (N_2202,N_1854,N_1863);
xor U2203 (N_2203,N_1606,N_1865);
or U2204 (N_2204,N_1798,N_1803);
nand U2205 (N_2205,N_1698,N_1629);
nand U2206 (N_2206,N_1709,N_1920);
nor U2207 (N_2207,N_1669,N_1860);
and U2208 (N_2208,N_1936,N_1946);
or U2209 (N_2209,N_1626,N_1820);
and U2210 (N_2210,N_1779,N_1947);
xnor U2211 (N_2211,N_1674,N_1597);
nand U2212 (N_2212,N_1893,N_1907);
nor U2213 (N_2213,N_1836,N_1846);
and U2214 (N_2214,N_1819,N_1543);
xor U2215 (N_2215,N_1502,N_1604);
nor U2216 (N_2216,N_1822,N_1693);
nand U2217 (N_2217,N_1755,N_1930);
or U2218 (N_2218,N_1879,N_1710);
xnor U2219 (N_2219,N_1970,N_1826);
nor U2220 (N_2220,N_1729,N_1576);
and U2221 (N_2221,N_1616,N_1763);
xor U2222 (N_2222,N_1814,N_1993);
nand U2223 (N_2223,N_1530,N_1958);
and U2224 (N_2224,N_1522,N_1852);
and U2225 (N_2225,N_1561,N_1639);
xnor U2226 (N_2226,N_1557,N_1918);
and U2227 (N_2227,N_1608,N_1940);
or U2228 (N_2228,N_1919,N_1785);
nand U2229 (N_2229,N_1969,N_1979);
xor U2230 (N_2230,N_1513,N_1533);
nor U2231 (N_2231,N_1656,N_1672);
xnor U2232 (N_2232,N_1675,N_1567);
or U2233 (N_2233,N_1905,N_1774);
xnor U2234 (N_2234,N_1896,N_1770);
nor U2235 (N_2235,N_1824,N_1886);
nor U2236 (N_2236,N_1900,N_1964);
xnor U2237 (N_2237,N_1908,N_1931);
nor U2238 (N_2238,N_1503,N_1910);
or U2239 (N_2239,N_1929,N_1986);
and U2240 (N_2240,N_1515,N_1775);
xor U2241 (N_2241,N_1548,N_1689);
and U2242 (N_2242,N_1642,N_1925);
and U2243 (N_2243,N_1818,N_1800);
and U2244 (N_2244,N_1734,N_1707);
and U2245 (N_2245,N_1664,N_1848);
or U2246 (N_2246,N_1565,N_1527);
and U2247 (N_2247,N_1614,N_1638);
xor U2248 (N_2248,N_1578,N_1862);
or U2249 (N_2249,N_1804,N_1812);
nor U2250 (N_2250,N_1625,N_1715);
and U2251 (N_2251,N_1995,N_1677);
nor U2252 (N_2252,N_1875,N_1986);
or U2253 (N_2253,N_1574,N_1784);
nor U2254 (N_2254,N_1656,N_1822);
xnor U2255 (N_2255,N_1855,N_1857);
xor U2256 (N_2256,N_1608,N_1600);
or U2257 (N_2257,N_1854,N_1789);
nor U2258 (N_2258,N_1659,N_1998);
or U2259 (N_2259,N_1837,N_1902);
nand U2260 (N_2260,N_1642,N_1777);
nor U2261 (N_2261,N_1758,N_1882);
and U2262 (N_2262,N_1910,N_1761);
and U2263 (N_2263,N_1827,N_1571);
xor U2264 (N_2264,N_1893,N_1760);
xor U2265 (N_2265,N_1944,N_1683);
nor U2266 (N_2266,N_1714,N_1766);
or U2267 (N_2267,N_1963,N_1697);
nand U2268 (N_2268,N_1883,N_1760);
nand U2269 (N_2269,N_1918,N_1721);
and U2270 (N_2270,N_1947,N_1961);
nor U2271 (N_2271,N_1579,N_1998);
nor U2272 (N_2272,N_1951,N_1854);
nor U2273 (N_2273,N_1803,N_1984);
and U2274 (N_2274,N_1974,N_1640);
xnor U2275 (N_2275,N_1727,N_1592);
nor U2276 (N_2276,N_1905,N_1894);
xor U2277 (N_2277,N_1902,N_1648);
xor U2278 (N_2278,N_1784,N_1653);
and U2279 (N_2279,N_1867,N_1745);
xnor U2280 (N_2280,N_1660,N_1630);
nand U2281 (N_2281,N_1976,N_1548);
nor U2282 (N_2282,N_1888,N_1855);
and U2283 (N_2283,N_1900,N_1937);
nor U2284 (N_2284,N_1796,N_1835);
nor U2285 (N_2285,N_1837,N_1923);
nand U2286 (N_2286,N_1621,N_1532);
nor U2287 (N_2287,N_1531,N_1703);
or U2288 (N_2288,N_1699,N_1767);
and U2289 (N_2289,N_1924,N_1700);
nor U2290 (N_2290,N_1781,N_1686);
nor U2291 (N_2291,N_1847,N_1654);
and U2292 (N_2292,N_1573,N_1733);
nor U2293 (N_2293,N_1722,N_1576);
nor U2294 (N_2294,N_1932,N_1829);
xor U2295 (N_2295,N_1819,N_1975);
nor U2296 (N_2296,N_1917,N_1503);
nor U2297 (N_2297,N_1640,N_1520);
or U2298 (N_2298,N_1888,N_1904);
nand U2299 (N_2299,N_1800,N_1860);
nor U2300 (N_2300,N_1551,N_1593);
xnor U2301 (N_2301,N_1874,N_1762);
xor U2302 (N_2302,N_1815,N_1977);
xnor U2303 (N_2303,N_1672,N_1903);
or U2304 (N_2304,N_1693,N_1953);
or U2305 (N_2305,N_1676,N_1943);
nand U2306 (N_2306,N_1925,N_1687);
or U2307 (N_2307,N_1576,N_1995);
or U2308 (N_2308,N_1719,N_1927);
or U2309 (N_2309,N_1738,N_1673);
nor U2310 (N_2310,N_1974,N_1589);
and U2311 (N_2311,N_1820,N_1592);
xnor U2312 (N_2312,N_1954,N_1631);
or U2313 (N_2313,N_1507,N_1970);
and U2314 (N_2314,N_1869,N_1631);
xor U2315 (N_2315,N_1530,N_1972);
xnor U2316 (N_2316,N_1716,N_1710);
nor U2317 (N_2317,N_1644,N_1985);
or U2318 (N_2318,N_1514,N_1632);
nand U2319 (N_2319,N_1803,N_1731);
and U2320 (N_2320,N_1650,N_1575);
xor U2321 (N_2321,N_1590,N_1638);
and U2322 (N_2322,N_1506,N_1942);
nand U2323 (N_2323,N_1744,N_1622);
and U2324 (N_2324,N_1583,N_1885);
and U2325 (N_2325,N_1790,N_1812);
nor U2326 (N_2326,N_1583,N_1685);
nand U2327 (N_2327,N_1563,N_1594);
or U2328 (N_2328,N_1785,N_1641);
nor U2329 (N_2329,N_1832,N_1907);
or U2330 (N_2330,N_1760,N_1658);
and U2331 (N_2331,N_1508,N_1576);
and U2332 (N_2332,N_1918,N_1818);
and U2333 (N_2333,N_1667,N_1943);
or U2334 (N_2334,N_1919,N_1562);
xor U2335 (N_2335,N_1590,N_1500);
or U2336 (N_2336,N_1783,N_1820);
nand U2337 (N_2337,N_1647,N_1727);
xnor U2338 (N_2338,N_1820,N_1550);
xor U2339 (N_2339,N_1516,N_1515);
xor U2340 (N_2340,N_1794,N_1993);
nand U2341 (N_2341,N_1893,N_1790);
or U2342 (N_2342,N_1707,N_1634);
nand U2343 (N_2343,N_1762,N_1934);
and U2344 (N_2344,N_1692,N_1705);
xnor U2345 (N_2345,N_1945,N_1667);
nor U2346 (N_2346,N_1853,N_1780);
and U2347 (N_2347,N_1515,N_1603);
and U2348 (N_2348,N_1537,N_1578);
nor U2349 (N_2349,N_1735,N_1521);
nor U2350 (N_2350,N_1771,N_1949);
and U2351 (N_2351,N_1690,N_1525);
nor U2352 (N_2352,N_1814,N_1944);
xor U2353 (N_2353,N_1666,N_1600);
and U2354 (N_2354,N_1537,N_1828);
nor U2355 (N_2355,N_1715,N_1703);
xnor U2356 (N_2356,N_1536,N_1527);
xnor U2357 (N_2357,N_1785,N_1956);
nor U2358 (N_2358,N_1714,N_1821);
and U2359 (N_2359,N_1563,N_1773);
or U2360 (N_2360,N_1871,N_1815);
nand U2361 (N_2361,N_1729,N_1553);
nand U2362 (N_2362,N_1785,N_1966);
xnor U2363 (N_2363,N_1564,N_1965);
nand U2364 (N_2364,N_1629,N_1942);
or U2365 (N_2365,N_1874,N_1608);
or U2366 (N_2366,N_1568,N_1601);
nor U2367 (N_2367,N_1962,N_1574);
or U2368 (N_2368,N_1956,N_1563);
nor U2369 (N_2369,N_1738,N_1944);
and U2370 (N_2370,N_1879,N_1778);
nor U2371 (N_2371,N_1623,N_1570);
and U2372 (N_2372,N_1726,N_1511);
nand U2373 (N_2373,N_1952,N_1755);
nor U2374 (N_2374,N_1674,N_1644);
xnor U2375 (N_2375,N_1990,N_1951);
xnor U2376 (N_2376,N_1598,N_1965);
xnor U2377 (N_2377,N_1897,N_1709);
nor U2378 (N_2378,N_1790,N_1664);
nor U2379 (N_2379,N_1762,N_1758);
xnor U2380 (N_2380,N_1779,N_1789);
nor U2381 (N_2381,N_1965,N_1616);
nand U2382 (N_2382,N_1974,N_1669);
and U2383 (N_2383,N_1505,N_1546);
nor U2384 (N_2384,N_1540,N_1860);
xor U2385 (N_2385,N_1697,N_1915);
xor U2386 (N_2386,N_1779,N_1734);
nor U2387 (N_2387,N_1934,N_1502);
or U2388 (N_2388,N_1972,N_1794);
and U2389 (N_2389,N_1527,N_1686);
and U2390 (N_2390,N_1741,N_1999);
and U2391 (N_2391,N_1555,N_1787);
xnor U2392 (N_2392,N_1726,N_1954);
nand U2393 (N_2393,N_1991,N_1509);
or U2394 (N_2394,N_1589,N_1967);
nor U2395 (N_2395,N_1772,N_1776);
or U2396 (N_2396,N_1655,N_1633);
or U2397 (N_2397,N_1862,N_1556);
or U2398 (N_2398,N_1579,N_1690);
and U2399 (N_2399,N_1732,N_1773);
or U2400 (N_2400,N_1882,N_1993);
xor U2401 (N_2401,N_1864,N_1508);
xnor U2402 (N_2402,N_1557,N_1533);
nand U2403 (N_2403,N_1712,N_1586);
nor U2404 (N_2404,N_1963,N_1507);
xor U2405 (N_2405,N_1871,N_1962);
nor U2406 (N_2406,N_1756,N_1840);
xnor U2407 (N_2407,N_1599,N_1801);
nor U2408 (N_2408,N_1983,N_1788);
xnor U2409 (N_2409,N_1654,N_1620);
and U2410 (N_2410,N_1988,N_1590);
and U2411 (N_2411,N_1651,N_1528);
nor U2412 (N_2412,N_1802,N_1510);
or U2413 (N_2413,N_1950,N_1562);
nor U2414 (N_2414,N_1912,N_1595);
and U2415 (N_2415,N_1865,N_1901);
xor U2416 (N_2416,N_1517,N_1864);
nand U2417 (N_2417,N_1720,N_1968);
nand U2418 (N_2418,N_1621,N_1552);
and U2419 (N_2419,N_1578,N_1805);
nand U2420 (N_2420,N_1723,N_1693);
nor U2421 (N_2421,N_1749,N_1655);
nor U2422 (N_2422,N_1706,N_1928);
or U2423 (N_2423,N_1553,N_1787);
and U2424 (N_2424,N_1963,N_1600);
or U2425 (N_2425,N_1919,N_1738);
nor U2426 (N_2426,N_1794,N_1891);
and U2427 (N_2427,N_1712,N_1715);
and U2428 (N_2428,N_1591,N_1594);
xor U2429 (N_2429,N_1699,N_1925);
or U2430 (N_2430,N_1796,N_1797);
nand U2431 (N_2431,N_1613,N_1507);
nor U2432 (N_2432,N_1911,N_1544);
nand U2433 (N_2433,N_1764,N_1612);
nor U2434 (N_2434,N_1581,N_1730);
and U2435 (N_2435,N_1680,N_1930);
and U2436 (N_2436,N_1534,N_1984);
or U2437 (N_2437,N_1937,N_1910);
and U2438 (N_2438,N_1697,N_1630);
or U2439 (N_2439,N_1586,N_1669);
nand U2440 (N_2440,N_1746,N_1567);
xnor U2441 (N_2441,N_1535,N_1668);
or U2442 (N_2442,N_1991,N_1760);
and U2443 (N_2443,N_1853,N_1590);
and U2444 (N_2444,N_1647,N_1953);
nand U2445 (N_2445,N_1779,N_1565);
xnor U2446 (N_2446,N_1792,N_1575);
and U2447 (N_2447,N_1718,N_1841);
xnor U2448 (N_2448,N_1852,N_1946);
or U2449 (N_2449,N_1527,N_1918);
nand U2450 (N_2450,N_1538,N_1515);
nand U2451 (N_2451,N_1580,N_1617);
and U2452 (N_2452,N_1595,N_1816);
and U2453 (N_2453,N_1676,N_1603);
xnor U2454 (N_2454,N_1630,N_1557);
and U2455 (N_2455,N_1564,N_1818);
nand U2456 (N_2456,N_1950,N_1556);
nor U2457 (N_2457,N_1854,N_1769);
nand U2458 (N_2458,N_1924,N_1614);
xor U2459 (N_2459,N_1827,N_1819);
xor U2460 (N_2460,N_1515,N_1989);
nand U2461 (N_2461,N_1910,N_1509);
or U2462 (N_2462,N_1883,N_1722);
or U2463 (N_2463,N_1563,N_1683);
and U2464 (N_2464,N_1664,N_1935);
and U2465 (N_2465,N_1689,N_1921);
nand U2466 (N_2466,N_1848,N_1750);
nor U2467 (N_2467,N_1548,N_1838);
or U2468 (N_2468,N_1758,N_1902);
xnor U2469 (N_2469,N_1792,N_1894);
and U2470 (N_2470,N_1958,N_1870);
or U2471 (N_2471,N_1823,N_1737);
and U2472 (N_2472,N_1583,N_1821);
nor U2473 (N_2473,N_1856,N_1503);
or U2474 (N_2474,N_1538,N_1886);
or U2475 (N_2475,N_1824,N_1667);
or U2476 (N_2476,N_1746,N_1976);
nand U2477 (N_2477,N_1795,N_1953);
xnor U2478 (N_2478,N_1809,N_1617);
nor U2479 (N_2479,N_1706,N_1716);
nand U2480 (N_2480,N_1752,N_1522);
nor U2481 (N_2481,N_1954,N_1623);
xor U2482 (N_2482,N_1802,N_1984);
nand U2483 (N_2483,N_1807,N_1912);
nor U2484 (N_2484,N_1599,N_1664);
or U2485 (N_2485,N_1767,N_1777);
and U2486 (N_2486,N_1782,N_1514);
and U2487 (N_2487,N_1539,N_1686);
or U2488 (N_2488,N_1739,N_1788);
xor U2489 (N_2489,N_1502,N_1540);
nand U2490 (N_2490,N_1942,N_1652);
nor U2491 (N_2491,N_1520,N_1744);
and U2492 (N_2492,N_1535,N_1576);
xor U2493 (N_2493,N_1546,N_1557);
or U2494 (N_2494,N_1785,N_1600);
nand U2495 (N_2495,N_1731,N_1671);
nor U2496 (N_2496,N_1699,N_1882);
xnor U2497 (N_2497,N_1989,N_1747);
nor U2498 (N_2498,N_1925,N_1700);
xor U2499 (N_2499,N_1999,N_1681);
nand U2500 (N_2500,N_2298,N_2252);
nor U2501 (N_2501,N_2367,N_2039);
or U2502 (N_2502,N_2406,N_2372);
nand U2503 (N_2503,N_2399,N_2014);
nand U2504 (N_2504,N_2151,N_2365);
xnor U2505 (N_2505,N_2186,N_2037);
and U2506 (N_2506,N_2294,N_2126);
nand U2507 (N_2507,N_2440,N_2047);
or U2508 (N_2508,N_2065,N_2046);
nor U2509 (N_2509,N_2192,N_2301);
xor U2510 (N_2510,N_2056,N_2246);
and U2511 (N_2511,N_2398,N_2305);
nor U2512 (N_2512,N_2110,N_2179);
nand U2513 (N_2513,N_2359,N_2084);
nor U2514 (N_2514,N_2468,N_2290);
nor U2515 (N_2515,N_2013,N_2419);
nand U2516 (N_2516,N_2401,N_2490);
nand U2517 (N_2517,N_2424,N_2346);
and U2518 (N_2518,N_2463,N_2445);
nand U2519 (N_2519,N_2420,N_2380);
and U2520 (N_2520,N_2122,N_2313);
or U2521 (N_2521,N_2432,N_2247);
nand U2522 (N_2522,N_2338,N_2370);
nor U2523 (N_2523,N_2194,N_2334);
or U2524 (N_2524,N_2384,N_2105);
nor U2525 (N_2525,N_2373,N_2091);
nor U2526 (N_2526,N_2415,N_2207);
nor U2527 (N_2527,N_2208,N_2141);
xor U2528 (N_2528,N_2352,N_2167);
or U2529 (N_2529,N_2456,N_2259);
nor U2530 (N_2530,N_2462,N_2072);
xnor U2531 (N_2531,N_2115,N_2342);
nand U2532 (N_2532,N_2286,N_2275);
nor U2533 (N_2533,N_2053,N_2035);
nor U2534 (N_2534,N_2009,N_2412);
xor U2535 (N_2535,N_2228,N_2098);
nand U2536 (N_2536,N_2332,N_2345);
nand U2537 (N_2537,N_2137,N_2357);
xor U2538 (N_2538,N_2333,N_2470);
and U2539 (N_2539,N_2184,N_2460);
xnor U2540 (N_2540,N_2066,N_2103);
nand U2541 (N_2541,N_2113,N_2466);
xnor U2542 (N_2542,N_2042,N_2389);
xor U2543 (N_2543,N_2385,N_2344);
or U2544 (N_2544,N_2237,N_2022);
nand U2545 (N_2545,N_2254,N_2457);
or U2546 (N_2546,N_2421,N_2293);
or U2547 (N_2547,N_2410,N_2443);
or U2548 (N_2548,N_2270,N_2128);
xor U2549 (N_2549,N_2317,N_2076);
nor U2550 (N_2550,N_2284,N_2494);
nor U2551 (N_2551,N_2364,N_2133);
xnor U2552 (N_2552,N_2161,N_2442);
and U2553 (N_2553,N_2086,N_2355);
nor U2554 (N_2554,N_2185,N_2243);
nor U2555 (N_2555,N_2465,N_2176);
nor U2556 (N_2556,N_2394,N_2255);
nor U2557 (N_2557,N_2267,N_2487);
xnor U2558 (N_2558,N_2145,N_2092);
nor U2559 (N_2559,N_2233,N_2132);
or U2560 (N_2560,N_2478,N_2016);
xnor U2561 (N_2561,N_2261,N_2429);
xor U2562 (N_2562,N_2172,N_2044);
nor U2563 (N_2563,N_2164,N_2127);
nor U2564 (N_2564,N_2190,N_2191);
xor U2565 (N_2565,N_2052,N_2241);
or U2566 (N_2566,N_2077,N_2390);
and U2567 (N_2567,N_2304,N_2337);
nor U2568 (N_2568,N_2257,N_2195);
nand U2569 (N_2569,N_2213,N_2393);
nand U2570 (N_2570,N_2150,N_2223);
xor U2571 (N_2571,N_2476,N_2276);
nand U2572 (N_2572,N_2116,N_2029);
nand U2573 (N_2573,N_2363,N_2239);
or U2574 (N_2574,N_2099,N_2388);
and U2575 (N_2575,N_2002,N_2483);
xor U2576 (N_2576,N_2263,N_2203);
or U2577 (N_2577,N_2413,N_2064);
nor U2578 (N_2578,N_2021,N_2378);
nand U2579 (N_2579,N_2278,N_2081);
nand U2580 (N_2580,N_2123,N_2454);
nor U2581 (N_2581,N_2031,N_2493);
nor U2582 (N_2582,N_2287,N_2376);
nand U2583 (N_2583,N_2019,N_2229);
and U2584 (N_2584,N_2451,N_2187);
xnor U2585 (N_2585,N_2196,N_2326);
nor U2586 (N_2586,N_2142,N_2330);
xnor U2587 (N_2587,N_2020,N_2093);
or U2588 (N_2588,N_2392,N_2461);
xnor U2589 (N_2589,N_2486,N_2422);
nand U2590 (N_2590,N_2168,N_2215);
xnor U2591 (N_2591,N_2260,N_2154);
nor U2592 (N_2592,N_2448,N_2446);
or U2593 (N_2593,N_2244,N_2004);
xor U2594 (N_2594,N_2489,N_2225);
or U2595 (N_2595,N_2467,N_2174);
nand U2596 (N_2596,N_2354,N_2049);
nand U2597 (N_2597,N_2234,N_2012);
and U2598 (N_2598,N_2006,N_2268);
nand U2599 (N_2599,N_2408,N_2315);
and U2600 (N_2600,N_2414,N_2158);
xor U2601 (N_2601,N_2235,N_2182);
nand U2602 (N_2602,N_2400,N_2003);
nor U2603 (N_2603,N_2485,N_2297);
and U2604 (N_2604,N_2499,N_2479);
nand U2605 (N_2605,N_2061,N_2481);
xor U2606 (N_2606,N_2480,N_2121);
and U2607 (N_2607,N_2095,N_2302);
nand U2608 (N_2608,N_2045,N_2030);
and U2609 (N_2609,N_2417,N_2189);
or U2610 (N_2610,N_2282,N_2271);
and U2611 (N_2611,N_2273,N_2048);
and U2612 (N_2612,N_2319,N_2375);
and U2613 (N_2613,N_2159,N_2202);
and U2614 (N_2614,N_2140,N_2070);
xnor U2615 (N_2615,N_2166,N_2368);
and U2616 (N_2616,N_2131,N_2078);
or U2617 (N_2617,N_2311,N_2124);
and U2618 (N_2618,N_2382,N_2032);
nand U2619 (N_2619,N_2114,N_2108);
xnor U2620 (N_2620,N_2232,N_2144);
or U2621 (N_2621,N_2227,N_2226);
or U2622 (N_2622,N_2308,N_2082);
and U2623 (N_2623,N_2007,N_2452);
or U2624 (N_2624,N_2079,N_2111);
xor U2625 (N_2625,N_2051,N_2430);
nor U2626 (N_2626,N_2216,N_2438);
nor U2627 (N_2627,N_2001,N_2075);
xor U2628 (N_2628,N_2265,N_2336);
nor U2629 (N_2629,N_2120,N_2100);
xor U2630 (N_2630,N_2102,N_2296);
nand U2631 (N_2631,N_2281,N_2057);
nor U2632 (N_2632,N_2221,N_2387);
nand U2633 (N_2633,N_2200,N_2143);
nor U2634 (N_2634,N_2283,N_2088);
nand U2635 (N_2635,N_2036,N_2224);
nor U2636 (N_2636,N_2374,N_2135);
xnor U2637 (N_2637,N_2397,N_2258);
or U2638 (N_2638,N_2183,N_2018);
and U2639 (N_2639,N_2104,N_2475);
nand U2640 (N_2640,N_2369,N_2096);
nand U2641 (N_2641,N_2193,N_2360);
nand U2642 (N_2642,N_2269,N_2175);
and U2643 (N_2643,N_2038,N_2222);
xnor U2644 (N_2644,N_2136,N_2146);
and U2645 (N_2645,N_2156,N_2165);
and U2646 (N_2646,N_2214,N_2469);
or U2647 (N_2647,N_2139,N_2251);
nor U2648 (N_2648,N_2325,N_2312);
xor U2649 (N_2649,N_2063,N_2425);
or U2650 (N_2650,N_2418,N_2059);
nor U2651 (N_2651,N_2211,N_2147);
nand U2652 (N_2652,N_2300,N_2000);
nand U2653 (N_2653,N_2205,N_2323);
nand U2654 (N_2654,N_2062,N_2027);
nand U2655 (N_2655,N_2130,N_2089);
or U2656 (N_2656,N_2043,N_2307);
and U2657 (N_2657,N_2427,N_2491);
nand U2658 (N_2658,N_2288,N_2238);
and U2659 (N_2659,N_2209,N_2178);
and U2660 (N_2660,N_2148,N_2231);
or U2661 (N_2661,N_2274,N_2160);
nand U2662 (N_2662,N_2118,N_2381);
or U2663 (N_2663,N_2033,N_2220);
xnor U2664 (N_2664,N_2498,N_2210);
and U2665 (N_2665,N_2107,N_2085);
nor U2666 (N_2666,N_2169,N_2152);
xor U2667 (N_2667,N_2264,N_2017);
and U2668 (N_2668,N_2010,N_2090);
and U2669 (N_2669,N_2201,N_2416);
and U2670 (N_2670,N_2248,N_2074);
nand U2671 (N_2671,N_2428,N_2157);
nor U2672 (N_2672,N_2155,N_2101);
nand U2673 (N_2673,N_2409,N_2492);
nor U2674 (N_2674,N_2383,N_2219);
xor U2675 (N_2675,N_2431,N_2453);
or U2676 (N_2676,N_2250,N_2071);
xnor U2677 (N_2677,N_2306,N_2005);
xor U2678 (N_2678,N_2181,N_2347);
and U2679 (N_2679,N_2285,N_2495);
nor U2680 (N_2680,N_2351,N_2015);
xnor U2681 (N_2681,N_2474,N_2329);
nand U2682 (N_2682,N_2358,N_2177);
and U2683 (N_2683,N_2441,N_2377);
or U2684 (N_2684,N_2386,N_2361);
or U2685 (N_2685,N_2058,N_2349);
nand U2686 (N_2686,N_2197,N_2112);
nor U2687 (N_2687,N_2435,N_2279);
and U2688 (N_2688,N_2437,N_2477);
xor U2689 (N_2689,N_2423,N_2362);
and U2690 (N_2690,N_2129,N_2055);
nand U2691 (N_2691,N_2069,N_2455);
and U2692 (N_2692,N_2180,N_2138);
and U2693 (N_2693,N_2087,N_2083);
nand U2694 (N_2694,N_2318,N_2280);
nand U2695 (N_2695,N_2371,N_2230);
or U2696 (N_2696,N_2067,N_2028);
nor U2697 (N_2697,N_2153,N_2447);
and U2698 (N_2698,N_2008,N_2343);
or U2699 (N_2699,N_2482,N_2391);
or U2700 (N_2700,N_2073,N_2188);
nor U2701 (N_2701,N_2405,N_2212);
xor U2702 (N_2702,N_2497,N_2149);
and U2703 (N_2703,N_2402,N_2291);
xnor U2704 (N_2704,N_2366,N_2034);
or U2705 (N_2705,N_2094,N_2316);
nand U2706 (N_2706,N_2080,N_2472);
nor U2707 (N_2707,N_2407,N_2041);
nand U2708 (N_2708,N_2170,N_2125);
and U2709 (N_2709,N_2218,N_2303);
nor U2710 (N_2710,N_2350,N_2068);
nor U2711 (N_2711,N_2198,N_2458);
or U2712 (N_2712,N_2436,N_2245);
xor U2713 (N_2713,N_2024,N_2289);
and U2714 (N_2714,N_2433,N_2050);
nor U2715 (N_2715,N_2162,N_2426);
nor U2716 (N_2716,N_2327,N_2025);
or U2717 (N_2717,N_2471,N_2320);
or U2718 (N_2718,N_2488,N_2411);
nand U2719 (N_2719,N_2339,N_2109);
and U2720 (N_2720,N_2444,N_2395);
nor U2721 (N_2721,N_2403,N_2292);
nor U2722 (N_2722,N_2404,N_2199);
xnor U2723 (N_2723,N_2464,N_2040);
or U2724 (N_2724,N_2117,N_2310);
and U2725 (N_2725,N_2272,N_2396);
or U2726 (N_2726,N_2353,N_2379);
or U2727 (N_2727,N_2295,N_2206);
xor U2728 (N_2728,N_2341,N_2256);
and U2729 (N_2729,N_2324,N_2011);
nand U2730 (N_2730,N_2484,N_2449);
or U2731 (N_2731,N_2262,N_2348);
xnor U2732 (N_2732,N_2277,N_2321);
nand U2733 (N_2733,N_2335,N_2328);
and U2734 (N_2734,N_2356,N_2473);
nand U2735 (N_2735,N_2119,N_2060);
nor U2736 (N_2736,N_2314,N_2459);
or U2737 (N_2737,N_2253,N_2439);
xnor U2738 (N_2738,N_2097,N_2054);
nor U2739 (N_2739,N_2331,N_2217);
or U2740 (N_2740,N_2299,N_2249);
and U2741 (N_2741,N_2026,N_2236);
nor U2742 (N_2742,N_2434,N_2204);
nand U2743 (N_2743,N_2340,N_2106);
nand U2744 (N_2744,N_2496,N_2309);
xnor U2745 (N_2745,N_2242,N_2171);
nor U2746 (N_2746,N_2173,N_2322);
nand U2747 (N_2747,N_2163,N_2450);
or U2748 (N_2748,N_2023,N_2134);
nor U2749 (N_2749,N_2266,N_2240);
xor U2750 (N_2750,N_2451,N_2360);
xnor U2751 (N_2751,N_2477,N_2135);
or U2752 (N_2752,N_2319,N_2108);
xor U2753 (N_2753,N_2033,N_2134);
nand U2754 (N_2754,N_2482,N_2009);
or U2755 (N_2755,N_2021,N_2046);
nand U2756 (N_2756,N_2458,N_2329);
nand U2757 (N_2757,N_2022,N_2321);
or U2758 (N_2758,N_2044,N_2321);
and U2759 (N_2759,N_2367,N_2107);
and U2760 (N_2760,N_2454,N_2465);
or U2761 (N_2761,N_2041,N_2385);
and U2762 (N_2762,N_2460,N_2099);
nand U2763 (N_2763,N_2346,N_2366);
nor U2764 (N_2764,N_2082,N_2331);
and U2765 (N_2765,N_2395,N_2059);
nor U2766 (N_2766,N_2471,N_2370);
nor U2767 (N_2767,N_2477,N_2211);
and U2768 (N_2768,N_2416,N_2144);
nand U2769 (N_2769,N_2157,N_2177);
or U2770 (N_2770,N_2140,N_2478);
nor U2771 (N_2771,N_2300,N_2134);
nand U2772 (N_2772,N_2263,N_2124);
xor U2773 (N_2773,N_2343,N_2435);
nor U2774 (N_2774,N_2084,N_2485);
and U2775 (N_2775,N_2150,N_2089);
or U2776 (N_2776,N_2306,N_2353);
xnor U2777 (N_2777,N_2031,N_2159);
nor U2778 (N_2778,N_2436,N_2431);
nor U2779 (N_2779,N_2486,N_2356);
or U2780 (N_2780,N_2108,N_2104);
and U2781 (N_2781,N_2423,N_2494);
xnor U2782 (N_2782,N_2268,N_2487);
xnor U2783 (N_2783,N_2205,N_2419);
or U2784 (N_2784,N_2136,N_2078);
xnor U2785 (N_2785,N_2057,N_2397);
nor U2786 (N_2786,N_2435,N_2401);
and U2787 (N_2787,N_2069,N_2260);
and U2788 (N_2788,N_2035,N_2403);
and U2789 (N_2789,N_2122,N_2351);
xor U2790 (N_2790,N_2089,N_2340);
nor U2791 (N_2791,N_2416,N_2021);
xor U2792 (N_2792,N_2195,N_2237);
nor U2793 (N_2793,N_2375,N_2249);
or U2794 (N_2794,N_2072,N_2005);
xor U2795 (N_2795,N_2048,N_2152);
nand U2796 (N_2796,N_2257,N_2492);
or U2797 (N_2797,N_2493,N_2386);
and U2798 (N_2798,N_2317,N_2044);
or U2799 (N_2799,N_2052,N_2118);
nand U2800 (N_2800,N_2434,N_2398);
and U2801 (N_2801,N_2372,N_2176);
and U2802 (N_2802,N_2274,N_2213);
or U2803 (N_2803,N_2331,N_2483);
nand U2804 (N_2804,N_2220,N_2285);
nor U2805 (N_2805,N_2060,N_2267);
nor U2806 (N_2806,N_2412,N_2157);
and U2807 (N_2807,N_2340,N_2137);
xor U2808 (N_2808,N_2062,N_2341);
xnor U2809 (N_2809,N_2383,N_2342);
xnor U2810 (N_2810,N_2246,N_2094);
and U2811 (N_2811,N_2319,N_2499);
and U2812 (N_2812,N_2304,N_2271);
and U2813 (N_2813,N_2329,N_2249);
nor U2814 (N_2814,N_2367,N_2479);
xnor U2815 (N_2815,N_2091,N_2124);
xnor U2816 (N_2816,N_2185,N_2271);
or U2817 (N_2817,N_2362,N_2034);
or U2818 (N_2818,N_2380,N_2415);
nor U2819 (N_2819,N_2449,N_2370);
nor U2820 (N_2820,N_2235,N_2365);
nand U2821 (N_2821,N_2261,N_2496);
or U2822 (N_2822,N_2362,N_2324);
nand U2823 (N_2823,N_2042,N_2151);
or U2824 (N_2824,N_2404,N_2304);
or U2825 (N_2825,N_2215,N_2471);
and U2826 (N_2826,N_2254,N_2165);
xor U2827 (N_2827,N_2281,N_2238);
nand U2828 (N_2828,N_2086,N_2269);
nand U2829 (N_2829,N_2385,N_2051);
and U2830 (N_2830,N_2359,N_2380);
nand U2831 (N_2831,N_2143,N_2142);
and U2832 (N_2832,N_2380,N_2480);
and U2833 (N_2833,N_2085,N_2024);
xor U2834 (N_2834,N_2431,N_2377);
and U2835 (N_2835,N_2443,N_2471);
xor U2836 (N_2836,N_2398,N_2228);
nor U2837 (N_2837,N_2119,N_2232);
xnor U2838 (N_2838,N_2150,N_2087);
nand U2839 (N_2839,N_2452,N_2223);
xor U2840 (N_2840,N_2241,N_2142);
xor U2841 (N_2841,N_2227,N_2456);
xnor U2842 (N_2842,N_2238,N_2030);
or U2843 (N_2843,N_2325,N_2273);
nor U2844 (N_2844,N_2076,N_2096);
xor U2845 (N_2845,N_2069,N_2164);
nor U2846 (N_2846,N_2487,N_2014);
nand U2847 (N_2847,N_2468,N_2325);
or U2848 (N_2848,N_2332,N_2212);
nand U2849 (N_2849,N_2294,N_2010);
or U2850 (N_2850,N_2043,N_2371);
and U2851 (N_2851,N_2318,N_2214);
nand U2852 (N_2852,N_2124,N_2008);
and U2853 (N_2853,N_2034,N_2436);
nand U2854 (N_2854,N_2385,N_2321);
and U2855 (N_2855,N_2162,N_2238);
and U2856 (N_2856,N_2489,N_2149);
nand U2857 (N_2857,N_2465,N_2439);
nor U2858 (N_2858,N_2014,N_2044);
or U2859 (N_2859,N_2025,N_2363);
nand U2860 (N_2860,N_2405,N_2025);
nand U2861 (N_2861,N_2214,N_2134);
xor U2862 (N_2862,N_2082,N_2033);
and U2863 (N_2863,N_2318,N_2186);
or U2864 (N_2864,N_2016,N_2379);
and U2865 (N_2865,N_2093,N_2415);
nand U2866 (N_2866,N_2213,N_2192);
nor U2867 (N_2867,N_2111,N_2276);
and U2868 (N_2868,N_2354,N_2265);
and U2869 (N_2869,N_2351,N_2059);
nand U2870 (N_2870,N_2064,N_2436);
xor U2871 (N_2871,N_2319,N_2429);
or U2872 (N_2872,N_2231,N_2377);
or U2873 (N_2873,N_2243,N_2453);
nand U2874 (N_2874,N_2473,N_2019);
or U2875 (N_2875,N_2217,N_2161);
xnor U2876 (N_2876,N_2496,N_2259);
nand U2877 (N_2877,N_2123,N_2457);
nor U2878 (N_2878,N_2400,N_2380);
xor U2879 (N_2879,N_2292,N_2253);
xnor U2880 (N_2880,N_2409,N_2457);
nand U2881 (N_2881,N_2097,N_2263);
nor U2882 (N_2882,N_2495,N_2385);
nor U2883 (N_2883,N_2213,N_2125);
and U2884 (N_2884,N_2289,N_2078);
nand U2885 (N_2885,N_2439,N_2355);
nand U2886 (N_2886,N_2327,N_2191);
nand U2887 (N_2887,N_2224,N_2458);
and U2888 (N_2888,N_2413,N_2083);
nor U2889 (N_2889,N_2235,N_2318);
or U2890 (N_2890,N_2016,N_2310);
nor U2891 (N_2891,N_2432,N_2137);
nand U2892 (N_2892,N_2016,N_2178);
and U2893 (N_2893,N_2174,N_2184);
and U2894 (N_2894,N_2158,N_2396);
or U2895 (N_2895,N_2288,N_2274);
nand U2896 (N_2896,N_2303,N_2222);
or U2897 (N_2897,N_2215,N_2490);
nand U2898 (N_2898,N_2298,N_2109);
nand U2899 (N_2899,N_2052,N_2381);
nor U2900 (N_2900,N_2495,N_2197);
nor U2901 (N_2901,N_2425,N_2465);
and U2902 (N_2902,N_2463,N_2055);
nand U2903 (N_2903,N_2033,N_2285);
or U2904 (N_2904,N_2304,N_2219);
nand U2905 (N_2905,N_2176,N_2081);
and U2906 (N_2906,N_2110,N_2030);
xnor U2907 (N_2907,N_2376,N_2411);
xor U2908 (N_2908,N_2179,N_2253);
xor U2909 (N_2909,N_2043,N_2299);
nand U2910 (N_2910,N_2268,N_2162);
xor U2911 (N_2911,N_2479,N_2005);
nor U2912 (N_2912,N_2011,N_2227);
xor U2913 (N_2913,N_2487,N_2182);
and U2914 (N_2914,N_2460,N_2323);
nand U2915 (N_2915,N_2039,N_2168);
nand U2916 (N_2916,N_2172,N_2349);
or U2917 (N_2917,N_2185,N_2352);
xnor U2918 (N_2918,N_2229,N_2287);
or U2919 (N_2919,N_2429,N_2118);
nor U2920 (N_2920,N_2018,N_2114);
xor U2921 (N_2921,N_2415,N_2015);
xor U2922 (N_2922,N_2183,N_2182);
nand U2923 (N_2923,N_2016,N_2222);
nor U2924 (N_2924,N_2356,N_2138);
and U2925 (N_2925,N_2210,N_2358);
and U2926 (N_2926,N_2045,N_2284);
nor U2927 (N_2927,N_2313,N_2469);
or U2928 (N_2928,N_2021,N_2476);
or U2929 (N_2929,N_2005,N_2249);
or U2930 (N_2930,N_2373,N_2451);
nor U2931 (N_2931,N_2252,N_2023);
nand U2932 (N_2932,N_2093,N_2079);
nand U2933 (N_2933,N_2354,N_2464);
and U2934 (N_2934,N_2387,N_2126);
nand U2935 (N_2935,N_2289,N_2019);
nor U2936 (N_2936,N_2010,N_2065);
xor U2937 (N_2937,N_2356,N_2477);
and U2938 (N_2938,N_2392,N_2356);
nand U2939 (N_2939,N_2109,N_2223);
and U2940 (N_2940,N_2065,N_2038);
nand U2941 (N_2941,N_2065,N_2386);
nor U2942 (N_2942,N_2392,N_2457);
xor U2943 (N_2943,N_2210,N_2493);
and U2944 (N_2944,N_2238,N_2475);
xnor U2945 (N_2945,N_2475,N_2205);
nor U2946 (N_2946,N_2368,N_2415);
xor U2947 (N_2947,N_2114,N_2315);
or U2948 (N_2948,N_2251,N_2220);
nor U2949 (N_2949,N_2464,N_2256);
and U2950 (N_2950,N_2457,N_2036);
or U2951 (N_2951,N_2302,N_2198);
xnor U2952 (N_2952,N_2287,N_2479);
nor U2953 (N_2953,N_2207,N_2381);
nand U2954 (N_2954,N_2432,N_2017);
and U2955 (N_2955,N_2039,N_2017);
or U2956 (N_2956,N_2198,N_2092);
nor U2957 (N_2957,N_2416,N_2205);
xor U2958 (N_2958,N_2357,N_2404);
or U2959 (N_2959,N_2403,N_2099);
and U2960 (N_2960,N_2396,N_2165);
and U2961 (N_2961,N_2146,N_2065);
or U2962 (N_2962,N_2131,N_2190);
xor U2963 (N_2963,N_2302,N_2393);
nor U2964 (N_2964,N_2489,N_2213);
nand U2965 (N_2965,N_2288,N_2246);
and U2966 (N_2966,N_2311,N_2412);
and U2967 (N_2967,N_2258,N_2126);
xor U2968 (N_2968,N_2246,N_2147);
and U2969 (N_2969,N_2083,N_2498);
xnor U2970 (N_2970,N_2214,N_2284);
or U2971 (N_2971,N_2068,N_2171);
xor U2972 (N_2972,N_2456,N_2388);
nor U2973 (N_2973,N_2252,N_2207);
nand U2974 (N_2974,N_2457,N_2407);
nand U2975 (N_2975,N_2451,N_2404);
or U2976 (N_2976,N_2224,N_2013);
xor U2977 (N_2977,N_2430,N_2251);
xnor U2978 (N_2978,N_2070,N_2466);
nand U2979 (N_2979,N_2089,N_2366);
or U2980 (N_2980,N_2453,N_2154);
and U2981 (N_2981,N_2271,N_2373);
nand U2982 (N_2982,N_2303,N_2162);
nand U2983 (N_2983,N_2017,N_2477);
and U2984 (N_2984,N_2265,N_2139);
nand U2985 (N_2985,N_2346,N_2089);
nor U2986 (N_2986,N_2077,N_2409);
nor U2987 (N_2987,N_2299,N_2082);
or U2988 (N_2988,N_2369,N_2408);
nor U2989 (N_2989,N_2286,N_2408);
nor U2990 (N_2990,N_2083,N_2462);
nand U2991 (N_2991,N_2299,N_2271);
or U2992 (N_2992,N_2022,N_2199);
nor U2993 (N_2993,N_2336,N_2046);
or U2994 (N_2994,N_2220,N_2087);
xor U2995 (N_2995,N_2285,N_2197);
xor U2996 (N_2996,N_2369,N_2058);
and U2997 (N_2997,N_2153,N_2169);
or U2998 (N_2998,N_2056,N_2269);
xnor U2999 (N_2999,N_2256,N_2401);
nand U3000 (N_3000,N_2640,N_2561);
or U3001 (N_3001,N_2839,N_2618);
xor U3002 (N_3002,N_2546,N_2917);
xor U3003 (N_3003,N_2620,N_2698);
and U3004 (N_3004,N_2852,N_2899);
and U3005 (N_3005,N_2908,N_2876);
xnor U3006 (N_3006,N_2748,N_2619);
nand U3007 (N_3007,N_2763,N_2842);
or U3008 (N_3008,N_2744,N_2802);
xor U3009 (N_3009,N_2527,N_2668);
xor U3010 (N_3010,N_2514,N_2736);
and U3011 (N_3011,N_2952,N_2968);
nor U3012 (N_3012,N_2568,N_2815);
xnor U3013 (N_3013,N_2935,N_2819);
nand U3014 (N_3014,N_2857,N_2879);
nor U3015 (N_3015,N_2881,N_2741);
and U3016 (N_3016,N_2642,N_2782);
nor U3017 (N_3017,N_2673,N_2610);
nand U3018 (N_3018,N_2700,N_2513);
xnor U3019 (N_3019,N_2954,N_2996);
and U3020 (N_3020,N_2577,N_2804);
nor U3021 (N_3021,N_2584,N_2504);
or U3022 (N_3022,N_2755,N_2833);
and U3023 (N_3023,N_2613,N_2501);
and U3024 (N_3024,N_2554,N_2516);
and U3025 (N_3025,N_2779,N_2647);
xnor U3026 (N_3026,N_2608,N_2630);
xor U3027 (N_3027,N_2683,N_2807);
xor U3028 (N_3028,N_2560,N_2578);
xor U3029 (N_3029,N_2787,N_2998);
xor U3030 (N_3030,N_2942,N_2667);
nor U3031 (N_3031,N_2880,N_2924);
nand U3032 (N_3032,N_2706,N_2559);
nand U3033 (N_3033,N_2891,N_2564);
and U3034 (N_3034,N_2987,N_2762);
and U3035 (N_3035,N_2540,N_2874);
xor U3036 (N_3036,N_2712,N_2536);
nor U3037 (N_3037,N_2701,N_2506);
nor U3038 (N_3038,N_2585,N_2720);
nand U3039 (N_3039,N_2580,N_2946);
nand U3040 (N_3040,N_2771,N_2709);
nand U3041 (N_3041,N_2750,N_2971);
and U3042 (N_3042,N_2726,N_2727);
nand U3043 (N_3043,N_2914,N_2983);
or U3044 (N_3044,N_2882,N_2962);
and U3045 (N_3045,N_2566,N_2686);
and U3046 (N_3046,N_2928,N_2558);
and U3047 (N_3047,N_2665,N_2752);
or U3048 (N_3048,N_2733,N_2766);
and U3049 (N_3049,N_2848,N_2943);
nor U3050 (N_3050,N_2838,N_2858);
nand U3051 (N_3051,N_2655,N_2767);
or U3052 (N_3052,N_2718,N_2722);
or U3053 (N_3053,N_2685,N_2747);
xnor U3054 (N_3054,N_2950,N_2934);
nand U3055 (N_3055,N_2575,N_2906);
xnor U3056 (N_3056,N_2789,N_2892);
xor U3057 (N_3057,N_2641,N_2598);
xnor U3058 (N_3058,N_2587,N_2932);
and U3059 (N_3059,N_2522,N_2623);
xnor U3060 (N_3060,N_2825,N_2740);
xnor U3061 (N_3061,N_2590,N_2854);
nand U3062 (N_3062,N_2520,N_2925);
nor U3063 (N_3063,N_2659,N_2860);
nand U3064 (N_3064,N_2688,N_2828);
or U3065 (N_3065,N_2916,N_2936);
or U3066 (N_3066,N_2687,N_2960);
xor U3067 (N_3067,N_2869,N_2864);
or U3068 (N_3068,N_2941,N_2978);
xor U3069 (N_3069,N_2672,N_2897);
and U3070 (N_3070,N_2510,N_2507);
nand U3071 (N_3071,N_2638,N_2657);
xnor U3072 (N_3072,N_2820,N_2915);
xnor U3073 (N_3073,N_2861,N_2565);
xor U3074 (N_3074,N_2602,N_2631);
and U3075 (N_3075,N_2739,N_2617);
nor U3076 (N_3076,N_2840,N_2656);
and U3077 (N_3077,N_2729,N_2624);
and U3078 (N_3078,N_2693,N_2576);
or U3079 (N_3079,N_2644,N_2535);
nor U3080 (N_3080,N_2889,N_2826);
nand U3081 (N_3081,N_2918,N_2518);
nor U3082 (N_3082,N_2877,N_2792);
xnor U3083 (N_3083,N_2749,N_2816);
or U3084 (N_3084,N_2615,N_2818);
nor U3085 (N_3085,N_2591,N_2929);
xnor U3086 (N_3086,N_2531,N_2616);
and U3087 (N_3087,N_2957,N_2886);
nand U3088 (N_3088,N_2949,N_2982);
and U3089 (N_3089,N_2539,N_2588);
nor U3090 (N_3090,N_2719,N_2837);
xor U3091 (N_3091,N_2959,N_2813);
nand U3092 (N_3092,N_2653,N_2545);
nor U3093 (N_3093,N_2601,N_2721);
and U3094 (N_3094,N_2902,N_2808);
nand U3095 (N_3095,N_2734,N_2732);
or U3096 (N_3096,N_2993,N_2984);
and U3097 (N_3097,N_2871,N_2500);
nor U3098 (N_3098,N_2851,N_2776);
and U3099 (N_3099,N_2538,N_2547);
and U3100 (N_3100,N_2937,N_2835);
xnor U3101 (N_3101,N_2788,N_2715);
or U3102 (N_3102,N_2626,N_2800);
or U3103 (N_3103,N_2682,N_2898);
or U3104 (N_3104,N_2745,N_2664);
nand U3105 (N_3105,N_2765,N_2542);
and U3106 (N_3106,N_2955,N_2533);
xor U3107 (N_3107,N_2684,N_2589);
nand U3108 (N_3108,N_2702,N_2853);
xor U3109 (N_3109,N_2903,N_2986);
nor U3110 (N_3110,N_2992,N_2883);
xnor U3111 (N_3111,N_2777,N_2743);
nand U3112 (N_3112,N_2637,N_2723);
xnor U3113 (N_3113,N_2563,N_2592);
and U3114 (N_3114,N_2660,N_2646);
or U3115 (N_3115,N_2738,N_2966);
nand U3116 (N_3116,N_2980,N_2594);
or U3117 (N_3117,N_2870,N_2574);
nand U3118 (N_3118,N_2939,N_2676);
or U3119 (N_3119,N_2969,N_2716);
xnor U3120 (N_3120,N_2856,N_2824);
and U3121 (N_3121,N_2521,N_2911);
and U3122 (N_3122,N_2836,N_2550);
or U3123 (N_3123,N_2849,N_2717);
nor U3124 (N_3124,N_2691,N_2821);
and U3125 (N_3125,N_2570,N_2710);
nand U3126 (N_3126,N_2703,N_2661);
xor U3127 (N_3127,N_2622,N_2629);
xnor U3128 (N_3128,N_2956,N_2525);
or U3129 (N_3129,N_2976,N_2675);
nand U3130 (N_3130,N_2707,N_2549);
and U3131 (N_3131,N_2798,N_2583);
nand U3132 (N_3132,N_2805,N_2769);
or U3133 (N_3133,N_2913,N_2582);
nor U3134 (N_3134,N_2964,N_2784);
or U3135 (N_3135,N_2865,N_2705);
and U3136 (N_3136,N_2600,N_2791);
and U3137 (N_3137,N_2552,N_2599);
nand U3138 (N_3138,N_2669,N_2991);
and U3139 (N_3139,N_2663,N_2572);
xnor U3140 (N_3140,N_2919,N_2519);
nor U3141 (N_3141,N_2888,N_2844);
or U3142 (N_3142,N_2632,N_2938);
or U3143 (N_3143,N_2556,N_2823);
xnor U3144 (N_3144,N_2873,N_2931);
nand U3145 (N_3145,N_2843,N_2887);
nand U3146 (N_3146,N_2772,N_2537);
nand U3147 (N_3147,N_2797,N_2728);
nand U3148 (N_3148,N_2811,N_2628);
nor U3149 (N_3149,N_2730,N_2812);
nand U3150 (N_3150,N_2958,N_2764);
or U3151 (N_3151,N_2773,N_2666);
or U3152 (N_3152,N_2737,N_2746);
nor U3153 (N_3153,N_2786,N_2847);
nor U3154 (N_3154,N_2948,N_2557);
nand U3155 (N_3155,N_2979,N_2544);
nand U3156 (N_3156,N_2759,N_2689);
and U3157 (N_3157,N_2830,N_2529);
nor U3158 (N_3158,N_2785,N_2990);
and U3159 (N_3159,N_2595,N_2562);
and U3160 (N_3160,N_2555,N_2526);
nor U3161 (N_3161,N_2794,N_2947);
xor U3162 (N_3162,N_2581,N_2645);
nor U3163 (N_3163,N_2895,N_2793);
and U3164 (N_3164,N_2944,N_2751);
nor U3165 (N_3165,N_2922,N_2674);
or U3166 (N_3166,N_2963,N_2855);
xor U3167 (N_3167,N_2708,N_2654);
or U3168 (N_3168,N_2995,N_2845);
and U3169 (N_3169,N_2896,N_2970);
nor U3170 (N_3170,N_2981,N_2834);
xor U3171 (N_3171,N_2593,N_2951);
nand U3172 (N_3172,N_2553,N_2977);
or U3173 (N_3173,N_2878,N_2651);
nand U3174 (N_3174,N_2909,N_2997);
nand U3175 (N_3175,N_2502,N_2671);
or U3176 (N_3176,N_2753,N_2774);
xnor U3177 (N_3177,N_2523,N_2639);
nor U3178 (N_3178,N_2863,N_2677);
or U3179 (N_3179,N_2894,N_2534);
xor U3180 (N_3180,N_2912,N_2961);
nor U3181 (N_3181,N_2515,N_2872);
and U3182 (N_3182,N_2757,N_2809);
nor U3183 (N_3183,N_2822,N_2636);
nand U3184 (N_3184,N_2670,N_2758);
nand U3185 (N_3185,N_2890,N_2790);
nand U3186 (N_3186,N_2953,N_2867);
nand U3187 (N_3187,N_2780,N_2796);
or U3188 (N_3188,N_2528,N_2586);
or U3189 (N_3189,N_2678,N_2841);
xor U3190 (N_3190,N_2596,N_2926);
nand U3191 (N_3191,N_2972,N_2868);
xnor U3192 (N_3192,N_2783,N_2754);
and U3193 (N_3193,N_2690,N_2567);
nand U3194 (N_3194,N_2633,N_2885);
or U3195 (N_3195,N_2635,N_2714);
nand U3196 (N_3196,N_2829,N_2781);
or U3197 (N_3197,N_2604,N_2904);
and U3198 (N_3198,N_2974,N_2650);
nand U3199 (N_3199,N_2508,N_2699);
or U3200 (N_3200,N_2579,N_2999);
nor U3201 (N_3201,N_2775,N_2967);
and U3202 (N_3202,N_2761,N_2503);
xor U3203 (N_3203,N_2731,N_2988);
xor U3204 (N_3204,N_2859,N_2512);
xnor U3205 (N_3205,N_2806,N_2921);
nand U3206 (N_3206,N_2910,N_2696);
and U3207 (N_3207,N_2524,N_2994);
nor U3208 (N_3208,N_2692,N_2541);
xnor U3209 (N_3209,N_2985,N_2923);
nor U3210 (N_3210,N_2900,N_2597);
and U3211 (N_3211,N_2517,N_2532);
xnor U3212 (N_3212,N_2905,N_2543);
and U3213 (N_3213,N_2801,N_2573);
nor U3214 (N_3214,N_2846,N_2569);
and U3215 (N_3215,N_2817,N_2827);
xnor U3216 (N_3216,N_2697,N_2606);
xor U3217 (N_3217,N_2933,N_2505);
and U3218 (N_3218,N_2901,N_2866);
xnor U3219 (N_3219,N_2814,N_2658);
or U3220 (N_3220,N_2875,N_2778);
or U3221 (N_3221,N_2530,N_2795);
nor U3222 (N_3222,N_2662,N_2605);
nand U3223 (N_3223,N_2803,N_2649);
nor U3224 (N_3224,N_2679,N_2551);
nor U3225 (N_3225,N_2725,N_2975);
xnor U3226 (N_3226,N_2832,N_2884);
nand U3227 (N_3227,N_2634,N_2627);
nor U3228 (N_3228,N_2927,N_2607);
or U3229 (N_3229,N_2648,N_2965);
xor U3230 (N_3230,N_2989,N_2930);
xnor U3231 (N_3231,N_2940,N_2509);
nand U3232 (N_3232,N_2694,N_2681);
or U3233 (N_3233,N_2511,N_2862);
nand U3234 (N_3234,N_2643,N_2614);
and U3235 (N_3235,N_2711,N_2742);
nor U3236 (N_3236,N_2611,N_2621);
and U3237 (N_3237,N_2735,N_2548);
or U3238 (N_3238,N_2652,N_2893);
nand U3239 (N_3239,N_2612,N_2907);
and U3240 (N_3240,N_2850,N_2973);
or U3241 (N_3241,N_2713,N_2704);
and U3242 (N_3242,N_2945,N_2680);
xnor U3243 (N_3243,N_2603,N_2770);
nor U3244 (N_3244,N_2920,N_2625);
xnor U3245 (N_3245,N_2831,N_2609);
xor U3246 (N_3246,N_2571,N_2799);
nand U3247 (N_3247,N_2756,N_2724);
or U3248 (N_3248,N_2760,N_2810);
xor U3249 (N_3249,N_2695,N_2768);
nand U3250 (N_3250,N_2943,N_2665);
nor U3251 (N_3251,N_2628,N_2977);
nor U3252 (N_3252,N_2796,N_2684);
or U3253 (N_3253,N_2789,N_2915);
and U3254 (N_3254,N_2544,N_2557);
nand U3255 (N_3255,N_2944,N_2971);
and U3256 (N_3256,N_2968,N_2551);
and U3257 (N_3257,N_2573,N_2551);
nand U3258 (N_3258,N_2691,N_2618);
xor U3259 (N_3259,N_2884,N_2654);
and U3260 (N_3260,N_2719,N_2988);
xor U3261 (N_3261,N_2549,N_2862);
nor U3262 (N_3262,N_2619,N_2638);
xnor U3263 (N_3263,N_2803,N_2597);
or U3264 (N_3264,N_2519,N_2545);
nor U3265 (N_3265,N_2974,N_2915);
nand U3266 (N_3266,N_2764,N_2983);
nor U3267 (N_3267,N_2918,N_2899);
xnor U3268 (N_3268,N_2741,N_2676);
nand U3269 (N_3269,N_2699,N_2812);
or U3270 (N_3270,N_2672,N_2583);
nor U3271 (N_3271,N_2545,N_2901);
xor U3272 (N_3272,N_2997,N_2769);
xnor U3273 (N_3273,N_2878,N_2772);
nor U3274 (N_3274,N_2694,N_2691);
or U3275 (N_3275,N_2623,N_2779);
nor U3276 (N_3276,N_2540,N_2904);
or U3277 (N_3277,N_2914,N_2845);
nor U3278 (N_3278,N_2599,N_2672);
and U3279 (N_3279,N_2795,N_2838);
nor U3280 (N_3280,N_2840,N_2977);
and U3281 (N_3281,N_2812,N_2957);
xor U3282 (N_3282,N_2547,N_2596);
and U3283 (N_3283,N_2886,N_2775);
and U3284 (N_3284,N_2810,N_2568);
nand U3285 (N_3285,N_2818,N_2577);
and U3286 (N_3286,N_2540,N_2650);
nand U3287 (N_3287,N_2931,N_2944);
nand U3288 (N_3288,N_2665,N_2813);
nor U3289 (N_3289,N_2739,N_2660);
nand U3290 (N_3290,N_2588,N_2938);
and U3291 (N_3291,N_2696,N_2928);
nand U3292 (N_3292,N_2595,N_2997);
xnor U3293 (N_3293,N_2971,N_2602);
or U3294 (N_3294,N_2749,N_2881);
or U3295 (N_3295,N_2938,N_2929);
nand U3296 (N_3296,N_2778,N_2733);
nand U3297 (N_3297,N_2640,N_2923);
xnor U3298 (N_3298,N_2784,N_2513);
xnor U3299 (N_3299,N_2807,N_2556);
nand U3300 (N_3300,N_2540,N_2960);
nand U3301 (N_3301,N_2618,N_2689);
nand U3302 (N_3302,N_2659,N_2832);
and U3303 (N_3303,N_2892,N_2632);
nor U3304 (N_3304,N_2797,N_2868);
nor U3305 (N_3305,N_2503,N_2722);
and U3306 (N_3306,N_2557,N_2928);
and U3307 (N_3307,N_2676,N_2589);
nor U3308 (N_3308,N_2534,N_2797);
xnor U3309 (N_3309,N_2759,N_2573);
nor U3310 (N_3310,N_2562,N_2614);
nand U3311 (N_3311,N_2760,N_2512);
xor U3312 (N_3312,N_2691,N_2852);
nand U3313 (N_3313,N_2651,N_2580);
and U3314 (N_3314,N_2584,N_2913);
and U3315 (N_3315,N_2643,N_2952);
nand U3316 (N_3316,N_2540,N_2796);
nor U3317 (N_3317,N_2884,N_2883);
xnor U3318 (N_3318,N_2740,N_2653);
or U3319 (N_3319,N_2680,N_2517);
nand U3320 (N_3320,N_2845,N_2896);
and U3321 (N_3321,N_2831,N_2723);
nand U3322 (N_3322,N_2759,N_2882);
nand U3323 (N_3323,N_2771,N_2910);
or U3324 (N_3324,N_2864,N_2632);
nor U3325 (N_3325,N_2732,N_2547);
and U3326 (N_3326,N_2897,N_2934);
nor U3327 (N_3327,N_2956,N_2734);
xnor U3328 (N_3328,N_2917,N_2762);
and U3329 (N_3329,N_2859,N_2692);
xnor U3330 (N_3330,N_2679,N_2824);
nand U3331 (N_3331,N_2903,N_2656);
or U3332 (N_3332,N_2981,N_2936);
nor U3333 (N_3333,N_2747,N_2882);
nor U3334 (N_3334,N_2574,N_2721);
or U3335 (N_3335,N_2528,N_2623);
or U3336 (N_3336,N_2767,N_2675);
nor U3337 (N_3337,N_2893,N_2900);
or U3338 (N_3338,N_2665,N_2737);
nor U3339 (N_3339,N_2525,N_2819);
nor U3340 (N_3340,N_2725,N_2963);
and U3341 (N_3341,N_2774,N_2640);
and U3342 (N_3342,N_2620,N_2548);
xnor U3343 (N_3343,N_2989,N_2540);
and U3344 (N_3344,N_2698,N_2623);
nor U3345 (N_3345,N_2667,N_2715);
or U3346 (N_3346,N_2672,N_2989);
and U3347 (N_3347,N_2976,N_2794);
and U3348 (N_3348,N_2963,N_2783);
xor U3349 (N_3349,N_2980,N_2884);
nand U3350 (N_3350,N_2616,N_2896);
nand U3351 (N_3351,N_2770,N_2586);
and U3352 (N_3352,N_2730,N_2814);
nor U3353 (N_3353,N_2721,N_2749);
nor U3354 (N_3354,N_2998,N_2751);
and U3355 (N_3355,N_2697,N_2532);
and U3356 (N_3356,N_2860,N_2945);
and U3357 (N_3357,N_2694,N_2577);
and U3358 (N_3358,N_2529,N_2581);
xnor U3359 (N_3359,N_2661,N_2898);
and U3360 (N_3360,N_2996,N_2960);
and U3361 (N_3361,N_2567,N_2529);
nor U3362 (N_3362,N_2695,N_2512);
and U3363 (N_3363,N_2966,N_2840);
nor U3364 (N_3364,N_2800,N_2525);
nor U3365 (N_3365,N_2833,N_2968);
xnor U3366 (N_3366,N_2987,N_2771);
or U3367 (N_3367,N_2758,N_2652);
and U3368 (N_3368,N_2805,N_2707);
and U3369 (N_3369,N_2610,N_2884);
xor U3370 (N_3370,N_2801,N_2969);
nor U3371 (N_3371,N_2520,N_2613);
nand U3372 (N_3372,N_2802,N_2970);
nor U3373 (N_3373,N_2851,N_2828);
nand U3374 (N_3374,N_2922,N_2819);
xnor U3375 (N_3375,N_2790,N_2758);
nor U3376 (N_3376,N_2718,N_2697);
and U3377 (N_3377,N_2669,N_2846);
or U3378 (N_3378,N_2760,N_2957);
nor U3379 (N_3379,N_2665,N_2942);
nor U3380 (N_3380,N_2826,N_2876);
xor U3381 (N_3381,N_2615,N_2786);
xnor U3382 (N_3382,N_2829,N_2635);
nor U3383 (N_3383,N_2728,N_2735);
and U3384 (N_3384,N_2509,N_2618);
xor U3385 (N_3385,N_2967,N_2746);
nor U3386 (N_3386,N_2573,N_2863);
nand U3387 (N_3387,N_2545,N_2840);
nor U3388 (N_3388,N_2719,N_2738);
xnor U3389 (N_3389,N_2942,N_2557);
and U3390 (N_3390,N_2997,N_2958);
or U3391 (N_3391,N_2651,N_2674);
and U3392 (N_3392,N_2672,N_2960);
xnor U3393 (N_3393,N_2574,N_2707);
nand U3394 (N_3394,N_2818,N_2819);
or U3395 (N_3395,N_2834,N_2924);
nand U3396 (N_3396,N_2687,N_2883);
nor U3397 (N_3397,N_2670,N_2937);
xnor U3398 (N_3398,N_2762,N_2555);
and U3399 (N_3399,N_2878,N_2779);
or U3400 (N_3400,N_2986,N_2724);
nand U3401 (N_3401,N_2639,N_2648);
nand U3402 (N_3402,N_2721,N_2850);
or U3403 (N_3403,N_2957,N_2775);
nor U3404 (N_3404,N_2774,N_2854);
xnor U3405 (N_3405,N_2682,N_2779);
or U3406 (N_3406,N_2755,N_2993);
and U3407 (N_3407,N_2642,N_2841);
and U3408 (N_3408,N_2550,N_2645);
and U3409 (N_3409,N_2615,N_2503);
xnor U3410 (N_3410,N_2889,N_2588);
nand U3411 (N_3411,N_2711,N_2688);
nor U3412 (N_3412,N_2581,N_2552);
and U3413 (N_3413,N_2947,N_2879);
nor U3414 (N_3414,N_2942,N_2642);
xnor U3415 (N_3415,N_2503,N_2594);
xnor U3416 (N_3416,N_2811,N_2502);
or U3417 (N_3417,N_2572,N_2617);
xor U3418 (N_3418,N_2732,N_2747);
nor U3419 (N_3419,N_2842,N_2520);
nor U3420 (N_3420,N_2758,N_2732);
xnor U3421 (N_3421,N_2771,N_2666);
xor U3422 (N_3422,N_2602,N_2997);
and U3423 (N_3423,N_2519,N_2998);
and U3424 (N_3424,N_2551,N_2630);
nand U3425 (N_3425,N_2961,N_2965);
xnor U3426 (N_3426,N_2677,N_2695);
nand U3427 (N_3427,N_2564,N_2859);
nand U3428 (N_3428,N_2691,N_2877);
or U3429 (N_3429,N_2882,N_2874);
xnor U3430 (N_3430,N_2601,N_2725);
nor U3431 (N_3431,N_2558,N_2986);
nand U3432 (N_3432,N_2693,N_2615);
xor U3433 (N_3433,N_2557,N_2589);
and U3434 (N_3434,N_2755,N_2554);
xor U3435 (N_3435,N_2723,N_2898);
and U3436 (N_3436,N_2748,N_2917);
nand U3437 (N_3437,N_2922,N_2779);
or U3438 (N_3438,N_2881,N_2893);
nand U3439 (N_3439,N_2701,N_2521);
xnor U3440 (N_3440,N_2616,N_2708);
or U3441 (N_3441,N_2683,N_2535);
nand U3442 (N_3442,N_2985,N_2676);
nand U3443 (N_3443,N_2555,N_2644);
nand U3444 (N_3444,N_2871,N_2649);
nand U3445 (N_3445,N_2753,N_2958);
xor U3446 (N_3446,N_2599,N_2681);
and U3447 (N_3447,N_2917,N_2622);
or U3448 (N_3448,N_2729,N_2875);
nand U3449 (N_3449,N_2887,N_2836);
xnor U3450 (N_3450,N_2614,N_2730);
xnor U3451 (N_3451,N_2788,N_2512);
or U3452 (N_3452,N_2937,N_2940);
and U3453 (N_3453,N_2620,N_2941);
or U3454 (N_3454,N_2987,N_2578);
or U3455 (N_3455,N_2857,N_2635);
and U3456 (N_3456,N_2602,N_2810);
and U3457 (N_3457,N_2754,N_2893);
and U3458 (N_3458,N_2730,N_2746);
nand U3459 (N_3459,N_2658,N_2936);
nand U3460 (N_3460,N_2629,N_2521);
or U3461 (N_3461,N_2629,N_2632);
or U3462 (N_3462,N_2677,N_2681);
and U3463 (N_3463,N_2806,N_2514);
nand U3464 (N_3464,N_2868,N_2788);
and U3465 (N_3465,N_2773,N_2921);
or U3466 (N_3466,N_2861,N_2825);
xnor U3467 (N_3467,N_2863,N_2682);
and U3468 (N_3468,N_2895,N_2745);
and U3469 (N_3469,N_2792,N_2924);
nor U3470 (N_3470,N_2899,N_2792);
and U3471 (N_3471,N_2654,N_2548);
nor U3472 (N_3472,N_2920,N_2610);
nor U3473 (N_3473,N_2965,N_2952);
nor U3474 (N_3474,N_2843,N_2757);
xor U3475 (N_3475,N_2745,N_2562);
nand U3476 (N_3476,N_2543,N_2652);
and U3477 (N_3477,N_2998,N_2563);
and U3478 (N_3478,N_2621,N_2688);
nand U3479 (N_3479,N_2629,N_2839);
nor U3480 (N_3480,N_2640,N_2703);
nand U3481 (N_3481,N_2533,N_2826);
and U3482 (N_3482,N_2781,N_2511);
nor U3483 (N_3483,N_2956,N_2630);
or U3484 (N_3484,N_2926,N_2552);
or U3485 (N_3485,N_2831,N_2980);
xor U3486 (N_3486,N_2907,N_2552);
or U3487 (N_3487,N_2665,N_2572);
and U3488 (N_3488,N_2640,N_2747);
and U3489 (N_3489,N_2796,N_2794);
or U3490 (N_3490,N_2610,N_2972);
or U3491 (N_3491,N_2811,N_2669);
and U3492 (N_3492,N_2693,N_2605);
xnor U3493 (N_3493,N_2982,N_2557);
or U3494 (N_3494,N_2548,N_2631);
and U3495 (N_3495,N_2757,N_2621);
nand U3496 (N_3496,N_2967,N_2841);
and U3497 (N_3497,N_2660,N_2778);
xnor U3498 (N_3498,N_2942,N_2539);
nand U3499 (N_3499,N_2842,N_2798);
and U3500 (N_3500,N_3309,N_3216);
or U3501 (N_3501,N_3006,N_3413);
and U3502 (N_3502,N_3240,N_3063);
nor U3503 (N_3503,N_3139,N_3062);
xnor U3504 (N_3504,N_3339,N_3440);
nand U3505 (N_3505,N_3369,N_3221);
or U3506 (N_3506,N_3347,N_3175);
xor U3507 (N_3507,N_3422,N_3459);
and U3508 (N_3508,N_3325,N_3072);
and U3509 (N_3509,N_3106,N_3035);
nand U3510 (N_3510,N_3020,N_3454);
or U3511 (N_3511,N_3248,N_3478);
and U3512 (N_3512,N_3277,N_3428);
nor U3513 (N_3513,N_3322,N_3361);
nand U3514 (N_3514,N_3242,N_3222);
xnor U3515 (N_3515,N_3269,N_3409);
or U3516 (N_3516,N_3193,N_3400);
or U3517 (N_3517,N_3229,N_3115);
nor U3518 (N_3518,N_3273,N_3394);
or U3519 (N_3519,N_3281,N_3226);
and U3520 (N_3520,N_3436,N_3206);
nor U3521 (N_3521,N_3233,N_3066);
nor U3522 (N_3522,N_3252,N_3326);
nand U3523 (N_3523,N_3195,N_3251);
nand U3524 (N_3524,N_3159,N_3158);
and U3525 (N_3525,N_3052,N_3191);
and U3526 (N_3526,N_3174,N_3276);
nand U3527 (N_3527,N_3462,N_3310);
nand U3528 (N_3528,N_3275,N_3085);
nand U3529 (N_3529,N_3403,N_3232);
nor U3530 (N_3530,N_3099,N_3386);
and U3531 (N_3531,N_3262,N_3101);
nand U3532 (N_3532,N_3435,N_3384);
xor U3533 (N_3533,N_3096,N_3170);
or U3534 (N_3534,N_3288,N_3267);
nor U3535 (N_3535,N_3113,N_3107);
nand U3536 (N_3536,N_3340,N_3258);
and U3537 (N_3537,N_3134,N_3357);
nand U3538 (N_3538,N_3137,N_3283);
xnor U3539 (N_3539,N_3482,N_3306);
nand U3540 (N_3540,N_3376,N_3131);
xor U3541 (N_3541,N_3238,N_3272);
xnor U3542 (N_3542,N_3122,N_3045);
and U3543 (N_3543,N_3025,N_3304);
xor U3544 (N_3544,N_3261,N_3093);
or U3545 (N_3545,N_3246,N_3147);
xor U3546 (N_3546,N_3321,N_3341);
nand U3547 (N_3547,N_3254,N_3377);
nor U3548 (N_3548,N_3203,N_3498);
nand U3549 (N_3549,N_3161,N_3287);
and U3550 (N_3550,N_3036,N_3418);
xnor U3551 (N_3551,N_3234,N_3366);
and U3552 (N_3552,N_3471,N_3406);
nand U3553 (N_3553,N_3064,N_3007);
or U3554 (N_3554,N_3235,N_3073);
xnor U3555 (N_3555,N_3399,N_3424);
and U3556 (N_3556,N_3303,N_3396);
or U3557 (N_3557,N_3003,N_3458);
and U3558 (N_3558,N_3358,N_3049);
or U3559 (N_3559,N_3327,N_3383);
and U3560 (N_3560,N_3059,N_3415);
and U3561 (N_3561,N_3264,N_3176);
or U3562 (N_3562,N_3363,N_3278);
nand U3563 (N_3563,N_3497,N_3213);
nand U3564 (N_3564,N_3127,N_3390);
nor U3565 (N_3565,N_3129,N_3402);
or U3566 (N_3566,N_3453,N_3004);
xnor U3567 (N_3567,N_3494,N_3198);
xor U3568 (N_3568,N_3112,N_3372);
and U3569 (N_3569,N_3490,N_3123);
nor U3570 (N_3570,N_3177,N_3168);
or U3571 (N_3571,N_3336,N_3393);
and U3572 (N_3572,N_3154,N_3451);
and U3573 (N_3573,N_3316,N_3280);
nor U3574 (N_3574,N_3499,N_3016);
nor U3575 (N_3575,N_3183,N_3128);
nor U3576 (N_3576,N_3373,N_3274);
or U3577 (N_3577,N_3169,N_3408);
nand U3578 (N_3578,N_3010,N_3385);
nor U3579 (N_3579,N_3181,N_3148);
nor U3580 (N_3580,N_3443,N_3038);
or U3581 (N_3581,N_3362,N_3382);
nor U3582 (N_3582,N_3136,N_3097);
or U3583 (N_3583,N_3445,N_3476);
xor U3584 (N_3584,N_3294,N_3268);
nand U3585 (N_3585,N_3237,N_3381);
nor U3586 (N_3586,N_3412,N_3313);
nor U3587 (N_3587,N_3114,N_3450);
and U3588 (N_3588,N_3444,N_3255);
nand U3589 (N_3589,N_3223,N_3087);
nor U3590 (N_3590,N_3411,N_3111);
nand U3591 (N_3591,N_3431,N_3419);
and U3592 (N_3592,N_3084,N_3370);
nor U3593 (N_3593,N_3051,N_3473);
nor U3594 (N_3594,N_3485,N_3282);
nand U3595 (N_3595,N_3076,N_3256);
or U3596 (N_3596,N_3236,N_3315);
nor U3597 (N_3597,N_3120,N_3050);
nand U3598 (N_3598,N_3253,N_3184);
or U3599 (N_3599,N_3019,N_3296);
and U3600 (N_3600,N_3047,N_3104);
nor U3601 (N_3601,N_3259,N_3053);
and U3602 (N_3602,N_3068,N_3230);
nor U3603 (N_3603,N_3439,N_3109);
xnor U3604 (N_3604,N_3164,N_3022);
xor U3605 (N_3605,N_3032,N_3046);
nand U3606 (N_3606,N_3429,N_3119);
and U3607 (N_3607,N_3080,N_3351);
xnor U3608 (N_3608,N_3426,N_3352);
nor U3609 (N_3609,N_3065,N_3416);
or U3610 (N_3610,N_3292,N_3491);
and U3611 (N_3611,N_3151,N_3487);
nand U3612 (N_3612,N_3000,N_3009);
nor U3613 (N_3613,N_3031,N_3495);
or U3614 (N_3614,N_3225,N_3037);
xnor U3615 (N_3615,N_3266,N_3295);
or U3616 (N_3616,N_3214,N_3124);
or U3617 (N_3617,N_3157,N_3026);
nand U3618 (N_3618,N_3320,N_3130);
xnor U3619 (N_3619,N_3297,N_3056);
and U3620 (N_3620,N_3388,N_3121);
nor U3621 (N_3621,N_3318,N_3142);
or U3622 (N_3622,N_3089,N_3227);
nor U3623 (N_3623,N_3263,N_3024);
nor U3624 (N_3624,N_3293,N_3144);
and U3625 (N_3625,N_3395,N_3241);
nor U3626 (N_3626,N_3329,N_3029);
xor U3627 (N_3627,N_3167,N_3185);
or U3628 (N_3628,N_3260,N_3171);
nor U3629 (N_3629,N_3102,N_3162);
nand U3630 (N_3630,N_3082,N_3015);
nor U3631 (N_3631,N_3011,N_3461);
nand U3632 (N_3632,N_3021,N_3217);
or U3633 (N_3633,N_3442,N_3243);
or U3634 (N_3634,N_3455,N_3150);
nor U3635 (N_3635,N_3166,N_3464);
or U3636 (N_3636,N_3218,N_3480);
xnor U3637 (N_3637,N_3279,N_3077);
or U3638 (N_3638,N_3187,N_3173);
or U3639 (N_3639,N_3379,N_3034);
nand U3640 (N_3640,N_3360,N_3474);
and U3641 (N_3641,N_3012,N_3135);
xnor U3642 (N_3642,N_3039,N_3219);
xor U3643 (N_3643,N_3014,N_3335);
or U3644 (N_3644,N_3190,N_3378);
xnor U3645 (N_3645,N_3479,N_3330);
or U3646 (N_3646,N_3323,N_3488);
nor U3647 (N_3647,N_3027,N_3475);
nor U3648 (N_3648,N_3465,N_3483);
nor U3649 (N_3649,N_3116,N_3407);
xor U3650 (N_3650,N_3250,N_3205);
xnor U3651 (N_3651,N_3457,N_3346);
xor U3652 (N_3652,N_3186,N_3091);
and U3653 (N_3653,N_3391,N_3138);
or U3654 (N_3654,N_3040,N_3299);
or U3655 (N_3655,N_3493,N_3140);
or U3656 (N_3656,N_3289,N_3300);
and U3657 (N_3657,N_3095,N_3212);
xnor U3658 (N_3658,N_3334,N_3333);
xor U3659 (N_3659,N_3331,N_3470);
nor U3660 (N_3660,N_3069,N_3200);
nor U3661 (N_3661,N_3404,N_3133);
and U3662 (N_3662,N_3055,N_3197);
nand U3663 (N_3663,N_3005,N_3088);
and U3664 (N_3664,N_3108,N_3496);
nand U3665 (N_3665,N_3152,N_3146);
nor U3666 (N_3666,N_3286,N_3305);
nor U3667 (N_3667,N_3054,N_3489);
nor U3668 (N_3668,N_3302,N_3224);
or U3669 (N_3669,N_3145,N_3466);
nand U3670 (N_3670,N_3434,N_3110);
xnor U3671 (N_3671,N_3058,N_3410);
or U3672 (N_3672,N_3201,N_3387);
nor U3673 (N_3673,N_3210,N_3421);
or U3674 (N_3674,N_3013,N_3389);
nor U3675 (N_3675,N_3332,N_3452);
or U3676 (N_3676,N_3239,N_3172);
xor U3677 (N_3677,N_3312,N_3420);
xor U3678 (N_3678,N_3002,N_3156);
nand U3679 (N_3679,N_3486,N_3061);
and U3680 (N_3680,N_3375,N_3467);
xor U3681 (N_3681,N_3118,N_3083);
or U3682 (N_3682,N_3060,N_3074);
and U3683 (N_3683,N_3041,N_3270);
and U3684 (N_3684,N_3290,N_3057);
nor U3685 (N_3685,N_3367,N_3307);
nand U3686 (N_3686,N_3477,N_3423);
nand U3687 (N_3687,N_3165,N_3067);
nor U3688 (N_3688,N_3414,N_3392);
xnor U3689 (N_3689,N_3196,N_3257);
xor U3690 (N_3690,N_3456,N_3079);
nor U3691 (N_3691,N_3324,N_3033);
and U3692 (N_3692,N_3208,N_3207);
and U3693 (N_3693,N_3141,N_3163);
or U3694 (N_3694,N_3350,N_3018);
nand U3695 (N_3695,N_3188,N_3160);
nand U3696 (N_3696,N_3228,N_3398);
nor U3697 (N_3697,N_3215,N_3365);
nand U3698 (N_3698,N_3460,N_3349);
or U3699 (N_3699,N_3245,N_3468);
and U3700 (N_3700,N_3086,N_3364);
and U3701 (N_3701,N_3182,N_3244);
nor U3702 (N_3702,N_3092,N_3204);
and U3703 (N_3703,N_3356,N_3094);
and U3704 (N_3704,N_3126,N_3354);
xor U3705 (N_3705,N_3078,N_3001);
nor U3706 (N_3706,N_3317,N_3397);
nor U3707 (N_3707,N_3328,N_3202);
nor U3708 (N_3708,N_3343,N_3374);
nor U3709 (N_3709,N_3359,N_3132);
xor U3710 (N_3710,N_3192,N_3153);
or U3711 (N_3711,N_3355,N_3023);
xnor U3712 (N_3712,N_3425,N_3117);
nand U3713 (N_3713,N_3211,N_3143);
or U3714 (N_3714,N_3247,N_3070);
or U3715 (N_3715,N_3199,N_3189);
nand U3716 (N_3716,N_3265,N_3401);
and U3717 (N_3717,N_3337,N_3433);
nand U3718 (N_3718,N_3342,N_3030);
xnor U3719 (N_3719,N_3285,N_3220);
nand U3720 (N_3720,N_3231,N_3371);
xor U3721 (N_3721,N_3448,N_3492);
xnor U3722 (N_3722,N_3284,N_3180);
and U3723 (N_3723,N_3155,N_3463);
and U3724 (N_3724,N_3353,N_3071);
or U3725 (N_3725,N_3469,N_3311);
xor U3726 (N_3726,N_3017,N_3048);
nand U3727 (N_3727,N_3446,N_3209);
nand U3728 (N_3728,N_3380,N_3432);
nand U3729 (N_3729,N_3178,N_3249);
and U3730 (N_3730,N_3368,N_3417);
or U3731 (N_3731,N_3298,N_3100);
xnor U3732 (N_3732,N_3179,N_3427);
nor U3733 (N_3733,N_3271,N_3044);
xnor U3734 (N_3734,N_3090,N_3314);
nor U3735 (N_3735,N_3344,N_3125);
or U3736 (N_3736,N_3438,N_3308);
nand U3737 (N_3737,N_3441,N_3042);
nor U3738 (N_3738,N_3405,N_3472);
xor U3739 (N_3739,N_3345,N_3301);
or U3740 (N_3740,N_3437,N_3103);
xor U3741 (N_3741,N_3481,N_3075);
nand U3742 (N_3742,N_3447,N_3449);
nor U3743 (N_3743,N_3430,N_3081);
nand U3744 (N_3744,N_3149,N_3338);
nor U3745 (N_3745,N_3348,N_3291);
and U3746 (N_3746,N_3484,N_3319);
or U3747 (N_3747,N_3105,N_3194);
nor U3748 (N_3748,N_3028,N_3043);
nand U3749 (N_3749,N_3098,N_3008);
and U3750 (N_3750,N_3366,N_3170);
nand U3751 (N_3751,N_3053,N_3383);
or U3752 (N_3752,N_3409,N_3372);
or U3753 (N_3753,N_3078,N_3461);
xnor U3754 (N_3754,N_3420,N_3104);
or U3755 (N_3755,N_3471,N_3205);
and U3756 (N_3756,N_3195,N_3220);
and U3757 (N_3757,N_3296,N_3120);
nand U3758 (N_3758,N_3014,N_3197);
and U3759 (N_3759,N_3118,N_3452);
or U3760 (N_3760,N_3193,N_3275);
xor U3761 (N_3761,N_3432,N_3315);
xnor U3762 (N_3762,N_3079,N_3441);
nand U3763 (N_3763,N_3240,N_3238);
or U3764 (N_3764,N_3182,N_3365);
nor U3765 (N_3765,N_3345,N_3381);
or U3766 (N_3766,N_3309,N_3370);
nand U3767 (N_3767,N_3350,N_3242);
nor U3768 (N_3768,N_3299,N_3317);
or U3769 (N_3769,N_3139,N_3436);
nor U3770 (N_3770,N_3409,N_3468);
and U3771 (N_3771,N_3192,N_3187);
or U3772 (N_3772,N_3481,N_3430);
and U3773 (N_3773,N_3293,N_3465);
or U3774 (N_3774,N_3466,N_3199);
or U3775 (N_3775,N_3451,N_3481);
xnor U3776 (N_3776,N_3457,N_3198);
nor U3777 (N_3777,N_3431,N_3234);
and U3778 (N_3778,N_3411,N_3019);
or U3779 (N_3779,N_3195,N_3078);
nor U3780 (N_3780,N_3134,N_3442);
or U3781 (N_3781,N_3215,N_3320);
nand U3782 (N_3782,N_3338,N_3470);
xnor U3783 (N_3783,N_3421,N_3147);
nand U3784 (N_3784,N_3056,N_3122);
xnor U3785 (N_3785,N_3455,N_3448);
xnor U3786 (N_3786,N_3106,N_3254);
nor U3787 (N_3787,N_3180,N_3351);
xor U3788 (N_3788,N_3303,N_3004);
nand U3789 (N_3789,N_3180,N_3039);
nor U3790 (N_3790,N_3329,N_3281);
nand U3791 (N_3791,N_3229,N_3379);
xor U3792 (N_3792,N_3003,N_3152);
nand U3793 (N_3793,N_3337,N_3368);
and U3794 (N_3794,N_3064,N_3214);
and U3795 (N_3795,N_3277,N_3409);
nand U3796 (N_3796,N_3346,N_3302);
nor U3797 (N_3797,N_3489,N_3388);
and U3798 (N_3798,N_3252,N_3223);
and U3799 (N_3799,N_3307,N_3132);
or U3800 (N_3800,N_3488,N_3389);
or U3801 (N_3801,N_3383,N_3221);
xnor U3802 (N_3802,N_3246,N_3090);
or U3803 (N_3803,N_3094,N_3449);
and U3804 (N_3804,N_3298,N_3188);
nand U3805 (N_3805,N_3380,N_3262);
nand U3806 (N_3806,N_3216,N_3193);
and U3807 (N_3807,N_3233,N_3111);
and U3808 (N_3808,N_3262,N_3076);
and U3809 (N_3809,N_3118,N_3156);
and U3810 (N_3810,N_3079,N_3476);
or U3811 (N_3811,N_3468,N_3097);
nand U3812 (N_3812,N_3499,N_3141);
nor U3813 (N_3813,N_3398,N_3084);
and U3814 (N_3814,N_3185,N_3420);
nand U3815 (N_3815,N_3211,N_3324);
or U3816 (N_3816,N_3246,N_3164);
nor U3817 (N_3817,N_3025,N_3195);
or U3818 (N_3818,N_3402,N_3218);
nand U3819 (N_3819,N_3268,N_3014);
xnor U3820 (N_3820,N_3063,N_3248);
xor U3821 (N_3821,N_3021,N_3202);
nand U3822 (N_3822,N_3296,N_3331);
nor U3823 (N_3823,N_3049,N_3475);
and U3824 (N_3824,N_3355,N_3178);
nand U3825 (N_3825,N_3367,N_3293);
nand U3826 (N_3826,N_3209,N_3399);
xnor U3827 (N_3827,N_3053,N_3003);
xnor U3828 (N_3828,N_3356,N_3478);
xor U3829 (N_3829,N_3099,N_3415);
nor U3830 (N_3830,N_3133,N_3330);
nand U3831 (N_3831,N_3010,N_3381);
and U3832 (N_3832,N_3320,N_3136);
and U3833 (N_3833,N_3120,N_3045);
or U3834 (N_3834,N_3220,N_3191);
xor U3835 (N_3835,N_3174,N_3141);
and U3836 (N_3836,N_3245,N_3102);
nor U3837 (N_3837,N_3034,N_3406);
nor U3838 (N_3838,N_3460,N_3404);
or U3839 (N_3839,N_3086,N_3262);
nand U3840 (N_3840,N_3410,N_3010);
nand U3841 (N_3841,N_3017,N_3397);
nor U3842 (N_3842,N_3267,N_3033);
nor U3843 (N_3843,N_3496,N_3287);
nand U3844 (N_3844,N_3209,N_3122);
xor U3845 (N_3845,N_3394,N_3012);
xor U3846 (N_3846,N_3408,N_3085);
and U3847 (N_3847,N_3228,N_3035);
and U3848 (N_3848,N_3112,N_3463);
or U3849 (N_3849,N_3088,N_3294);
nand U3850 (N_3850,N_3463,N_3021);
xor U3851 (N_3851,N_3446,N_3447);
nand U3852 (N_3852,N_3055,N_3136);
nand U3853 (N_3853,N_3280,N_3021);
and U3854 (N_3854,N_3241,N_3433);
xnor U3855 (N_3855,N_3444,N_3376);
nand U3856 (N_3856,N_3312,N_3337);
and U3857 (N_3857,N_3338,N_3148);
nand U3858 (N_3858,N_3232,N_3197);
nor U3859 (N_3859,N_3469,N_3112);
xor U3860 (N_3860,N_3184,N_3114);
nor U3861 (N_3861,N_3003,N_3325);
xor U3862 (N_3862,N_3189,N_3142);
nor U3863 (N_3863,N_3072,N_3175);
and U3864 (N_3864,N_3098,N_3417);
or U3865 (N_3865,N_3443,N_3272);
xor U3866 (N_3866,N_3229,N_3064);
and U3867 (N_3867,N_3438,N_3006);
nor U3868 (N_3868,N_3460,N_3137);
nand U3869 (N_3869,N_3240,N_3408);
and U3870 (N_3870,N_3093,N_3258);
nor U3871 (N_3871,N_3401,N_3055);
xor U3872 (N_3872,N_3315,N_3074);
xnor U3873 (N_3873,N_3411,N_3029);
xnor U3874 (N_3874,N_3310,N_3212);
nand U3875 (N_3875,N_3360,N_3077);
xor U3876 (N_3876,N_3268,N_3187);
and U3877 (N_3877,N_3155,N_3058);
nand U3878 (N_3878,N_3429,N_3445);
and U3879 (N_3879,N_3019,N_3034);
or U3880 (N_3880,N_3022,N_3292);
or U3881 (N_3881,N_3205,N_3299);
nor U3882 (N_3882,N_3201,N_3284);
xor U3883 (N_3883,N_3389,N_3045);
xnor U3884 (N_3884,N_3282,N_3280);
xor U3885 (N_3885,N_3154,N_3322);
or U3886 (N_3886,N_3282,N_3456);
xnor U3887 (N_3887,N_3398,N_3140);
and U3888 (N_3888,N_3346,N_3364);
or U3889 (N_3889,N_3461,N_3085);
nor U3890 (N_3890,N_3313,N_3474);
nor U3891 (N_3891,N_3312,N_3498);
nand U3892 (N_3892,N_3209,N_3200);
nor U3893 (N_3893,N_3370,N_3228);
or U3894 (N_3894,N_3143,N_3040);
and U3895 (N_3895,N_3183,N_3029);
nor U3896 (N_3896,N_3379,N_3211);
xor U3897 (N_3897,N_3003,N_3089);
or U3898 (N_3898,N_3022,N_3191);
or U3899 (N_3899,N_3394,N_3366);
or U3900 (N_3900,N_3228,N_3103);
xor U3901 (N_3901,N_3282,N_3429);
nand U3902 (N_3902,N_3286,N_3142);
nand U3903 (N_3903,N_3256,N_3058);
xor U3904 (N_3904,N_3491,N_3053);
nand U3905 (N_3905,N_3483,N_3267);
or U3906 (N_3906,N_3103,N_3385);
and U3907 (N_3907,N_3170,N_3430);
and U3908 (N_3908,N_3179,N_3430);
nand U3909 (N_3909,N_3388,N_3166);
nand U3910 (N_3910,N_3255,N_3244);
or U3911 (N_3911,N_3128,N_3008);
xor U3912 (N_3912,N_3485,N_3358);
xor U3913 (N_3913,N_3175,N_3180);
nor U3914 (N_3914,N_3359,N_3271);
or U3915 (N_3915,N_3097,N_3096);
or U3916 (N_3916,N_3408,N_3178);
nor U3917 (N_3917,N_3179,N_3242);
or U3918 (N_3918,N_3405,N_3183);
and U3919 (N_3919,N_3480,N_3044);
nor U3920 (N_3920,N_3388,N_3353);
nand U3921 (N_3921,N_3364,N_3434);
nor U3922 (N_3922,N_3375,N_3148);
or U3923 (N_3923,N_3446,N_3164);
xnor U3924 (N_3924,N_3091,N_3131);
and U3925 (N_3925,N_3288,N_3414);
nor U3926 (N_3926,N_3375,N_3064);
and U3927 (N_3927,N_3380,N_3498);
or U3928 (N_3928,N_3128,N_3226);
nand U3929 (N_3929,N_3203,N_3102);
xor U3930 (N_3930,N_3284,N_3043);
xnor U3931 (N_3931,N_3476,N_3395);
xnor U3932 (N_3932,N_3226,N_3451);
nand U3933 (N_3933,N_3226,N_3159);
and U3934 (N_3934,N_3220,N_3084);
nor U3935 (N_3935,N_3461,N_3340);
nand U3936 (N_3936,N_3218,N_3315);
nand U3937 (N_3937,N_3405,N_3195);
nor U3938 (N_3938,N_3255,N_3383);
nand U3939 (N_3939,N_3366,N_3095);
or U3940 (N_3940,N_3474,N_3384);
nor U3941 (N_3941,N_3357,N_3229);
xnor U3942 (N_3942,N_3365,N_3276);
xnor U3943 (N_3943,N_3411,N_3077);
nor U3944 (N_3944,N_3344,N_3221);
and U3945 (N_3945,N_3055,N_3190);
nand U3946 (N_3946,N_3318,N_3489);
nor U3947 (N_3947,N_3400,N_3440);
or U3948 (N_3948,N_3236,N_3009);
and U3949 (N_3949,N_3366,N_3105);
nand U3950 (N_3950,N_3258,N_3167);
nor U3951 (N_3951,N_3175,N_3413);
nor U3952 (N_3952,N_3404,N_3137);
xnor U3953 (N_3953,N_3124,N_3142);
and U3954 (N_3954,N_3105,N_3349);
xor U3955 (N_3955,N_3050,N_3125);
nand U3956 (N_3956,N_3313,N_3355);
nor U3957 (N_3957,N_3124,N_3259);
or U3958 (N_3958,N_3347,N_3004);
nor U3959 (N_3959,N_3351,N_3134);
or U3960 (N_3960,N_3105,N_3458);
nor U3961 (N_3961,N_3356,N_3104);
or U3962 (N_3962,N_3416,N_3368);
xnor U3963 (N_3963,N_3394,N_3407);
or U3964 (N_3964,N_3124,N_3381);
and U3965 (N_3965,N_3349,N_3302);
nand U3966 (N_3966,N_3084,N_3435);
nor U3967 (N_3967,N_3088,N_3260);
nand U3968 (N_3968,N_3014,N_3168);
nor U3969 (N_3969,N_3313,N_3337);
nor U3970 (N_3970,N_3076,N_3041);
and U3971 (N_3971,N_3106,N_3319);
nand U3972 (N_3972,N_3099,N_3192);
xnor U3973 (N_3973,N_3008,N_3402);
xor U3974 (N_3974,N_3054,N_3009);
and U3975 (N_3975,N_3215,N_3003);
or U3976 (N_3976,N_3059,N_3353);
nand U3977 (N_3977,N_3063,N_3465);
xor U3978 (N_3978,N_3303,N_3411);
or U3979 (N_3979,N_3115,N_3373);
and U3980 (N_3980,N_3306,N_3095);
nand U3981 (N_3981,N_3036,N_3379);
nor U3982 (N_3982,N_3087,N_3352);
and U3983 (N_3983,N_3195,N_3095);
nor U3984 (N_3984,N_3436,N_3086);
nor U3985 (N_3985,N_3057,N_3473);
nor U3986 (N_3986,N_3278,N_3181);
nor U3987 (N_3987,N_3019,N_3480);
and U3988 (N_3988,N_3496,N_3331);
nor U3989 (N_3989,N_3320,N_3313);
and U3990 (N_3990,N_3146,N_3293);
nor U3991 (N_3991,N_3252,N_3109);
xor U3992 (N_3992,N_3031,N_3180);
or U3993 (N_3993,N_3021,N_3166);
or U3994 (N_3994,N_3121,N_3185);
or U3995 (N_3995,N_3444,N_3397);
xnor U3996 (N_3996,N_3455,N_3035);
or U3997 (N_3997,N_3480,N_3272);
and U3998 (N_3998,N_3264,N_3361);
or U3999 (N_3999,N_3236,N_3470);
xnor U4000 (N_4000,N_3648,N_3908);
xor U4001 (N_4001,N_3567,N_3954);
xor U4002 (N_4002,N_3946,N_3762);
or U4003 (N_4003,N_3530,N_3957);
or U4004 (N_4004,N_3594,N_3851);
nand U4005 (N_4005,N_3756,N_3660);
or U4006 (N_4006,N_3965,N_3532);
or U4007 (N_4007,N_3739,N_3736);
xnor U4008 (N_4008,N_3573,N_3525);
or U4009 (N_4009,N_3933,N_3841);
nand U4010 (N_4010,N_3990,N_3794);
xnor U4011 (N_4011,N_3628,N_3776);
nand U4012 (N_4012,N_3615,N_3845);
and U4013 (N_4013,N_3602,N_3672);
xor U4014 (N_4014,N_3562,N_3669);
xnor U4015 (N_4015,N_3824,N_3925);
xor U4016 (N_4016,N_3880,N_3759);
xor U4017 (N_4017,N_3597,N_3639);
xor U4018 (N_4018,N_3766,N_3898);
nand U4019 (N_4019,N_3775,N_3840);
and U4020 (N_4020,N_3867,N_3976);
nand U4021 (N_4021,N_3600,N_3553);
nor U4022 (N_4022,N_3797,N_3924);
and U4023 (N_4023,N_3773,N_3588);
xnor U4024 (N_4024,N_3504,N_3813);
or U4025 (N_4025,N_3650,N_3698);
and U4026 (N_4026,N_3838,N_3630);
nand U4027 (N_4027,N_3901,N_3595);
nor U4028 (N_4028,N_3966,N_3564);
nor U4029 (N_4029,N_3655,N_3877);
and U4030 (N_4030,N_3651,N_3677);
nor U4031 (N_4031,N_3528,N_3599);
and U4032 (N_4032,N_3844,N_3605);
xnor U4033 (N_4033,N_3832,N_3506);
xor U4034 (N_4034,N_3685,N_3806);
nor U4035 (N_4035,N_3747,N_3757);
and U4036 (N_4036,N_3787,N_3996);
xnor U4037 (N_4037,N_3916,N_3695);
or U4038 (N_4038,N_3603,N_3612);
or U4039 (N_4039,N_3548,N_3661);
and U4040 (N_4040,N_3937,N_3812);
nor U4041 (N_4041,N_3883,N_3549);
and U4042 (N_4042,N_3590,N_3904);
or U4043 (N_4043,N_3755,N_3589);
xor U4044 (N_4044,N_3778,N_3860);
and U4045 (N_4045,N_3729,N_3936);
nor U4046 (N_4046,N_3905,N_3953);
and U4047 (N_4047,N_3679,N_3551);
nand U4048 (N_4048,N_3952,N_3823);
xnor U4049 (N_4049,N_3740,N_3702);
and U4050 (N_4050,N_3720,N_3791);
nand U4051 (N_4051,N_3945,N_3703);
or U4052 (N_4052,N_3738,N_3746);
xnor U4053 (N_4053,N_3897,N_3899);
nor U4054 (N_4054,N_3529,N_3558);
nand U4055 (N_4055,N_3886,N_3550);
nor U4056 (N_4056,N_3938,N_3843);
xor U4057 (N_4057,N_3503,N_3539);
xor U4058 (N_4058,N_3725,N_3818);
nor U4059 (N_4059,N_3917,N_3792);
and U4060 (N_4060,N_3790,N_3948);
xor U4061 (N_4061,N_3994,N_3986);
and U4062 (N_4062,N_3663,N_3930);
nor U4063 (N_4063,N_3998,N_3693);
xor U4064 (N_4064,N_3638,N_3714);
nand U4065 (N_4065,N_3682,N_3799);
and U4066 (N_4066,N_3890,N_3934);
nand U4067 (N_4067,N_3804,N_3942);
nor U4068 (N_4068,N_3712,N_3560);
and U4069 (N_4069,N_3967,N_3878);
xor U4070 (N_4070,N_3859,N_3795);
nor U4071 (N_4071,N_3970,N_3817);
or U4072 (N_4072,N_3857,N_3542);
or U4073 (N_4073,N_3516,N_3983);
nand U4074 (N_4074,N_3944,N_3742);
or U4075 (N_4075,N_3989,N_3834);
and U4076 (N_4076,N_3500,N_3671);
or U4077 (N_4077,N_3535,N_3544);
nand U4078 (N_4078,N_3999,N_3598);
nor U4079 (N_4079,N_3931,N_3502);
and U4080 (N_4080,N_3670,N_3637);
xor U4081 (N_4081,N_3950,N_3825);
nand U4082 (N_4082,N_3918,N_3984);
nand U4083 (N_4083,N_3912,N_3520);
and U4084 (N_4084,N_3808,N_3760);
or U4085 (N_4085,N_3675,N_3853);
and U4086 (N_4086,N_3872,N_3708);
xor U4087 (N_4087,N_3764,N_3837);
nor U4088 (N_4088,N_3568,N_3796);
nor U4089 (N_4089,N_3518,N_3765);
xor U4090 (N_4090,N_3889,N_3507);
or U4091 (N_4091,N_3659,N_3616);
xor U4092 (N_4092,N_3971,N_3586);
nor U4093 (N_4093,N_3839,N_3955);
and U4094 (N_4094,N_3910,N_3995);
xor U4095 (N_4095,N_3624,N_3537);
or U4096 (N_4096,N_3761,N_3949);
nor U4097 (N_4097,N_3533,N_3514);
nand U4098 (N_4098,N_3563,N_3977);
nor U4099 (N_4099,N_3610,N_3782);
nand U4100 (N_4100,N_3814,N_3634);
nor U4101 (N_4101,N_3617,N_3858);
nor U4102 (N_4102,N_3830,N_3831);
or U4103 (N_4103,N_3727,N_3960);
nor U4104 (N_4104,N_3958,N_3571);
xnor U4105 (N_4105,N_3884,N_3801);
and U4106 (N_4106,N_3927,N_3632);
nor U4107 (N_4107,N_3572,N_3678);
nand U4108 (N_4108,N_3515,N_3710);
or U4109 (N_4109,N_3730,N_3940);
nand U4110 (N_4110,N_3694,N_3688);
nor U4111 (N_4111,N_3517,N_3654);
xor U4112 (N_4112,N_3674,N_3613);
and U4113 (N_4113,N_3980,N_3723);
nand U4114 (N_4114,N_3829,N_3821);
nand U4115 (N_4115,N_3767,N_3956);
or U4116 (N_4116,N_3754,N_3541);
xor U4117 (N_4117,N_3676,N_3644);
or U4118 (N_4118,N_3850,N_3581);
or U4119 (N_4119,N_3777,N_3784);
and U4120 (N_4120,N_3854,N_3869);
and U4121 (N_4121,N_3815,N_3785);
and U4122 (N_4122,N_3547,N_3704);
or U4123 (N_4123,N_3735,N_3882);
and U4124 (N_4124,N_3578,N_3749);
and U4125 (N_4125,N_3522,N_3943);
xnor U4126 (N_4126,N_3716,N_3923);
nand U4127 (N_4127,N_3719,N_3750);
xor U4128 (N_4128,N_3583,N_3875);
nor U4129 (N_4129,N_3896,N_3501);
nor U4130 (N_4130,N_3763,N_3584);
or U4131 (N_4131,N_3687,N_3577);
xnor U4132 (N_4132,N_3892,N_3647);
xor U4133 (N_4133,N_3932,N_3789);
nor U4134 (N_4134,N_3665,N_3513);
or U4135 (N_4135,N_3524,N_3546);
nand U4136 (N_4136,N_3592,N_3512);
or U4137 (N_4137,N_3689,N_3874);
nand U4138 (N_4138,N_3575,N_3987);
or U4139 (N_4139,N_3900,N_3914);
nor U4140 (N_4140,N_3523,N_3696);
xnor U4141 (N_4141,N_3629,N_3633);
xnor U4142 (N_4142,N_3935,N_3623);
or U4143 (N_4143,N_3582,N_3656);
or U4144 (N_4144,N_3711,N_3591);
nor U4145 (N_4145,N_3626,N_3643);
nor U4146 (N_4146,N_3893,N_3508);
nor U4147 (N_4147,N_3873,N_3627);
nor U4148 (N_4148,N_3680,N_3636);
xor U4149 (N_4149,N_3731,N_3961);
and U4150 (N_4150,N_3555,N_3536);
and U4151 (N_4151,N_3732,N_3673);
nor U4152 (N_4152,N_3509,N_3635);
xnor U4153 (N_4153,N_3733,N_3565);
nor U4154 (N_4154,N_3863,N_3652);
and U4155 (N_4155,N_3649,N_3741);
nand U4156 (N_4156,N_3803,N_3768);
or U4157 (N_4157,N_3705,N_3753);
xnor U4158 (N_4158,N_3646,N_3601);
and U4159 (N_4159,N_3653,N_3540);
xnor U4160 (N_4160,N_3667,N_3622);
nor U4161 (N_4161,N_3527,N_3822);
nand U4162 (N_4162,N_3992,N_3511);
nor U4163 (N_4163,N_3793,N_3666);
xor U4164 (N_4164,N_3557,N_3816);
nor U4165 (N_4165,N_3751,N_3915);
or U4166 (N_4166,N_3788,N_3922);
nand U4167 (N_4167,N_3852,N_3706);
xor U4168 (N_4168,N_3566,N_3798);
or U4169 (N_4169,N_3964,N_3774);
nor U4170 (N_4170,N_3724,N_3713);
nand U4171 (N_4171,N_3833,N_3781);
or U4172 (N_4172,N_3895,N_3941);
nand U4173 (N_4173,N_3861,N_3826);
xor U4174 (N_4174,N_3979,N_3668);
nor U4175 (N_4175,N_3836,N_3748);
nand U4176 (N_4176,N_3929,N_3690);
nand U4177 (N_4177,N_3607,N_3543);
and U4178 (N_4178,N_3614,N_3819);
nor U4179 (N_4179,N_3593,N_3870);
xor U4180 (N_4180,N_3631,N_3981);
or U4181 (N_4181,N_3576,N_3664);
xor U4182 (N_4182,N_3856,N_3700);
and U4183 (N_4183,N_3692,N_3887);
or U4184 (N_4184,N_3920,N_3973);
and U4185 (N_4185,N_3888,N_3894);
xnor U4186 (N_4186,N_3985,N_3618);
and U4187 (N_4187,N_3596,N_3745);
or U4188 (N_4188,N_3909,N_3570);
or U4189 (N_4189,N_3807,N_3828);
and U4190 (N_4190,N_3526,N_3835);
and U4191 (N_4191,N_3662,N_3969);
or U4192 (N_4192,N_3734,N_3913);
and U4193 (N_4193,N_3805,N_3951);
nand U4194 (N_4194,N_3531,N_3993);
or U4195 (N_4195,N_3538,N_3921);
or U4196 (N_4196,N_3606,N_3902);
nand U4197 (N_4197,N_3876,N_3972);
nor U4198 (N_4198,N_3962,N_3519);
nor U4199 (N_4199,N_3718,N_3800);
xnor U4200 (N_4200,N_3691,N_3772);
xor U4201 (N_4201,N_3619,N_3848);
nand U4202 (N_4202,N_3928,N_3871);
xnor U4203 (N_4203,N_3620,N_3657);
nand U4204 (N_4204,N_3786,N_3642);
nor U4205 (N_4205,N_3744,N_3699);
nor U4206 (N_4206,N_3847,N_3997);
or U4207 (N_4207,N_3580,N_3988);
xor U4208 (N_4208,N_3554,N_3585);
nor U4209 (N_4209,N_3810,N_3947);
and U4210 (N_4210,N_3780,N_3842);
xor U4211 (N_4211,N_3545,N_3771);
and U4212 (N_4212,N_3697,N_3820);
nand U4213 (N_4213,N_3802,N_3811);
or U4214 (N_4214,N_3604,N_3879);
or U4215 (N_4215,N_3722,N_3556);
nand U4216 (N_4216,N_3641,N_3683);
or U4217 (N_4217,N_3728,N_3737);
nor U4218 (N_4218,N_3868,N_3906);
nand U4219 (N_4219,N_3919,N_3521);
nor U4220 (N_4220,N_3758,N_3574);
or U4221 (N_4221,N_3505,N_3959);
or U4222 (N_4222,N_3645,N_3552);
and U4223 (N_4223,N_3939,N_3849);
nand U4224 (N_4224,N_3864,N_3701);
and U4225 (N_4225,N_3559,N_3686);
nor U4226 (N_4226,N_3911,N_3621);
xor U4227 (N_4227,N_3783,N_3681);
nor U4228 (N_4228,N_3926,N_3561);
or U4229 (N_4229,N_3963,N_3866);
xnor U4230 (N_4230,N_3534,N_3510);
nand U4231 (N_4231,N_3770,N_3975);
and U4232 (N_4232,N_3717,N_3968);
nand U4233 (N_4233,N_3809,N_3743);
nor U4234 (N_4234,N_3881,N_3769);
nor U4235 (N_4235,N_3991,N_3569);
or U4236 (N_4236,N_3625,N_3846);
or U4237 (N_4237,N_3903,N_3611);
nor U4238 (N_4238,N_3891,N_3579);
and U4239 (N_4239,N_3608,N_3752);
xor U4240 (N_4240,N_3721,N_3855);
or U4241 (N_4241,N_3726,N_3885);
and U4242 (N_4242,N_3640,N_3658);
nand U4243 (N_4243,N_3715,N_3779);
and U4244 (N_4244,N_3587,N_3978);
nand U4245 (N_4245,N_3709,N_3974);
and U4246 (N_4246,N_3609,N_3907);
nand U4247 (N_4247,N_3827,N_3707);
nor U4248 (N_4248,N_3982,N_3684);
nand U4249 (N_4249,N_3865,N_3862);
nor U4250 (N_4250,N_3832,N_3544);
and U4251 (N_4251,N_3537,N_3589);
nor U4252 (N_4252,N_3971,N_3941);
and U4253 (N_4253,N_3625,N_3521);
and U4254 (N_4254,N_3549,N_3652);
or U4255 (N_4255,N_3647,N_3677);
nor U4256 (N_4256,N_3993,N_3695);
xor U4257 (N_4257,N_3920,N_3764);
xor U4258 (N_4258,N_3658,N_3988);
nand U4259 (N_4259,N_3954,N_3883);
and U4260 (N_4260,N_3903,N_3999);
nand U4261 (N_4261,N_3914,N_3587);
or U4262 (N_4262,N_3643,N_3809);
or U4263 (N_4263,N_3525,N_3775);
and U4264 (N_4264,N_3540,N_3692);
nor U4265 (N_4265,N_3570,N_3507);
nor U4266 (N_4266,N_3681,N_3903);
or U4267 (N_4267,N_3687,N_3905);
nand U4268 (N_4268,N_3548,N_3550);
nor U4269 (N_4269,N_3638,N_3645);
or U4270 (N_4270,N_3778,N_3558);
nand U4271 (N_4271,N_3738,N_3880);
nand U4272 (N_4272,N_3904,N_3658);
xor U4273 (N_4273,N_3548,N_3651);
nand U4274 (N_4274,N_3921,N_3586);
nor U4275 (N_4275,N_3746,N_3857);
xnor U4276 (N_4276,N_3902,N_3689);
or U4277 (N_4277,N_3618,N_3706);
and U4278 (N_4278,N_3654,N_3981);
or U4279 (N_4279,N_3880,N_3775);
and U4280 (N_4280,N_3845,N_3781);
nor U4281 (N_4281,N_3541,N_3523);
nor U4282 (N_4282,N_3638,N_3979);
nand U4283 (N_4283,N_3596,N_3705);
nand U4284 (N_4284,N_3640,N_3956);
nand U4285 (N_4285,N_3564,N_3567);
nor U4286 (N_4286,N_3604,N_3852);
and U4287 (N_4287,N_3657,N_3622);
or U4288 (N_4288,N_3688,N_3663);
and U4289 (N_4289,N_3604,N_3580);
nor U4290 (N_4290,N_3805,N_3665);
or U4291 (N_4291,N_3810,N_3640);
nand U4292 (N_4292,N_3569,N_3549);
nand U4293 (N_4293,N_3640,N_3597);
xnor U4294 (N_4294,N_3856,N_3802);
or U4295 (N_4295,N_3551,N_3938);
and U4296 (N_4296,N_3881,N_3795);
nand U4297 (N_4297,N_3656,N_3947);
nor U4298 (N_4298,N_3795,N_3899);
nor U4299 (N_4299,N_3890,N_3788);
nand U4300 (N_4300,N_3597,N_3913);
nor U4301 (N_4301,N_3718,N_3733);
and U4302 (N_4302,N_3547,N_3710);
nand U4303 (N_4303,N_3965,N_3630);
xor U4304 (N_4304,N_3833,N_3783);
or U4305 (N_4305,N_3661,N_3874);
nor U4306 (N_4306,N_3810,N_3906);
nor U4307 (N_4307,N_3814,N_3917);
or U4308 (N_4308,N_3666,N_3984);
nand U4309 (N_4309,N_3722,N_3862);
xnor U4310 (N_4310,N_3700,N_3807);
or U4311 (N_4311,N_3954,N_3775);
nand U4312 (N_4312,N_3571,N_3774);
nor U4313 (N_4313,N_3649,N_3681);
nand U4314 (N_4314,N_3615,N_3738);
nor U4315 (N_4315,N_3891,N_3792);
xnor U4316 (N_4316,N_3860,N_3616);
nand U4317 (N_4317,N_3565,N_3822);
nor U4318 (N_4318,N_3595,N_3678);
or U4319 (N_4319,N_3621,N_3519);
nor U4320 (N_4320,N_3942,N_3843);
xor U4321 (N_4321,N_3968,N_3842);
nor U4322 (N_4322,N_3838,N_3972);
xnor U4323 (N_4323,N_3604,N_3743);
xor U4324 (N_4324,N_3593,N_3958);
xnor U4325 (N_4325,N_3939,N_3539);
and U4326 (N_4326,N_3676,N_3753);
xnor U4327 (N_4327,N_3693,N_3858);
xnor U4328 (N_4328,N_3822,N_3770);
nor U4329 (N_4329,N_3692,N_3991);
xnor U4330 (N_4330,N_3944,N_3744);
nand U4331 (N_4331,N_3701,N_3911);
nand U4332 (N_4332,N_3660,N_3979);
nor U4333 (N_4333,N_3517,N_3581);
xnor U4334 (N_4334,N_3680,N_3686);
nand U4335 (N_4335,N_3828,N_3604);
nor U4336 (N_4336,N_3568,N_3752);
xnor U4337 (N_4337,N_3812,N_3710);
nor U4338 (N_4338,N_3557,N_3669);
or U4339 (N_4339,N_3844,N_3823);
xor U4340 (N_4340,N_3522,N_3675);
xnor U4341 (N_4341,N_3969,N_3591);
xnor U4342 (N_4342,N_3694,N_3525);
nor U4343 (N_4343,N_3881,N_3957);
xnor U4344 (N_4344,N_3821,N_3981);
nor U4345 (N_4345,N_3703,N_3908);
or U4346 (N_4346,N_3937,N_3599);
nor U4347 (N_4347,N_3511,N_3838);
and U4348 (N_4348,N_3591,N_3997);
and U4349 (N_4349,N_3756,N_3859);
and U4350 (N_4350,N_3552,N_3536);
nor U4351 (N_4351,N_3551,N_3788);
nor U4352 (N_4352,N_3712,N_3877);
nand U4353 (N_4353,N_3512,N_3721);
or U4354 (N_4354,N_3661,N_3681);
nor U4355 (N_4355,N_3877,N_3805);
or U4356 (N_4356,N_3626,N_3864);
nor U4357 (N_4357,N_3918,N_3559);
and U4358 (N_4358,N_3647,N_3978);
nor U4359 (N_4359,N_3642,N_3577);
nand U4360 (N_4360,N_3705,N_3713);
and U4361 (N_4361,N_3829,N_3688);
xor U4362 (N_4362,N_3812,N_3854);
or U4363 (N_4363,N_3503,N_3796);
nor U4364 (N_4364,N_3688,N_3590);
nor U4365 (N_4365,N_3740,N_3898);
or U4366 (N_4366,N_3775,N_3949);
xnor U4367 (N_4367,N_3831,N_3782);
xor U4368 (N_4368,N_3876,N_3984);
xnor U4369 (N_4369,N_3703,N_3570);
xor U4370 (N_4370,N_3661,N_3914);
nand U4371 (N_4371,N_3899,N_3952);
nor U4372 (N_4372,N_3588,N_3852);
nand U4373 (N_4373,N_3769,N_3680);
and U4374 (N_4374,N_3668,N_3618);
nand U4375 (N_4375,N_3528,N_3600);
nor U4376 (N_4376,N_3783,N_3663);
or U4377 (N_4377,N_3663,N_3881);
nor U4378 (N_4378,N_3781,N_3742);
or U4379 (N_4379,N_3550,N_3804);
nand U4380 (N_4380,N_3744,N_3516);
nand U4381 (N_4381,N_3897,N_3680);
and U4382 (N_4382,N_3907,N_3898);
or U4383 (N_4383,N_3744,N_3610);
xnor U4384 (N_4384,N_3654,N_3562);
xor U4385 (N_4385,N_3855,N_3720);
xor U4386 (N_4386,N_3697,N_3500);
and U4387 (N_4387,N_3850,N_3640);
nand U4388 (N_4388,N_3897,N_3729);
nand U4389 (N_4389,N_3551,N_3944);
nand U4390 (N_4390,N_3567,N_3772);
and U4391 (N_4391,N_3602,N_3770);
nand U4392 (N_4392,N_3795,N_3606);
xnor U4393 (N_4393,N_3926,N_3521);
nand U4394 (N_4394,N_3845,N_3924);
xnor U4395 (N_4395,N_3707,N_3634);
and U4396 (N_4396,N_3913,N_3629);
nor U4397 (N_4397,N_3879,N_3717);
nand U4398 (N_4398,N_3724,N_3866);
and U4399 (N_4399,N_3912,N_3877);
and U4400 (N_4400,N_3736,N_3572);
xor U4401 (N_4401,N_3537,N_3999);
and U4402 (N_4402,N_3770,N_3625);
xnor U4403 (N_4403,N_3767,N_3828);
nor U4404 (N_4404,N_3586,N_3917);
and U4405 (N_4405,N_3724,N_3710);
xor U4406 (N_4406,N_3884,N_3804);
nand U4407 (N_4407,N_3613,N_3660);
and U4408 (N_4408,N_3692,N_3726);
or U4409 (N_4409,N_3981,N_3716);
nor U4410 (N_4410,N_3979,N_3914);
xor U4411 (N_4411,N_3526,N_3553);
nor U4412 (N_4412,N_3633,N_3935);
xor U4413 (N_4413,N_3932,N_3793);
and U4414 (N_4414,N_3907,N_3788);
nand U4415 (N_4415,N_3583,N_3926);
or U4416 (N_4416,N_3738,N_3529);
xnor U4417 (N_4417,N_3771,N_3637);
or U4418 (N_4418,N_3690,N_3512);
nor U4419 (N_4419,N_3690,N_3806);
nor U4420 (N_4420,N_3857,N_3507);
nand U4421 (N_4421,N_3765,N_3647);
nand U4422 (N_4422,N_3615,N_3746);
nor U4423 (N_4423,N_3836,N_3574);
or U4424 (N_4424,N_3990,N_3636);
and U4425 (N_4425,N_3619,N_3917);
and U4426 (N_4426,N_3993,N_3518);
or U4427 (N_4427,N_3787,N_3714);
and U4428 (N_4428,N_3717,N_3585);
or U4429 (N_4429,N_3525,N_3973);
or U4430 (N_4430,N_3680,N_3532);
nor U4431 (N_4431,N_3932,N_3828);
xnor U4432 (N_4432,N_3600,N_3508);
and U4433 (N_4433,N_3913,N_3904);
nor U4434 (N_4434,N_3873,N_3636);
nand U4435 (N_4435,N_3961,N_3868);
xor U4436 (N_4436,N_3574,N_3623);
nor U4437 (N_4437,N_3565,N_3930);
xnor U4438 (N_4438,N_3664,N_3659);
or U4439 (N_4439,N_3704,N_3894);
nand U4440 (N_4440,N_3698,N_3640);
and U4441 (N_4441,N_3743,N_3925);
xor U4442 (N_4442,N_3735,N_3840);
nor U4443 (N_4443,N_3978,N_3996);
or U4444 (N_4444,N_3973,N_3922);
and U4445 (N_4445,N_3507,N_3772);
or U4446 (N_4446,N_3855,N_3744);
nor U4447 (N_4447,N_3653,N_3671);
xor U4448 (N_4448,N_3702,N_3953);
and U4449 (N_4449,N_3856,N_3814);
nand U4450 (N_4450,N_3665,N_3992);
nor U4451 (N_4451,N_3744,N_3614);
or U4452 (N_4452,N_3873,N_3668);
nor U4453 (N_4453,N_3542,N_3562);
nand U4454 (N_4454,N_3868,N_3620);
nand U4455 (N_4455,N_3614,N_3501);
xor U4456 (N_4456,N_3795,N_3613);
xnor U4457 (N_4457,N_3742,N_3536);
or U4458 (N_4458,N_3663,N_3907);
xor U4459 (N_4459,N_3601,N_3653);
and U4460 (N_4460,N_3662,N_3888);
nand U4461 (N_4461,N_3754,N_3547);
nand U4462 (N_4462,N_3564,N_3628);
xor U4463 (N_4463,N_3896,N_3888);
nand U4464 (N_4464,N_3883,N_3724);
xor U4465 (N_4465,N_3644,N_3981);
nand U4466 (N_4466,N_3913,N_3869);
xor U4467 (N_4467,N_3541,N_3681);
nand U4468 (N_4468,N_3993,N_3542);
and U4469 (N_4469,N_3772,N_3824);
or U4470 (N_4470,N_3620,N_3591);
and U4471 (N_4471,N_3792,N_3863);
nand U4472 (N_4472,N_3943,N_3714);
and U4473 (N_4473,N_3647,N_3693);
xor U4474 (N_4474,N_3711,N_3787);
or U4475 (N_4475,N_3681,N_3990);
nor U4476 (N_4476,N_3985,N_3581);
and U4477 (N_4477,N_3798,N_3502);
nand U4478 (N_4478,N_3737,N_3864);
and U4479 (N_4479,N_3978,N_3970);
and U4480 (N_4480,N_3515,N_3871);
or U4481 (N_4481,N_3549,N_3603);
nand U4482 (N_4482,N_3618,N_3773);
and U4483 (N_4483,N_3907,N_3514);
xor U4484 (N_4484,N_3615,N_3529);
or U4485 (N_4485,N_3543,N_3684);
or U4486 (N_4486,N_3838,N_3706);
or U4487 (N_4487,N_3882,N_3843);
and U4488 (N_4488,N_3765,N_3925);
nand U4489 (N_4489,N_3693,N_3561);
and U4490 (N_4490,N_3995,N_3920);
nor U4491 (N_4491,N_3518,N_3510);
nor U4492 (N_4492,N_3763,N_3721);
nand U4493 (N_4493,N_3510,N_3788);
and U4494 (N_4494,N_3593,N_3582);
xor U4495 (N_4495,N_3535,N_3565);
nor U4496 (N_4496,N_3552,N_3980);
and U4497 (N_4497,N_3937,N_3930);
nor U4498 (N_4498,N_3986,N_3666);
or U4499 (N_4499,N_3898,N_3972);
nor U4500 (N_4500,N_4393,N_4220);
nor U4501 (N_4501,N_4051,N_4428);
and U4502 (N_4502,N_4484,N_4367);
and U4503 (N_4503,N_4158,N_4398);
or U4504 (N_4504,N_4238,N_4360);
or U4505 (N_4505,N_4138,N_4109);
xor U4506 (N_4506,N_4422,N_4200);
nand U4507 (N_4507,N_4432,N_4154);
xnor U4508 (N_4508,N_4479,N_4172);
and U4509 (N_4509,N_4232,N_4358);
xor U4510 (N_4510,N_4499,N_4298);
xor U4511 (N_4511,N_4126,N_4108);
or U4512 (N_4512,N_4343,N_4076);
nor U4513 (N_4513,N_4205,N_4122);
nand U4514 (N_4514,N_4282,N_4046);
xor U4515 (N_4515,N_4020,N_4347);
or U4516 (N_4516,N_4447,N_4204);
xor U4517 (N_4517,N_4181,N_4057);
and U4518 (N_4518,N_4225,N_4178);
xor U4519 (N_4519,N_4330,N_4470);
or U4520 (N_4520,N_4169,N_4216);
nor U4521 (N_4521,N_4354,N_4237);
xor U4522 (N_4522,N_4086,N_4176);
nand U4523 (N_4523,N_4319,N_4023);
nor U4524 (N_4524,N_4124,N_4287);
nand U4525 (N_4525,N_4437,N_4102);
nand U4526 (N_4526,N_4105,N_4257);
xnor U4527 (N_4527,N_4445,N_4440);
nor U4528 (N_4528,N_4083,N_4413);
nand U4529 (N_4529,N_4435,N_4091);
or U4530 (N_4530,N_4261,N_4151);
and U4531 (N_4531,N_4338,N_4009);
and U4532 (N_4532,N_4424,N_4116);
nand U4533 (N_4533,N_4193,N_4117);
nor U4534 (N_4534,N_4025,N_4164);
or U4535 (N_4535,N_4133,N_4002);
and U4536 (N_4536,N_4192,N_4431);
xor U4537 (N_4537,N_4494,N_4007);
or U4538 (N_4538,N_4317,N_4034);
nand U4539 (N_4539,N_4455,N_4197);
or U4540 (N_4540,N_4452,N_4331);
xnor U4541 (N_4541,N_4371,N_4297);
and U4542 (N_4542,N_4386,N_4453);
or U4543 (N_4543,N_4092,N_4352);
xnor U4544 (N_4544,N_4483,N_4449);
nand U4545 (N_4545,N_4219,N_4035);
xor U4546 (N_4546,N_4241,N_4326);
nor U4547 (N_4547,N_4161,N_4230);
or U4548 (N_4548,N_4471,N_4361);
nand U4549 (N_4549,N_4210,N_4269);
and U4550 (N_4550,N_4231,N_4212);
nor U4551 (N_4551,N_4396,N_4142);
nand U4552 (N_4552,N_4356,N_4295);
nand U4553 (N_4553,N_4429,N_4341);
and U4554 (N_4554,N_4156,N_4081);
and U4555 (N_4555,N_4168,N_4072);
nor U4556 (N_4556,N_4497,N_4469);
nand U4557 (N_4557,N_4467,N_4421);
nor U4558 (N_4558,N_4337,N_4388);
nand U4559 (N_4559,N_4253,N_4475);
nand U4560 (N_4560,N_4378,N_4407);
nor U4561 (N_4561,N_4476,N_4387);
nor U4562 (N_4562,N_4120,N_4084);
xnor U4563 (N_4563,N_4087,N_4148);
nor U4564 (N_4564,N_4442,N_4404);
nand U4565 (N_4565,N_4325,N_4199);
and U4566 (N_4566,N_4420,N_4304);
and U4567 (N_4567,N_4480,N_4082);
nor U4568 (N_4568,N_4278,N_4111);
nand U4569 (N_4569,N_4362,N_4094);
and U4570 (N_4570,N_4474,N_4121);
xnor U4571 (N_4571,N_4183,N_4136);
and U4572 (N_4572,N_4370,N_4299);
xor U4573 (N_4573,N_4018,N_4332);
nor U4574 (N_4574,N_4281,N_4245);
xnor U4575 (N_4575,N_4415,N_4090);
xor U4576 (N_4576,N_4139,N_4208);
nand U4577 (N_4577,N_4194,N_4173);
or U4578 (N_4578,N_4485,N_4242);
or U4579 (N_4579,N_4477,N_4016);
and U4580 (N_4580,N_4067,N_4384);
nor U4581 (N_4581,N_4265,N_4079);
or U4582 (N_4582,N_4180,N_4272);
or U4583 (N_4583,N_4191,N_4135);
xor U4584 (N_4584,N_4436,N_4328);
nor U4585 (N_4585,N_4275,N_4163);
or U4586 (N_4586,N_4236,N_4008);
nor U4587 (N_4587,N_4377,N_4303);
xor U4588 (N_4588,N_4374,N_4159);
nor U4589 (N_4589,N_4305,N_4464);
nand U4590 (N_4590,N_4403,N_4300);
nand U4591 (N_4591,N_4426,N_4399);
or U4592 (N_4592,N_4088,N_4149);
and U4593 (N_4593,N_4335,N_4053);
or U4594 (N_4594,N_4036,N_4410);
nor U4595 (N_4595,N_4492,N_4198);
nand U4596 (N_4596,N_4277,N_4400);
xnor U4597 (N_4597,N_4414,N_4038);
and U4598 (N_4598,N_4250,N_4114);
nor U4599 (N_4599,N_4177,N_4292);
nand U4600 (N_4600,N_4058,N_4248);
nand U4601 (N_4601,N_4486,N_4215);
nand U4602 (N_4602,N_4255,N_4301);
xnor U4603 (N_4603,N_4000,N_4376);
xnor U4604 (N_4604,N_4129,N_4221);
xor U4605 (N_4605,N_4329,N_4234);
nor U4606 (N_4606,N_4307,N_4383);
nor U4607 (N_4607,N_4206,N_4373);
xnor U4608 (N_4608,N_4350,N_4014);
nand U4609 (N_4609,N_4382,N_4030);
or U4610 (N_4610,N_4165,N_4381);
xnor U4611 (N_4611,N_4458,N_4359);
and U4612 (N_4612,N_4095,N_4048);
or U4613 (N_4613,N_4351,N_4251);
nor U4614 (N_4614,N_4478,N_4070);
nor U4615 (N_4615,N_4260,N_4003);
or U4616 (N_4616,N_4147,N_4213);
and U4617 (N_4617,N_4267,N_4185);
or U4618 (N_4618,N_4227,N_4033);
and U4619 (N_4619,N_4071,N_4152);
xor U4620 (N_4620,N_4011,N_4170);
or U4621 (N_4621,N_4355,N_4296);
xor U4622 (N_4622,N_4107,N_4392);
xor U4623 (N_4623,N_4468,N_4451);
nand U4624 (N_4624,N_4247,N_4055);
nor U4625 (N_4625,N_4043,N_4283);
and U4626 (N_4626,N_4327,N_4363);
xnor U4627 (N_4627,N_4150,N_4119);
xor U4628 (N_4628,N_4130,N_4271);
and U4629 (N_4629,N_4203,N_4425);
nand U4630 (N_4630,N_4324,N_4141);
nand U4631 (N_4631,N_4256,N_4005);
and U4632 (N_4632,N_4409,N_4320);
xnor U4633 (N_4633,N_4228,N_4032);
or U4634 (N_4634,N_4379,N_4021);
and U4635 (N_4635,N_4321,N_4184);
xor U4636 (N_4636,N_4293,N_4490);
nor U4637 (N_4637,N_4202,N_4101);
nor U4638 (N_4638,N_4353,N_4457);
or U4639 (N_4639,N_4438,N_4397);
xnor U4640 (N_4640,N_4103,N_4244);
and U4641 (N_4641,N_4187,N_4050);
xor U4642 (N_4642,N_4259,N_4294);
and U4643 (N_4643,N_4391,N_4024);
nor U4644 (N_4644,N_4174,N_4439);
nor U4645 (N_4645,N_4040,N_4039);
and U4646 (N_4646,N_4380,N_4276);
xnor U4647 (N_4647,N_4450,N_4308);
xor U4648 (N_4648,N_4186,N_4411);
nor U4649 (N_4649,N_4104,N_4270);
or U4650 (N_4650,N_4306,N_4062);
nor U4651 (N_4651,N_4207,N_4465);
xor U4652 (N_4652,N_4446,N_4226);
nand U4653 (N_4653,N_4162,N_4113);
and U4654 (N_4654,N_4097,N_4430);
nor U4655 (N_4655,N_4229,N_4418);
nand U4656 (N_4656,N_4029,N_4128);
nand U4657 (N_4657,N_4498,N_4179);
and U4658 (N_4658,N_4013,N_4123);
or U4659 (N_4659,N_4235,N_4290);
nand U4660 (N_4660,N_4146,N_4074);
or U4661 (N_4661,N_4357,N_4315);
xnor U4662 (N_4662,N_4110,N_4372);
and U4663 (N_4663,N_4314,N_4077);
and U4664 (N_4664,N_4054,N_4375);
and U4665 (N_4665,N_4167,N_4118);
nor U4666 (N_4666,N_4263,N_4243);
or U4667 (N_4667,N_4273,N_4309);
or U4668 (N_4668,N_4344,N_4322);
nand U4669 (N_4669,N_4157,N_4311);
nand U4670 (N_4670,N_4448,N_4280);
xor U4671 (N_4671,N_4209,N_4010);
and U4672 (N_4672,N_4427,N_4318);
xnor U4673 (N_4673,N_4342,N_4027);
nor U4674 (N_4674,N_4346,N_4078);
nand U4675 (N_4675,N_4454,N_4482);
xor U4676 (N_4676,N_4065,N_4390);
and U4677 (N_4677,N_4489,N_4394);
xnor U4678 (N_4678,N_4182,N_4288);
and U4679 (N_4679,N_4160,N_4252);
xor U4680 (N_4680,N_4064,N_4015);
and U4681 (N_4681,N_4481,N_4348);
nor U4682 (N_4682,N_4196,N_4461);
nand U4683 (N_4683,N_4045,N_4313);
nor U4684 (N_4684,N_4444,N_4166);
nor U4685 (N_4685,N_4060,N_4417);
nor U4686 (N_4686,N_4402,N_4408);
nor U4687 (N_4687,N_4333,N_4127);
nand U4688 (N_4688,N_4153,N_4125);
and U4689 (N_4689,N_4443,N_4068);
and U4690 (N_4690,N_4369,N_4496);
and U4691 (N_4691,N_4291,N_4339);
or U4692 (N_4692,N_4223,N_4217);
xnor U4693 (N_4693,N_4144,N_4066);
or U4694 (N_4694,N_4044,N_4279);
xor U4695 (N_4695,N_4052,N_4385);
or U4696 (N_4696,N_4047,N_4462);
or U4697 (N_4697,N_4340,N_4175);
and U4698 (N_4698,N_4365,N_4017);
nand U4699 (N_4699,N_4345,N_4246);
or U4700 (N_4700,N_4006,N_4137);
nand U4701 (N_4701,N_4089,N_4389);
nand U4702 (N_4702,N_4233,N_4222);
nor U4703 (N_4703,N_4423,N_4211);
nand U4704 (N_4704,N_4249,N_4466);
xnor U4705 (N_4705,N_4495,N_4266);
nor U4706 (N_4706,N_4224,N_4366);
nand U4707 (N_4707,N_4488,N_4093);
nor U4708 (N_4708,N_4310,N_4132);
xnor U4709 (N_4709,N_4099,N_4028);
nor U4710 (N_4710,N_4491,N_4069);
nand U4711 (N_4711,N_4075,N_4368);
xor U4712 (N_4712,N_4019,N_4131);
or U4713 (N_4713,N_4412,N_4406);
xnor U4714 (N_4714,N_4349,N_4312);
nand U4715 (N_4715,N_4098,N_4364);
and U4716 (N_4716,N_4188,N_4268);
nand U4717 (N_4717,N_4195,N_4112);
and U4718 (N_4718,N_4472,N_4115);
nand U4719 (N_4719,N_4493,N_4323);
xor U4720 (N_4720,N_4037,N_4316);
or U4721 (N_4721,N_4096,N_4134);
and U4722 (N_4722,N_4004,N_4031);
or U4723 (N_4723,N_4285,N_4042);
xnor U4724 (N_4724,N_4258,N_4106);
nor U4725 (N_4725,N_4080,N_4459);
xnor U4726 (N_4726,N_4145,N_4218);
or U4727 (N_4727,N_4254,N_4143);
or U4728 (N_4728,N_4262,N_4473);
nor U4729 (N_4729,N_4140,N_4155);
nand U4730 (N_4730,N_4487,N_4100);
nor U4731 (N_4731,N_4022,N_4401);
nor U4732 (N_4732,N_4416,N_4171);
and U4733 (N_4733,N_4012,N_4336);
nand U4734 (N_4734,N_4460,N_4049);
nand U4735 (N_4735,N_4302,N_4056);
xnor U4736 (N_4736,N_4190,N_4214);
nand U4737 (N_4737,N_4073,N_4441);
nor U4738 (N_4738,N_4433,N_4405);
nand U4739 (N_4739,N_4274,N_4239);
xnor U4740 (N_4740,N_4286,N_4434);
nor U4741 (N_4741,N_4240,N_4419);
xor U4742 (N_4742,N_4201,N_4334);
or U4743 (N_4743,N_4063,N_4041);
nor U4744 (N_4744,N_4284,N_4061);
nor U4745 (N_4745,N_4289,N_4395);
or U4746 (N_4746,N_4001,N_4189);
xor U4747 (N_4747,N_4026,N_4463);
nor U4748 (N_4748,N_4264,N_4456);
xnor U4749 (N_4749,N_4085,N_4059);
nand U4750 (N_4750,N_4316,N_4269);
nand U4751 (N_4751,N_4066,N_4448);
xor U4752 (N_4752,N_4320,N_4215);
xor U4753 (N_4753,N_4270,N_4471);
nor U4754 (N_4754,N_4010,N_4397);
nor U4755 (N_4755,N_4156,N_4398);
nand U4756 (N_4756,N_4167,N_4484);
nor U4757 (N_4757,N_4055,N_4160);
nand U4758 (N_4758,N_4472,N_4360);
nand U4759 (N_4759,N_4494,N_4189);
or U4760 (N_4760,N_4414,N_4165);
nand U4761 (N_4761,N_4349,N_4059);
xnor U4762 (N_4762,N_4030,N_4410);
or U4763 (N_4763,N_4483,N_4369);
and U4764 (N_4764,N_4160,N_4320);
nor U4765 (N_4765,N_4396,N_4105);
or U4766 (N_4766,N_4017,N_4454);
xnor U4767 (N_4767,N_4424,N_4320);
and U4768 (N_4768,N_4102,N_4315);
and U4769 (N_4769,N_4009,N_4408);
xnor U4770 (N_4770,N_4264,N_4008);
and U4771 (N_4771,N_4403,N_4011);
xor U4772 (N_4772,N_4179,N_4385);
and U4773 (N_4773,N_4400,N_4061);
and U4774 (N_4774,N_4163,N_4207);
and U4775 (N_4775,N_4410,N_4346);
or U4776 (N_4776,N_4091,N_4169);
xnor U4777 (N_4777,N_4141,N_4182);
xnor U4778 (N_4778,N_4469,N_4182);
nor U4779 (N_4779,N_4201,N_4475);
or U4780 (N_4780,N_4465,N_4024);
nand U4781 (N_4781,N_4108,N_4339);
nor U4782 (N_4782,N_4396,N_4420);
or U4783 (N_4783,N_4307,N_4298);
nand U4784 (N_4784,N_4259,N_4000);
or U4785 (N_4785,N_4443,N_4280);
or U4786 (N_4786,N_4334,N_4117);
nand U4787 (N_4787,N_4278,N_4357);
xor U4788 (N_4788,N_4402,N_4051);
xor U4789 (N_4789,N_4218,N_4260);
nor U4790 (N_4790,N_4257,N_4018);
xor U4791 (N_4791,N_4179,N_4455);
nand U4792 (N_4792,N_4343,N_4017);
nand U4793 (N_4793,N_4333,N_4418);
and U4794 (N_4794,N_4111,N_4138);
xor U4795 (N_4795,N_4496,N_4175);
and U4796 (N_4796,N_4435,N_4020);
nor U4797 (N_4797,N_4113,N_4376);
and U4798 (N_4798,N_4262,N_4011);
or U4799 (N_4799,N_4201,N_4422);
nor U4800 (N_4800,N_4229,N_4048);
nor U4801 (N_4801,N_4303,N_4211);
nor U4802 (N_4802,N_4405,N_4037);
nor U4803 (N_4803,N_4333,N_4197);
xor U4804 (N_4804,N_4017,N_4239);
or U4805 (N_4805,N_4280,N_4145);
nand U4806 (N_4806,N_4329,N_4451);
or U4807 (N_4807,N_4189,N_4449);
and U4808 (N_4808,N_4359,N_4168);
xor U4809 (N_4809,N_4176,N_4309);
and U4810 (N_4810,N_4079,N_4133);
nor U4811 (N_4811,N_4040,N_4404);
and U4812 (N_4812,N_4237,N_4022);
xnor U4813 (N_4813,N_4271,N_4151);
xnor U4814 (N_4814,N_4285,N_4187);
xor U4815 (N_4815,N_4475,N_4353);
nand U4816 (N_4816,N_4381,N_4074);
xor U4817 (N_4817,N_4499,N_4282);
nor U4818 (N_4818,N_4275,N_4463);
nand U4819 (N_4819,N_4314,N_4138);
nand U4820 (N_4820,N_4361,N_4331);
nor U4821 (N_4821,N_4313,N_4350);
nor U4822 (N_4822,N_4458,N_4181);
or U4823 (N_4823,N_4497,N_4174);
and U4824 (N_4824,N_4060,N_4281);
nor U4825 (N_4825,N_4251,N_4316);
xor U4826 (N_4826,N_4479,N_4239);
nor U4827 (N_4827,N_4036,N_4207);
or U4828 (N_4828,N_4322,N_4057);
and U4829 (N_4829,N_4005,N_4224);
nor U4830 (N_4830,N_4140,N_4480);
or U4831 (N_4831,N_4489,N_4470);
and U4832 (N_4832,N_4412,N_4446);
or U4833 (N_4833,N_4261,N_4292);
nand U4834 (N_4834,N_4218,N_4076);
and U4835 (N_4835,N_4062,N_4213);
or U4836 (N_4836,N_4108,N_4235);
nand U4837 (N_4837,N_4449,N_4325);
xnor U4838 (N_4838,N_4342,N_4154);
and U4839 (N_4839,N_4092,N_4188);
nand U4840 (N_4840,N_4364,N_4141);
nand U4841 (N_4841,N_4463,N_4446);
or U4842 (N_4842,N_4143,N_4084);
nor U4843 (N_4843,N_4217,N_4187);
or U4844 (N_4844,N_4056,N_4063);
nand U4845 (N_4845,N_4252,N_4182);
and U4846 (N_4846,N_4051,N_4330);
nor U4847 (N_4847,N_4112,N_4355);
and U4848 (N_4848,N_4382,N_4015);
xnor U4849 (N_4849,N_4404,N_4233);
nand U4850 (N_4850,N_4049,N_4297);
xnor U4851 (N_4851,N_4186,N_4158);
nand U4852 (N_4852,N_4072,N_4035);
nor U4853 (N_4853,N_4007,N_4227);
xor U4854 (N_4854,N_4128,N_4007);
and U4855 (N_4855,N_4134,N_4148);
nor U4856 (N_4856,N_4238,N_4289);
nand U4857 (N_4857,N_4097,N_4004);
xnor U4858 (N_4858,N_4486,N_4356);
nor U4859 (N_4859,N_4029,N_4028);
nor U4860 (N_4860,N_4117,N_4079);
or U4861 (N_4861,N_4423,N_4377);
xnor U4862 (N_4862,N_4292,N_4231);
nor U4863 (N_4863,N_4379,N_4052);
nor U4864 (N_4864,N_4209,N_4185);
and U4865 (N_4865,N_4208,N_4220);
or U4866 (N_4866,N_4010,N_4126);
and U4867 (N_4867,N_4247,N_4051);
nor U4868 (N_4868,N_4219,N_4303);
xor U4869 (N_4869,N_4170,N_4463);
or U4870 (N_4870,N_4243,N_4375);
and U4871 (N_4871,N_4370,N_4367);
or U4872 (N_4872,N_4490,N_4147);
nor U4873 (N_4873,N_4117,N_4003);
xor U4874 (N_4874,N_4173,N_4349);
xor U4875 (N_4875,N_4123,N_4038);
nor U4876 (N_4876,N_4401,N_4229);
and U4877 (N_4877,N_4099,N_4380);
nor U4878 (N_4878,N_4330,N_4225);
xor U4879 (N_4879,N_4215,N_4459);
nor U4880 (N_4880,N_4453,N_4199);
and U4881 (N_4881,N_4193,N_4251);
xor U4882 (N_4882,N_4119,N_4275);
xnor U4883 (N_4883,N_4248,N_4243);
or U4884 (N_4884,N_4282,N_4271);
nor U4885 (N_4885,N_4332,N_4360);
or U4886 (N_4886,N_4208,N_4076);
nand U4887 (N_4887,N_4182,N_4016);
and U4888 (N_4888,N_4012,N_4075);
and U4889 (N_4889,N_4115,N_4199);
and U4890 (N_4890,N_4211,N_4457);
xnor U4891 (N_4891,N_4317,N_4486);
and U4892 (N_4892,N_4467,N_4197);
or U4893 (N_4893,N_4291,N_4262);
xor U4894 (N_4894,N_4366,N_4499);
and U4895 (N_4895,N_4010,N_4013);
xor U4896 (N_4896,N_4384,N_4126);
nand U4897 (N_4897,N_4228,N_4036);
and U4898 (N_4898,N_4496,N_4023);
nor U4899 (N_4899,N_4448,N_4300);
xor U4900 (N_4900,N_4131,N_4204);
xor U4901 (N_4901,N_4397,N_4399);
nor U4902 (N_4902,N_4352,N_4084);
and U4903 (N_4903,N_4336,N_4010);
nor U4904 (N_4904,N_4089,N_4136);
and U4905 (N_4905,N_4360,N_4364);
and U4906 (N_4906,N_4221,N_4116);
xor U4907 (N_4907,N_4067,N_4182);
and U4908 (N_4908,N_4370,N_4337);
or U4909 (N_4909,N_4226,N_4067);
nand U4910 (N_4910,N_4486,N_4146);
xor U4911 (N_4911,N_4191,N_4249);
nor U4912 (N_4912,N_4320,N_4300);
or U4913 (N_4913,N_4065,N_4345);
nand U4914 (N_4914,N_4023,N_4080);
xnor U4915 (N_4915,N_4075,N_4424);
and U4916 (N_4916,N_4167,N_4389);
nand U4917 (N_4917,N_4370,N_4386);
and U4918 (N_4918,N_4373,N_4312);
xnor U4919 (N_4919,N_4311,N_4447);
xnor U4920 (N_4920,N_4165,N_4480);
or U4921 (N_4921,N_4137,N_4439);
and U4922 (N_4922,N_4007,N_4451);
nor U4923 (N_4923,N_4011,N_4413);
or U4924 (N_4924,N_4240,N_4077);
xor U4925 (N_4925,N_4492,N_4412);
nor U4926 (N_4926,N_4005,N_4315);
or U4927 (N_4927,N_4460,N_4173);
or U4928 (N_4928,N_4003,N_4005);
nor U4929 (N_4929,N_4407,N_4291);
xor U4930 (N_4930,N_4049,N_4394);
or U4931 (N_4931,N_4466,N_4487);
nor U4932 (N_4932,N_4466,N_4259);
xor U4933 (N_4933,N_4253,N_4177);
nor U4934 (N_4934,N_4169,N_4238);
or U4935 (N_4935,N_4178,N_4402);
nand U4936 (N_4936,N_4430,N_4393);
nor U4937 (N_4937,N_4301,N_4405);
xnor U4938 (N_4938,N_4413,N_4342);
or U4939 (N_4939,N_4044,N_4348);
or U4940 (N_4940,N_4014,N_4423);
and U4941 (N_4941,N_4316,N_4322);
nor U4942 (N_4942,N_4305,N_4443);
nor U4943 (N_4943,N_4001,N_4482);
nand U4944 (N_4944,N_4152,N_4197);
xnor U4945 (N_4945,N_4143,N_4064);
nor U4946 (N_4946,N_4338,N_4369);
or U4947 (N_4947,N_4104,N_4395);
or U4948 (N_4948,N_4139,N_4474);
or U4949 (N_4949,N_4294,N_4013);
and U4950 (N_4950,N_4024,N_4109);
xnor U4951 (N_4951,N_4255,N_4421);
and U4952 (N_4952,N_4275,N_4482);
nand U4953 (N_4953,N_4132,N_4217);
and U4954 (N_4954,N_4375,N_4492);
and U4955 (N_4955,N_4242,N_4162);
or U4956 (N_4956,N_4307,N_4095);
nor U4957 (N_4957,N_4157,N_4142);
or U4958 (N_4958,N_4248,N_4223);
or U4959 (N_4959,N_4062,N_4096);
nand U4960 (N_4960,N_4101,N_4410);
and U4961 (N_4961,N_4175,N_4217);
or U4962 (N_4962,N_4184,N_4035);
nor U4963 (N_4963,N_4338,N_4381);
nand U4964 (N_4964,N_4242,N_4413);
nand U4965 (N_4965,N_4393,N_4308);
xor U4966 (N_4966,N_4124,N_4334);
and U4967 (N_4967,N_4232,N_4092);
and U4968 (N_4968,N_4391,N_4051);
nand U4969 (N_4969,N_4128,N_4009);
nand U4970 (N_4970,N_4124,N_4022);
nand U4971 (N_4971,N_4272,N_4260);
nor U4972 (N_4972,N_4345,N_4382);
nor U4973 (N_4973,N_4440,N_4413);
or U4974 (N_4974,N_4268,N_4273);
xnor U4975 (N_4975,N_4383,N_4332);
xnor U4976 (N_4976,N_4290,N_4295);
xor U4977 (N_4977,N_4090,N_4131);
nand U4978 (N_4978,N_4076,N_4382);
nand U4979 (N_4979,N_4199,N_4039);
and U4980 (N_4980,N_4006,N_4251);
nor U4981 (N_4981,N_4316,N_4401);
xor U4982 (N_4982,N_4355,N_4009);
nand U4983 (N_4983,N_4346,N_4090);
nand U4984 (N_4984,N_4370,N_4381);
or U4985 (N_4985,N_4269,N_4209);
xnor U4986 (N_4986,N_4333,N_4284);
or U4987 (N_4987,N_4437,N_4192);
nor U4988 (N_4988,N_4476,N_4181);
nand U4989 (N_4989,N_4199,N_4180);
nand U4990 (N_4990,N_4487,N_4249);
and U4991 (N_4991,N_4441,N_4223);
and U4992 (N_4992,N_4250,N_4177);
or U4993 (N_4993,N_4040,N_4065);
nand U4994 (N_4994,N_4279,N_4416);
or U4995 (N_4995,N_4355,N_4136);
xnor U4996 (N_4996,N_4353,N_4304);
nor U4997 (N_4997,N_4474,N_4291);
and U4998 (N_4998,N_4042,N_4173);
or U4999 (N_4999,N_4188,N_4418);
and U5000 (N_5000,N_4569,N_4872);
nor U5001 (N_5001,N_4884,N_4821);
and U5002 (N_5002,N_4779,N_4896);
and U5003 (N_5003,N_4502,N_4622);
and U5004 (N_5004,N_4618,N_4905);
or U5005 (N_5005,N_4591,N_4557);
xor U5006 (N_5006,N_4841,N_4715);
nand U5007 (N_5007,N_4750,N_4631);
and U5008 (N_5008,N_4547,N_4735);
and U5009 (N_5009,N_4994,N_4516);
or U5010 (N_5010,N_4555,N_4558);
xnor U5011 (N_5011,N_4966,N_4991);
nor U5012 (N_5012,N_4962,N_4679);
and U5013 (N_5013,N_4746,N_4827);
nor U5014 (N_5014,N_4568,N_4504);
or U5015 (N_5015,N_4640,N_4623);
and U5016 (N_5016,N_4916,N_4990);
nand U5017 (N_5017,N_4778,N_4908);
nand U5018 (N_5018,N_4927,N_4606);
xnor U5019 (N_5019,N_4721,N_4712);
or U5020 (N_5020,N_4535,N_4984);
or U5021 (N_5021,N_4789,N_4621);
xnor U5022 (N_5022,N_4782,N_4880);
nor U5023 (N_5023,N_4726,N_4707);
xor U5024 (N_5024,N_4744,N_4545);
xor U5025 (N_5025,N_4722,N_4594);
or U5026 (N_5026,N_4826,N_4706);
xor U5027 (N_5027,N_4894,N_4743);
or U5028 (N_5028,N_4694,N_4757);
and U5029 (N_5029,N_4633,N_4992);
and U5030 (N_5030,N_4663,N_4929);
nand U5031 (N_5031,N_4532,N_4548);
nand U5032 (N_5032,N_4736,N_4833);
or U5033 (N_5033,N_4592,N_4509);
and U5034 (N_5034,N_4940,N_4514);
xor U5035 (N_5035,N_4745,N_4812);
or U5036 (N_5036,N_4588,N_4834);
nand U5037 (N_5037,N_4832,N_4564);
nor U5038 (N_5038,N_4787,N_4944);
nand U5039 (N_5039,N_4956,N_4703);
nand U5040 (N_5040,N_4737,N_4854);
or U5041 (N_5041,N_4711,N_4612);
xor U5042 (N_5042,N_4919,N_4915);
or U5043 (N_5043,N_4921,N_4772);
xnor U5044 (N_5044,N_4856,N_4732);
xnor U5045 (N_5045,N_4644,N_4760);
and U5046 (N_5046,N_4552,N_4646);
nor U5047 (N_5047,N_4936,N_4730);
or U5048 (N_5048,N_4563,N_4906);
nand U5049 (N_5049,N_4723,N_4943);
nand U5050 (N_5050,N_4926,N_4878);
and U5051 (N_5051,N_4501,N_4598);
nand U5052 (N_5052,N_4651,N_4574);
nand U5053 (N_5053,N_4752,N_4813);
and U5054 (N_5054,N_4815,N_4965);
or U5055 (N_5055,N_4979,N_4754);
and U5056 (N_5056,N_4907,N_4783);
nand U5057 (N_5057,N_4843,N_4603);
and U5058 (N_5058,N_4800,N_4851);
or U5059 (N_5059,N_4868,N_4579);
nand U5060 (N_5060,N_4852,N_4751);
nor U5061 (N_5061,N_4912,N_4528);
nor U5062 (N_5062,N_4611,N_4625);
and U5063 (N_5063,N_4533,N_4677);
or U5064 (N_5064,N_4734,N_4823);
and U5065 (N_5065,N_4518,N_4928);
and U5066 (N_5066,N_4945,N_4570);
and U5067 (N_5067,N_4550,N_4520);
and U5068 (N_5068,N_4681,N_4902);
xor U5069 (N_5069,N_4777,N_4881);
or U5070 (N_5070,N_4600,N_4567);
or U5071 (N_5071,N_4871,N_4521);
and U5072 (N_5072,N_4537,N_4585);
xor U5073 (N_5073,N_4627,N_4889);
or U5074 (N_5074,N_4717,N_4553);
nand U5075 (N_5075,N_4804,N_4785);
or U5076 (N_5076,N_4828,N_4716);
nand U5077 (N_5077,N_4937,N_4686);
and U5078 (N_5078,N_4581,N_4769);
nor U5079 (N_5079,N_4576,N_4503);
and U5080 (N_5080,N_4835,N_4885);
or U5081 (N_5081,N_4909,N_4764);
nand U5082 (N_5082,N_4903,N_4875);
and U5083 (N_5083,N_4948,N_4659);
nand U5084 (N_5084,N_4605,N_4808);
xor U5085 (N_5085,N_4977,N_4859);
or U5086 (N_5086,N_4914,N_4634);
or U5087 (N_5087,N_4515,N_4952);
nand U5088 (N_5088,N_4650,N_4687);
or U5089 (N_5089,N_4556,N_4742);
nor U5090 (N_5090,N_4930,N_4980);
xnor U5091 (N_5091,N_4900,N_4655);
nand U5092 (N_5092,N_4680,N_4572);
nand U5093 (N_5093,N_4628,N_4607);
nand U5094 (N_5094,N_4954,N_4517);
or U5095 (N_5095,N_4788,N_4719);
or U5096 (N_5096,N_4829,N_4850);
or U5097 (N_5097,N_4709,N_4697);
nor U5098 (N_5098,N_4846,N_4784);
nor U5099 (N_5099,N_4874,N_4791);
nand U5100 (N_5100,N_4656,N_4869);
or U5101 (N_5101,N_4961,N_4725);
nand U5102 (N_5102,N_4675,N_4566);
or U5103 (N_5103,N_4780,N_4773);
and U5104 (N_5104,N_4806,N_4708);
xnor U5105 (N_5105,N_4848,N_4538);
nor U5106 (N_5106,N_4599,N_4849);
or U5107 (N_5107,N_4797,N_4892);
xnor U5108 (N_5108,N_4536,N_4822);
or U5109 (N_5109,N_4638,N_4972);
and U5110 (N_5110,N_4811,N_4768);
or U5111 (N_5111,N_4584,N_4602);
xnor U5112 (N_5112,N_4761,N_4989);
nor U5113 (N_5113,N_4705,N_4786);
or U5114 (N_5114,N_4692,N_4809);
nor U5115 (N_5115,N_4624,N_4647);
and U5116 (N_5116,N_4910,N_4898);
nor U5117 (N_5117,N_4951,N_4941);
nand U5118 (N_5118,N_4747,N_4616);
and U5119 (N_5119,N_4855,N_4560);
or U5120 (N_5120,N_4601,N_4890);
or U5121 (N_5121,N_4924,N_4974);
nand U5122 (N_5122,N_4817,N_4544);
xor U5123 (N_5123,N_4571,N_4530);
or U5124 (N_5124,N_4527,N_4895);
xor U5125 (N_5125,N_4740,N_4939);
xnor U5126 (N_5126,N_4957,N_4559);
and U5127 (N_5127,N_4587,N_4993);
and U5128 (N_5128,N_4700,N_4714);
nand U5129 (N_5129,N_4513,N_4604);
and U5130 (N_5130,N_4645,N_4987);
or U5131 (N_5131,N_4887,N_4891);
and U5132 (N_5132,N_4539,N_4934);
nor U5133 (N_5133,N_4731,N_4920);
nor U5134 (N_5134,N_4767,N_4864);
or U5135 (N_5135,N_4801,N_4917);
xor U5136 (N_5136,N_4653,N_4798);
nand U5137 (N_5137,N_4583,N_4531);
xor U5138 (N_5138,N_4582,N_4971);
or U5139 (N_5139,N_4978,N_4674);
and U5140 (N_5140,N_4888,N_4728);
and U5141 (N_5141,N_4727,N_4932);
and U5142 (N_5142,N_4877,N_4613);
xor U5143 (N_5143,N_4771,N_4540);
nand U5144 (N_5144,N_4673,N_4671);
xor U5145 (N_5145,N_4549,N_4969);
nor U5146 (N_5146,N_4642,N_4672);
or U5147 (N_5147,N_4718,N_4838);
or U5148 (N_5148,N_4586,N_4844);
or U5149 (N_5149,N_4814,N_4762);
xnor U5150 (N_5150,N_4876,N_4639);
nor U5151 (N_5151,N_4997,N_4949);
or U5152 (N_5152,N_4635,N_4589);
and U5153 (N_5153,N_4577,N_4842);
nand U5154 (N_5154,N_4933,N_4820);
xnor U5155 (N_5155,N_4938,N_4996);
or U5156 (N_5156,N_4565,N_4657);
nor U5157 (N_5157,N_4925,N_4981);
xnor U5158 (N_5158,N_4665,N_4510);
and U5159 (N_5159,N_4955,N_4867);
and U5160 (N_5160,N_4873,N_4830);
xor U5161 (N_5161,N_4755,N_4632);
nand U5162 (N_5162,N_4541,N_4649);
or U5163 (N_5163,N_4946,N_4614);
nor U5164 (N_5164,N_4702,N_4662);
and U5165 (N_5165,N_4683,N_4654);
or U5166 (N_5166,N_4523,N_4652);
and U5167 (N_5167,N_4695,N_4668);
and U5168 (N_5168,N_4561,N_4629);
or U5169 (N_5169,N_4950,N_4865);
nand U5170 (N_5170,N_4790,N_4774);
nor U5171 (N_5171,N_4836,N_4696);
nor U5172 (N_5172,N_4999,N_4542);
nor U5173 (N_5173,N_4882,N_4562);
and U5174 (N_5174,N_4897,N_4636);
xor U5175 (N_5175,N_4983,N_4546);
nor U5176 (N_5176,N_4637,N_4597);
or U5177 (N_5177,N_4698,N_4682);
or U5178 (N_5178,N_4796,N_4879);
nand U5179 (N_5179,N_4522,N_4626);
and U5180 (N_5180,N_4739,N_4839);
or U5181 (N_5181,N_4641,N_4947);
xor U5182 (N_5182,N_4741,N_4967);
or U5183 (N_5183,N_4866,N_4863);
and U5184 (N_5184,N_4664,N_4781);
and U5185 (N_5185,N_4923,N_4942);
and U5186 (N_5186,N_4704,N_4505);
nand U5187 (N_5187,N_4795,N_4935);
and U5188 (N_5188,N_4543,N_4960);
nor U5189 (N_5189,N_4525,N_4508);
nand U5190 (N_5190,N_4985,N_4615);
nor U5191 (N_5191,N_4753,N_4918);
nand U5192 (N_5192,N_4710,N_4660);
xnor U5193 (N_5193,N_4529,N_4578);
nor U5194 (N_5194,N_4963,N_4775);
xnor U5195 (N_5195,N_4959,N_4630);
nand U5196 (N_5196,N_4699,N_4853);
xnor U5197 (N_5197,N_4575,N_4911);
xor U5198 (N_5198,N_4810,N_4860);
nor U5199 (N_5199,N_4619,N_4676);
nand U5200 (N_5200,N_4685,N_4512);
xor U5201 (N_5201,N_4968,N_4904);
nor U5202 (N_5202,N_4975,N_4701);
nor U5203 (N_5203,N_4958,N_4986);
and U5204 (N_5204,N_4953,N_4667);
nand U5205 (N_5205,N_4748,N_4617);
or U5206 (N_5206,N_4690,N_4551);
xor U5207 (N_5207,N_4913,N_4688);
or U5208 (N_5208,N_4973,N_4661);
and U5209 (N_5209,N_4770,N_4643);
or U5210 (N_5210,N_4759,N_4609);
nor U5211 (N_5211,N_4595,N_4608);
nor U5212 (N_5212,N_4519,N_4610);
nor U5213 (N_5213,N_4901,N_4729);
nor U5214 (N_5214,N_4893,N_4763);
nor U5215 (N_5215,N_4511,N_4819);
and U5216 (N_5216,N_4678,N_4824);
and U5217 (N_5217,N_4976,N_4837);
and U5218 (N_5218,N_4794,N_4807);
nand U5219 (N_5219,N_4816,N_4862);
or U5220 (N_5220,N_4720,N_4766);
nor U5221 (N_5221,N_4818,N_4803);
nand U5222 (N_5222,N_4666,N_4931);
and U5223 (N_5223,N_4506,N_4886);
and U5224 (N_5224,N_4669,N_4593);
and U5225 (N_5225,N_4713,N_4870);
xor U5226 (N_5226,N_4857,N_4684);
xnor U5227 (N_5227,N_4799,N_4825);
xnor U5228 (N_5228,N_4995,N_4765);
nand U5229 (N_5229,N_4861,N_4507);
and U5230 (N_5230,N_4524,N_4590);
xnor U5231 (N_5231,N_4749,N_4964);
nor U5232 (N_5232,N_4596,N_4738);
and U5233 (N_5233,N_4802,N_4776);
nand U5234 (N_5234,N_4756,N_4793);
nor U5235 (N_5235,N_4982,N_4580);
nand U5236 (N_5236,N_4847,N_4526);
nand U5237 (N_5237,N_4648,N_4554);
and U5238 (N_5238,N_4831,N_4970);
and U5239 (N_5239,N_4500,N_4840);
nor U5240 (N_5240,N_4922,N_4534);
nand U5241 (N_5241,N_4670,N_4805);
nor U5242 (N_5242,N_4689,N_4998);
nor U5243 (N_5243,N_4691,N_4620);
and U5244 (N_5244,N_4899,N_4733);
or U5245 (N_5245,N_4573,N_4792);
xnor U5246 (N_5246,N_4988,N_4658);
nand U5247 (N_5247,N_4724,N_4758);
xnor U5248 (N_5248,N_4858,N_4845);
or U5249 (N_5249,N_4883,N_4693);
nand U5250 (N_5250,N_4881,N_4773);
xnor U5251 (N_5251,N_4755,N_4731);
xor U5252 (N_5252,N_4525,N_4768);
nor U5253 (N_5253,N_4816,N_4961);
and U5254 (N_5254,N_4712,N_4528);
nor U5255 (N_5255,N_4982,N_4989);
and U5256 (N_5256,N_4514,N_4741);
nand U5257 (N_5257,N_4516,N_4870);
nand U5258 (N_5258,N_4554,N_4743);
nor U5259 (N_5259,N_4594,N_4654);
nand U5260 (N_5260,N_4690,N_4700);
xor U5261 (N_5261,N_4692,N_4745);
nor U5262 (N_5262,N_4907,N_4586);
nor U5263 (N_5263,N_4521,N_4873);
and U5264 (N_5264,N_4769,N_4507);
nor U5265 (N_5265,N_4906,N_4801);
nor U5266 (N_5266,N_4918,N_4890);
nor U5267 (N_5267,N_4997,N_4959);
nor U5268 (N_5268,N_4880,N_4721);
and U5269 (N_5269,N_4876,N_4589);
nor U5270 (N_5270,N_4851,N_4725);
nor U5271 (N_5271,N_4612,N_4691);
or U5272 (N_5272,N_4843,N_4594);
and U5273 (N_5273,N_4685,N_4977);
or U5274 (N_5274,N_4815,N_4999);
nor U5275 (N_5275,N_4844,N_4712);
nand U5276 (N_5276,N_4544,N_4919);
and U5277 (N_5277,N_4625,N_4699);
or U5278 (N_5278,N_4834,N_4958);
or U5279 (N_5279,N_4915,N_4746);
nand U5280 (N_5280,N_4520,N_4868);
or U5281 (N_5281,N_4781,N_4806);
nor U5282 (N_5282,N_4764,N_4538);
nand U5283 (N_5283,N_4750,N_4533);
nand U5284 (N_5284,N_4700,N_4650);
nand U5285 (N_5285,N_4796,N_4831);
nor U5286 (N_5286,N_4808,N_4571);
or U5287 (N_5287,N_4957,N_4977);
nand U5288 (N_5288,N_4777,N_4814);
nand U5289 (N_5289,N_4867,N_4513);
or U5290 (N_5290,N_4520,N_4584);
xnor U5291 (N_5291,N_4922,N_4946);
or U5292 (N_5292,N_4664,N_4918);
nor U5293 (N_5293,N_4805,N_4795);
xnor U5294 (N_5294,N_4556,N_4932);
nor U5295 (N_5295,N_4588,N_4727);
xor U5296 (N_5296,N_4750,N_4996);
nand U5297 (N_5297,N_4994,N_4951);
or U5298 (N_5298,N_4634,N_4797);
nand U5299 (N_5299,N_4735,N_4910);
xor U5300 (N_5300,N_4834,N_4727);
and U5301 (N_5301,N_4500,N_4950);
or U5302 (N_5302,N_4703,N_4783);
xor U5303 (N_5303,N_4874,N_4998);
xor U5304 (N_5304,N_4507,N_4939);
nor U5305 (N_5305,N_4581,N_4949);
xor U5306 (N_5306,N_4756,N_4518);
or U5307 (N_5307,N_4787,N_4672);
xor U5308 (N_5308,N_4952,N_4798);
nand U5309 (N_5309,N_4553,N_4922);
nor U5310 (N_5310,N_4813,N_4586);
nor U5311 (N_5311,N_4832,N_4833);
or U5312 (N_5312,N_4530,N_4636);
or U5313 (N_5313,N_4697,N_4586);
nand U5314 (N_5314,N_4708,N_4863);
nor U5315 (N_5315,N_4796,N_4704);
nor U5316 (N_5316,N_4999,N_4755);
nor U5317 (N_5317,N_4623,N_4680);
nand U5318 (N_5318,N_4725,N_4678);
nor U5319 (N_5319,N_4886,N_4809);
nor U5320 (N_5320,N_4865,N_4878);
nor U5321 (N_5321,N_4760,N_4935);
nor U5322 (N_5322,N_4813,N_4692);
and U5323 (N_5323,N_4577,N_4963);
nand U5324 (N_5324,N_4868,N_4965);
and U5325 (N_5325,N_4533,N_4870);
nor U5326 (N_5326,N_4714,N_4567);
xnor U5327 (N_5327,N_4563,N_4771);
xnor U5328 (N_5328,N_4808,N_4599);
or U5329 (N_5329,N_4827,N_4529);
and U5330 (N_5330,N_4931,N_4733);
and U5331 (N_5331,N_4612,N_4975);
or U5332 (N_5332,N_4722,N_4590);
or U5333 (N_5333,N_4526,N_4923);
nand U5334 (N_5334,N_4984,N_4544);
or U5335 (N_5335,N_4660,N_4667);
xnor U5336 (N_5336,N_4973,N_4682);
nor U5337 (N_5337,N_4657,N_4531);
nor U5338 (N_5338,N_4783,N_4776);
and U5339 (N_5339,N_4775,N_4647);
and U5340 (N_5340,N_4940,N_4885);
xor U5341 (N_5341,N_4592,N_4873);
xor U5342 (N_5342,N_4608,N_4714);
nand U5343 (N_5343,N_4748,N_4760);
nor U5344 (N_5344,N_4689,N_4611);
nor U5345 (N_5345,N_4675,N_4632);
and U5346 (N_5346,N_4697,N_4656);
nand U5347 (N_5347,N_4605,N_4765);
nand U5348 (N_5348,N_4797,N_4849);
and U5349 (N_5349,N_4874,N_4527);
and U5350 (N_5350,N_4789,N_4874);
xor U5351 (N_5351,N_4926,N_4876);
nor U5352 (N_5352,N_4766,N_4844);
nand U5353 (N_5353,N_4733,N_4563);
nand U5354 (N_5354,N_4896,N_4518);
nand U5355 (N_5355,N_4705,N_4611);
xnor U5356 (N_5356,N_4872,N_4984);
nor U5357 (N_5357,N_4991,N_4760);
or U5358 (N_5358,N_4561,N_4757);
nand U5359 (N_5359,N_4548,N_4914);
nand U5360 (N_5360,N_4890,N_4835);
xnor U5361 (N_5361,N_4501,N_4627);
and U5362 (N_5362,N_4569,N_4889);
or U5363 (N_5363,N_4694,N_4543);
nand U5364 (N_5364,N_4512,N_4975);
or U5365 (N_5365,N_4678,N_4796);
and U5366 (N_5366,N_4510,N_4764);
or U5367 (N_5367,N_4835,N_4831);
nand U5368 (N_5368,N_4687,N_4822);
nor U5369 (N_5369,N_4960,N_4930);
and U5370 (N_5370,N_4824,N_4749);
and U5371 (N_5371,N_4856,N_4938);
nand U5372 (N_5372,N_4574,N_4845);
nand U5373 (N_5373,N_4850,N_4726);
nor U5374 (N_5374,N_4736,N_4797);
nor U5375 (N_5375,N_4695,N_4950);
xnor U5376 (N_5376,N_4812,N_4624);
or U5377 (N_5377,N_4836,N_4600);
and U5378 (N_5378,N_4731,N_4790);
nand U5379 (N_5379,N_4902,N_4957);
nor U5380 (N_5380,N_4982,N_4591);
nand U5381 (N_5381,N_4752,N_4695);
nor U5382 (N_5382,N_4747,N_4787);
nor U5383 (N_5383,N_4954,N_4673);
nor U5384 (N_5384,N_4677,N_4973);
nor U5385 (N_5385,N_4979,N_4749);
nor U5386 (N_5386,N_4845,N_4510);
nand U5387 (N_5387,N_4874,N_4971);
or U5388 (N_5388,N_4564,N_4864);
or U5389 (N_5389,N_4660,N_4592);
xor U5390 (N_5390,N_4934,N_4675);
and U5391 (N_5391,N_4857,N_4703);
and U5392 (N_5392,N_4575,N_4839);
or U5393 (N_5393,N_4533,N_4608);
and U5394 (N_5394,N_4530,N_4561);
xnor U5395 (N_5395,N_4959,N_4846);
xor U5396 (N_5396,N_4721,N_4964);
xnor U5397 (N_5397,N_4737,N_4968);
or U5398 (N_5398,N_4982,N_4883);
or U5399 (N_5399,N_4796,N_4657);
nand U5400 (N_5400,N_4777,N_4710);
and U5401 (N_5401,N_4787,N_4517);
nand U5402 (N_5402,N_4896,N_4884);
nor U5403 (N_5403,N_4635,N_4945);
and U5404 (N_5404,N_4593,N_4655);
xnor U5405 (N_5405,N_4565,N_4568);
xnor U5406 (N_5406,N_4500,N_4771);
nand U5407 (N_5407,N_4698,N_4811);
nand U5408 (N_5408,N_4541,N_4859);
xor U5409 (N_5409,N_4608,N_4840);
xnor U5410 (N_5410,N_4744,N_4658);
nand U5411 (N_5411,N_4938,N_4837);
and U5412 (N_5412,N_4845,N_4649);
and U5413 (N_5413,N_4611,N_4899);
nor U5414 (N_5414,N_4791,N_4767);
nand U5415 (N_5415,N_4519,N_4722);
nand U5416 (N_5416,N_4685,N_4766);
or U5417 (N_5417,N_4832,N_4512);
nand U5418 (N_5418,N_4732,N_4575);
or U5419 (N_5419,N_4965,N_4711);
xnor U5420 (N_5420,N_4926,N_4977);
or U5421 (N_5421,N_4987,N_4978);
nor U5422 (N_5422,N_4544,N_4949);
and U5423 (N_5423,N_4609,N_4804);
or U5424 (N_5424,N_4852,N_4660);
nor U5425 (N_5425,N_4636,N_4943);
nand U5426 (N_5426,N_4846,N_4841);
or U5427 (N_5427,N_4903,N_4669);
xnor U5428 (N_5428,N_4900,N_4511);
xnor U5429 (N_5429,N_4935,N_4712);
or U5430 (N_5430,N_4956,N_4603);
xnor U5431 (N_5431,N_4687,N_4864);
and U5432 (N_5432,N_4633,N_4838);
or U5433 (N_5433,N_4541,N_4750);
nand U5434 (N_5434,N_4865,N_4634);
xnor U5435 (N_5435,N_4559,N_4811);
nor U5436 (N_5436,N_4857,N_4647);
nand U5437 (N_5437,N_4999,N_4916);
nor U5438 (N_5438,N_4713,N_4782);
nor U5439 (N_5439,N_4918,N_4795);
nand U5440 (N_5440,N_4986,N_4585);
or U5441 (N_5441,N_4661,N_4663);
nand U5442 (N_5442,N_4823,N_4867);
nor U5443 (N_5443,N_4866,N_4506);
xnor U5444 (N_5444,N_4750,N_4517);
nand U5445 (N_5445,N_4668,N_4827);
nor U5446 (N_5446,N_4559,N_4680);
and U5447 (N_5447,N_4884,N_4680);
or U5448 (N_5448,N_4604,N_4795);
and U5449 (N_5449,N_4509,N_4958);
and U5450 (N_5450,N_4944,N_4894);
xnor U5451 (N_5451,N_4681,N_4856);
or U5452 (N_5452,N_4825,N_4809);
nand U5453 (N_5453,N_4749,N_4848);
nand U5454 (N_5454,N_4786,N_4782);
and U5455 (N_5455,N_4511,N_4642);
or U5456 (N_5456,N_4870,N_4667);
xor U5457 (N_5457,N_4668,N_4984);
xor U5458 (N_5458,N_4872,N_4525);
or U5459 (N_5459,N_4667,N_4935);
or U5460 (N_5460,N_4781,N_4549);
or U5461 (N_5461,N_4695,N_4924);
xor U5462 (N_5462,N_4679,N_4515);
and U5463 (N_5463,N_4617,N_4540);
xnor U5464 (N_5464,N_4648,N_4680);
xor U5465 (N_5465,N_4666,N_4972);
or U5466 (N_5466,N_4667,N_4886);
nand U5467 (N_5467,N_4631,N_4562);
nand U5468 (N_5468,N_4807,N_4791);
xnor U5469 (N_5469,N_4813,N_4637);
nor U5470 (N_5470,N_4984,N_4930);
xor U5471 (N_5471,N_4542,N_4968);
nand U5472 (N_5472,N_4815,N_4980);
nor U5473 (N_5473,N_4580,N_4636);
nor U5474 (N_5474,N_4908,N_4789);
xor U5475 (N_5475,N_4564,N_4571);
nand U5476 (N_5476,N_4930,N_4894);
or U5477 (N_5477,N_4784,N_4965);
nor U5478 (N_5478,N_4779,N_4719);
nand U5479 (N_5479,N_4515,N_4625);
and U5480 (N_5480,N_4892,N_4944);
nor U5481 (N_5481,N_4649,N_4545);
xnor U5482 (N_5482,N_4895,N_4606);
xnor U5483 (N_5483,N_4779,N_4723);
or U5484 (N_5484,N_4565,N_4718);
nand U5485 (N_5485,N_4974,N_4591);
and U5486 (N_5486,N_4760,N_4761);
nand U5487 (N_5487,N_4753,N_4846);
xor U5488 (N_5488,N_4782,N_4528);
and U5489 (N_5489,N_4685,N_4981);
or U5490 (N_5490,N_4687,N_4660);
xnor U5491 (N_5491,N_4666,N_4709);
or U5492 (N_5492,N_4690,N_4889);
nand U5493 (N_5493,N_4797,N_4836);
and U5494 (N_5494,N_4884,N_4618);
nand U5495 (N_5495,N_4565,N_4766);
nand U5496 (N_5496,N_4545,N_4880);
or U5497 (N_5497,N_4632,N_4703);
nor U5498 (N_5498,N_4526,N_4828);
xnor U5499 (N_5499,N_4812,N_4876);
xnor U5500 (N_5500,N_5399,N_5119);
xor U5501 (N_5501,N_5162,N_5247);
and U5502 (N_5502,N_5023,N_5005);
xor U5503 (N_5503,N_5236,N_5206);
and U5504 (N_5504,N_5418,N_5033);
or U5505 (N_5505,N_5228,N_5131);
and U5506 (N_5506,N_5483,N_5268);
or U5507 (N_5507,N_5179,N_5043);
xor U5508 (N_5508,N_5322,N_5342);
xor U5509 (N_5509,N_5030,N_5263);
or U5510 (N_5510,N_5024,N_5360);
xor U5511 (N_5511,N_5185,N_5385);
or U5512 (N_5512,N_5312,N_5411);
nor U5513 (N_5513,N_5029,N_5413);
nand U5514 (N_5514,N_5383,N_5090);
and U5515 (N_5515,N_5428,N_5197);
or U5516 (N_5516,N_5126,N_5157);
xor U5517 (N_5517,N_5477,N_5438);
xor U5518 (N_5518,N_5432,N_5401);
xor U5519 (N_5519,N_5310,N_5417);
and U5520 (N_5520,N_5335,N_5020);
and U5521 (N_5521,N_5051,N_5192);
nand U5522 (N_5522,N_5077,N_5094);
or U5523 (N_5523,N_5098,N_5294);
or U5524 (N_5524,N_5371,N_5173);
or U5525 (N_5525,N_5048,N_5277);
or U5526 (N_5526,N_5425,N_5265);
nor U5527 (N_5527,N_5042,N_5149);
and U5528 (N_5528,N_5164,N_5245);
or U5529 (N_5529,N_5424,N_5221);
xor U5530 (N_5530,N_5158,N_5150);
and U5531 (N_5531,N_5229,N_5469);
and U5532 (N_5532,N_5456,N_5317);
or U5533 (N_5533,N_5487,N_5292);
and U5534 (N_5534,N_5073,N_5085);
or U5535 (N_5535,N_5047,N_5414);
xor U5536 (N_5536,N_5255,N_5121);
nand U5537 (N_5537,N_5234,N_5110);
or U5538 (N_5538,N_5352,N_5395);
xor U5539 (N_5539,N_5130,N_5106);
nor U5540 (N_5540,N_5052,N_5137);
and U5541 (N_5541,N_5187,N_5481);
nand U5542 (N_5542,N_5099,N_5434);
nand U5543 (N_5543,N_5114,N_5128);
nand U5544 (N_5544,N_5316,N_5061);
or U5545 (N_5545,N_5233,N_5348);
or U5546 (N_5546,N_5058,N_5412);
and U5547 (N_5547,N_5012,N_5146);
nand U5548 (N_5548,N_5186,N_5189);
or U5549 (N_5549,N_5443,N_5261);
or U5550 (N_5550,N_5135,N_5408);
xnor U5551 (N_5551,N_5423,N_5472);
or U5552 (N_5552,N_5046,N_5065);
xnor U5553 (N_5553,N_5470,N_5168);
or U5554 (N_5554,N_5444,N_5172);
nor U5555 (N_5555,N_5270,N_5184);
or U5556 (N_5556,N_5323,N_5384);
and U5557 (N_5557,N_5156,N_5226);
nor U5558 (N_5558,N_5392,N_5279);
xor U5559 (N_5559,N_5325,N_5321);
or U5560 (N_5560,N_5416,N_5116);
nor U5561 (N_5561,N_5243,N_5252);
xnor U5562 (N_5562,N_5393,N_5183);
xnor U5563 (N_5563,N_5091,N_5223);
and U5564 (N_5564,N_5057,N_5374);
and U5565 (N_5565,N_5329,N_5377);
and U5566 (N_5566,N_5108,N_5286);
xnor U5567 (N_5567,N_5476,N_5458);
and U5568 (N_5568,N_5295,N_5246);
xor U5569 (N_5569,N_5217,N_5080);
nor U5570 (N_5570,N_5358,N_5003);
nand U5571 (N_5571,N_5264,N_5153);
nor U5572 (N_5572,N_5349,N_5367);
or U5573 (N_5573,N_5039,N_5141);
nor U5574 (N_5574,N_5390,N_5379);
nand U5575 (N_5575,N_5288,N_5134);
or U5576 (N_5576,N_5467,N_5147);
or U5577 (N_5577,N_5207,N_5339);
xnor U5578 (N_5578,N_5350,N_5307);
nor U5579 (N_5579,N_5016,N_5182);
nor U5580 (N_5580,N_5239,N_5262);
and U5581 (N_5581,N_5082,N_5407);
and U5582 (N_5582,N_5142,N_5375);
xnor U5583 (N_5583,N_5070,N_5124);
xnor U5584 (N_5584,N_5087,N_5143);
or U5585 (N_5585,N_5249,N_5465);
nand U5586 (N_5586,N_5256,N_5449);
nand U5587 (N_5587,N_5370,N_5151);
and U5588 (N_5588,N_5479,N_5118);
xor U5589 (N_5589,N_5439,N_5355);
nand U5590 (N_5590,N_5362,N_5364);
or U5591 (N_5591,N_5299,N_5170);
nor U5592 (N_5592,N_5345,N_5426);
and U5593 (N_5593,N_5209,N_5171);
nor U5594 (N_5594,N_5204,N_5492);
or U5595 (N_5595,N_5244,N_5014);
xor U5596 (N_5596,N_5400,N_5336);
or U5597 (N_5597,N_5471,N_5049);
nor U5598 (N_5598,N_5420,N_5177);
xor U5599 (N_5599,N_5037,N_5340);
and U5600 (N_5600,N_5160,N_5290);
and U5601 (N_5601,N_5260,N_5457);
and U5602 (N_5602,N_5232,N_5396);
xnor U5603 (N_5603,N_5495,N_5344);
and U5604 (N_5604,N_5356,N_5284);
or U5605 (N_5605,N_5027,N_5011);
nand U5606 (N_5606,N_5123,N_5405);
or U5607 (N_5607,N_5103,N_5190);
nor U5608 (N_5608,N_5442,N_5009);
xor U5609 (N_5609,N_5044,N_5437);
nor U5610 (N_5610,N_5213,N_5330);
and U5611 (N_5611,N_5218,N_5025);
xnor U5612 (N_5612,N_5293,N_5369);
xor U5613 (N_5613,N_5271,N_5493);
or U5614 (N_5614,N_5034,N_5155);
nand U5615 (N_5615,N_5254,N_5165);
xor U5616 (N_5616,N_5109,N_5205);
nor U5617 (N_5617,N_5161,N_5274);
and U5618 (N_5618,N_5409,N_5459);
and U5619 (N_5619,N_5386,N_5282);
nand U5620 (N_5620,N_5445,N_5306);
nand U5621 (N_5621,N_5196,N_5113);
xnor U5622 (N_5622,N_5333,N_5188);
and U5623 (N_5623,N_5002,N_5427);
nand U5624 (N_5624,N_5068,N_5231);
and U5625 (N_5625,N_5324,N_5431);
or U5626 (N_5626,N_5104,N_5494);
xor U5627 (N_5627,N_5127,N_5117);
nand U5628 (N_5628,N_5314,N_5337);
and U5629 (N_5629,N_5305,N_5199);
nor U5630 (N_5630,N_5320,N_5269);
and U5631 (N_5631,N_5166,N_5436);
nor U5632 (N_5632,N_5328,N_5391);
and U5633 (N_5633,N_5019,N_5338);
or U5634 (N_5634,N_5191,N_5403);
nor U5635 (N_5635,N_5429,N_5266);
and U5636 (N_5636,N_5140,N_5482);
or U5637 (N_5637,N_5415,N_5010);
nor U5638 (N_5638,N_5389,N_5353);
and U5639 (N_5639,N_5067,N_5222);
nand U5640 (N_5640,N_5347,N_5300);
or U5641 (N_5641,N_5219,N_5096);
and U5642 (N_5642,N_5253,N_5346);
and U5643 (N_5643,N_5304,N_5394);
nand U5644 (N_5644,N_5071,N_5296);
and U5645 (N_5645,N_5132,N_5035);
or U5646 (N_5646,N_5298,N_5129);
and U5647 (N_5647,N_5361,N_5214);
nand U5648 (N_5648,N_5276,N_5022);
nor U5649 (N_5649,N_5251,N_5489);
xor U5650 (N_5650,N_5063,N_5194);
nor U5651 (N_5651,N_5102,N_5241);
or U5652 (N_5652,N_5101,N_5363);
nor U5653 (N_5653,N_5380,N_5210);
nor U5654 (N_5654,N_5062,N_5138);
nor U5655 (N_5655,N_5453,N_5499);
xor U5656 (N_5656,N_5258,N_5032);
nand U5657 (N_5657,N_5435,N_5167);
nor U5658 (N_5658,N_5451,N_5097);
and U5659 (N_5659,N_5287,N_5498);
xor U5660 (N_5660,N_5275,N_5125);
xor U5661 (N_5661,N_5064,N_5332);
and U5662 (N_5662,N_5454,N_5488);
and U5663 (N_5663,N_5175,N_5208);
and U5664 (N_5664,N_5159,N_5406);
or U5665 (N_5665,N_5163,N_5053);
nor U5666 (N_5666,N_5050,N_5017);
and U5667 (N_5667,N_5475,N_5169);
xor U5668 (N_5668,N_5297,N_5216);
nor U5669 (N_5669,N_5054,N_5315);
nor U5670 (N_5670,N_5013,N_5368);
nand U5671 (N_5671,N_5404,N_5031);
and U5672 (N_5672,N_5351,N_5319);
nand U5673 (N_5673,N_5430,N_5088);
nand U5674 (N_5674,N_5478,N_5397);
xnor U5675 (N_5675,N_5318,N_5302);
xnor U5676 (N_5676,N_5308,N_5285);
and U5677 (N_5677,N_5388,N_5281);
nand U5678 (N_5678,N_5200,N_5086);
and U5679 (N_5679,N_5001,N_5026);
xnor U5680 (N_5680,N_5484,N_5485);
or U5681 (N_5681,N_5291,N_5235);
nand U5682 (N_5682,N_5278,N_5497);
and U5683 (N_5683,N_5468,N_5331);
nor U5684 (N_5684,N_5075,N_5133);
or U5685 (N_5685,N_5452,N_5076);
nor U5686 (N_5686,N_5084,N_5461);
xor U5687 (N_5687,N_5107,N_5301);
or U5688 (N_5688,N_5230,N_5100);
or U5689 (N_5689,N_5176,N_5004);
xor U5690 (N_5690,N_5450,N_5083);
or U5691 (N_5691,N_5440,N_5242);
nand U5692 (N_5692,N_5365,N_5227);
nor U5693 (N_5693,N_5145,N_5174);
or U5694 (N_5694,N_5419,N_5008);
nor U5695 (N_5695,N_5382,N_5040);
nor U5696 (N_5696,N_5466,N_5021);
xnor U5697 (N_5697,N_5378,N_5248);
and U5698 (N_5698,N_5203,N_5343);
and U5699 (N_5699,N_5448,N_5366);
or U5700 (N_5700,N_5092,N_5240);
and U5701 (N_5701,N_5066,N_5491);
and U5702 (N_5702,N_5387,N_5211);
nand U5703 (N_5703,N_5373,N_5225);
xnor U5704 (N_5704,N_5000,N_5462);
or U5705 (N_5705,N_5273,N_5069);
and U5706 (N_5706,N_5354,N_5480);
xnor U5707 (N_5707,N_5224,N_5148);
or U5708 (N_5708,N_5036,N_5309);
xnor U5709 (N_5709,N_5311,N_5376);
or U5710 (N_5710,N_5015,N_5074);
nor U5711 (N_5711,N_5327,N_5144);
xor U5712 (N_5712,N_5154,N_5152);
nor U5713 (N_5713,N_5326,N_5357);
and U5714 (N_5714,N_5056,N_5112);
nand U5715 (N_5715,N_5195,N_5402);
nand U5716 (N_5716,N_5055,N_5202);
xor U5717 (N_5717,N_5267,N_5115);
or U5718 (N_5718,N_5095,N_5398);
and U5719 (N_5719,N_5093,N_5028);
and U5720 (N_5720,N_5089,N_5136);
nor U5721 (N_5721,N_5441,N_5060);
or U5722 (N_5722,N_5410,N_5198);
nor U5723 (N_5723,N_5111,N_5359);
xnor U5724 (N_5724,N_5180,N_5490);
nand U5725 (N_5725,N_5045,N_5341);
nand U5726 (N_5726,N_5238,N_5072);
nand U5727 (N_5727,N_5496,N_5259);
nand U5728 (N_5728,N_5422,N_5006);
xnor U5729 (N_5729,N_5193,N_5455);
or U5730 (N_5730,N_5059,N_5460);
and U5731 (N_5731,N_5303,N_5433);
xnor U5732 (N_5732,N_5122,N_5220);
xor U5733 (N_5733,N_5081,N_5041);
or U5734 (N_5734,N_5473,N_5381);
or U5735 (N_5735,N_5257,N_5105);
and U5736 (N_5736,N_5421,N_5486);
nor U5737 (N_5737,N_5139,N_5272);
nor U5738 (N_5738,N_5078,N_5446);
or U5739 (N_5739,N_5212,N_5447);
nand U5740 (N_5740,N_5283,N_5463);
xnor U5741 (N_5741,N_5215,N_5201);
nor U5742 (N_5742,N_5178,N_5120);
nand U5743 (N_5743,N_5038,N_5464);
nor U5744 (N_5744,N_5280,N_5181);
nor U5745 (N_5745,N_5334,N_5018);
nor U5746 (N_5746,N_5250,N_5372);
nand U5747 (N_5747,N_5007,N_5079);
nand U5748 (N_5748,N_5289,N_5313);
nor U5749 (N_5749,N_5474,N_5237);
xnor U5750 (N_5750,N_5151,N_5276);
nand U5751 (N_5751,N_5220,N_5367);
and U5752 (N_5752,N_5408,N_5110);
nand U5753 (N_5753,N_5039,N_5358);
xnor U5754 (N_5754,N_5189,N_5337);
nand U5755 (N_5755,N_5021,N_5248);
nand U5756 (N_5756,N_5477,N_5008);
nand U5757 (N_5757,N_5436,N_5217);
or U5758 (N_5758,N_5108,N_5344);
nand U5759 (N_5759,N_5430,N_5148);
or U5760 (N_5760,N_5318,N_5451);
xnor U5761 (N_5761,N_5365,N_5027);
nand U5762 (N_5762,N_5456,N_5381);
nand U5763 (N_5763,N_5179,N_5481);
xnor U5764 (N_5764,N_5315,N_5299);
and U5765 (N_5765,N_5356,N_5162);
xnor U5766 (N_5766,N_5272,N_5011);
nand U5767 (N_5767,N_5066,N_5227);
or U5768 (N_5768,N_5264,N_5129);
nand U5769 (N_5769,N_5343,N_5067);
and U5770 (N_5770,N_5423,N_5494);
nor U5771 (N_5771,N_5340,N_5000);
xor U5772 (N_5772,N_5410,N_5196);
and U5773 (N_5773,N_5068,N_5494);
and U5774 (N_5774,N_5073,N_5352);
and U5775 (N_5775,N_5279,N_5012);
or U5776 (N_5776,N_5384,N_5079);
and U5777 (N_5777,N_5110,N_5354);
nor U5778 (N_5778,N_5326,N_5241);
or U5779 (N_5779,N_5114,N_5009);
and U5780 (N_5780,N_5261,N_5351);
xnor U5781 (N_5781,N_5153,N_5327);
xnor U5782 (N_5782,N_5144,N_5157);
xnor U5783 (N_5783,N_5376,N_5157);
or U5784 (N_5784,N_5281,N_5003);
nor U5785 (N_5785,N_5284,N_5148);
or U5786 (N_5786,N_5476,N_5408);
nand U5787 (N_5787,N_5431,N_5153);
nand U5788 (N_5788,N_5291,N_5287);
and U5789 (N_5789,N_5142,N_5030);
nor U5790 (N_5790,N_5063,N_5494);
and U5791 (N_5791,N_5026,N_5432);
or U5792 (N_5792,N_5003,N_5309);
or U5793 (N_5793,N_5413,N_5449);
nand U5794 (N_5794,N_5176,N_5006);
xnor U5795 (N_5795,N_5179,N_5036);
nand U5796 (N_5796,N_5461,N_5116);
nor U5797 (N_5797,N_5349,N_5255);
xor U5798 (N_5798,N_5494,N_5035);
nor U5799 (N_5799,N_5057,N_5133);
nor U5800 (N_5800,N_5489,N_5342);
nor U5801 (N_5801,N_5318,N_5360);
and U5802 (N_5802,N_5332,N_5404);
nand U5803 (N_5803,N_5475,N_5194);
nand U5804 (N_5804,N_5251,N_5227);
xnor U5805 (N_5805,N_5031,N_5054);
xnor U5806 (N_5806,N_5194,N_5444);
xnor U5807 (N_5807,N_5375,N_5262);
nand U5808 (N_5808,N_5377,N_5022);
or U5809 (N_5809,N_5332,N_5475);
nand U5810 (N_5810,N_5103,N_5266);
xnor U5811 (N_5811,N_5384,N_5198);
nor U5812 (N_5812,N_5363,N_5380);
nand U5813 (N_5813,N_5389,N_5275);
nand U5814 (N_5814,N_5349,N_5392);
nand U5815 (N_5815,N_5401,N_5068);
and U5816 (N_5816,N_5064,N_5201);
nor U5817 (N_5817,N_5076,N_5430);
and U5818 (N_5818,N_5375,N_5134);
and U5819 (N_5819,N_5319,N_5065);
and U5820 (N_5820,N_5413,N_5118);
xnor U5821 (N_5821,N_5322,N_5191);
nand U5822 (N_5822,N_5022,N_5071);
or U5823 (N_5823,N_5080,N_5284);
xor U5824 (N_5824,N_5238,N_5255);
or U5825 (N_5825,N_5112,N_5172);
nor U5826 (N_5826,N_5450,N_5487);
or U5827 (N_5827,N_5159,N_5426);
xor U5828 (N_5828,N_5430,N_5403);
nand U5829 (N_5829,N_5114,N_5443);
or U5830 (N_5830,N_5308,N_5437);
nand U5831 (N_5831,N_5288,N_5234);
or U5832 (N_5832,N_5126,N_5487);
or U5833 (N_5833,N_5352,N_5103);
nand U5834 (N_5834,N_5193,N_5057);
or U5835 (N_5835,N_5283,N_5105);
nor U5836 (N_5836,N_5176,N_5150);
xnor U5837 (N_5837,N_5393,N_5005);
or U5838 (N_5838,N_5161,N_5458);
nor U5839 (N_5839,N_5375,N_5091);
xor U5840 (N_5840,N_5249,N_5024);
nor U5841 (N_5841,N_5039,N_5357);
nand U5842 (N_5842,N_5012,N_5191);
xor U5843 (N_5843,N_5028,N_5342);
nor U5844 (N_5844,N_5070,N_5110);
or U5845 (N_5845,N_5175,N_5394);
nor U5846 (N_5846,N_5208,N_5460);
nand U5847 (N_5847,N_5138,N_5195);
or U5848 (N_5848,N_5059,N_5332);
nand U5849 (N_5849,N_5269,N_5434);
or U5850 (N_5850,N_5337,N_5265);
or U5851 (N_5851,N_5110,N_5121);
and U5852 (N_5852,N_5013,N_5203);
xnor U5853 (N_5853,N_5272,N_5120);
or U5854 (N_5854,N_5012,N_5078);
or U5855 (N_5855,N_5369,N_5333);
nand U5856 (N_5856,N_5123,N_5332);
nor U5857 (N_5857,N_5157,N_5271);
nor U5858 (N_5858,N_5383,N_5130);
nor U5859 (N_5859,N_5437,N_5045);
nand U5860 (N_5860,N_5194,N_5472);
or U5861 (N_5861,N_5420,N_5296);
nor U5862 (N_5862,N_5150,N_5160);
and U5863 (N_5863,N_5465,N_5144);
nor U5864 (N_5864,N_5079,N_5068);
and U5865 (N_5865,N_5241,N_5344);
and U5866 (N_5866,N_5129,N_5293);
nor U5867 (N_5867,N_5322,N_5326);
xor U5868 (N_5868,N_5266,N_5469);
xor U5869 (N_5869,N_5183,N_5290);
xor U5870 (N_5870,N_5091,N_5271);
xor U5871 (N_5871,N_5382,N_5475);
xor U5872 (N_5872,N_5426,N_5074);
xnor U5873 (N_5873,N_5364,N_5310);
and U5874 (N_5874,N_5412,N_5144);
nand U5875 (N_5875,N_5389,N_5479);
and U5876 (N_5876,N_5007,N_5005);
and U5877 (N_5877,N_5180,N_5474);
nor U5878 (N_5878,N_5345,N_5177);
xnor U5879 (N_5879,N_5397,N_5166);
and U5880 (N_5880,N_5315,N_5321);
nand U5881 (N_5881,N_5497,N_5477);
nor U5882 (N_5882,N_5019,N_5129);
and U5883 (N_5883,N_5408,N_5096);
or U5884 (N_5884,N_5198,N_5393);
or U5885 (N_5885,N_5243,N_5450);
xnor U5886 (N_5886,N_5025,N_5129);
nor U5887 (N_5887,N_5308,N_5341);
or U5888 (N_5888,N_5450,N_5095);
or U5889 (N_5889,N_5211,N_5011);
or U5890 (N_5890,N_5401,N_5405);
and U5891 (N_5891,N_5093,N_5190);
nor U5892 (N_5892,N_5399,N_5290);
nand U5893 (N_5893,N_5378,N_5188);
nand U5894 (N_5894,N_5039,N_5415);
nor U5895 (N_5895,N_5212,N_5316);
and U5896 (N_5896,N_5152,N_5135);
xor U5897 (N_5897,N_5172,N_5347);
nand U5898 (N_5898,N_5137,N_5179);
xor U5899 (N_5899,N_5366,N_5320);
and U5900 (N_5900,N_5176,N_5033);
or U5901 (N_5901,N_5084,N_5490);
or U5902 (N_5902,N_5068,N_5080);
nor U5903 (N_5903,N_5488,N_5199);
nand U5904 (N_5904,N_5151,N_5133);
nor U5905 (N_5905,N_5374,N_5478);
nor U5906 (N_5906,N_5354,N_5478);
or U5907 (N_5907,N_5371,N_5166);
nand U5908 (N_5908,N_5298,N_5238);
xor U5909 (N_5909,N_5238,N_5350);
or U5910 (N_5910,N_5463,N_5418);
xnor U5911 (N_5911,N_5033,N_5402);
and U5912 (N_5912,N_5193,N_5291);
nor U5913 (N_5913,N_5294,N_5085);
or U5914 (N_5914,N_5119,N_5247);
nor U5915 (N_5915,N_5197,N_5291);
nor U5916 (N_5916,N_5378,N_5327);
xor U5917 (N_5917,N_5315,N_5025);
xnor U5918 (N_5918,N_5285,N_5088);
nor U5919 (N_5919,N_5098,N_5238);
or U5920 (N_5920,N_5408,N_5130);
or U5921 (N_5921,N_5090,N_5117);
nor U5922 (N_5922,N_5171,N_5442);
nor U5923 (N_5923,N_5080,N_5129);
xor U5924 (N_5924,N_5216,N_5015);
nand U5925 (N_5925,N_5480,N_5438);
or U5926 (N_5926,N_5149,N_5116);
and U5927 (N_5927,N_5384,N_5316);
xor U5928 (N_5928,N_5010,N_5193);
or U5929 (N_5929,N_5005,N_5315);
nor U5930 (N_5930,N_5182,N_5228);
and U5931 (N_5931,N_5137,N_5427);
or U5932 (N_5932,N_5202,N_5289);
and U5933 (N_5933,N_5090,N_5024);
xnor U5934 (N_5934,N_5077,N_5180);
nor U5935 (N_5935,N_5052,N_5158);
or U5936 (N_5936,N_5037,N_5178);
nor U5937 (N_5937,N_5254,N_5185);
xnor U5938 (N_5938,N_5429,N_5188);
nand U5939 (N_5939,N_5128,N_5366);
nor U5940 (N_5940,N_5290,N_5056);
and U5941 (N_5941,N_5424,N_5482);
nand U5942 (N_5942,N_5235,N_5394);
nand U5943 (N_5943,N_5225,N_5348);
or U5944 (N_5944,N_5261,N_5296);
or U5945 (N_5945,N_5394,N_5408);
and U5946 (N_5946,N_5148,N_5344);
nor U5947 (N_5947,N_5217,N_5311);
and U5948 (N_5948,N_5237,N_5166);
and U5949 (N_5949,N_5093,N_5416);
nor U5950 (N_5950,N_5227,N_5483);
nand U5951 (N_5951,N_5278,N_5130);
or U5952 (N_5952,N_5323,N_5280);
nand U5953 (N_5953,N_5267,N_5140);
xnor U5954 (N_5954,N_5415,N_5371);
and U5955 (N_5955,N_5037,N_5357);
or U5956 (N_5956,N_5201,N_5308);
or U5957 (N_5957,N_5281,N_5475);
and U5958 (N_5958,N_5309,N_5108);
or U5959 (N_5959,N_5431,N_5132);
nor U5960 (N_5960,N_5059,N_5407);
or U5961 (N_5961,N_5233,N_5082);
or U5962 (N_5962,N_5058,N_5101);
nor U5963 (N_5963,N_5182,N_5330);
nand U5964 (N_5964,N_5077,N_5329);
nand U5965 (N_5965,N_5467,N_5127);
nand U5966 (N_5966,N_5143,N_5115);
nand U5967 (N_5967,N_5265,N_5210);
nor U5968 (N_5968,N_5037,N_5375);
or U5969 (N_5969,N_5084,N_5472);
nand U5970 (N_5970,N_5108,N_5310);
xor U5971 (N_5971,N_5193,N_5459);
or U5972 (N_5972,N_5053,N_5285);
xnor U5973 (N_5973,N_5107,N_5207);
nor U5974 (N_5974,N_5346,N_5304);
nand U5975 (N_5975,N_5460,N_5471);
or U5976 (N_5976,N_5274,N_5458);
or U5977 (N_5977,N_5495,N_5315);
nor U5978 (N_5978,N_5051,N_5332);
nand U5979 (N_5979,N_5272,N_5256);
xor U5980 (N_5980,N_5052,N_5468);
xor U5981 (N_5981,N_5016,N_5478);
xnor U5982 (N_5982,N_5092,N_5023);
and U5983 (N_5983,N_5056,N_5253);
or U5984 (N_5984,N_5045,N_5199);
xnor U5985 (N_5985,N_5325,N_5186);
and U5986 (N_5986,N_5217,N_5172);
or U5987 (N_5987,N_5231,N_5151);
and U5988 (N_5988,N_5190,N_5281);
or U5989 (N_5989,N_5132,N_5264);
nor U5990 (N_5990,N_5276,N_5472);
nand U5991 (N_5991,N_5453,N_5120);
nand U5992 (N_5992,N_5037,N_5006);
xor U5993 (N_5993,N_5257,N_5358);
xor U5994 (N_5994,N_5376,N_5307);
xor U5995 (N_5995,N_5015,N_5039);
nor U5996 (N_5996,N_5293,N_5421);
xor U5997 (N_5997,N_5430,N_5044);
and U5998 (N_5998,N_5271,N_5402);
xnor U5999 (N_5999,N_5219,N_5148);
xor U6000 (N_6000,N_5542,N_5985);
xnor U6001 (N_6001,N_5883,N_5510);
xor U6002 (N_6002,N_5680,N_5647);
or U6003 (N_6003,N_5891,N_5743);
or U6004 (N_6004,N_5689,N_5988);
nor U6005 (N_6005,N_5601,N_5912);
nor U6006 (N_6006,N_5771,N_5563);
nand U6007 (N_6007,N_5640,N_5678);
and U6008 (N_6008,N_5858,N_5502);
and U6009 (N_6009,N_5557,N_5942);
xor U6010 (N_6010,N_5862,N_5797);
xnor U6011 (N_6011,N_5749,N_5781);
nand U6012 (N_6012,N_5984,N_5931);
and U6013 (N_6013,N_5802,N_5685);
and U6014 (N_6014,N_5614,N_5994);
xnor U6015 (N_6015,N_5998,N_5583);
nand U6016 (N_6016,N_5661,N_5795);
or U6017 (N_6017,N_5559,N_5698);
and U6018 (N_6018,N_5898,N_5788);
xnor U6019 (N_6019,N_5881,N_5709);
nor U6020 (N_6020,N_5700,N_5990);
nor U6021 (N_6021,N_5848,N_5969);
nor U6022 (N_6022,N_5522,N_5579);
nor U6023 (N_6023,N_5565,N_5524);
xnor U6024 (N_6024,N_5547,N_5977);
or U6025 (N_6025,N_5983,N_5777);
nand U6026 (N_6026,N_5918,N_5784);
xnor U6027 (N_6027,N_5529,N_5809);
and U6028 (N_6028,N_5785,N_5548);
or U6029 (N_6029,N_5663,N_5625);
nor U6030 (N_6030,N_5901,N_5842);
nand U6031 (N_6031,N_5699,N_5531);
xnor U6032 (N_6032,N_5824,N_5748);
nor U6033 (N_6033,N_5896,N_5948);
nor U6034 (N_6034,N_5925,N_5854);
nor U6035 (N_6035,N_5533,N_5880);
and U6036 (N_6036,N_5799,N_5725);
nand U6037 (N_6037,N_5742,N_5708);
nand U6038 (N_6038,N_5882,N_5782);
nand U6039 (N_6039,N_5778,N_5947);
xor U6040 (N_6040,N_5550,N_5933);
nor U6041 (N_6041,N_5597,N_5960);
and U6042 (N_6042,N_5512,N_5551);
xnor U6043 (N_6043,N_5852,N_5786);
or U6044 (N_6044,N_5779,N_5595);
nand U6045 (N_6045,N_5909,N_5615);
or U6046 (N_6046,N_5902,N_5835);
nor U6047 (N_6047,N_5818,N_5554);
nor U6048 (N_6048,N_5707,N_5874);
xnor U6049 (N_6049,N_5635,N_5847);
or U6050 (N_6050,N_5576,N_5613);
nand U6051 (N_6051,N_5666,N_5841);
nor U6052 (N_6052,N_5861,N_5922);
nor U6053 (N_6053,N_5754,N_5889);
xnor U6054 (N_6054,N_5975,N_5617);
or U6055 (N_6055,N_5683,N_5571);
or U6056 (N_6056,N_5637,N_5538);
or U6057 (N_6057,N_5812,N_5721);
or U6058 (N_6058,N_5506,N_5758);
and U6059 (N_6059,N_5991,N_5671);
nor U6060 (N_6060,N_5591,N_5829);
or U6061 (N_6061,N_5611,N_5935);
nand U6062 (N_6062,N_5703,N_5753);
and U6063 (N_6063,N_5780,N_5575);
nand U6064 (N_6064,N_5927,N_5573);
or U6065 (N_6065,N_5993,N_5610);
nor U6066 (N_6066,N_5627,N_5745);
nand U6067 (N_6067,N_5688,N_5772);
nor U6068 (N_6068,N_5769,N_5641);
nand U6069 (N_6069,N_5978,N_5855);
or U6070 (N_6070,N_5783,N_5820);
nand U6071 (N_6071,N_5645,N_5500);
nand U6072 (N_6072,N_5945,N_5530);
nor U6073 (N_6073,N_5845,N_5732);
nand U6074 (N_6074,N_5713,N_5814);
xnor U6075 (N_6075,N_5821,N_5652);
or U6076 (N_6076,N_5885,N_5787);
xor U6077 (N_6077,N_5875,N_5757);
xor U6078 (N_6078,N_5908,N_5914);
or U6079 (N_6079,N_5919,N_5718);
nor U6080 (N_6080,N_5599,N_5904);
nor U6081 (N_6081,N_5892,N_5752);
and U6082 (N_6082,N_5553,N_5924);
and U6083 (N_6083,N_5884,N_5876);
nand U6084 (N_6084,N_5936,N_5793);
and U6085 (N_6085,N_5744,N_5995);
and U6086 (N_6086,N_5537,N_5646);
and U6087 (N_6087,N_5629,N_5832);
nand U6088 (N_6088,N_5727,N_5955);
xnor U6089 (N_6089,N_5677,N_5593);
nor U6090 (N_6090,N_5711,N_5943);
nand U6091 (N_6091,N_5710,N_5886);
xor U6092 (N_6092,N_5736,N_5837);
and U6093 (N_6093,N_5655,N_5839);
or U6094 (N_6094,N_5740,N_5910);
nand U6095 (N_6095,N_5923,N_5584);
nor U6096 (N_6096,N_5650,N_5932);
xnor U6097 (N_6097,N_5967,N_5660);
xnor U6098 (N_6098,N_5776,N_5792);
xor U6099 (N_6099,N_5750,N_5761);
xor U6100 (N_6100,N_5760,N_5705);
nand U6101 (N_6101,N_5735,N_5774);
and U6102 (N_6102,N_5501,N_5695);
and U6103 (N_6103,N_5964,N_5622);
nand U6104 (N_6104,N_5519,N_5656);
nor U6105 (N_6105,N_5878,N_5746);
nand U6106 (N_6106,N_5976,N_5632);
nor U6107 (N_6107,N_5897,N_5596);
nor U6108 (N_6108,N_5694,N_5653);
or U6109 (N_6109,N_5903,N_5556);
xnor U6110 (N_6110,N_5719,N_5668);
or U6111 (N_6111,N_5962,N_5911);
nand U6112 (N_6112,N_5589,N_5765);
or U6113 (N_6113,N_5968,N_5941);
or U6114 (N_6114,N_5633,N_5569);
or U6115 (N_6115,N_5965,N_5838);
and U6116 (N_6116,N_5631,N_5513);
and U6117 (N_6117,N_5527,N_5895);
or U6118 (N_6118,N_5654,N_5686);
or U6119 (N_6119,N_5853,N_5980);
xor U6120 (N_6120,N_5828,N_5630);
nand U6121 (N_6121,N_5605,N_5626);
xnor U6122 (N_6122,N_5731,N_5511);
or U6123 (N_6123,N_5581,N_5851);
and U6124 (N_6124,N_5900,N_5602);
xnor U6125 (N_6125,N_5939,N_5737);
nor U6126 (N_6126,N_5940,N_5715);
and U6127 (N_6127,N_5712,N_5831);
nand U6128 (N_6128,N_5866,N_5893);
nor U6129 (N_6129,N_5937,N_5956);
or U6130 (N_6130,N_5649,N_5726);
or U6131 (N_6131,N_5616,N_5679);
and U6132 (N_6132,N_5864,N_5982);
nor U6133 (N_6133,N_5672,N_5681);
and U6134 (N_6134,N_5815,N_5578);
nand U6135 (N_6135,N_5624,N_5766);
nand U6136 (N_6136,N_5598,N_5791);
nor U6137 (N_6137,N_5534,N_5620);
nand U6138 (N_6138,N_5996,N_5526);
or U6139 (N_6139,N_5844,N_5926);
nor U6140 (N_6140,N_5734,N_5634);
and U6141 (N_6141,N_5850,N_5642);
or U6142 (N_6142,N_5849,N_5860);
nand U6143 (N_6143,N_5716,N_5808);
xor U6144 (N_6144,N_5644,N_5585);
and U6145 (N_6145,N_5868,N_5805);
xor U6146 (N_6146,N_5971,N_5833);
xor U6147 (N_6147,N_5768,N_5528);
and U6148 (N_6148,N_5676,N_5545);
or U6149 (N_6149,N_5609,N_5747);
or U6150 (N_6150,N_5917,N_5890);
or U6151 (N_6151,N_5669,N_5561);
or U6152 (N_6152,N_5973,N_5907);
and U6153 (N_6153,N_5504,N_5894);
or U6154 (N_6154,N_5773,N_5603);
and U6155 (N_6155,N_5525,N_5899);
xnor U6156 (N_6156,N_5834,N_5755);
xnor U6157 (N_6157,N_5830,N_5934);
or U6158 (N_6158,N_5639,N_5566);
nand U6159 (N_6159,N_5577,N_5564);
and U6160 (N_6160,N_5558,N_5836);
nor U6161 (N_6161,N_5872,N_5863);
nand U6162 (N_6162,N_5658,N_5612);
and U6163 (N_6163,N_5873,N_5811);
nand U6164 (N_6164,N_5540,N_5913);
nor U6165 (N_6165,N_5801,N_5509);
nor U6166 (N_6166,N_5870,N_5920);
nand U6167 (N_6167,N_5789,N_5687);
nor U6168 (N_6168,N_5505,N_5588);
nand U6169 (N_6169,N_5944,N_5972);
nand U6170 (N_6170,N_5767,N_5827);
nor U6171 (N_6171,N_5701,N_5572);
or U6172 (N_6172,N_5692,N_5515);
or U6173 (N_6173,N_5549,N_5704);
nor U6174 (N_6174,N_5775,N_5670);
or U6175 (N_6175,N_5921,N_5816);
or U6176 (N_6176,N_5963,N_5702);
xor U6177 (N_6177,N_5543,N_5722);
nor U6178 (N_6178,N_5696,N_5987);
nor U6179 (N_6179,N_5518,N_5877);
or U6180 (N_6180,N_5974,N_5954);
nand U6181 (N_6181,N_5667,N_5733);
and U6182 (N_6182,N_5590,N_5636);
nor U6183 (N_6183,N_5682,N_5800);
xnor U6184 (N_6184,N_5567,N_5856);
nor U6185 (N_6185,N_5706,N_5915);
nand U6186 (N_6186,N_5621,N_5807);
and U6187 (N_6187,N_5693,N_5790);
nor U6188 (N_6188,N_5675,N_5763);
or U6189 (N_6189,N_5981,N_5587);
xor U6190 (N_6190,N_5989,N_5532);
nand U6191 (N_6191,N_5846,N_5979);
or U6192 (N_6192,N_5729,N_5888);
and U6193 (N_6193,N_5720,N_5796);
nand U6194 (N_6194,N_5997,N_5823);
or U6195 (N_6195,N_5651,N_5826);
nor U6196 (N_6196,N_5552,N_5517);
and U6197 (N_6197,N_5813,N_5717);
or U6198 (N_6198,N_5619,N_5929);
xnor U6199 (N_6199,N_5887,N_5546);
or U6200 (N_6200,N_5560,N_5536);
nor U6201 (N_6201,N_5516,N_5810);
nor U6202 (N_6202,N_5674,N_5673);
xnor U6203 (N_6203,N_5503,N_5822);
or U6204 (N_6204,N_5999,N_5952);
xnor U6205 (N_6205,N_5508,N_5643);
nor U6206 (N_6206,N_5957,N_5825);
and U6207 (N_6207,N_5867,N_5865);
and U6208 (N_6208,N_5580,N_5770);
nand U6209 (N_6209,N_5574,N_5840);
xor U6210 (N_6210,N_5523,N_5623);
xor U6211 (N_6211,N_5930,N_5664);
or U6212 (N_6212,N_5756,N_5728);
or U6213 (N_6213,N_5938,N_5628);
and U6214 (N_6214,N_5905,N_5638);
xnor U6215 (N_6215,N_5544,N_5986);
xnor U6216 (N_6216,N_5568,N_5879);
and U6217 (N_6217,N_5950,N_5521);
and U6218 (N_6218,N_5662,N_5586);
and U6219 (N_6219,N_5541,N_5871);
or U6220 (N_6220,N_5859,N_5764);
xnor U6221 (N_6221,N_5738,N_5659);
nand U6222 (N_6222,N_5804,N_5514);
nor U6223 (N_6223,N_5958,N_5966);
nand U6224 (N_6224,N_5684,N_5592);
and U6225 (N_6225,N_5507,N_5697);
and U6226 (N_6226,N_5739,N_5535);
and U6227 (N_6227,N_5946,N_5562);
xor U6228 (N_6228,N_5843,N_5714);
nor U6229 (N_6229,N_5906,N_5723);
and U6230 (N_6230,N_5657,N_5690);
nand U6231 (N_6231,N_5600,N_5606);
and U6232 (N_6232,N_5992,N_5665);
nor U6233 (N_6233,N_5691,N_5970);
or U6234 (N_6234,N_5869,N_5570);
nand U6235 (N_6235,N_5594,N_5959);
and U6236 (N_6236,N_5741,N_5857);
nand U6237 (N_6237,N_5539,N_5604);
xnor U6238 (N_6238,N_5961,N_5817);
xnor U6239 (N_6239,N_5618,N_5648);
nand U6240 (N_6240,N_5928,N_5520);
nand U6241 (N_6241,N_5806,N_5762);
xnor U6242 (N_6242,N_5951,N_5751);
nor U6243 (N_6243,N_5949,N_5607);
xor U6244 (N_6244,N_5759,N_5803);
and U6245 (N_6245,N_5724,N_5819);
nand U6246 (N_6246,N_5794,N_5730);
nor U6247 (N_6247,N_5916,N_5555);
and U6248 (N_6248,N_5953,N_5582);
xor U6249 (N_6249,N_5608,N_5798);
nand U6250 (N_6250,N_5798,N_5750);
and U6251 (N_6251,N_5643,N_5749);
nor U6252 (N_6252,N_5540,N_5606);
nand U6253 (N_6253,N_5745,N_5952);
nand U6254 (N_6254,N_5510,N_5693);
xor U6255 (N_6255,N_5695,N_5542);
or U6256 (N_6256,N_5643,N_5688);
nand U6257 (N_6257,N_5768,N_5994);
and U6258 (N_6258,N_5614,N_5738);
or U6259 (N_6259,N_5978,N_5864);
nor U6260 (N_6260,N_5831,N_5997);
xor U6261 (N_6261,N_5804,N_5724);
nand U6262 (N_6262,N_5555,N_5960);
or U6263 (N_6263,N_5704,N_5867);
and U6264 (N_6264,N_5896,N_5529);
or U6265 (N_6265,N_5712,N_5770);
nand U6266 (N_6266,N_5828,N_5998);
nand U6267 (N_6267,N_5786,N_5531);
nand U6268 (N_6268,N_5959,N_5538);
or U6269 (N_6269,N_5714,N_5899);
nor U6270 (N_6270,N_5956,N_5878);
and U6271 (N_6271,N_5901,N_5827);
xor U6272 (N_6272,N_5518,N_5629);
and U6273 (N_6273,N_5757,N_5677);
nor U6274 (N_6274,N_5769,N_5982);
nor U6275 (N_6275,N_5771,N_5869);
xor U6276 (N_6276,N_5671,N_5807);
or U6277 (N_6277,N_5763,N_5950);
and U6278 (N_6278,N_5751,N_5845);
xnor U6279 (N_6279,N_5724,N_5764);
xor U6280 (N_6280,N_5675,N_5717);
nor U6281 (N_6281,N_5574,N_5800);
or U6282 (N_6282,N_5586,N_5599);
nor U6283 (N_6283,N_5905,N_5680);
nor U6284 (N_6284,N_5980,N_5921);
or U6285 (N_6285,N_5828,N_5875);
and U6286 (N_6286,N_5709,N_5965);
nand U6287 (N_6287,N_5703,N_5891);
xor U6288 (N_6288,N_5963,N_5690);
xor U6289 (N_6289,N_5690,N_5512);
or U6290 (N_6290,N_5965,N_5598);
or U6291 (N_6291,N_5760,N_5636);
xor U6292 (N_6292,N_5538,N_5524);
and U6293 (N_6293,N_5848,N_5715);
nand U6294 (N_6294,N_5800,N_5783);
xor U6295 (N_6295,N_5756,N_5570);
nor U6296 (N_6296,N_5743,N_5659);
and U6297 (N_6297,N_5927,N_5939);
and U6298 (N_6298,N_5782,N_5970);
nand U6299 (N_6299,N_5570,N_5819);
or U6300 (N_6300,N_5599,N_5676);
and U6301 (N_6301,N_5828,N_5751);
nand U6302 (N_6302,N_5699,N_5822);
xor U6303 (N_6303,N_5976,N_5731);
nor U6304 (N_6304,N_5690,N_5554);
nor U6305 (N_6305,N_5759,N_5578);
nor U6306 (N_6306,N_5775,N_5843);
nand U6307 (N_6307,N_5512,N_5794);
and U6308 (N_6308,N_5825,N_5567);
or U6309 (N_6309,N_5831,N_5858);
and U6310 (N_6310,N_5786,N_5773);
xor U6311 (N_6311,N_5948,N_5520);
nand U6312 (N_6312,N_5806,N_5825);
nand U6313 (N_6313,N_5700,N_5780);
or U6314 (N_6314,N_5510,N_5821);
nor U6315 (N_6315,N_5957,N_5533);
xor U6316 (N_6316,N_5632,N_5578);
xor U6317 (N_6317,N_5561,N_5689);
and U6318 (N_6318,N_5998,N_5506);
nor U6319 (N_6319,N_5507,N_5687);
xor U6320 (N_6320,N_5647,N_5602);
xnor U6321 (N_6321,N_5620,N_5858);
and U6322 (N_6322,N_5868,N_5833);
nor U6323 (N_6323,N_5551,N_5511);
nand U6324 (N_6324,N_5837,N_5615);
and U6325 (N_6325,N_5582,N_5700);
nor U6326 (N_6326,N_5984,N_5934);
or U6327 (N_6327,N_5600,N_5522);
nand U6328 (N_6328,N_5508,N_5757);
xor U6329 (N_6329,N_5850,N_5926);
nor U6330 (N_6330,N_5628,N_5826);
xor U6331 (N_6331,N_5952,N_5878);
nor U6332 (N_6332,N_5902,N_5863);
and U6333 (N_6333,N_5688,N_5840);
or U6334 (N_6334,N_5988,N_5573);
nand U6335 (N_6335,N_5840,N_5673);
nor U6336 (N_6336,N_5937,N_5640);
xor U6337 (N_6337,N_5721,N_5750);
or U6338 (N_6338,N_5655,N_5797);
nand U6339 (N_6339,N_5714,N_5915);
or U6340 (N_6340,N_5521,N_5571);
and U6341 (N_6341,N_5562,N_5853);
nand U6342 (N_6342,N_5900,N_5559);
nor U6343 (N_6343,N_5520,N_5910);
nor U6344 (N_6344,N_5697,N_5621);
or U6345 (N_6345,N_5687,N_5697);
nand U6346 (N_6346,N_5579,N_5703);
and U6347 (N_6347,N_5548,N_5997);
and U6348 (N_6348,N_5528,N_5556);
xor U6349 (N_6349,N_5511,N_5522);
nor U6350 (N_6350,N_5705,N_5964);
nand U6351 (N_6351,N_5602,N_5807);
nor U6352 (N_6352,N_5803,N_5823);
nand U6353 (N_6353,N_5757,N_5936);
and U6354 (N_6354,N_5968,N_5582);
nor U6355 (N_6355,N_5633,N_5590);
or U6356 (N_6356,N_5682,N_5962);
nor U6357 (N_6357,N_5598,N_5644);
and U6358 (N_6358,N_5676,N_5945);
nor U6359 (N_6359,N_5581,N_5601);
and U6360 (N_6360,N_5946,N_5650);
and U6361 (N_6361,N_5866,N_5731);
or U6362 (N_6362,N_5644,N_5880);
xor U6363 (N_6363,N_5767,N_5678);
and U6364 (N_6364,N_5615,N_5815);
nand U6365 (N_6365,N_5728,N_5532);
xnor U6366 (N_6366,N_5859,N_5793);
and U6367 (N_6367,N_5894,N_5631);
xor U6368 (N_6368,N_5948,N_5967);
or U6369 (N_6369,N_5557,N_5884);
or U6370 (N_6370,N_5949,N_5723);
and U6371 (N_6371,N_5834,N_5519);
or U6372 (N_6372,N_5582,N_5642);
or U6373 (N_6373,N_5901,N_5810);
or U6374 (N_6374,N_5852,N_5873);
or U6375 (N_6375,N_5676,N_5828);
or U6376 (N_6376,N_5572,N_5726);
nor U6377 (N_6377,N_5877,N_5555);
nand U6378 (N_6378,N_5697,N_5974);
nor U6379 (N_6379,N_5675,N_5780);
and U6380 (N_6380,N_5524,N_5902);
or U6381 (N_6381,N_5534,N_5664);
xnor U6382 (N_6382,N_5764,N_5741);
xor U6383 (N_6383,N_5672,N_5627);
or U6384 (N_6384,N_5965,N_5572);
or U6385 (N_6385,N_5893,N_5904);
and U6386 (N_6386,N_5669,N_5926);
nor U6387 (N_6387,N_5614,N_5885);
or U6388 (N_6388,N_5925,N_5915);
nor U6389 (N_6389,N_5552,N_5874);
nand U6390 (N_6390,N_5980,N_5670);
nor U6391 (N_6391,N_5938,N_5648);
and U6392 (N_6392,N_5516,N_5859);
xor U6393 (N_6393,N_5535,N_5642);
and U6394 (N_6394,N_5525,N_5763);
and U6395 (N_6395,N_5726,N_5667);
nand U6396 (N_6396,N_5879,N_5688);
nand U6397 (N_6397,N_5871,N_5761);
and U6398 (N_6398,N_5570,N_5581);
and U6399 (N_6399,N_5734,N_5802);
nor U6400 (N_6400,N_5931,N_5671);
xnor U6401 (N_6401,N_5948,N_5587);
and U6402 (N_6402,N_5985,N_5690);
xnor U6403 (N_6403,N_5934,N_5877);
nor U6404 (N_6404,N_5597,N_5849);
and U6405 (N_6405,N_5750,N_5937);
xor U6406 (N_6406,N_5917,N_5744);
nand U6407 (N_6407,N_5659,N_5877);
and U6408 (N_6408,N_5711,N_5739);
nor U6409 (N_6409,N_5515,N_5769);
xor U6410 (N_6410,N_5574,N_5774);
xor U6411 (N_6411,N_5713,N_5673);
xor U6412 (N_6412,N_5716,N_5694);
or U6413 (N_6413,N_5925,N_5514);
nor U6414 (N_6414,N_5567,N_5848);
nor U6415 (N_6415,N_5821,N_5912);
nor U6416 (N_6416,N_5843,N_5792);
xnor U6417 (N_6417,N_5618,N_5511);
or U6418 (N_6418,N_5922,N_5690);
or U6419 (N_6419,N_5693,N_5872);
xnor U6420 (N_6420,N_5510,N_5664);
and U6421 (N_6421,N_5512,N_5593);
nor U6422 (N_6422,N_5730,N_5571);
nor U6423 (N_6423,N_5912,N_5537);
and U6424 (N_6424,N_5873,N_5712);
nand U6425 (N_6425,N_5720,N_5578);
and U6426 (N_6426,N_5777,N_5526);
nand U6427 (N_6427,N_5653,N_5610);
nand U6428 (N_6428,N_5835,N_5520);
and U6429 (N_6429,N_5580,N_5992);
nand U6430 (N_6430,N_5555,N_5649);
and U6431 (N_6431,N_5973,N_5763);
and U6432 (N_6432,N_5641,N_5772);
xor U6433 (N_6433,N_5646,N_5718);
xnor U6434 (N_6434,N_5830,N_5928);
nor U6435 (N_6435,N_5907,N_5728);
or U6436 (N_6436,N_5990,N_5580);
or U6437 (N_6437,N_5577,N_5551);
xor U6438 (N_6438,N_5570,N_5500);
xnor U6439 (N_6439,N_5542,N_5713);
nand U6440 (N_6440,N_5715,N_5684);
nand U6441 (N_6441,N_5753,N_5897);
xor U6442 (N_6442,N_5809,N_5741);
and U6443 (N_6443,N_5688,N_5868);
nor U6444 (N_6444,N_5774,N_5562);
and U6445 (N_6445,N_5830,N_5601);
or U6446 (N_6446,N_5801,N_5790);
xnor U6447 (N_6447,N_5928,N_5936);
nor U6448 (N_6448,N_5536,N_5844);
xnor U6449 (N_6449,N_5549,N_5716);
xnor U6450 (N_6450,N_5844,N_5794);
nand U6451 (N_6451,N_5870,N_5676);
or U6452 (N_6452,N_5669,N_5672);
or U6453 (N_6453,N_5878,N_5644);
nand U6454 (N_6454,N_5584,N_5933);
nand U6455 (N_6455,N_5743,N_5593);
and U6456 (N_6456,N_5757,N_5995);
xor U6457 (N_6457,N_5857,N_5626);
nand U6458 (N_6458,N_5693,N_5871);
xor U6459 (N_6459,N_5563,N_5619);
and U6460 (N_6460,N_5909,N_5814);
or U6461 (N_6461,N_5512,N_5975);
nor U6462 (N_6462,N_5998,N_5700);
or U6463 (N_6463,N_5816,N_5682);
and U6464 (N_6464,N_5859,N_5657);
and U6465 (N_6465,N_5998,N_5590);
or U6466 (N_6466,N_5914,N_5864);
nor U6467 (N_6467,N_5567,N_5766);
or U6468 (N_6468,N_5577,N_5642);
and U6469 (N_6469,N_5502,N_5956);
nor U6470 (N_6470,N_5601,N_5660);
or U6471 (N_6471,N_5626,N_5661);
nor U6472 (N_6472,N_5656,N_5555);
and U6473 (N_6473,N_5875,N_5657);
nand U6474 (N_6474,N_5636,N_5543);
nor U6475 (N_6475,N_5984,N_5935);
nor U6476 (N_6476,N_5713,N_5541);
xnor U6477 (N_6477,N_5887,N_5617);
nor U6478 (N_6478,N_5859,N_5986);
and U6479 (N_6479,N_5581,N_5852);
nor U6480 (N_6480,N_5793,N_5598);
xnor U6481 (N_6481,N_5717,N_5953);
and U6482 (N_6482,N_5714,N_5845);
nor U6483 (N_6483,N_5753,N_5860);
or U6484 (N_6484,N_5637,N_5527);
xor U6485 (N_6485,N_5810,N_5980);
xor U6486 (N_6486,N_5778,N_5579);
nor U6487 (N_6487,N_5614,N_5513);
nor U6488 (N_6488,N_5889,N_5560);
and U6489 (N_6489,N_5593,N_5964);
xor U6490 (N_6490,N_5502,N_5809);
xor U6491 (N_6491,N_5747,N_5773);
nor U6492 (N_6492,N_5940,N_5501);
and U6493 (N_6493,N_5919,N_5849);
nand U6494 (N_6494,N_5610,N_5698);
xnor U6495 (N_6495,N_5762,N_5679);
or U6496 (N_6496,N_5620,N_5992);
nor U6497 (N_6497,N_5681,N_5750);
xor U6498 (N_6498,N_5904,N_5815);
nand U6499 (N_6499,N_5987,N_5945);
or U6500 (N_6500,N_6399,N_6075);
or U6501 (N_6501,N_6062,N_6108);
nand U6502 (N_6502,N_6230,N_6289);
nor U6503 (N_6503,N_6394,N_6268);
nand U6504 (N_6504,N_6372,N_6170);
nor U6505 (N_6505,N_6460,N_6453);
or U6506 (N_6506,N_6214,N_6169);
xnor U6507 (N_6507,N_6208,N_6336);
nand U6508 (N_6508,N_6191,N_6386);
nand U6509 (N_6509,N_6311,N_6498);
nand U6510 (N_6510,N_6163,N_6225);
and U6511 (N_6511,N_6217,N_6109);
nor U6512 (N_6512,N_6390,N_6067);
nor U6513 (N_6513,N_6165,N_6402);
and U6514 (N_6514,N_6448,N_6167);
nand U6515 (N_6515,N_6081,N_6377);
xor U6516 (N_6516,N_6398,N_6361);
nand U6517 (N_6517,N_6428,N_6357);
and U6518 (N_6518,N_6072,N_6138);
xnor U6519 (N_6519,N_6292,N_6481);
nand U6520 (N_6520,N_6478,N_6100);
or U6521 (N_6521,N_6181,N_6029);
or U6522 (N_6522,N_6309,N_6203);
or U6523 (N_6523,N_6254,N_6299);
xnor U6524 (N_6524,N_6199,N_6294);
xor U6525 (N_6525,N_6044,N_6452);
nand U6526 (N_6526,N_6284,N_6272);
nor U6527 (N_6527,N_6126,N_6008);
nor U6528 (N_6528,N_6283,N_6241);
and U6529 (N_6529,N_6302,N_6330);
and U6530 (N_6530,N_6485,N_6031);
nor U6531 (N_6531,N_6094,N_6347);
nand U6532 (N_6532,N_6133,N_6378);
nor U6533 (N_6533,N_6216,N_6016);
or U6534 (N_6534,N_6425,N_6183);
and U6535 (N_6535,N_6000,N_6104);
nor U6536 (N_6536,N_6212,N_6195);
xor U6537 (N_6537,N_6366,N_6397);
xor U6538 (N_6538,N_6451,N_6429);
nand U6539 (N_6539,N_6455,N_6221);
or U6540 (N_6540,N_6479,N_6105);
xnor U6541 (N_6541,N_6407,N_6079);
or U6542 (N_6542,N_6381,N_6318);
and U6543 (N_6543,N_6352,N_6269);
nand U6544 (N_6544,N_6063,N_6237);
or U6545 (N_6545,N_6238,N_6266);
or U6546 (N_6546,N_6112,N_6490);
nor U6547 (N_6547,N_6280,N_6323);
or U6548 (N_6548,N_6045,N_6436);
nand U6549 (N_6549,N_6279,N_6161);
or U6550 (N_6550,N_6246,N_6441);
and U6551 (N_6551,N_6058,N_6140);
nand U6552 (N_6552,N_6431,N_6022);
and U6553 (N_6553,N_6004,N_6301);
nor U6554 (N_6554,N_6445,N_6009);
or U6555 (N_6555,N_6414,N_6190);
and U6556 (N_6556,N_6337,N_6365);
and U6557 (N_6557,N_6276,N_6349);
nor U6558 (N_6558,N_6278,N_6093);
nand U6559 (N_6559,N_6229,N_6019);
xnor U6560 (N_6560,N_6182,N_6202);
xor U6561 (N_6561,N_6400,N_6052);
xor U6562 (N_6562,N_6111,N_6099);
or U6563 (N_6563,N_6113,N_6091);
or U6564 (N_6564,N_6332,N_6185);
and U6565 (N_6565,N_6495,N_6007);
nor U6566 (N_6566,N_6355,N_6486);
or U6567 (N_6567,N_6257,N_6427);
nor U6568 (N_6568,N_6315,N_6059);
nor U6569 (N_6569,N_6175,N_6442);
xor U6570 (N_6570,N_6321,N_6494);
or U6571 (N_6571,N_6340,N_6408);
nor U6572 (N_6572,N_6032,N_6382);
or U6573 (N_6573,N_6440,N_6159);
or U6574 (N_6574,N_6085,N_6135);
nand U6575 (N_6575,N_6086,N_6303);
or U6576 (N_6576,N_6128,N_6092);
nor U6577 (N_6577,N_6261,N_6350);
and U6578 (N_6578,N_6069,N_6136);
nor U6579 (N_6579,N_6065,N_6437);
nand U6580 (N_6580,N_6252,N_6018);
or U6581 (N_6581,N_6348,N_6375);
and U6582 (N_6582,N_6376,N_6148);
xor U6583 (N_6583,N_6173,N_6373);
nand U6584 (N_6584,N_6057,N_6468);
nor U6585 (N_6585,N_6459,N_6014);
xor U6586 (N_6586,N_6040,N_6047);
nand U6587 (N_6587,N_6061,N_6172);
and U6588 (N_6588,N_6450,N_6464);
nor U6589 (N_6589,N_6147,N_6404);
nor U6590 (N_6590,N_6473,N_6034);
and U6591 (N_6591,N_6213,N_6189);
nor U6592 (N_6592,N_6243,N_6412);
or U6593 (N_6593,N_6358,N_6168);
nor U6594 (N_6594,N_6090,N_6041);
nor U6595 (N_6595,N_6205,N_6291);
nand U6596 (N_6596,N_6070,N_6393);
or U6597 (N_6597,N_6368,N_6083);
nand U6598 (N_6598,N_6155,N_6433);
or U6599 (N_6599,N_6290,N_6422);
nor U6600 (N_6600,N_6298,N_6120);
nand U6601 (N_6601,N_6035,N_6462);
nand U6602 (N_6602,N_6258,N_6286);
or U6603 (N_6603,N_6364,N_6074);
xnor U6604 (N_6604,N_6265,N_6322);
or U6605 (N_6605,N_6320,N_6435);
and U6606 (N_6606,N_6124,N_6327);
xor U6607 (N_6607,N_6098,N_6219);
nor U6608 (N_6608,N_6475,N_6248);
xnor U6609 (N_6609,N_6305,N_6097);
nand U6610 (N_6610,N_6446,N_6489);
nand U6611 (N_6611,N_6162,N_6021);
nor U6612 (N_6612,N_6256,N_6369);
or U6613 (N_6613,N_6415,N_6343);
xnor U6614 (N_6614,N_6483,N_6263);
or U6615 (N_6615,N_6253,N_6068);
nor U6616 (N_6616,N_6324,N_6417);
and U6617 (N_6617,N_6432,N_6293);
nand U6618 (N_6618,N_6260,N_6288);
or U6619 (N_6619,N_6020,N_6131);
and U6620 (N_6620,N_6444,N_6331);
and U6621 (N_6621,N_6244,N_6472);
nand U6622 (N_6622,N_6319,N_6117);
nor U6623 (N_6623,N_6026,N_6344);
or U6624 (N_6624,N_6192,N_6329);
xnor U6625 (N_6625,N_6151,N_6024);
or U6626 (N_6626,N_6235,N_6210);
or U6627 (N_6627,N_6046,N_6143);
xnor U6628 (N_6628,N_6082,N_6411);
and U6629 (N_6629,N_6177,N_6122);
nor U6630 (N_6630,N_6346,N_6033);
or U6631 (N_6631,N_6255,N_6011);
or U6632 (N_6632,N_6048,N_6179);
nor U6633 (N_6633,N_6297,N_6410);
and U6634 (N_6634,N_6304,N_6461);
nand U6635 (N_6635,N_6234,N_6198);
xnor U6636 (N_6636,N_6457,N_6454);
nand U6637 (N_6637,N_6465,N_6353);
nand U6638 (N_6638,N_6474,N_6188);
and U6639 (N_6639,N_6132,N_6012);
nand U6640 (N_6640,N_6363,N_6267);
and U6641 (N_6641,N_6102,N_6273);
xor U6642 (N_6642,N_6326,N_6150);
xor U6643 (N_6643,N_6264,N_6333);
nor U6644 (N_6644,N_6447,N_6028);
or U6645 (N_6645,N_6206,N_6222);
and U6646 (N_6646,N_6129,N_6227);
and U6647 (N_6647,N_6491,N_6077);
or U6648 (N_6648,N_6002,N_6418);
and U6649 (N_6649,N_6017,N_6054);
or U6650 (N_6650,N_6317,N_6088);
and U6651 (N_6651,N_6335,N_6209);
xnor U6652 (N_6652,N_6421,N_6476);
nand U6653 (N_6653,N_6039,N_6463);
nand U6654 (N_6654,N_6371,N_6419);
nand U6655 (N_6655,N_6119,N_6171);
and U6656 (N_6656,N_6449,N_6275);
nand U6657 (N_6657,N_6114,N_6466);
or U6658 (N_6658,N_6379,N_6184);
nor U6659 (N_6659,N_6027,N_6176);
or U6660 (N_6660,N_6064,N_6080);
or U6661 (N_6661,N_6125,N_6409);
nand U6662 (N_6662,N_6477,N_6240);
nor U6663 (N_6663,N_6197,N_6313);
nand U6664 (N_6664,N_6001,N_6383);
nand U6665 (N_6665,N_6359,N_6285);
nand U6666 (N_6666,N_6201,N_6174);
nand U6667 (N_6667,N_6438,N_6010);
xnor U6668 (N_6668,N_6307,N_6396);
or U6669 (N_6669,N_6356,N_6277);
nand U6670 (N_6670,N_6430,N_6043);
xor U6671 (N_6671,N_6308,N_6089);
or U6672 (N_6672,N_6499,N_6193);
xnor U6673 (N_6673,N_6149,N_6194);
or U6674 (N_6674,N_6233,N_6484);
or U6675 (N_6675,N_6084,N_6127);
nand U6676 (N_6676,N_6496,N_6416);
nand U6677 (N_6677,N_6424,N_6367);
nand U6678 (N_6678,N_6005,N_6003);
and U6679 (N_6679,N_6134,N_6154);
xor U6680 (N_6680,N_6116,N_6239);
xnor U6681 (N_6681,N_6316,N_6049);
or U6682 (N_6682,N_6187,N_6482);
or U6683 (N_6683,N_6076,N_6232);
xor U6684 (N_6684,N_6456,N_6137);
and U6685 (N_6685,N_6078,N_6118);
nor U6686 (N_6686,N_6443,N_6110);
or U6687 (N_6687,N_6095,N_6388);
nor U6688 (N_6688,N_6215,N_6360);
xor U6689 (N_6689,N_6270,N_6392);
nand U6690 (N_6690,N_6351,N_6306);
nand U6691 (N_6691,N_6186,N_6287);
nand U6692 (N_6692,N_6025,N_6488);
nand U6693 (N_6693,N_6471,N_6341);
nand U6694 (N_6694,N_6247,N_6497);
or U6695 (N_6695,N_6158,N_6030);
nand U6696 (N_6696,N_6385,N_6242);
xnor U6697 (N_6697,N_6345,N_6395);
or U6698 (N_6698,N_6434,N_6180);
and U6699 (N_6699,N_6226,N_6493);
xor U6700 (N_6700,N_6339,N_6224);
nor U6701 (N_6701,N_6271,N_6391);
nor U6702 (N_6702,N_6439,N_6259);
nand U6703 (N_6703,N_6156,N_6338);
nand U6704 (N_6704,N_6055,N_6142);
or U6705 (N_6705,N_6312,N_6071);
or U6706 (N_6706,N_6211,N_6152);
nand U6707 (N_6707,N_6228,N_6096);
nand U6708 (N_6708,N_6387,N_6066);
nand U6709 (N_6709,N_6139,N_6153);
nand U6710 (N_6710,N_6141,N_6042);
and U6711 (N_6711,N_6051,N_6250);
or U6712 (N_6712,N_6374,N_6207);
and U6713 (N_6713,N_6458,N_6370);
nand U6714 (N_6714,N_6023,N_6231);
nor U6715 (N_6715,N_6121,N_6115);
and U6716 (N_6716,N_6362,N_6300);
nand U6717 (N_6717,N_6013,N_6492);
or U6718 (N_6718,N_6123,N_6406);
and U6719 (N_6719,N_6145,N_6087);
or U6720 (N_6720,N_6281,N_6314);
nor U6721 (N_6721,N_6144,N_6384);
and U6722 (N_6722,N_6470,N_6296);
nand U6723 (N_6723,N_6334,N_6251);
nor U6724 (N_6724,N_6423,N_6380);
and U6725 (N_6725,N_6420,N_6295);
xor U6726 (N_6726,N_6403,N_6200);
and U6727 (N_6727,N_6467,N_6354);
and U6728 (N_6728,N_6166,N_6325);
xor U6729 (N_6729,N_6157,N_6160);
and U6730 (N_6730,N_6274,N_6178);
nand U6731 (N_6731,N_6015,N_6037);
nand U6732 (N_6732,N_6164,N_6328);
nor U6733 (N_6733,N_6282,N_6060);
nor U6734 (N_6734,N_6073,N_6107);
nand U6735 (N_6735,N_6101,N_6196);
nand U6736 (N_6736,N_6006,N_6310);
and U6737 (N_6737,N_6223,N_6218);
xnor U6738 (N_6738,N_6038,N_6220);
xor U6739 (N_6739,N_6405,N_6401);
xor U6740 (N_6740,N_6245,N_6249);
or U6741 (N_6741,N_6036,N_6262);
nand U6742 (N_6742,N_6050,N_6236);
xnor U6743 (N_6743,N_6480,N_6204);
nand U6744 (N_6744,N_6146,N_6103);
and U6745 (N_6745,N_6342,N_6469);
or U6746 (N_6746,N_6413,N_6106);
xnor U6747 (N_6747,N_6053,N_6426);
xnor U6748 (N_6748,N_6389,N_6130);
or U6749 (N_6749,N_6487,N_6056);
xor U6750 (N_6750,N_6290,N_6077);
xnor U6751 (N_6751,N_6068,N_6094);
nor U6752 (N_6752,N_6318,N_6087);
or U6753 (N_6753,N_6085,N_6325);
and U6754 (N_6754,N_6080,N_6450);
xor U6755 (N_6755,N_6127,N_6454);
nand U6756 (N_6756,N_6478,N_6206);
nor U6757 (N_6757,N_6060,N_6336);
and U6758 (N_6758,N_6102,N_6001);
and U6759 (N_6759,N_6489,N_6244);
nor U6760 (N_6760,N_6325,N_6041);
xor U6761 (N_6761,N_6162,N_6325);
and U6762 (N_6762,N_6011,N_6100);
xor U6763 (N_6763,N_6335,N_6256);
or U6764 (N_6764,N_6271,N_6101);
nand U6765 (N_6765,N_6232,N_6039);
xor U6766 (N_6766,N_6447,N_6041);
nor U6767 (N_6767,N_6276,N_6160);
and U6768 (N_6768,N_6363,N_6166);
and U6769 (N_6769,N_6048,N_6111);
nor U6770 (N_6770,N_6200,N_6492);
xor U6771 (N_6771,N_6286,N_6115);
or U6772 (N_6772,N_6270,N_6379);
xnor U6773 (N_6773,N_6357,N_6001);
and U6774 (N_6774,N_6023,N_6064);
or U6775 (N_6775,N_6327,N_6261);
nand U6776 (N_6776,N_6148,N_6462);
nor U6777 (N_6777,N_6118,N_6291);
or U6778 (N_6778,N_6333,N_6078);
and U6779 (N_6779,N_6009,N_6150);
or U6780 (N_6780,N_6333,N_6349);
or U6781 (N_6781,N_6396,N_6447);
and U6782 (N_6782,N_6023,N_6082);
nand U6783 (N_6783,N_6250,N_6392);
or U6784 (N_6784,N_6161,N_6281);
nand U6785 (N_6785,N_6445,N_6198);
nor U6786 (N_6786,N_6491,N_6140);
or U6787 (N_6787,N_6389,N_6252);
and U6788 (N_6788,N_6491,N_6128);
or U6789 (N_6789,N_6406,N_6079);
xnor U6790 (N_6790,N_6287,N_6300);
and U6791 (N_6791,N_6439,N_6288);
or U6792 (N_6792,N_6216,N_6368);
nor U6793 (N_6793,N_6100,N_6206);
and U6794 (N_6794,N_6091,N_6363);
or U6795 (N_6795,N_6312,N_6079);
and U6796 (N_6796,N_6285,N_6156);
and U6797 (N_6797,N_6087,N_6023);
and U6798 (N_6798,N_6499,N_6466);
nor U6799 (N_6799,N_6058,N_6339);
nand U6800 (N_6800,N_6149,N_6219);
and U6801 (N_6801,N_6086,N_6202);
or U6802 (N_6802,N_6101,N_6089);
xor U6803 (N_6803,N_6346,N_6266);
and U6804 (N_6804,N_6489,N_6079);
and U6805 (N_6805,N_6176,N_6308);
and U6806 (N_6806,N_6288,N_6356);
and U6807 (N_6807,N_6263,N_6200);
xnor U6808 (N_6808,N_6130,N_6098);
nor U6809 (N_6809,N_6214,N_6315);
xor U6810 (N_6810,N_6145,N_6386);
nand U6811 (N_6811,N_6096,N_6246);
xor U6812 (N_6812,N_6351,N_6041);
nor U6813 (N_6813,N_6170,N_6299);
and U6814 (N_6814,N_6246,N_6036);
xor U6815 (N_6815,N_6339,N_6018);
nor U6816 (N_6816,N_6153,N_6435);
and U6817 (N_6817,N_6481,N_6149);
nor U6818 (N_6818,N_6131,N_6022);
nand U6819 (N_6819,N_6102,N_6465);
nand U6820 (N_6820,N_6172,N_6119);
and U6821 (N_6821,N_6170,N_6234);
nand U6822 (N_6822,N_6403,N_6112);
nand U6823 (N_6823,N_6044,N_6445);
or U6824 (N_6824,N_6263,N_6154);
and U6825 (N_6825,N_6326,N_6496);
nand U6826 (N_6826,N_6316,N_6439);
nor U6827 (N_6827,N_6315,N_6279);
xnor U6828 (N_6828,N_6077,N_6386);
nor U6829 (N_6829,N_6345,N_6226);
xnor U6830 (N_6830,N_6072,N_6002);
xor U6831 (N_6831,N_6052,N_6367);
nor U6832 (N_6832,N_6330,N_6292);
or U6833 (N_6833,N_6086,N_6203);
nand U6834 (N_6834,N_6468,N_6117);
xor U6835 (N_6835,N_6133,N_6027);
nor U6836 (N_6836,N_6339,N_6485);
xor U6837 (N_6837,N_6007,N_6312);
nor U6838 (N_6838,N_6176,N_6245);
nor U6839 (N_6839,N_6193,N_6047);
nand U6840 (N_6840,N_6381,N_6009);
or U6841 (N_6841,N_6369,N_6040);
nand U6842 (N_6842,N_6288,N_6228);
xnor U6843 (N_6843,N_6327,N_6051);
nor U6844 (N_6844,N_6493,N_6240);
and U6845 (N_6845,N_6433,N_6252);
xnor U6846 (N_6846,N_6482,N_6420);
or U6847 (N_6847,N_6085,N_6186);
nor U6848 (N_6848,N_6446,N_6328);
nor U6849 (N_6849,N_6370,N_6068);
or U6850 (N_6850,N_6140,N_6270);
nor U6851 (N_6851,N_6385,N_6347);
and U6852 (N_6852,N_6197,N_6294);
nand U6853 (N_6853,N_6227,N_6278);
or U6854 (N_6854,N_6270,N_6028);
and U6855 (N_6855,N_6125,N_6230);
or U6856 (N_6856,N_6108,N_6306);
nor U6857 (N_6857,N_6330,N_6129);
and U6858 (N_6858,N_6381,N_6473);
or U6859 (N_6859,N_6052,N_6297);
xor U6860 (N_6860,N_6234,N_6159);
nor U6861 (N_6861,N_6196,N_6106);
nor U6862 (N_6862,N_6380,N_6116);
xnor U6863 (N_6863,N_6484,N_6049);
nor U6864 (N_6864,N_6288,N_6480);
nor U6865 (N_6865,N_6486,N_6211);
or U6866 (N_6866,N_6024,N_6393);
or U6867 (N_6867,N_6341,N_6225);
nor U6868 (N_6868,N_6306,N_6041);
and U6869 (N_6869,N_6322,N_6090);
or U6870 (N_6870,N_6083,N_6242);
and U6871 (N_6871,N_6284,N_6172);
or U6872 (N_6872,N_6136,N_6440);
xor U6873 (N_6873,N_6081,N_6133);
and U6874 (N_6874,N_6360,N_6165);
nand U6875 (N_6875,N_6129,N_6428);
xnor U6876 (N_6876,N_6370,N_6081);
nor U6877 (N_6877,N_6407,N_6192);
nor U6878 (N_6878,N_6150,N_6069);
xor U6879 (N_6879,N_6242,N_6188);
and U6880 (N_6880,N_6081,N_6251);
xor U6881 (N_6881,N_6295,N_6403);
nand U6882 (N_6882,N_6452,N_6367);
or U6883 (N_6883,N_6051,N_6167);
nor U6884 (N_6884,N_6400,N_6209);
nor U6885 (N_6885,N_6419,N_6139);
nor U6886 (N_6886,N_6097,N_6471);
or U6887 (N_6887,N_6426,N_6068);
nand U6888 (N_6888,N_6210,N_6139);
nor U6889 (N_6889,N_6474,N_6431);
xor U6890 (N_6890,N_6165,N_6374);
nand U6891 (N_6891,N_6146,N_6400);
or U6892 (N_6892,N_6418,N_6145);
xor U6893 (N_6893,N_6482,N_6278);
nand U6894 (N_6894,N_6312,N_6352);
nor U6895 (N_6895,N_6076,N_6344);
xnor U6896 (N_6896,N_6245,N_6229);
or U6897 (N_6897,N_6459,N_6496);
xor U6898 (N_6898,N_6189,N_6101);
nor U6899 (N_6899,N_6107,N_6368);
xnor U6900 (N_6900,N_6479,N_6037);
or U6901 (N_6901,N_6035,N_6166);
nor U6902 (N_6902,N_6367,N_6200);
xnor U6903 (N_6903,N_6377,N_6169);
nand U6904 (N_6904,N_6201,N_6034);
nand U6905 (N_6905,N_6499,N_6266);
nor U6906 (N_6906,N_6336,N_6070);
nand U6907 (N_6907,N_6153,N_6378);
nor U6908 (N_6908,N_6108,N_6109);
and U6909 (N_6909,N_6242,N_6252);
and U6910 (N_6910,N_6439,N_6005);
xnor U6911 (N_6911,N_6293,N_6093);
nor U6912 (N_6912,N_6224,N_6209);
nor U6913 (N_6913,N_6261,N_6053);
or U6914 (N_6914,N_6258,N_6078);
xnor U6915 (N_6915,N_6325,N_6392);
or U6916 (N_6916,N_6304,N_6438);
or U6917 (N_6917,N_6467,N_6410);
nor U6918 (N_6918,N_6154,N_6433);
xnor U6919 (N_6919,N_6285,N_6478);
xnor U6920 (N_6920,N_6094,N_6328);
and U6921 (N_6921,N_6380,N_6399);
xnor U6922 (N_6922,N_6389,N_6459);
nand U6923 (N_6923,N_6241,N_6192);
xor U6924 (N_6924,N_6021,N_6001);
and U6925 (N_6925,N_6242,N_6165);
nor U6926 (N_6926,N_6457,N_6496);
and U6927 (N_6927,N_6082,N_6395);
nand U6928 (N_6928,N_6007,N_6470);
nand U6929 (N_6929,N_6321,N_6492);
nor U6930 (N_6930,N_6072,N_6207);
and U6931 (N_6931,N_6224,N_6327);
nor U6932 (N_6932,N_6084,N_6294);
nand U6933 (N_6933,N_6405,N_6449);
nand U6934 (N_6934,N_6216,N_6453);
nor U6935 (N_6935,N_6412,N_6268);
and U6936 (N_6936,N_6306,N_6173);
and U6937 (N_6937,N_6045,N_6263);
nor U6938 (N_6938,N_6378,N_6092);
nor U6939 (N_6939,N_6213,N_6182);
and U6940 (N_6940,N_6285,N_6243);
nor U6941 (N_6941,N_6268,N_6484);
nand U6942 (N_6942,N_6074,N_6145);
and U6943 (N_6943,N_6062,N_6337);
nor U6944 (N_6944,N_6313,N_6250);
xor U6945 (N_6945,N_6124,N_6133);
xor U6946 (N_6946,N_6287,N_6083);
nor U6947 (N_6947,N_6281,N_6179);
nand U6948 (N_6948,N_6437,N_6198);
and U6949 (N_6949,N_6492,N_6402);
nand U6950 (N_6950,N_6384,N_6427);
xnor U6951 (N_6951,N_6435,N_6164);
nand U6952 (N_6952,N_6104,N_6139);
or U6953 (N_6953,N_6049,N_6264);
nand U6954 (N_6954,N_6288,N_6103);
or U6955 (N_6955,N_6318,N_6354);
and U6956 (N_6956,N_6336,N_6186);
xnor U6957 (N_6957,N_6037,N_6218);
and U6958 (N_6958,N_6374,N_6277);
nor U6959 (N_6959,N_6087,N_6436);
nor U6960 (N_6960,N_6402,N_6272);
nor U6961 (N_6961,N_6486,N_6417);
nand U6962 (N_6962,N_6027,N_6066);
nand U6963 (N_6963,N_6012,N_6207);
or U6964 (N_6964,N_6175,N_6282);
nor U6965 (N_6965,N_6034,N_6414);
and U6966 (N_6966,N_6458,N_6373);
nand U6967 (N_6967,N_6220,N_6198);
nand U6968 (N_6968,N_6111,N_6325);
or U6969 (N_6969,N_6357,N_6115);
nand U6970 (N_6970,N_6261,N_6459);
and U6971 (N_6971,N_6203,N_6424);
and U6972 (N_6972,N_6053,N_6067);
and U6973 (N_6973,N_6200,N_6150);
xor U6974 (N_6974,N_6218,N_6498);
xnor U6975 (N_6975,N_6246,N_6489);
and U6976 (N_6976,N_6084,N_6374);
or U6977 (N_6977,N_6475,N_6160);
nand U6978 (N_6978,N_6483,N_6059);
xor U6979 (N_6979,N_6371,N_6012);
and U6980 (N_6980,N_6186,N_6381);
nand U6981 (N_6981,N_6453,N_6309);
nor U6982 (N_6982,N_6327,N_6245);
nand U6983 (N_6983,N_6199,N_6159);
and U6984 (N_6984,N_6415,N_6013);
or U6985 (N_6985,N_6320,N_6042);
and U6986 (N_6986,N_6097,N_6463);
or U6987 (N_6987,N_6033,N_6450);
nand U6988 (N_6988,N_6458,N_6355);
xnor U6989 (N_6989,N_6011,N_6450);
nand U6990 (N_6990,N_6368,N_6386);
xor U6991 (N_6991,N_6316,N_6083);
nor U6992 (N_6992,N_6271,N_6165);
and U6993 (N_6993,N_6382,N_6344);
nand U6994 (N_6994,N_6324,N_6052);
nor U6995 (N_6995,N_6259,N_6451);
or U6996 (N_6996,N_6121,N_6338);
and U6997 (N_6997,N_6468,N_6050);
and U6998 (N_6998,N_6366,N_6384);
xor U6999 (N_6999,N_6278,N_6095);
or U7000 (N_7000,N_6603,N_6869);
nand U7001 (N_7001,N_6846,N_6651);
and U7002 (N_7002,N_6828,N_6920);
and U7003 (N_7003,N_6726,N_6527);
nor U7004 (N_7004,N_6643,N_6905);
or U7005 (N_7005,N_6542,N_6978);
and U7006 (N_7006,N_6964,N_6916);
and U7007 (N_7007,N_6953,N_6788);
and U7008 (N_7008,N_6656,N_6973);
nor U7009 (N_7009,N_6545,N_6895);
nor U7010 (N_7010,N_6647,N_6981);
and U7011 (N_7011,N_6983,N_6810);
nand U7012 (N_7012,N_6717,N_6673);
nor U7013 (N_7013,N_6640,N_6525);
xnor U7014 (N_7014,N_6849,N_6989);
nand U7015 (N_7015,N_6734,N_6712);
nand U7016 (N_7016,N_6519,N_6777);
nand U7017 (N_7017,N_6757,N_6735);
nand U7018 (N_7018,N_6744,N_6679);
xnor U7019 (N_7019,N_6610,N_6677);
nor U7020 (N_7020,N_6618,N_6960);
and U7021 (N_7021,N_6838,N_6991);
xnor U7022 (N_7022,N_6945,N_6512);
nor U7023 (N_7023,N_6613,N_6641);
xnor U7024 (N_7024,N_6601,N_6770);
or U7025 (N_7025,N_6936,N_6522);
and U7026 (N_7026,N_6820,N_6795);
nor U7027 (N_7027,N_6886,N_6521);
or U7028 (N_7028,N_6811,N_6959);
nand U7029 (N_7029,N_6866,N_6763);
nor U7030 (N_7030,N_6695,N_6766);
xor U7031 (N_7031,N_6719,N_6848);
or U7032 (N_7032,N_6706,N_6546);
nand U7033 (N_7033,N_6721,N_6705);
nand U7034 (N_7034,N_6865,N_6885);
xor U7035 (N_7035,N_6720,N_6691);
xor U7036 (N_7036,N_6906,N_6778);
xor U7037 (N_7037,N_6535,N_6617);
nand U7038 (N_7038,N_6898,N_6941);
xor U7039 (N_7039,N_6834,N_6997);
nor U7040 (N_7040,N_6662,N_6680);
xnor U7041 (N_7041,N_6952,N_6919);
and U7042 (N_7042,N_6711,N_6917);
and U7043 (N_7043,N_6854,N_6665);
and U7044 (N_7044,N_6914,N_6873);
xor U7045 (N_7045,N_6551,N_6876);
and U7046 (N_7046,N_6929,N_6541);
nor U7047 (N_7047,N_6681,N_6765);
or U7048 (N_7048,N_6709,N_6903);
nor U7049 (N_7049,N_6825,N_6670);
and U7050 (N_7050,N_6716,N_6697);
xnor U7051 (N_7051,N_6867,N_6547);
xnor U7052 (N_7052,N_6657,N_6708);
nand U7053 (N_7053,N_6794,N_6597);
xnor U7054 (N_7054,N_6500,N_6600);
nor U7055 (N_7055,N_6782,N_6713);
or U7056 (N_7056,N_6570,N_6502);
nor U7057 (N_7057,N_6791,N_6571);
xnor U7058 (N_7058,N_6683,N_6559);
nor U7059 (N_7059,N_6769,N_6950);
xnor U7060 (N_7060,N_6969,N_6528);
nor U7061 (N_7061,N_6893,N_6944);
or U7062 (N_7062,N_6655,N_6624);
xnor U7063 (N_7063,N_6847,N_6799);
xor U7064 (N_7064,N_6575,N_6574);
nor U7065 (N_7065,N_6607,N_6890);
xor U7066 (N_7066,N_6646,N_6913);
and U7067 (N_7067,N_6722,N_6773);
and U7068 (N_7068,N_6622,N_6856);
nor U7069 (N_7069,N_6555,N_6779);
nand U7070 (N_7070,N_6988,N_6619);
xor U7071 (N_7071,N_6623,N_6503);
and U7072 (N_7072,N_6628,N_6768);
xnor U7073 (N_7073,N_6684,N_6654);
nor U7074 (N_7074,N_6967,N_6675);
nor U7075 (N_7075,N_6910,N_6669);
and U7076 (N_7076,N_6784,N_6518);
and U7077 (N_7077,N_6809,N_6668);
nand U7078 (N_7078,N_6862,N_6948);
nor U7079 (N_7079,N_6605,N_6998);
nor U7080 (N_7080,N_6614,N_6676);
or U7081 (N_7081,N_6965,N_6639);
nor U7082 (N_7082,N_6537,N_6790);
nand U7083 (N_7083,N_6753,N_6818);
nand U7084 (N_7084,N_6560,N_6736);
nor U7085 (N_7085,N_6933,N_6842);
xnor U7086 (N_7086,N_6700,N_6805);
and U7087 (N_7087,N_6531,N_6501);
nor U7088 (N_7088,N_6858,N_6615);
nand U7089 (N_7089,N_6850,N_6634);
nor U7090 (N_7090,N_6658,N_6844);
nand U7091 (N_7091,N_6909,N_6694);
xor U7092 (N_7092,N_6632,N_6940);
nand U7093 (N_7093,N_6772,N_6589);
and U7094 (N_7094,N_6663,N_6751);
nor U7095 (N_7095,N_6802,N_6693);
xnor U7096 (N_7096,N_6598,N_6715);
and U7097 (N_7097,N_6852,N_6934);
nand U7098 (N_7098,N_6892,N_6793);
or U7099 (N_7099,N_6888,N_6976);
nand U7100 (N_7100,N_6999,N_6509);
and U7101 (N_7101,N_6671,N_6556);
and U7102 (N_7102,N_6985,N_6733);
or U7103 (N_7103,N_6723,N_6877);
nor U7104 (N_7104,N_6748,N_6591);
xor U7105 (N_7105,N_6776,N_6907);
or U7106 (N_7106,N_6739,N_6507);
nand U7107 (N_7107,N_6760,N_6819);
xnor U7108 (N_7108,N_6650,N_6644);
or U7109 (N_7109,N_6621,N_6666);
nand U7110 (N_7110,N_6743,N_6841);
nor U7111 (N_7111,N_6817,N_6826);
nor U7112 (N_7112,N_6821,N_6963);
or U7113 (N_7113,N_6516,N_6652);
or U7114 (N_7114,N_6863,N_6786);
nor U7115 (N_7115,N_6755,N_6642);
and U7116 (N_7116,N_6543,N_6911);
xnor U7117 (N_7117,N_6878,N_6980);
and U7118 (N_7118,N_6554,N_6504);
nand U7119 (N_7119,N_6874,N_6861);
and U7120 (N_7120,N_6704,N_6583);
xor U7121 (N_7121,N_6979,N_6803);
and U7122 (N_7122,N_6882,N_6538);
or U7123 (N_7123,N_6667,N_6703);
nor U7124 (N_7124,N_6664,N_6569);
and U7125 (N_7125,N_6958,N_6520);
nand U7126 (N_7126,N_6742,N_6781);
nand U7127 (N_7127,N_6792,N_6517);
nor U7128 (N_7128,N_6899,N_6774);
and U7129 (N_7129,N_6672,N_6629);
or U7130 (N_7130,N_6686,N_6835);
xnor U7131 (N_7131,N_6824,N_6645);
nor U7132 (N_7132,N_6692,N_6937);
nor U7133 (N_7133,N_6827,N_6785);
or U7134 (N_7134,N_6689,N_6891);
xor U7135 (N_7135,N_6922,N_6631);
and U7136 (N_7136,N_6729,N_6630);
xnor U7137 (N_7137,N_6996,N_6956);
and U7138 (N_7138,N_6581,N_6690);
nand U7139 (N_7139,N_6699,N_6946);
nand U7140 (N_7140,N_6602,N_6864);
xnor U7141 (N_7141,N_6771,N_6539);
or U7142 (N_7142,N_6740,N_6764);
nand U7143 (N_7143,N_6725,N_6800);
xor U7144 (N_7144,N_6612,N_6579);
and U7145 (N_7145,N_6568,N_6935);
nand U7146 (N_7146,N_6883,N_6586);
and U7147 (N_7147,N_6696,N_6900);
or U7148 (N_7148,N_6975,N_6831);
nor U7149 (N_7149,N_6633,N_6566);
nor U7150 (N_7150,N_6808,N_6884);
nor U7151 (N_7151,N_6599,N_6904);
nor U7152 (N_7152,N_6529,N_6839);
nor U7153 (N_7153,N_6947,N_6731);
xor U7154 (N_7154,N_6972,N_6797);
nand U7155 (N_7155,N_6759,N_6505);
and U7156 (N_7156,N_6833,N_6747);
xnor U7157 (N_7157,N_6783,N_6550);
and U7158 (N_7158,N_6932,N_6995);
nand U7159 (N_7159,N_6648,N_6807);
or U7160 (N_7160,N_6564,N_6889);
or U7161 (N_7161,N_6840,N_6659);
nor U7162 (N_7162,N_6636,N_6604);
and U7163 (N_7163,N_6752,N_6620);
and U7164 (N_7164,N_6710,N_6548);
nand U7165 (N_7165,N_6931,N_6737);
nor U7166 (N_7166,N_6804,N_6506);
nand U7167 (N_7167,N_6993,N_6741);
xor U7168 (N_7168,N_6860,N_6596);
xor U7169 (N_7169,N_6724,N_6962);
nor U7170 (N_7170,N_6511,N_6971);
nand U7171 (N_7171,N_6609,N_6930);
xor U7172 (N_7172,N_6585,N_6749);
and U7173 (N_7173,N_6961,N_6822);
nand U7174 (N_7174,N_6510,N_6576);
xnor U7175 (N_7175,N_6938,N_6851);
xor U7176 (N_7176,N_6837,N_6756);
nand U7177 (N_7177,N_6966,N_6870);
xnor U7178 (N_7178,N_6801,N_6557);
and U7179 (N_7179,N_6578,N_6813);
nor U7180 (N_7180,N_6608,N_6942);
nand U7181 (N_7181,N_6682,N_6762);
and U7182 (N_7182,N_6881,N_6532);
or U7183 (N_7183,N_6754,N_6887);
or U7184 (N_7184,N_6515,N_6698);
and U7185 (N_7185,N_6927,N_6982);
and U7186 (N_7186,N_6926,N_6540);
and U7187 (N_7187,N_6745,N_6590);
nand U7188 (N_7188,N_6836,N_6627);
or U7189 (N_7189,N_6635,N_6787);
and U7190 (N_7190,N_6812,N_6879);
xnor U7191 (N_7191,N_6685,N_6949);
xnor U7192 (N_7192,N_6707,N_6625);
and U7193 (N_7193,N_6580,N_6536);
nand U7194 (N_7194,N_6990,N_6688);
or U7195 (N_7195,N_6746,N_6616);
xnor U7196 (N_7196,N_6855,N_6514);
or U7197 (N_7197,N_6524,N_6814);
nor U7198 (N_7198,N_6552,N_6563);
nor U7199 (N_7199,N_6859,N_6565);
nand U7200 (N_7200,N_6678,N_6951);
and U7201 (N_7201,N_6761,N_6939);
xnor U7202 (N_7202,N_6798,N_6845);
nand U7203 (N_7203,N_6830,N_6880);
nor U7204 (N_7204,N_6718,N_6796);
nor U7205 (N_7205,N_6611,N_6829);
and U7206 (N_7206,N_6606,N_6894);
nor U7207 (N_7207,N_6549,N_6558);
or U7208 (N_7208,N_6918,N_6595);
xor U7209 (N_7209,N_6815,N_6573);
and U7210 (N_7210,N_6533,N_6513);
nor U7211 (N_7211,N_6584,N_6572);
and U7212 (N_7212,N_6653,N_6561);
nand U7213 (N_7213,N_6730,N_6832);
nand U7214 (N_7214,N_6701,N_6994);
or U7215 (N_7215,N_6732,N_6902);
xnor U7216 (N_7216,N_6928,N_6577);
nand U7217 (N_7217,N_6530,N_6915);
and U7218 (N_7218,N_6875,N_6534);
xor U7219 (N_7219,N_6857,N_6526);
and U7220 (N_7220,N_6775,N_6508);
and U7221 (N_7221,N_6553,N_6871);
xnor U7222 (N_7222,N_6823,N_6780);
or U7223 (N_7223,N_6660,N_6955);
xor U7224 (N_7224,N_6587,N_6853);
nand U7225 (N_7225,N_6649,N_6702);
or U7226 (N_7226,N_6789,N_6957);
and U7227 (N_7227,N_6714,N_6974);
and U7228 (N_7228,N_6843,N_6727);
xnor U7229 (N_7229,N_6968,N_6872);
nor U7230 (N_7230,N_6562,N_6588);
xor U7231 (N_7231,N_6592,N_6901);
or U7232 (N_7232,N_6896,N_6924);
nand U7233 (N_7233,N_6816,N_6970);
xnor U7234 (N_7234,N_6674,N_6925);
or U7235 (N_7235,N_6921,N_6544);
nand U7236 (N_7236,N_6912,N_6567);
nand U7237 (N_7237,N_6767,N_6992);
and U7238 (N_7238,N_6593,N_6908);
or U7239 (N_7239,N_6758,N_6986);
or U7240 (N_7240,N_6661,N_6687);
or U7241 (N_7241,N_6977,N_6738);
nor U7242 (N_7242,N_6728,N_6806);
xor U7243 (N_7243,N_6638,N_6984);
and U7244 (N_7244,N_6868,N_6626);
and U7245 (N_7245,N_6582,N_6594);
and U7246 (N_7246,N_6897,N_6954);
nand U7247 (N_7247,N_6637,N_6923);
or U7248 (N_7248,N_6750,N_6943);
or U7249 (N_7249,N_6523,N_6987);
nor U7250 (N_7250,N_6953,N_6658);
or U7251 (N_7251,N_6517,N_6726);
xnor U7252 (N_7252,N_6955,N_6932);
or U7253 (N_7253,N_6822,N_6686);
and U7254 (N_7254,N_6996,N_6877);
xnor U7255 (N_7255,N_6578,N_6971);
xnor U7256 (N_7256,N_6974,N_6804);
and U7257 (N_7257,N_6538,N_6983);
nand U7258 (N_7258,N_6906,N_6946);
xor U7259 (N_7259,N_6622,N_6964);
and U7260 (N_7260,N_6737,N_6888);
nor U7261 (N_7261,N_6839,N_6991);
xor U7262 (N_7262,N_6973,N_6881);
or U7263 (N_7263,N_6651,N_6758);
xnor U7264 (N_7264,N_6820,N_6946);
nor U7265 (N_7265,N_6554,N_6660);
or U7266 (N_7266,N_6608,N_6627);
nor U7267 (N_7267,N_6535,N_6943);
and U7268 (N_7268,N_6982,N_6646);
and U7269 (N_7269,N_6948,N_6782);
and U7270 (N_7270,N_6755,N_6623);
nand U7271 (N_7271,N_6801,N_6799);
nand U7272 (N_7272,N_6586,N_6911);
or U7273 (N_7273,N_6715,N_6656);
nand U7274 (N_7274,N_6904,N_6817);
or U7275 (N_7275,N_6845,N_6649);
or U7276 (N_7276,N_6720,N_6714);
nand U7277 (N_7277,N_6788,N_6884);
xor U7278 (N_7278,N_6760,N_6515);
or U7279 (N_7279,N_6521,N_6854);
xnor U7280 (N_7280,N_6990,N_6649);
nand U7281 (N_7281,N_6847,N_6521);
or U7282 (N_7282,N_6627,N_6624);
nor U7283 (N_7283,N_6654,N_6895);
or U7284 (N_7284,N_6542,N_6806);
and U7285 (N_7285,N_6581,N_6995);
or U7286 (N_7286,N_6652,N_6986);
xnor U7287 (N_7287,N_6732,N_6944);
or U7288 (N_7288,N_6695,N_6737);
nor U7289 (N_7289,N_6810,N_6760);
nor U7290 (N_7290,N_6812,N_6760);
nand U7291 (N_7291,N_6531,N_6951);
or U7292 (N_7292,N_6576,N_6847);
and U7293 (N_7293,N_6866,N_6760);
nor U7294 (N_7294,N_6989,N_6767);
and U7295 (N_7295,N_6851,N_6904);
or U7296 (N_7296,N_6735,N_6900);
nand U7297 (N_7297,N_6924,N_6968);
and U7298 (N_7298,N_6516,N_6697);
nor U7299 (N_7299,N_6569,N_6502);
nor U7300 (N_7300,N_6914,N_6954);
xor U7301 (N_7301,N_6778,N_6803);
xnor U7302 (N_7302,N_6862,N_6966);
nor U7303 (N_7303,N_6519,N_6845);
and U7304 (N_7304,N_6749,N_6859);
or U7305 (N_7305,N_6768,N_6763);
or U7306 (N_7306,N_6745,N_6862);
and U7307 (N_7307,N_6909,N_6742);
or U7308 (N_7308,N_6508,N_6744);
and U7309 (N_7309,N_6800,N_6966);
or U7310 (N_7310,N_6575,N_6688);
nor U7311 (N_7311,N_6877,N_6981);
xor U7312 (N_7312,N_6587,N_6699);
nor U7313 (N_7313,N_6566,N_6653);
xnor U7314 (N_7314,N_6555,N_6580);
xor U7315 (N_7315,N_6874,N_6700);
or U7316 (N_7316,N_6540,N_6826);
and U7317 (N_7317,N_6633,N_6594);
and U7318 (N_7318,N_6584,N_6543);
nor U7319 (N_7319,N_6742,N_6838);
nand U7320 (N_7320,N_6881,N_6521);
or U7321 (N_7321,N_6792,N_6998);
nor U7322 (N_7322,N_6556,N_6886);
nor U7323 (N_7323,N_6912,N_6701);
and U7324 (N_7324,N_6533,N_6793);
nand U7325 (N_7325,N_6534,N_6919);
or U7326 (N_7326,N_6610,N_6944);
xor U7327 (N_7327,N_6834,N_6819);
and U7328 (N_7328,N_6863,N_6603);
xnor U7329 (N_7329,N_6821,N_6912);
nor U7330 (N_7330,N_6906,N_6805);
and U7331 (N_7331,N_6943,N_6749);
xnor U7332 (N_7332,N_6825,N_6520);
and U7333 (N_7333,N_6579,N_6627);
xnor U7334 (N_7334,N_6618,N_6836);
xnor U7335 (N_7335,N_6781,N_6626);
and U7336 (N_7336,N_6520,N_6614);
or U7337 (N_7337,N_6782,N_6813);
nor U7338 (N_7338,N_6603,N_6818);
or U7339 (N_7339,N_6571,N_6972);
nand U7340 (N_7340,N_6952,N_6740);
nand U7341 (N_7341,N_6545,N_6675);
nor U7342 (N_7342,N_6892,N_6840);
xor U7343 (N_7343,N_6526,N_6930);
nor U7344 (N_7344,N_6936,N_6928);
nor U7345 (N_7345,N_6970,N_6857);
and U7346 (N_7346,N_6675,N_6942);
xor U7347 (N_7347,N_6658,N_6819);
nand U7348 (N_7348,N_6946,N_6903);
nand U7349 (N_7349,N_6769,N_6696);
xnor U7350 (N_7350,N_6555,N_6583);
nand U7351 (N_7351,N_6605,N_6521);
nor U7352 (N_7352,N_6539,N_6816);
nor U7353 (N_7353,N_6556,N_6548);
and U7354 (N_7354,N_6592,N_6668);
xnor U7355 (N_7355,N_6822,N_6681);
nor U7356 (N_7356,N_6897,N_6623);
and U7357 (N_7357,N_6903,N_6583);
nor U7358 (N_7358,N_6507,N_6872);
xor U7359 (N_7359,N_6643,N_6595);
nor U7360 (N_7360,N_6800,N_6753);
and U7361 (N_7361,N_6530,N_6770);
or U7362 (N_7362,N_6762,N_6959);
and U7363 (N_7363,N_6986,N_6795);
xor U7364 (N_7364,N_6578,N_6848);
and U7365 (N_7365,N_6808,N_6933);
or U7366 (N_7366,N_6931,N_6860);
xnor U7367 (N_7367,N_6545,N_6871);
nor U7368 (N_7368,N_6823,N_6840);
nor U7369 (N_7369,N_6895,N_6928);
xnor U7370 (N_7370,N_6777,N_6629);
nor U7371 (N_7371,N_6883,N_6743);
xor U7372 (N_7372,N_6841,N_6599);
xor U7373 (N_7373,N_6902,N_6589);
nand U7374 (N_7374,N_6602,N_6662);
and U7375 (N_7375,N_6531,N_6827);
nor U7376 (N_7376,N_6593,N_6866);
nor U7377 (N_7377,N_6649,N_6792);
and U7378 (N_7378,N_6562,N_6587);
or U7379 (N_7379,N_6777,N_6724);
and U7380 (N_7380,N_6989,N_6938);
and U7381 (N_7381,N_6692,N_6816);
nand U7382 (N_7382,N_6598,N_6968);
nor U7383 (N_7383,N_6980,N_6611);
nand U7384 (N_7384,N_6666,N_6706);
and U7385 (N_7385,N_6526,N_6582);
nand U7386 (N_7386,N_6995,N_6545);
nor U7387 (N_7387,N_6803,N_6522);
and U7388 (N_7388,N_6586,N_6518);
nand U7389 (N_7389,N_6832,N_6983);
nand U7390 (N_7390,N_6574,N_6855);
nor U7391 (N_7391,N_6948,N_6827);
and U7392 (N_7392,N_6811,N_6759);
nand U7393 (N_7393,N_6945,N_6778);
or U7394 (N_7394,N_6510,N_6737);
xnor U7395 (N_7395,N_6506,N_6831);
nand U7396 (N_7396,N_6598,N_6704);
or U7397 (N_7397,N_6594,N_6770);
xnor U7398 (N_7398,N_6734,N_6908);
nor U7399 (N_7399,N_6583,N_6525);
or U7400 (N_7400,N_6777,N_6640);
and U7401 (N_7401,N_6943,N_6568);
nor U7402 (N_7402,N_6769,N_6704);
and U7403 (N_7403,N_6522,N_6854);
nand U7404 (N_7404,N_6738,N_6567);
or U7405 (N_7405,N_6683,N_6661);
nor U7406 (N_7406,N_6558,N_6979);
nand U7407 (N_7407,N_6641,N_6887);
or U7408 (N_7408,N_6621,N_6940);
xor U7409 (N_7409,N_6698,N_6635);
nor U7410 (N_7410,N_6688,N_6950);
nor U7411 (N_7411,N_6826,N_6755);
or U7412 (N_7412,N_6948,N_6922);
and U7413 (N_7413,N_6611,N_6961);
nand U7414 (N_7414,N_6650,N_6624);
and U7415 (N_7415,N_6992,N_6877);
nand U7416 (N_7416,N_6626,N_6516);
xnor U7417 (N_7417,N_6702,N_6966);
nor U7418 (N_7418,N_6713,N_6578);
nand U7419 (N_7419,N_6592,N_6547);
nand U7420 (N_7420,N_6929,N_6890);
xor U7421 (N_7421,N_6805,N_6547);
nor U7422 (N_7422,N_6765,N_6507);
nor U7423 (N_7423,N_6507,N_6782);
nor U7424 (N_7424,N_6813,N_6779);
xor U7425 (N_7425,N_6824,N_6668);
and U7426 (N_7426,N_6688,N_6881);
nand U7427 (N_7427,N_6846,N_6533);
xnor U7428 (N_7428,N_6726,N_6561);
or U7429 (N_7429,N_6845,N_6531);
nor U7430 (N_7430,N_6587,N_6532);
nor U7431 (N_7431,N_6967,N_6855);
and U7432 (N_7432,N_6752,N_6898);
and U7433 (N_7433,N_6703,N_6610);
nor U7434 (N_7434,N_6540,N_6727);
nor U7435 (N_7435,N_6615,N_6773);
nor U7436 (N_7436,N_6633,N_6671);
and U7437 (N_7437,N_6637,N_6730);
and U7438 (N_7438,N_6657,N_6555);
or U7439 (N_7439,N_6844,N_6879);
nor U7440 (N_7440,N_6655,N_6956);
xnor U7441 (N_7441,N_6515,N_6637);
or U7442 (N_7442,N_6530,N_6682);
and U7443 (N_7443,N_6944,N_6772);
and U7444 (N_7444,N_6897,N_6537);
nand U7445 (N_7445,N_6843,N_6812);
xor U7446 (N_7446,N_6779,N_6689);
xor U7447 (N_7447,N_6755,N_6943);
xor U7448 (N_7448,N_6565,N_6973);
nand U7449 (N_7449,N_6876,N_6792);
nor U7450 (N_7450,N_6685,N_6852);
or U7451 (N_7451,N_6889,N_6671);
nor U7452 (N_7452,N_6841,N_6766);
and U7453 (N_7453,N_6875,N_6987);
or U7454 (N_7454,N_6736,N_6950);
nor U7455 (N_7455,N_6883,N_6874);
and U7456 (N_7456,N_6972,N_6766);
nand U7457 (N_7457,N_6920,N_6989);
or U7458 (N_7458,N_6939,N_6777);
xnor U7459 (N_7459,N_6521,N_6936);
or U7460 (N_7460,N_6915,N_6565);
nor U7461 (N_7461,N_6902,N_6616);
and U7462 (N_7462,N_6655,N_6925);
or U7463 (N_7463,N_6887,N_6791);
and U7464 (N_7464,N_6686,N_6636);
nand U7465 (N_7465,N_6517,N_6522);
nand U7466 (N_7466,N_6752,N_6687);
nor U7467 (N_7467,N_6736,N_6826);
nor U7468 (N_7468,N_6602,N_6913);
or U7469 (N_7469,N_6607,N_6598);
nand U7470 (N_7470,N_6985,N_6945);
and U7471 (N_7471,N_6515,N_6998);
nand U7472 (N_7472,N_6865,N_6799);
nor U7473 (N_7473,N_6853,N_6966);
nand U7474 (N_7474,N_6599,N_6674);
nand U7475 (N_7475,N_6686,N_6921);
and U7476 (N_7476,N_6672,N_6867);
or U7477 (N_7477,N_6601,N_6872);
nor U7478 (N_7478,N_6806,N_6910);
nor U7479 (N_7479,N_6950,N_6549);
xor U7480 (N_7480,N_6721,N_6757);
and U7481 (N_7481,N_6558,N_6723);
xor U7482 (N_7482,N_6779,N_6907);
nand U7483 (N_7483,N_6852,N_6786);
nand U7484 (N_7484,N_6754,N_6910);
nor U7485 (N_7485,N_6564,N_6755);
or U7486 (N_7486,N_6572,N_6741);
and U7487 (N_7487,N_6632,N_6541);
and U7488 (N_7488,N_6806,N_6608);
xor U7489 (N_7489,N_6992,N_6589);
or U7490 (N_7490,N_6989,N_6559);
and U7491 (N_7491,N_6863,N_6598);
and U7492 (N_7492,N_6569,N_6601);
xnor U7493 (N_7493,N_6737,N_6939);
nor U7494 (N_7494,N_6538,N_6750);
xnor U7495 (N_7495,N_6591,N_6886);
or U7496 (N_7496,N_6595,N_6600);
and U7497 (N_7497,N_6959,N_6829);
and U7498 (N_7498,N_6622,N_6510);
nor U7499 (N_7499,N_6599,N_6748);
or U7500 (N_7500,N_7329,N_7420);
xnor U7501 (N_7501,N_7181,N_7139);
xnor U7502 (N_7502,N_7410,N_7497);
nand U7503 (N_7503,N_7268,N_7218);
and U7504 (N_7504,N_7494,N_7109);
nand U7505 (N_7505,N_7026,N_7284);
and U7506 (N_7506,N_7168,N_7438);
nand U7507 (N_7507,N_7290,N_7093);
xor U7508 (N_7508,N_7396,N_7449);
and U7509 (N_7509,N_7165,N_7355);
and U7510 (N_7510,N_7309,N_7276);
or U7511 (N_7511,N_7246,N_7205);
xor U7512 (N_7512,N_7445,N_7281);
xnor U7513 (N_7513,N_7316,N_7404);
and U7514 (N_7514,N_7248,N_7365);
nor U7515 (N_7515,N_7388,N_7482);
xnor U7516 (N_7516,N_7473,N_7015);
or U7517 (N_7517,N_7024,N_7237);
nor U7518 (N_7518,N_7287,N_7389);
and U7519 (N_7519,N_7000,N_7079);
or U7520 (N_7520,N_7417,N_7346);
nand U7521 (N_7521,N_7002,N_7190);
or U7522 (N_7522,N_7282,N_7435);
nand U7523 (N_7523,N_7127,N_7354);
nor U7524 (N_7524,N_7209,N_7336);
xnor U7525 (N_7525,N_7129,N_7498);
or U7526 (N_7526,N_7451,N_7308);
xnor U7527 (N_7527,N_7489,N_7342);
nand U7528 (N_7528,N_7334,N_7300);
nor U7529 (N_7529,N_7448,N_7469);
xnor U7530 (N_7530,N_7226,N_7235);
nand U7531 (N_7531,N_7245,N_7422);
xnor U7532 (N_7532,N_7278,N_7499);
nand U7533 (N_7533,N_7458,N_7399);
nor U7534 (N_7534,N_7359,N_7080);
nand U7535 (N_7535,N_7151,N_7046);
nand U7536 (N_7536,N_7124,N_7020);
or U7537 (N_7537,N_7186,N_7317);
nand U7538 (N_7538,N_7102,N_7457);
nand U7539 (N_7539,N_7207,N_7242);
and U7540 (N_7540,N_7006,N_7108);
xnor U7541 (N_7541,N_7089,N_7176);
or U7542 (N_7542,N_7374,N_7173);
xor U7543 (N_7543,N_7141,N_7042);
nor U7544 (N_7544,N_7189,N_7369);
nand U7545 (N_7545,N_7311,N_7440);
nand U7546 (N_7546,N_7164,N_7286);
or U7547 (N_7547,N_7312,N_7363);
nand U7548 (N_7548,N_7357,N_7013);
and U7549 (N_7549,N_7328,N_7044);
and U7550 (N_7550,N_7283,N_7279);
nand U7551 (N_7551,N_7107,N_7257);
nor U7552 (N_7552,N_7122,N_7274);
nor U7553 (N_7553,N_7091,N_7398);
or U7554 (N_7554,N_7431,N_7188);
nand U7555 (N_7555,N_7111,N_7126);
nor U7556 (N_7556,N_7432,N_7266);
or U7557 (N_7557,N_7063,N_7385);
nand U7558 (N_7558,N_7381,N_7053);
nor U7559 (N_7559,N_7455,N_7050);
xor U7560 (N_7560,N_7210,N_7043);
nor U7561 (N_7561,N_7201,N_7123);
and U7562 (N_7562,N_7153,N_7215);
nor U7563 (N_7563,N_7045,N_7411);
xnor U7564 (N_7564,N_7016,N_7262);
nand U7565 (N_7565,N_7267,N_7480);
nor U7566 (N_7566,N_7345,N_7040);
nor U7567 (N_7567,N_7027,N_7409);
or U7568 (N_7568,N_7038,N_7170);
nor U7569 (N_7569,N_7113,N_7330);
xnor U7570 (N_7570,N_7104,N_7012);
nor U7571 (N_7571,N_7483,N_7082);
nand U7572 (N_7572,N_7474,N_7072);
and U7573 (N_7573,N_7003,N_7150);
nor U7574 (N_7574,N_7019,N_7460);
and U7575 (N_7575,N_7228,N_7137);
and U7576 (N_7576,N_7280,N_7251);
nor U7577 (N_7577,N_7001,N_7378);
nor U7578 (N_7578,N_7264,N_7037);
and U7579 (N_7579,N_7491,N_7018);
xnor U7580 (N_7580,N_7254,N_7293);
nor U7581 (N_7581,N_7277,N_7306);
or U7582 (N_7582,N_7064,N_7232);
and U7583 (N_7583,N_7061,N_7412);
nor U7584 (N_7584,N_7339,N_7128);
and U7585 (N_7585,N_7476,N_7493);
nor U7586 (N_7586,N_7322,N_7094);
xnor U7587 (N_7587,N_7444,N_7343);
or U7588 (N_7588,N_7252,N_7405);
nand U7589 (N_7589,N_7090,N_7169);
nand U7590 (N_7590,N_7041,N_7115);
xor U7591 (N_7591,N_7211,N_7352);
or U7592 (N_7592,N_7022,N_7059);
nand U7593 (N_7593,N_7350,N_7275);
nand U7594 (N_7594,N_7301,N_7477);
and U7595 (N_7595,N_7179,N_7010);
xnor U7596 (N_7596,N_7307,N_7233);
or U7597 (N_7597,N_7344,N_7028);
xor U7598 (N_7598,N_7361,N_7486);
nor U7599 (N_7599,N_7305,N_7120);
nand U7600 (N_7600,N_7341,N_7263);
nand U7601 (N_7601,N_7400,N_7145);
xor U7602 (N_7602,N_7078,N_7056);
or U7603 (N_7603,N_7394,N_7291);
nor U7604 (N_7604,N_7067,N_7005);
or U7605 (N_7605,N_7429,N_7348);
and U7606 (N_7606,N_7244,N_7017);
or U7607 (N_7607,N_7464,N_7426);
xnor U7608 (N_7608,N_7321,N_7324);
or U7609 (N_7609,N_7358,N_7478);
and U7610 (N_7610,N_7269,N_7335);
nor U7611 (N_7611,N_7118,N_7265);
xnor U7612 (N_7612,N_7202,N_7456);
nand U7613 (N_7613,N_7163,N_7199);
and U7614 (N_7614,N_7391,N_7007);
and U7615 (N_7615,N_7051,N_7062);
nor U7616 (N_7616,N_7192,N_7453);
or U7617 (N_7617,N_7468,N_7416);
nand U7618 (N_7618,N_7360,N_7241);
xor U7619 (N_7619,N_7171,N_7260);
xor U7620 (N_7620,N_7092,N_7304);
and U7621 (N_7621,N_7386,N_7152);
nand U7622 (N_7622,N_7368,N_7114);
nand U7623 (N_7623,N_7234,N_7178);
xor U7624 (N_7624,N_7140,N_7406);
xor U7625 (N_7625,N_7213,N_7187);
or U7626 (N_7626,N_7049,N_7194);
or U7627 (N_7627,N_7162,N_7481);
xnor U7628 (N_7628,N_7098,N_7434);
or U7629 (N_7629,N_7177,N_7105);
nor U7630 (N_7630,N_7297,N_7052);
or U7631 (N_7631,N_7096,N_7214);
nand U7632 (N_7632,N_7161,N_7069);
and U7633 (N_7633,N_7184,N_7351);
nor U7634 (N_7634,N_7087,N_7095);
or U7635 (N_7635,N_7239,N_7475);
nor U7636 (N_7636,N_7462,N_7238);
nand U7637 (N_7637,N_7356,N_7261);
nor U7638 (N_7638,N_7054,N_7097);
nor U7639 (N_7639,N_7414,N_7172);
nor U7640 (N_7640,N_7379,N_7047);
xor U7641 (N_7641,N_7048,N_7193);
nand U7642 (N_7642,N_7395,N_7138);
and U7643 (N_7643,N_7110,N_7326);
or U7644 (N_7644,N_7073,N_7294);
and U7645 (N_7645,N_7272,N_7011);
nand U7646 (N_7646,N_7160,N_7415);
xnor U7647 (N_7647,N_7101,N_7025);
xor U7648 (N_7648,N_7479,N_7229);
xnor U7649 (N_7649,N_7144,N_7470);
nand U7650 (N_7650,N_7467,N_7472);
and U7651 (N_7651,N_7250,N_7222);
or U7652 (N_7652,N_7454,N_7292);
or U7653 (N_7653,N_7366,N_7196);
nor U7654 (N_7654,N_7488,N_7407);
and U7655 (N_7655,N_7303,N_7384);
and U7656 (N_7656,N_7197,N_7117);
xor U7657 (N_7657,N_7157,N_7195);
xor U7658 (N_7658,N_7459,N_7296);
xnor U7659 (N_7659,N_7208,N_7231);
nor U7660 (N_7660,N_7134,N_7077);
xor U7661 (N_7661,N_7495,N_7247);
or U7662 (N_7662,N_7143,N_7375);
or U7663 (N_7663,N_7450,N_7034);
or U7664 (N_7664,N_7014,N_7065);
or U7665 (N_7665,N_7319,N_7402);
nand U7666 (N_7666,N_7299,N_7273);
or U7667 (N_7667,N_7058,N_7349);
or U7668 (N_7668,N_7112,N_7135);
nand U7669 (N_7669,N_7206,N_7039);
nand U7670 (N_7670,N_7223,N_7332);
nor U7671 (N_7671,N_7433,N_7008);
xor U7672 (N_7672,N_7447,N_7023);
nor U7673 (N_7673,N_7200,N_7382);
nand U7674 (N_7674,N_7131,N_7183);
xor U7675 (N_7675,N_7310,N_7066);
and U7676 (N_7676,N_7076,N_7325);
or U7677 (N_7677,N_7367,N_7485);
nor U7678 (N_7678,N_7413,N_7372);
nor U7679 (N_7679,N_7340,N_7156);
and U7680 (N_7680,N_7377,N_7383);
nand U7681 (N_7681,N_7259,N_7146);
nor U7682 (N_7682,N_7337,N_7032);
nand U7683 (N_7683,N_7390,N_7106);
xnor U7684 (N_7684,N_7333,N_7217);
nand U7685 (N_7685,N_7258,N_7130);
nand U7686 (N_7686,N_7083,N_7148);
nor U7687 (N_7687,N_7204,N_7371);
or U7688 (N_7688,N_7031,N_7216);
xnor U7689 (N_7689,N_7219,N_7256);
and U7690 (N_7690,N_7203,N_7227);
and U7691 (N_7691,N_7180,N_7155);
nor U7692 (N_7692,N_7033,N_7387);
or U7693 (N_7693,N_7253,N_7119);
nor U7694 (N_7694,N_7225,N_7428);
and U7695 (N_7695,N_7174,N_7376);
and U7696 (N_7696,N_7315,N_7136);
and U7697 (N_7697,N_7085,N_7182);
or U7698 (N_7698,N_7461,N_7465);
nor U7699 (N_7699,N_7471,N_7380);
xor U7700 (N_7700,N_7185,N_7298);
and U7701 (N_7701,N_7125,N_7313);
nand U7702 (N_7702,N_7484,N_7021);
nand U7703 (N_7703,N_7175,N_7392);
xnor U7704 (N_7704,N_7198,N_7060);
and U7705 (N_7705,N_7220,N_7030);
nand U7706 (N_7706,N_7166,N_7236);
nor U7707 (N_7707,N_7347,N_7487);
nand U7708 (N_7708,N_7295,N_7167);
and U7709 (N_7709,N_7353,N_7421);
nor U7710 (N_7710,N_7423,N_7436);
nor U7711 (N_7711,N_7318,N_7191);
nor U7712 (N_7712,N_7029,N_7442);
nor U7713 (N_7713,N_7224,N_7133);
nor U7714 (N_7714,N_7249,N_7323);
xnor U7715 (N_7715,N_7075,N_7441);
xor U7716 (N_7716,N_7397,N_7289);
and U7717 (N_7717,N_7320,N_7086);
nor U7718 (N_7718,N_7240,N_7418);
nand U7719 (N_7719,N_7285,N_7009);
xor U7720 (N_7720,N_7147,N_7364);
nor U7721 (N_7721,N_7370,N_7103);
xor U7722 (N_7722,N_7338,N_7419);
and U7723 (N_7723,N_7427,N_7255);
nor U7724 (N_7724,N_7425,N_7437);
xor U7725 (N_7725,N_7142,N_7463);
nand U7726 (N_7726,N_7439,N_7154);
and U7727 (N_7727,N_7212,N_7466);
xnor U7728 (N_7728,N_7403,N_7496);
and U7729 (N_7729,N_7068,N_7158);
or U7730 (N_7730,N_7132,N_7159);
nor U7731 (N_7731,N_7004,N_7452);
nand U7732 (N_7732,N_7221,N_7100);
xnor U7733 (N_7733,N_7074,N_7036);
and U7734 (N_7734,N_7084,N_7035);
and U7735 (N_7735,N_7492,N_7331);
or U7736 (N_7736,N_7446,N_7071);
or U7737 (N_7737,N_7055,N_7314);
or U7738 (N_7738,N_7430,N_7401);
or U7739 (N_7739,N_7424,N_7302);
or U7740 (N_7740,N_7393,N_7099);
xnor U7741 (N_7741,N_7373,N_7408);
nor U7742 (N_7742,N_7327,N_7270);
or U7743 (N_7743,N_7230,N_7362);
and U7744 (N_7744,N_7116,N_7271);
or U7745 (N_7745,N_7088,N_7070);
nand U7746 (N_7746,N_7149,N_7288);
nand U7747 (N_7747,N_7243,N_7443);
nor U7748 (N_7748,N_7490,N_7057);
nor U7749 (N_7749,N_7121,N_7081);
or U7750 (N_7750,N_7411,N_7451);
xor U7751 (N_7751,N_7238,N_7363);
nand U7752 (N_7752,N_7398,N_7115);
nand U7753 (N_7753,N_7363,N_7146);
xnor U7754 (N_7754,N_7015,N_7178);
or U7755 (N_7755,N_7050,N_7325);
and U7756 (N_7756,N_7156,N_7255);
nand U7757 (N_7757,N_7442,N_7261);
and U7758 (N_7758,N_7074,N_7461);
nor U7759 (N_7759,N_7411,N_7171);
or U7760 (N_7760,N_7476,N_7270);
xor U7761 (N_7761,N_7219,N_7457);
or U7762 (N_7762,N_7308,N_7140);
and U7763 (N_7763,N_7315,N_7468);
nor U7764 (N_7764,N_7183,N_7210);
nand U7765 (N_7765,N_7024,N_7329);
xor U7766 (N_7766,N_7192,N_7268);
xor U7767 (N_7767,N_7208,N_7293);
or U7768 (N_7768,N_7415,N_7455);
and U7769 (N_7769,N_7317,N_7316);
and U7770 (N_7770,N_7381,N_7399);
or U7771 (N_7771,N_7278,N_7029);
nand U7772 (N_7772,N_7072,N_7270);
nor U7773 (N_7773,N_7100,N_7184);
xor U7774 (N_7774,N_7151,N_7358);
nor U7775 (N_7775,N_7020,N_7161);
xor U7776 (N_7776,N_7027,N_7066);
nor U7777 (N_7777,N_7200,N_7408);
nand U7778 (N_7778,N_7399,N_7453);
nand U7779 (N_7779,N_7132,N_7332);
or U7780 (N_7780,N_7026,N_7206);
nor U7781 (N_7781,N_7428,N_7459);
and U7782 (N_7782,N_7348,N_7382);
and U7783 (N_7783,N_7312,N_7341);
nor U7784 (N_7784,N_7085,N_7202);
and U7785 (N_7785,N_7308,N_7045);
nand U7786 (N_7786,N_7398,N_7408);
nand U7787 (N_7787,N_7197,N_7359);
nand U7788 (N_7788,N_7007,N_7296);
and U7789 (N_7789,N_7085,N_7268);
and U7790 (N_7790,N_7174,N_7147);
xor U7791 (N_7791,N_7020,N_7295);
or U7792 (N_7792,N_7153,N_7271);
and U7793 (N_7793,N_7288,N_7073);
nor U7794 (N_7794,N_7433,N_7450);
or U7795 (N_7795,N_7090,N_7371);
xor U7796 (N_7796,N_7148,N_7103);
and U7797 (N_7797,N_7218,N_7328);
nand U7798 (N_7798,N_7027,N_7160);
and U7799 (N_7799,N_7492,N_7008);
or U7800 (N_7800,N_7470,N_7450);
xor U7801 (N_7801,N_7140,N_7489);
xor U7802 (N_7802,N_7258,N_7455);
and U7803 (N_7803,N_7065,N_7178);
or U7804 (N_7804,N_7118,N_7214);
and U7805 (N_7805,N_7292,N_7357);
and U7806 (N_7806,N_7284,N_7016);
nor U7807 (N_7807,N_7498,N_7153);
nand U7808 (N_7808,N_7455,N_7316);
xnor U7809 (N_7809,N_7242,N_7173);
or U7810 (N_7810,N_7374,N_7264);
nor U7811 (N_7811,N_7015,N_7333);
and U7812 (N_7812,N_7150,N_7246);
xnor U7813 (N_7813,N_7341,N_7202);
nand U7814 (N_7814,N_7248,N_7122);
or U7815 (N_7815,N_7316,N_7111);
xnor U7816 (N_7816,N_7377,N_7189);
or U7817 (N_7817,N_7250,N_7131);
or U7818 (N_7818,N_7167,N_7144);
or U7819 (N_7819,N_7165,N_7327);
or U7820 (N_7820,N_7437,N_7320);
and U7821 (N_7821,N_7120,N_7284);
and U7822 (N_7822,N_7150,N_7345);
nand U7823 (N_7823,N_7199,N_7250);
xor U7824 (N_7824,N_7163,N_7368);
and U7825 (N_7825,N_7369,N_7321);
or U7826 (N_7826,N_7335,N_7091);
and U7827 (N_7827,N_7084,N_7425);
nand U7828 (N_7828,N_7069,N_7257);
or U7829 (N_7829,N_7407,N_7239);
or U7830 (N_7830,N_7035,N_7354);
nand U7831 (N_7831,N_7461,N_7479);
or U7832 (N_7832,N_7374,N_7081);
nand U7833 (N_7833,N_7113,N_7028);
nand U7834 (N_7834,N_7348,N_7065);
nand U7835 (N_7835,N_7158,N_7132);
or U7836 (N_7836,N_7338,N_7475);
xor U7837 (N_7837,N_7075,N_7469);
xor U7838 (N_7838,N_7408,N_7379);
nor U7839 (N_7839,N_7202,N_7323);
nor U7840 (N_7840,N_7432,N_7265);
or U7841 (N_7841,N_7289,N_7446);
nand U7842 (N_7842,N_7229,N_7253);
or U7843 (N_7843,N_7085,N_7423);
xnor U7844 (N_7844,N_7254,N_7497);
or U7845 (N_7845,N_7280,N_7453);
xor U7846 (N_7846,N_7123,N_7214);
or U7847 (N_7847,N_7109,N_7015);
nand U7848 (N_7848,N_7105,N_7338);
or U7849 (N_7849,N_7154,N_7428);
nor U7850 (N_7850,N_7014,N_7259);
nor U7851 (N_7851,N_7490,N_7012);
and U7852 (N_7852,N_7196,N_7356);
nand U7853 (N_7853,N_7389,N_7129);
or U7854 (N_7854,N_7137,N_7424);
nand U7855 (N_7855,N_7283,N_7202);
nor U7856 (N_7856,N_7289,N_7432);
and U7857 (N_7857,N_7411,N_7035);
and U7858 (N_7858,N_7293,N_7101);
and U7859 (N_7859,N_7197,N_7450);
or U7860 (N_7860,N_7329,N_7423);
xor U7861 (N_7861,N_7099,N_7280);
and U7862 (N_7862,N_7468,N_7383);
and U7863 (N_7863,N_7351,N_7333);
nand U7864 (N_7864,N_7238,N_7441);
or U7865 (N_7865,N_7407,N_7153);
or U7866 (N_7866,N_7038,N_7270);
nand U7867 (N_7867,N_7149,N_7233);
and U7868 (N_7868,N_7215,N_7309);
or U7869 (N_7869,N_7205,N_7092);
xnor U7870 (N_7870,N_7302,N_7452);
nor U7871 (N_7871,N_7492,N_7239);
and U7872 (N_7872,N_7175,N_7292);
xnor U7873 (N_7873,N_7248,N_7398);
xnor U7874 (N_7874,N_7486,N_7418);
nand U7875 (N_7875,N_7072,N_7191);
nand U7876 (N_7876,N_7014,N_7472);
or U7877 (N_7877,N_7422,N_7348);
xnor U7878 (N_7878,N_7235,N_7400);
xor U7879 (N_7879,N_7002,N_7123);
nand U7880 (N_7880,N_7414,N_7393);
and U7881 (N_7881,N_7035,N_7124);
and U7882 (N_7882,N_7411,N_7414);
nand U7883 (N_7883,N_7475,N_7479);
and U7884 (N_7884,N_7071,N_7063);
or U7885 (N_7885,N_7362,N_7374);
nand U7886 (N_7886,N_7432,N_7023);
xnor U7887 (N_7887,N_7023,N_7487);
or U7888 (N_7888,N_7328,N_7007);
and U7889 (N_7889,N_7050,N_7394);
nand U7890 (N_7890,N_7477,N_7300);
or U7891 (N_7891,N_7322,N_7102);
and U7892 (N_7892,N_7354,N_7162);
xnor U7893 (N_7893,N_7396,N_7024);
or U7894 (N_7894,N_7141,N_7372);
xor U7895 (N_7895,N_7456,N_7037);
or U7896 (N_7896,N_7269,N_7143);
xor U7897 (N_7897,N_7299,N_7244);
nand U7898 (N_7898,N_7086,N_7401);
or U7899 (N_7899,N_7308,N_7182);
or U7900 (N_7900,N_7071,N_7194);
xor U7901 (N_7901,N_7157,N_7174);
or U7902 (N_7902,N_7266,N_7186);
xnor U7903 (N_7903,N_7175,N_7491);
xor U7904 (N_7904,N_7134,N_7231);
and U7905 (N_7905,N_7127,N_7496);
xnor U7906 (N_7906,N_7244,N_7438);
xor U7907 (N_7907,N_7055,N_7340);
or U7908 (N_7908,N_7031,N_7257);
nor U7909 (N_7909,N_7288,N_7032);
and U7910 (N_7910,N_7347,N_7112);
or U7911 (N_7911,N_7043,N_7285);
nor U7912 (N_7912,N_7285,N_7155);
and U7913 (N_7913,N_7292,N_7006);
nor U7914 (N_7914,N_7033,N_7200);
nor U7915 (N_7915,N_7369,N_7018);
nand U7916 (N_7916,N_7447,N_7126);
nand U7917 (N_7917,N_7317,N_7161);
or U7918 (N_7918,N_7404,N_7066);
xor U7919 (N_7919,N_7107,N_7308);
nand U7920 (N_7920,N_7462,N_7174);
nor U7921 (N_7921,N_7308,N_7411);
or U7922 (N_7922,N_7318,N_7181);
nand U7923 (N_7923,N_7128,N_7429);
nand U7924 (N_7924,N_7226,N_7269);
nand U7925 (N_7925,N_7495,N_7017);
nand U7926 (N_7926,N_7424,N_7356);
or U7927 (N_7927,N_7039,N_7095);
xor U7928 (N_7928,N_7251,N_7134);
nand U7929 (N_7929,N_7199,N_7025);
and U7930 (N_7930,N_7375,N_7425);
or U7931 (N_7931,N_7447,N_7075);
and U7932 (N_7932,N_7299,N_7147);
nand U7933 (N_7933,N_7209,N_7070);
nand U7934 (N_7934,N_7117,N_7030);
nor U7935 (N_7935,N_7288,N_7499);
and U7936 (N_7936,N_7280,N_7061);
and U7937 (N_7937,N_7235,N_7205);
or U7938 (N_7938,N_7176,N_7477);
nor U7939 (N_7939,N_7320,N_7058);
and U7940 (N_7940,N_7010,N_7308);
nand U7941 (N_7941,N_7199,N_7379);
and U7942 (N_7942,N_7052,N_7090);
nor U7943 (N_7943,N_7197,N_7447);
nand U7944 (N_7944,N_7180,N_7019);
nand U7945 (N_7945,N_7324,N_7101);
nor U7946 (N_7946,N_7190,N_7299);
and U7947 (N_7947,N_7246,N_7051);
or U7948 (N_7948,N_7184,N_7362);
xor U7949 (N_7949,N_7277,N_7097);
nor U7950 (N_7950,N_7251,N_7392);
and U7951 (N_7951,N_7464,N_7225);
xnor U7952 (N_7952,N_7355,N_7397);
xor U7953 (N_7953,N_7194,N_7164);
and U7954 (N_7954,N_7297,N_7181);
xnor U7955 (N_7955,N_7437,N_7106);
nor U7956 (N_7956,N_7332,N_7456);
nor U7957 (N_7957,N_7160,N_7069);
or U7958 (N_7958,N_7346,N_7045);
xor U7959 (N_7959,N_7148,N_7468);
or U7960 (N_7960,N_7030,N_7397);
nand U7961 (N_7961,N_7488,N_7333);
nor U7962 (N_7962,N_7262,N_7462);
nor U7963 (N_7963,N_7109,N_7452);
and U7964 (N_7964,N_7147,N_7088);
xnor U7965 (N_7965,N_7293,N_7490);
or U7966 (N_7966,N_7481,N_7466);
nand U7967 (N_7967,N_7295,N_7035);
and U7968 (N_7968,N_7265,N_7239);
or U7969 (N_7969,N_7051,N_7443);
nand U7970 (N_7970,N_7088,N_7309);
or U7971 (N_7971,N_7413,N_7109);
and U7972 (N_7972,N_7439,N_7362);
nor U7973 (N_7973,N_7461,N_7270);
or U7974 (N_7974,N_7013,N_7127);
and U7975 (N_7975,N_7385,N_7217);
nand U7976 (N_7976,N_7371,N_7096);
or U7977 (N_7977,N_7071,N_7092);
and U7978 (N_7978,N_7415,N_7412);
nand U7979 (N_7979,N_7098,N_7429);
xor U7980 (N_7980,N_7445,N_7094);
or U7981 (N_7981,N_7155,N_7403);
nor U7982 (N_7982,N_7066,N_7121);
nand U7983 (N_7983,N_7049,N_7094);
or U7984 (N_7984,N_7332,N_7285);
xnor U7985 (N_7985,N_7103,N_7185);
and U7986 (N_7986,N_7341,N_7207);
or U7987 (N_7987,N_7076,N_7369);
or U7988 (N_7988,N_7124,N_7492);
or U7989 (N_7989,N_7306,N_7088);
nand U7990 (N_7990,N_7179,N_7421);
xor U7991 (N_7991,N_7383,N_7424);
xnor U7992 (N_7992,N_7274,N_7227);
and U7993 (N_7993,N_7084,N_7434);
nand U7994 (N_7994,N_7430,N_7492);
nand U7995 (N_7995,N_7053,N_7010);
nand U7996 (N_7996,N_7213,N_7225);
or U7997 (N_7997,N_7403,N_7179);
or U7998 (N_7998,N_7387,N_7381);
or U7999 (N_7999,N_7214,N_7428);
and U8000 (N_8000,N_7590,N_7938);
nand U8001 (N_8001,N_7867,N_7976);
nand U8002 (N_8002,N_7956,N_7954);
nor U8003 (N_8003,N_7663,N_7715);
and U8004 (N_8004,N_7631,N_7640);
xor U8005 (N_8005,N_7769,N_7842);
or U8006 (N_8006,N_7818,N_7877);
xor U8007 (N_8007,N_7849,N_7983);
nand U8008 (N_8008,N_7764,N_7721);
nor U8009 (N_8009,N_7655,N_7755);
xor U8010 (N_8010,N_7667,N_7757);
xnor U8011 (N_8011,N_7793,N_7767);
and U8012 (N_8012,N_7947,N_7795);
nand U8013 (N_8013,N_7624,N_7873);
xor U8014 (N_8014,N_7942,N_7791);
or U8015 (N_8015,N_7718,N_7882);
nand U8016 (N_8016,N_7776,N_7933);
and U8017 (N_8017,N_7523,N_7888);
xor U8018 (N_8018,N_7589,N_7991);
xor U8019 (N_8019,N_7846,N_7747);
or U8020 (N_8020,N_7814,N_7593);
nand U8021 (N_8021,N_7709,N_7733);
nor U8022 (N_8022,N_7910,N_7837);
or U8023 (N_8023,N_7774,N_7836);
nor U8024 (N_8024,N_7899,N_7690);
xnor U8025 (N_8025,N_7832,N_7978);
and U8026 (N_8026,N_7746,N_7719);
or U8027 (N_8027,N_7519,N_7967);
xnor U8028 (N_8028,N_7966,N_7940);
or U8029 (N_8029,N_7710,N_7621);
xor U8030 (N_8030,N_7905,N_7854);
xor U8031 (N_8031,N_7839,N_7527);
and U8032 (N_8032,N_7704,N_7762);
and U8033 (N_8033,N_7861,N_7745);
or U8034 (N_8034,N_7508,N_7807);
nand U8035 (N_8035,N_7516,N_7602);
or U8036 (N_8036,N_7581,N_7619);
xnor U8037 (N_8037,N_7911,N_7939);
nand U8038 (N_8038,N_7985,N_7772);
and U8039 (N_8039,N_7789,N_7734);
xnor U8040 (N_8040,N_7633,N_7657);
or U8041 (N_8041,N_7731,N_7565);
nand U8042 (N_8042,N_7951,N_7792);
or U8043 (N_8043,N_7923,N_7890);
xnor U8044 (N_8044,N_7968,N_7986);
xor U8045 (N_8045,N_7670,N_7622);
and U8046 (N_8046,N_7521,N_7994);
xor U8047 (N_8047,N_7564,N_7863);
nand U8048 (N_8048,N_7726,N_7920);
or U8049 (N_8049,N_7703,N_7828);
nor U8050 (N_8050,N_7771,N_7594);
nor U8051 (N_8051,N_7889,N_7765);
and U8052 (N_8052,N_7809,N_7981);
xnor U8053 (N_8053,N_7833,N_7572);
or U8054 (N_8054,N_7558,N_7618);
or U8055 (N_8055,N_7610,N_7936);
nor U8056 (N_8056,N_7801,N_7740);
nor U8057 (N_8057,N_7777,N_7872);
or U8058 (N_8058,N_7608,N_7559);
nor U8059 (N_8059,N_7768,N_7579);
nand U8060 (N_8060,N_7959,N_7636);
nand U8061 (N_8061,N_7672,N_7742);
nor U8062 (N_8062,N_7871,N_7826);
or U8063 (N_8063,N_7666,N_7961);
and U8064 (N_8064,N_7835,N_7680);
xor U8065 (N_8065,N_7563,N_7783);
or U8066 (N_8066,N_7847,N_7605);
xnor U8067 (N_8067,N_7674,N_7834);
nand U8068 (N_8068,N_7857,N_7571);
and U8069 (N_8069,N_7713,N_7596);
or U8070 (N_8070,N_7517,N_7796);
and U8071 (N_8071,N_7993,N_7798);
and U8072 (N_8072,N_7843,N_7884);
nor U8073 (N_8073,N_7611,N_7706);
or U8074 (N_8074,N_7858,N_7931);
or U8075 (N_8075,N_7570,N_7525);
nor U8076 (N_8076,N_7896,N_7658);
or U8077 (N_8077,N_7566,N_7584);
nand U8078 (N_8078,N_7827,N_7720);
xor U8079 (N_8079,N_7530,N_7965);
nand U8080 (N_8080,N_7944,N_7599);
and U8081 (N_8081,N_7567,N_7819);
xor U8082 (N_8082,N_7695,N_7630);
or U8083 (N_8083,N_7930,N_7901);
or U8084 (N_8084,N_7506,N_7536);
nand U8085 (N_8085,N_7803,N_7885);
and U8086 (N_8086,N_7908,N_7925);
and U8087 (N_8087,N_7752,N_7600);
xnor U8088 (N_8088,N_7543,N_7679);
and U8089 (N_8089,N_7788,N_7504);
nand U8090 (N_8090,N_7948,N_7500);
nor U8091 (N_8091,N_7648,N_7637);
xnor U8092 (N_8092,N_7779,N_7784);
and U8093 (N_8093,N_7775,N_7649);
or U8094 (N_8094,N_7917,N_7675);
nor U8095 (N_8095,N_7964,N_7886);
nor U8096 (N_8096,N_7802,N_7627);
and U8097 (N_8097,N_7513,N_7879);
nor U8098 (N_8098,N_7741,N_7972);
nand U8099 (N_8099,N_7759,N_7805);
nor U8100 (N_8100,N_7941,N_7705);
xnor U8101 (N_8101,N_7787,N_7639);
nand U8102 (N_8102,N_7794,N_7856);
nor U8103 (N_8103,N_7524,N_7989);
and U8104 (N_8104,N_7824,N_7617);
nand U8105 (N_8105,N_7573,N_7505);
xor U8106 (N_8106,N_7613,N_7817);
nor U8107 (N_8107,N_7894,N_7945);
or U8108 (N_8108,N_7660,N_7628);
or U8109 (N_8109,N_7934,N_7603);
nor U8110 (N_8110,N_7971,N_7816);
or U8111 (N_8111,N_7669,N_7546);
nor U8112 (N_8112,N_7661,N_7987);
xnor U8113 (N_8113,N_7575,N_7864);
or U8114 (N_8114,N_7756,N_7708);
and U8115 (N_8115,N_7682,N_7641);
xnor U8116 (N_8116,N_7743,N_7691);
nor U8117 (N_8117,N_7897,N_7969);
nor U8118 (N_8118,N_7912,N_7970);
nand U8119 (N_8119,N_7509,N_7620);
xor U8120 (N_8120,N_7738,N_7852);
and U8121 (N_8121,N_7712,N_7963);
nand U8122 (N_8122,N_7609,N_7693);
or U8123 (N_8123,N_7697,N_7552);
or U8124 (N_8124,N_7548,N_7568);
and U8125 (N_8125,N_7545,N_7725);
or U8126 (N_8126,N_7977,N_7561);
and U8127 (N_8127,N_7550,N_7980);
and U8128 (N_8128,N_7999,N_7585);
nand U8129 (N_8129,N_7612,N_7821);
nor U8130 (N_8130,N_7623,N_7902);
nand U8131 (N_8131,N_7766,N_7577);
or U8132 (N_8132,N_7651,N_7730);
and U8133 (N_8133,N_7689,N_7683);
or U8134 (N_8134,N_7601,N_7534);
and U8135 (N_8135,N_7647,N_7522);
nand U8136 (N_8136,N_7662,N_7732);
or U8137 (N_8137,N_7866,N_7526);
nand U8138 (N_8138,N_7898,N_7644);
xor U8139 (N_8139,N_7781,N_7786);
or U8140 (N_8140,N_7937,N_7869);
or U8141 (N_8141,N_7900,N_7825);
and U8142 (N_8142,N_7549,N_7702);
nor U8143 (N_8143,N_7727,N_7996);
nor U8144 (N_8144,N_7553,N_7915);
nor U8145 (N_8145,N_7955,N_7583);
xnor U8146 (N_8146,N_7950,N_7728);
xor U8147 (N_8147,N_7514,N_7698);
nor U8148 (N_8148,N_7876,N_7904);
and U8149 (N_8149,N_7962,N_7533);
or U8150 (N_8150,N_7770,N_7973);
xor U8151 (N_8151,N_7541,N_7532);
nand U8152 (N_8152,N_7810,N_7754);
and U8153 (N_8153,N_7737,N_7952);
or U8154 (N_8154,N_7848,N_7539);
or U8155 (N_8155,N_7806,N_7595);
nand U8156 (N_8156,N_7652,N_7537);
xor U8157 (N_8157,N_7699,N_7927);
or U8158 (N_8158,N_7960,N_7850);
nor U8159 (N_8159,N_7574,N_7748);
nand U8160 (N_8160,N_7614,N_7928);
nand U8161 (N_8161,N_7701,N_7520);
and U8162 (N_8162,N_7913,N_7685);
nand U8163 (N_8163,N_7700,N_7844);
nand U8164 (N_8164,N_7782,N_7638);
or U8165 (N_8165,N_7780,N_7665);
and U8166 (N_8166,N_7625,N_7760);
nand U8167 (N_8167,N_7909,N_7949);
nand U8168 (N_8168,N_7653,N_7813);
nor U8169 (N_8169,N_7929,N_7831);
xnor U8170 (N_8170,N_7946,N_7507);
nor U8171 (N_8171,N_7607,N_7671);
or U8172 (N_8172,N_7684,N_7544);
xor U8173 (N_8173,N_7606,N_7840);
xor U8174 (N_8174,N_7643,N_7722);
nor U8175 (N_8175,N_7724,N_7569);
nand U8176 (N_8176,N_7749,N_7763);
and U8177 (N_8177,N_7554,N_7845);
nor U8178 (N_8178,N_7736,N_7812);
xor U8179 (N_8179,N_7502,N_7739);
nand U8180 (N_8180,N_7984,N_7865);
nor U8181 (N_8181,N_7855,N_7868);
and U8182 (N_8182,N_7676,N_7935);
nor U8183 (N_8183,N_7578,N_7587);
and U8184 (N_8184,N_7518,N_7645);
nand U8185 (N_8185,N_7556,N_7510);
and U8186 (N_8186,N_7893,N_7677);
nand U8187 (N_8187,N_7932,N_7642);
xnor U8188 (N_8188,N_7503,N_7841);
or U8189 (N_8189,N_7535,N_7668);
or U8190 (N_8190,N_7907,N_7922);
and U8191 (N_8191,N_7529,N_7903);
nor U8192 (N_8192,N_7778,N_7988);
xor U8193 (N_8193,N_7598,N_7918);
nor U8194 (N_8194,N_7597,N_7875);
nand U8195 (N_8195,N_7582,N_7696);
nand U8196 (N_8196,N_7853,N_7632);
nor U8197 (N_8197,N_7678,N_7878);
nor U8198 (N_8198,N_7943,N_7634);
nand U8199 (N_8199,N_7735,N_7799);
nor U8200 (N_8200,N_7591,N_7838);
xor U8201 (N_8201,N_7975,N_7751);
xnor U8202 (N_8202,N_7895,N_7982);
xnor U8203 (N_8203,N_7512,N_7820);
xor U8204 (N_8204,N_7790,N_7919);
and U8205 (N_8205,N_7880,N_7773);
and U8206 (N_8206,N_7870,N_7729);
or U8207 (N_8207,N_7542,N_7629);
nand U8208 (N_8208,N_7881,N_7750);
and U8209 (N_8209,N_7635,N_7822);
or U8210 (N_8210,N_7892,N_7815);
or U8211 (N_8211,N_7753,N_7830);
and U8212 (N_8212,N_7992,N_7707);
or U8213 (N_8213,N_7758,N_7654);
nor U8214 (N_8214,N_7859,N_7562);
and U8215 (N_8215,N_7906,N_7586);
xnor U8216 (N_8216,N_7615,N_7538);
and U8217 (N_8217,N_7531,N_7688);
or U8218 (N_8218,N_7501,N_7659);
xor U8219 (N_8219,N_7547,N_7997);
nand U8220 (N_8220,N_7604,N_7511);
nand U8221 (N_8221,N_7916,N_7811);
and U8222 (N_8222,N_7953,N_7592);
and U8223 (N_8223,N_7694,N_7860);
xor U8224 (N_8224,N_7711,N_7580);
nand U8225 (N_8225,N_7560,N_7540);
or U8226 (N_8226,N_7829,N_7656);
xnor U8227 (N_8227,N_7926,N_7998);
or U8228 (N_8228,N_7874,N_7797);
nor U8229 (N_8229,N_7515,N_7979);
or U8230 (N_8230,N_7804,N_7761);
and U8231 (N_8231,N_7958,N_7555);
xnor U8232 (N_8232,N_7914,N_7716);
nand U8233 (N_8233,N_7551,N_7692);
nor U8234 (N_8234,N_7650,N_7616);
and U8235 (N_8235,N_7990,N_7924);
and U8236 (N_8236,N_7557,N_7887);
or U8237 (N_8237,N_7681,N_7808);
nor U8238 (N_8238,N_7528,N_7687);
nor U8239 (N_8239,N_7664,N_7785);
and U8240 (N_8240,N_7576,N_7957);
nand U8241 (N_8241,N_7921,N_7588);
nand U8242 (N_8242,N_7862,N_7995);
and U8243 (N_8243,N_7891,N_7851);
and U8244 (N_8244,N_7800,N_7717);
nand U8245 (N_8245,N_7883,N_7673);
xor U8246 (N_8246,N_7714,N_7823);
or U8247 (N_8247,N_7974,N_7626);
nor U8248 (N_8248,N_7723,N_7646);
nand U8249 (N_8249,N_7686,N_7744);
nand U8250 (N_8250,N_7511,N_7682);
and U8251 (N_8251,N_7828,N_7707);
or U8252 (N_8252,N_7770,N_7778);
or U8253 (N_8253,N_7936,N_7836);
and U8254 (N_8254,N_7802,N_7513);
and U8255 (N_8255,N_7796,N_7700);
and U8256 (N_8256,N_7650,N_7530);
nand U8257 (N_8257,N_7644,N_7548);
or U8258 (N_8258,N_7871,N_7947);
or U8259 (N_8259,N_7906,N_7991);
nor U8260 (N_8260,N_7782,N_7957);
nand U8261 (N_8261,N_7860,N_7645);
or U8262 (N_8262,N_7649,N_7923);
nand U8263 (N_8263,N_7599,N_7897);
and U8264 (N_8264,N_7885,N_7836);
xnor U8265 (N_8265,N_7674,N_7887);
and U8266 (N_8266,N_7658,N_7824);
nor U8267 (N_8267,N_7937,N_7729);
and U8268 (N_8268,N_7872,N_7613);
nor U8269 (N_8269,N_7593,N_7953);
and U8270 (N_8270,N_7790,N_7622);
and U8271 (N_8271,N_7988,N_7726);
nor U8272 (N_8272,N_7932,N_7902);
nand U8273 (N_8273,N_7676,N_7647);
nand U8274 (N_8274,N_7905,N_7945);
and U8275 (N_8275,N_7769,N_7977);
or U8276 (N_8276,N_7840,N_7949);
nand U8277 (N_8277,N_7961,N_7918);
or U8278 (N_8278,N_7785,N_7688);
nand U8279 (N_8279,N_7802,N_7685);
xnor U8280 (N_8280,N_7889,N_7523);
xor U8281 (N_8281,N_7603,N_7604);
xor U8282 (N_8282,N_7920,N_7851);
xnor U8283 (N_8283,N_7728,N_7734);
xor U8284 (N_8284,N_7780,N_7762);
nand U8285 (N_8285,N_7966,N_7683);
or U8286 (N_8286,N_7511,N_7555);
or U8287 (N_8287,N_7765,N_7639);
and U8288 (N_8288,N_7872,N_7507);
and U8289 (N_8289,N_7759,N_7828);
or U8290 (N_8290,N_7801,N_7614);
or U8291 (N_8291,N_7770,N_7848);
or U8292 (N_8292,N_7975,N_7998);
xnor U8293 (N_8293,N_7786,N_7771);
nand U8294 (N_8294,N_7699,N_7667);
nor U8295 (N_8295,N_7874,N_7951);
nand U8296 (N_8296,N_7566,N_7793);
or U8297 (N_8297,N_7622,N_7811);
nand U8298 (N_8298,N_7960,N_7657);
and U8299 (N_8299,N_7594,N_7508);
nand U8300 (N_8300,N_7662,N_7602);
and U8301 (N_8301,N_7838,N_7906);
xor U8302 (N_8302,N_7974,N_7519);
nand U8303 (N_8303,N_7638,N_7701);
nor U8304 (N_8304,N_7965,N_7516);
and U8305 (N_8305,N_7954,N_7672);
nor U8306 (N_8306,N_7785,N_7783);
nand U8307 (N_8307,N_7693,N_7734);
and U8308 (N_8308,N_7607,N_7603);
nand U8309 (N_8309,N_7984,N_7942);
nor U8310 (N_8310,N_7764,N_7819);
nor U8311 (N_8311,N_7859,N_7839);
or U8312 (N_8312,N_7747,N_7775);
nand U8313 (N_8313,N_7739,N_7837);
nand U8314 (N_8314,N_7580,N_7862);
and U8315 (N_8315,N_7821,N_7723);
and U8316 (N_8316,N_7650,N_7615);
or U8317 (N_8317,N_7903,N_7914);
xor U8318 (N_8318,N_7514,N_7897);
or U8319 (N_8319,N_7556,N_7939);
xnor U8320 (N_8320,N_7642,N_7535);
nor U8321 (N_8321,N_7596,N_7944);
and U8322 (N_8322,N_7741,N_7577);
xor U8323 (N_8323,N_7668,N_7685);
nor U8324 (N_8324,N_7756,N_7591);
xnor U8325 (N_8325,N_7506,N_7930);
or U8326 (N_8326,N_7901,N_7882);
nor U8327 (N_8327,N_7964,N_7576);
and U8328 (N_8328,N_7710,N_7945);
nand U8329 (N_8329,N_7663,N_7714);
nand U8330 (N_8330,N_7609,N_7998);
xor U8331 (N_8331,N_7997,N_7706);
and U8332 (N_8332,N_7727,N_7896);
and U8333 (N_8333,N_7815,N_7502);
nor U8334 (N_8334,N_7979,N_7543);
or U8335 (N_8335,N_7904,N_7839);
nor U8336 (N_8336,N_7768,N_7701);
xor U8337 (N_8337,N_7990,N_7712);
xnor U8338 (N_8338,N_7549,N_7874);
or U8339 (N_8339,N_7900,N_7946);
xnor U8340 (N_8340,N_7912,N_7952);
and U8341 (N_8341,N_7728,N_7629);
nor U8342 (N_8342,N_7677,N_7694);
nor U8343 (N_8343,N_7820,N_7825);
xor U8344 (N_8344,N_7850,N_7847);
and U8345 (N_8345,N_7657,N_7700);
nor U8346 (N_8346,N_7616,N_7870);
xor U8347 (N_8347,N_7625,N_7587);
nand U8348 (N_8348,N_7927,N_7873);
or U8349 (N_8349,N_7638,N_7786);
or U8350 (N_8350,N_7622,N_7626);
xnor U8351 (N_8351,N_7970,N_7836);
nor U8352 (N_8352,N_7809,N_7579);
and U8353 (N_8353,N_7611,N_7916);
and U8354 (N_8354,N_7892,N_7603);
or U8355 (N_8355,N_7530,N_7660);
xor U8356 (N_8356,N_7775,N_7612);
and U8357 (N_8357,N_7505,N_7937);
and U8358 (N_8358,N_7630,N_7756);
nand U8359 (N_8359,N_7990,N_7628);
or U8360 (N_8360,N_7878,N_7668);
xnor U8361 (N_8361,N_7522,N_7550);
nand U8362 (N_8362,N_7967,N_7708);
nor U8363 (N_8363,N_7999,N_7837);
nor U8364 (N_8364,N_7819,N_7957);
xnor U8365 (N_8365,N_7545,N_7514);
xor U8366 (N_8366,N_7569,N_7835);
nand U8367 (N_8367,N_7691,N_7931);
and U8368 (N_8368,N_7709,N_7885);
nor U8369 (N_8369,N_7569,N_7580);
nor U8370 (N_8370,N_7606,N_7749);
or U8371 (N_8371,N_7580,N_7825);
nor U8372 (N_8372,N_7632,N_7925);
and U8373 (N_8373,N_7708,N_7931);
and U8374 (N_8374,N_7547,N_7959);
nor U8375 (N_8375,N_7567,N_7859);
xnor U8376 (N_8376,N_7702,N_7853);
xnor U8377 (N_8377,N_7979,N_7535);
xnor U8378 (N_8378,N_7719,N_7841);
or U8379 (N_8379,N_7713,N_7914);
and U8380 (N_8380,N_7750,N_7520);
and U8381 (N_8381,N_7588,N_7990);
nor U8382 (N_8382,N_7550,N_7868);
xor U8383 (N_8383,N_7604,N_7795);
nand U8384 (N_8384,N_7547,N_7893);
nand U8385 (N_8385,N_7725,N_7944);
nand U8386 (N_8386,N_7768,N_7658);
nor U8387 (N_8387,N_7810,N_7932);
nor U8388 (N_8388,N_7992,N_7791);
nor U8389 (N_8389,N_7681,N_7834);
xnor U8390 (N_8390,N_7811,N_7703);
and U8391 (N_8391,N_7956,N_7668);
nor U8392 (N_8392,N_7572,N_7590);
and U8393 (N_8393,N_7806,N_7849);
and U8394 (N_8394,N_7970,N_7732);
or U8395 (N_8395,N_7849,N_7900);
xor U8396 (N_8396,N_7696,N_7909);
and U8397 (N_8397,N_7712,N_7680);
or U8398 (N_8398,N_7517,N_7837);
xnor U8399 (N_8399,N_7674,N_7675);
or U8400 (N_8400,N_7510,N_7985);
xor U8401 (N_8401,N_7622,N_7697);
and U8402 (N_8402,N_7745,N_7708);
nand U8403 (N_8403,N_7674,N_7740);
or U8404 (N_8404,N_7732,N_7535);
and U8405 (N_8405,N_7871,N_7847);
xnor U8406 (N_8406,N_7682,N_7959);
and U8407 (N_8407,N_7569,N_7908);
nand U8408 (N_8408,N_7741,N_7734);
and U8409 (N_8409,N_7949,N_7851);
or U8410 (N_8410,N_7911,N_7589);
nand U8411 (N_8411,N_7918,N_7683);
and U8412 (N_8412,N_7724,N_7557);
or U8413 (N_8413,N_7704,N_7565);
xnor U8414 (N_8414,N_7968,N_7948);
nor U8415 (N_8415,N_7672,N_7503);
nand U8416 (N_8416,N_7527,N_7548);
or U8417 (N_8417,N_7847,N_7500);
or U8418 (N_8418,N_7891,N_7721);
or U8419 (N_8419,N_7523,N_7697);
nand U8420 (N_8420,N_7921,N_7764);
xnor U8421 (N_8421,N_7530,N_7647);
xnor U8422 (N_8422,N_7739,N_7552);
nand U8423 (N_8423,N_7542,N_7724);
and U8424 (N_8424,N_7706,N_7549);
xnor U8425 (N_8425,N_7510,N_7592);
xor U8426 (N_8426,N_7594,N_7722);
or U8427 (N_8427,N_7527,N_7896);
nor U8428 (N_8428,N_7860,N_7782);
or U8429 (N_8429,N_7733,N_7741);
and U8430 (N_8430,N_7771,N_7607);
nor U8431 (N_8431,N_7941,N_7816);
nand U8432 (N_8432,N_7673,N_7644);
and U8433 (N_8433,N_7673,N_7554);
nor U8434 (N_8434,N_7679,N_7985);
xor U8435 (N_8435,N_7962,N_7614);
nand U8436 (N_8436,N_7810,N_7667);
xor U8437 (N_8437,N_7691,N_7850);
and U8438 (N_8438,N_7717,N_7932);
or U8439 (N_8439,N_7665,N_7520);
or U8440 (N_8440,N_7997,N_7515);
and U8441 (N_8441,N_7509,N_7694);
or U8442 (N_8442,N_7521,N_7731);
nor U8443 (N_8443,N_7851,N_7914);
nor U8444 (N_8444,N_7774,N_7748);
or U8445 (N_8445,N_7955,N_7724);
or U8446 (N_8446,N_7852,N_7776);
xor U8447 (N_8447,N_7635,N_7808);
nand U8448 (N_8448,N_7703,N_7535);
or U8449 (N_8449,N_7602,N_7556);
and U8450 (N_8450,N_7814,N_7664);
nor U8451 (N_8451,N_7549,N_7537);
nand U8452 (N_8452,N_7889,N_7966);
nor U8453 (N_8453,N_7978,N_7625);
or U8454 (N_8454,N_7585,N_7747);
nand U8455 (N_8455,N_7983,N_7679);
or U8456 (N_8456,N_7773,N_7541);
nor U8457 (N_8457,N_7913,N_7681);
nor U8458 (N_8458,N_7626,N_7866);
xnor U8459 (N_8459,N_7864,N_7942);
nor U8460 (N_8460,N_7927,N_7833);
nand U8461 (N_8461,N_7669,N_7694);
and U8462 (N_8462,N_7949,N_7567);
xor U8463 (N_8463,N_7634,N_7599);
and U8464 (N_8464,N_7650,N_7980);
nor U8465 (N_8465,N_7590,N_7727);
xor U8466 (N_8466,N_7817,N_7766);
or U8467 (N_8467,N_7686,N_7962);
nand U8468 (N_8468,N_7885,N_7845);
nor U8469 (N_8469,N_7884,N_7964);
nand U8470 (N_8470,N_7690,N_7858);
nand U8471 (N_8471,N_7878,N_7727);
or U8472 (N_8472,N_7678,N_7570);
xor U8473 (N_8473,N_7646,N_7996);
or U8474 (N_8474,N_7751,N_7741);
and U8475 (N_8475,N_7920,N_7841);
or U8476 (N_8476,N_7856,N_7718);
nand U8477 (N_8477,N_7945,N_7760);
nand U8478 (N_8478,N_7894,N_7521);
or U8479 (N_8479,N_7882,N_7535);
and U8480 (N_8480,N_7917,N_7866);
nand U8481 (N_8481,N_7523,N_7977);
nor U8482 (N_8482,N_7761,N_7676);
and U8483 (N_8483,N_7651,N_7737);
and U8484 (N_8484,N_7683,N_7735);
or U8485 (N_8485,N_7680,N_7890);
nor U8486 (N_8486,N_7655,N_7897);
or U8487 (N_8487,N_7870,N_7785);
nor U8488 (N_8488,N_7978,N_7805);
nor U8489 (N_8489,N_7505,N_7978);
xnor U8490 (N_8490,N_7925,N_7688);
xor U8491 (N_8491,N_7903,N_7525);
nor U8492 (N_8492,N_7987,N_7925);
nand U8493 (N_8493,N_7957,N_7898);
nand U8494 (N_8494,N_7819,N_7853);
xnor U8495 (N_8495,N_7526,N_7736);
xnor U8496 (N_8496,N_7748,N_7698);
and U8497 (N_8497,N_7503,N_7559);
xnor U8498 (N_8498,N_7643,N_7588);
nor U8499 (N_8499,N_7862,N_7718);
xnor U8500 (N_8500,N_8185,N_8391);
or U8501 (N_8501,N_8280,N_8113);
or U8502 (N_8502,N_8061,N_8382);
nand U8503 (N_8503,N_8116,N_8101);
xnor U8504 (N_8504,N_8444,N_8056);
nand U8505 (N_8505,N_8152,N_8432);
nor U8506 (N_8506,N_8484,N_8016);
nand U8507 (N_8507,N_8012,N_8017);
xnor U8508 (N_8508,N_8239,N_8314);
xnor U8509 (N_8509,N_8203,N_8440);
and U8510 (N_8510,N_8347,N_8478);
xnor U8511 (N_8511,N_8163,N_8335);
or U8512 (N_8512,N_8408,N_8452);
nand U8513 (N_8513,N_8127,N_8243);
and U8514 (N_8514,N_8054,N_8349);
xnor U8515 (N_8515,N_8147,N_8206);
or U8516 (N_8516,N_8260,N_8044);
nor U8517 (N_8517,N_8342,N_8262);
xor U8518 (N_8518,N_8164,N_8160);
or U8519 (N_8519,N_8247,N_8242);
nor U8520 (N_8520,N_8167,N_8186);
and U8521 (N_8521,N_8060,N_8098);
nand U8522 (N_8522,N_8304,N_8482);
or U8523 (N_8523,N_8006,N_8305);
nor U8524 (N_8524,N_8213,N_8040);
nor U8525 (N_8525,N_8316,N_8465);
nand U8526 (N_8526,N_8226,N_8339);
xor U8527 (N_8527,N_8337,N_8192);
and U8528 (N_8528,N_8086,N_8177);
and U8529 (N_8529,N_8139,N_8053);
nor U8530 (N_8530,N_8464,N_8197);
nor U8531 (N_8531,N_8151,N_8324);
nor U8532 (N_8532,N_8145,N_8463);
and U8533 (N_8533,N_8428,N_8067);
nor U8534 (N_8534,N_8183,N_8115);
nand U8535 (N_8535,N_8495,N_8011);
xor U8536 (N_8536,N_8446,N_8377);
xor U8537 (N_8537,N_8393,N_8355);
or U8538 (N_8538,N_8050,N_8274);
xnor U8539 (N_8539,N_8368,N_8422);
nor U8540 (N_8540,N_8244,N_8130);
nor U8541 (N_8541,N_8443,N_8078);
and U8542 (N_8542,N_8299,N_8180);
or U8543 (N_8543,N_8483,N_8229);
or U8544 (N_8544,N_8387,N_8404);
xor U8545 (N_8545,N_8051,N_8319);
nand U8546 (N_8546,N_8133,N_8036);
and U8547 (N_8547,N_8198,N_8204);
xnor U8548 (N_8548,N_8003,N_8459);
nor U8549 (N_8549,N_8137,N_8271);
xor U8550 (N_8550,N_8158,N_8207);
or U8551 (N_8551,N_8202,N_8336);
nand U8552 (N_8552,N_8072,N_8140);
or U8553 (N_8553,N_8296,N_8048);
xnor U8554 (N_8554,N_8331,N_8175);
nand U8555 (N_8555,N_8058,N_8248);
nor U8556 (N_8556,N_8380,N_8475);
nor U8557 (N_8557,N_8272,N_8093);
xor U8558 (N_8558,N_8128,N_8302);
nor U8559 (N_8559,N_8491,N_8153);
nand U8560 (N_8560,N_8227,N_8090);
nor U8561 (N_8561,N_8341,N_8450);
and U8562 (N_8562,N_8104,N_8497);
and U8563 (N_8563,N_8317,N_8245);
and U8564 (N_8564,N_8170,N_8343);
nand U8565 (N_8565,N_8265,N_8405);
and U8566 (N_8566,N_8390,N_8166);
nand U8567 (N_8567,N_8474,N_8263);
nor U8568 (N_8568,N_8083,N_8320);
xor U8569 (N_8569,N_8400,N_8254);
and U8570 (N_8570,N_8370,N_8020);
nand U8571 (N_8571,N_8079,N_8470);
nand U8572 (N_8572,N_8217,N_8126);
nand U8573 (N_8573,N_8389,N_8436);
xor U8574 (N_8574,N_8410,N_8286);
and U8575 (N_8575,N_8407,N_8315);
nand U8576 (N_8576,N_8434,N_8066);
nor U8577 (N_8577,N_8398,N_8330);
or U8578 (N_8578,N_8125,N_8381);
nor U8579 (N_8579,N_8477,N_8426);
nand U8580 (N_8580,N_8451,N_8224);
nand U8581 (N_8581,N_8418,N_8350);
or U8582 (N_8582,N_8414,N_8258);
and U8583 (N_8583,N_8176,N_8211);
or U8584 (N_8584,N_8494,N_8385);
xnor U8585 (N_8585,N_8279,N_8237);
or U8586 (N_8586,N_8310,N_8362);
or U8587 (N_8587,N_8069,N_8073);
nand U8588 (N_8588,N_8216,N_8332);
nor U8589 (N_8589,N_8291,N_8082);
and U8590 (N_8590,N_8027,N_8225);
or U8591 (N_8591,N_8124,N_8384);
nand U8592 (N_8592,N_8222,N_8046);
nand U8593 (N_8593,N_8107,N_8029);
nand U8594 (N_8594,N_8295,N_8089);
xnor U8595 (N_8595,N_8136,N_8270);
xor U8596 (N_8596,N_8156,N_8037);
and U8597 (N_8597,N_8032,N_8498);
xor U8598 (N_8598,N_8181,N_8255);
and U8599 (N_8599,N_8000,N_8193);
or U8600 (N_8600,N_8018,N_8297);
or U8601 (N_8601,N_8005,N_8490);
xor U8602 (N_8602,N_8019,N_8218);
or U8603 (N_8603,N_8357,N_8257);
or U8604 (N_8604,N_8448,N_8120);
nand U8605 (N_8605,N_8150,N_8173);
xnor U8606 (N_8606,N_8488,N_8352);
nand U8607 (N_8607,N_8172,N_8038);
nand U8608 (N_8608,N_8154,N_8111);
xnor U8609 (N_8609,N_8236,N_8187);
nor U8610 (N_8610,N_8306,N_8009);
xor U8611 (N_8611,N_8201,N_8025);
and U8612 (N_8612,N_8273,N_8161);
and U8613 (N_8613,N_8420,N_8290);
nor U8614 (N_8614,N_8182,N_8219);
nand U8615 (N_8615,N_8416,N_8402);
nand U8616 (N_8616,N_8269,N_8162);
nor U8617 (N_8617,N_8059,N_8303);
nor U8618 (N_8618,N_8472,N_8447);
or U8619 (N_8619,N_8344,N_8076);
nor U8620 (N_8620,N_8462,N_8194);
nor U8621 (N_8621,N_8435,N_8052);
and U8622 (N_8622,N_8184,N_8430);
nor U8623 (N_8623,N_8351,N_8442);
and U8624 (N_8624,N_8460,N_8031);
nor U8625 (N_8625,N_8417,N_8205);
nand U8626 (N_8626,N_8132,N_8449);
xnor U8627 (N_8627,N_8469,N_8250);
nand U8628 (N_8628,N_8041,N_8424);
nand U8629 (N_8629,N_8092,N_8441);
and U8630 (N_8630,N_8015,N_8109);
or U8631 (N_8631,N_8007,N_8088);
nor U8632 (N_8632,N_8457,N_8293);
and U8633 (N_8633,N_8148,N_8345);
nor U8634 (N_8634,N_8325,N_8021);
nand U8635 (N_8635,N_8308,N_8221);
or U8636 (N_8636,N_8371,N_8013);
nand U8637 (N_8637,N_8171,N_8396);
nand U8638 (N_8638,N_8010,N_8057);
or U8639 (N_8639,N_8231,N_8008);
xnor U8640 (N_8640,N_8481,N_8375);
xnor U8641 (N_8641,N_8433,N_8334);
xnor U8642 (N_8642,N_8085,N_8112);
and U8643 (N_8643,N_8095,N_8118);
nor U8644 (N_8644,N_8300,N_8261);
nand U8645 (N_8645,N_8063,N_8196);
xor U8646 (N_8646,N_8264,N_8356);
or U8647 (N_8647,N_8365,N_8281);
or U8648 (N_8648,N_8071,N_8080);
and U8649 (N_8649,N_8397,N_8283);
nand U8650 (N_8650,N_8394,N_8045);
and U8651 (N_8651,N_8493,N_8249);
nor U8652 (N_8652,N_8168,N_8354);
or U8653 (N_8653,N_8106,N_8142);
nor U8654 (N_8654,N_8346,N_8077);
xor U8655 (N_8655,N_8340,N_8146);
and U8656 (N_8656,N_8253,N_8240);
or U8657 (N_8657,N_8372,N_8131);
or U8658 (N_8658,N_8144,N_8277);
and U8659 (N_8659,N_8466,N_8359);
xnor U8660 (N_8660,N_8411,N_8323);
or U8661 (N_8661,N_8333,N_8395);
xnor U8662 (N_8662,N_8454,N_8055);
nor U8663 (N_8663,N_8287,N_8232);
and U8664 (N_8664,N_8386,N_8409);
xnor U8665 (N_8665,N_8406,N_8214);
nor U8666 (N_8666,N_8366,N_8476);
or U8667 (N_8667,N_8313,N_8030);
or U8668 (N_8668,N_8373,N_8292);
and U8669 (N_8669,N_8473,N_8022);
nor U8670 (N_8670,N_8421,N_8049);
xor U8671 (N_8671,N_8311,N_8135);
and U8672 (N_8672,N_8376,N_8399);
xor U8673 (N_8673,N_8122,N_8097);
nor U8674 (N_8674,N_8075,N_8276);
nor U8675 (N_8675,N_8275,N_8492);
nor U8676 (N_8676,N_8412,N_8246);
or U8677 (N_8677,N_8178,N_8487);
and U8678 (N_8678,N_8094,N_8278);
nor U8679 (N_8679,N_8378,N_8119);
xnor U8680 (N_8680,N_8438,N_8121);
nor U8681 (N_8681,N_8208,N_8065);
nand U8682 (N_8682,N_8110,N_8348);
and U8683 (N_8683,N_8403,N_8001);
nand U8684 (N_8684,N_8179,N_8468);
nor U8685 (N_8685,N_8195,N_8100);
nor U8686 (N_8686,N_8230,N_8228);
xor U8687 (N_8687,N_8445,N_8458);
xnor U8688 (N_8688,N_8379,N_8363);
nand U8689 (N_8689,N_8499,N_8456);
nor U8690 (N_8690,N_8423,N_8134);
xor U8691 (N_8691,N_8024,N_8014);
nor U8692 (N_8692,N_8087,N_8401);
nand U8693 (N_8693,N_8096,N_8070);
and U8694 (N_8694,N_8210,N_8062);
or U8695 (N_8695,N_8322,N_8453);
xnor U8696 (N_8696,N_8425,N_8353);
nand U8697 (N_8697,N_8431,N_8383);
or U8698 (N_8698,N_8103,N_8266);
or U8699 (N_8699,N_8212,N_8068);
and U8700 (N_8700,N_8200,N_8486);
or U8701 (N_8701,N_8461,N_8294);
xor U8702 (N_8702,N_8329,N_8489);
and U8703 (N_8703,N_8108,N_8091);
xnor U8704 (N_8704,N_8233,N_8105);
or U8705 (N_8705,N_8471,N_8026);
or U8706 (N_8706,N_8485,N_8074);
nand U8707 (N_8707,N_8039,N_8157);
nand U8708 (N_8708,N_8215,N_8259);
or U8709 (N_8709,N_8419,N_8223);
or U8710 (N_8710,N_8149,N_8043);
nor U8711 (N_8711,N_8155,N_8251);
nor U8712 (N_8712,N_8437,N_8338);
nor U8713 (N_8713,N_8190,N_8189);
nor U8714 (N_8714,N_8252,N_8129);
or U8715 (N_8715,N_8023,N_8004);
or U8716 (N_8716,N_8326,N_8256);
nor U8717 (N_8717,N_8084,N_8288);
or U8718 (N_8718,N_8364,N_8321);
xor U8719 (N_8719,N_8455,N_8141);
or U8720 (N_8720,N_8268,N_8479);
nand U8721 (N_8721,N_8028,N_8312);
or U8722 (N_8722,N_8099,N_8327);
nor U8723 (N_8723,N_8360,N_8174);
xnor U8724 (N_8724,N_8358,N_8439);
xnor U8725 (N_8725,N_8123,N_8429);
or U8726 (N_8726,N_8102,N_8143);
or U8727 (N_8727,N_8367,N_8307);
or U8728 (N_8728,N_8035,N_8427);
or U8729 (N_8729,N_8267,N_8361);
xnor U8730 (N_8730,N_8159,N_8169);
xor U8731 (N_8731,N_8081,N_8238);
or U8732 (N_8732,N_8392,N_8220);
and U8733 (N_8733,N_8165,N_8064);
or U8734 (N_8734,N_8042,N_8234);
xnor U8735 (N_8735,N_8309,N_8033);
or U8736 (N_8736,N_8415,N_8114);
nand U8737 (N_8737,N_8138,N_8285);
xor U8738 (N_8738,N_8235,N_8369);
or U8739 (N_8739,N_8241,N_8199);
xor U8740 (N_8740,N_8117,N_8002);
nor U8741 (N_8741,N_8047,N_8318);
and U8742 (N_8742,N_8467,N_8298);
nand U8743 (N_8743,N_8282,N_8289);
xor U8744 (N_8744,N_8328,N_8413);
or U8745 (N_8745,N_8480,N_8388);
and U8746 (N_8746,N_8209,N_8374);
and U8747 (N_8747,N_8284,N_8034);
or U8748 (N_8748,N_8496,N_8191);
xor U8749 (N_8749,N_8301,N_8188);
and U8750 (N_8750,N_8355,N_8157);
nand U8751 (N_8751,N_8156,N_8366);
xnor U8752 (N_8752,N_8144,N_8173);
nand U8753 (N_8753,N_8442,N_8017);
or U8754 (N_8754,N_8251,N_8259);
xor U8755 (N_8755,N_8032,N_8422);
or U8756 (N_8756,N_8048,N_8274);
and U8757 (N_8757,N_8262,N_8034);
nand U8758 (N_8758,N_8303,N_8116);
xnor U8759 (N_8759,N_8251,N_8234);
or U8760 (N_8760,N_8384,N_8326);
xnor U8761 (N_8761,N_8261,N_8450);
nand U8762 (N_8762,N_8042,N_8006);
nor U8763 (N_8763,N_8484,N_8209);
and U8764 (N_8764,N_8207,N_8423);
and U8765 (N_8765,N_8259,N_8065);
nand U8766 (N_8766,N_8292,N_8283);
or U8767 (N_8767,N_8294,N_8317);
or U8768 (N_8768,N_8008,N_8016);
xor U8769 (N_8769,N_8379,N_8358);
nor U8770 (N_8770,N_8291,N_8205);
xor U8771 (N_8771,N_8104,N_8182);
xor U8772 (N_8772,N_8239,N_8218);
and U8773 (N_8773,N_8202,N_8210);
nor U8774 (N_8774,N_8099,N_8170);
nand U8775 (N_8775,N_8325,N_8113);
or U8776 (N_8776,N_8109,N_8445);
and U8777 (N_8777,N_8271,N_8216);
or U8778 (N_8778,N_8370,N_8457);
and U8779 (N_8779,N_8408,N_8490);
nor U8780 (N_8780,N_8424,N_8499);
xnor U8781 (N_8781,N_8117,N_8438);
xnor U8782 (N_8782,N_8101,N_8176);
xor U8783 (N_8783,N_8175,N_8492);
and U8784 (N_8784,N_8181,N_8457);
nor U8785 (N_8785,N_8176,N_8112);
and U8786 (N_8786,N_8102,N_8267);
xnor U8787 (N_8787,N_8054,N_8072);
nor U8788 (N_8788,N_8006,N_8455);
or U8789 (N_8789,N_8490,N_8338);
or U8790 (N_8790,N_8424,N_8298);
or U8791 (N_8791,N_8293,N_8196);
nor U8792 (N_8792,N_8336,N_8345);
or U8793 (N_8793,N_8349,N_8421);
nand U8794 (N_8794,N_8042,N_8267);
and U8795 (N_8795,N_8153,N_8192);
xnor U8796 (N_8796,N_8390,N_8011);
and U8797 (N_8797,N_8421,N_8385);
xnor U8798 (N_8798,N_8180,N_8416);
nor U8799 (N_8799,N_8329,N_8062);
xnor U8800 (N_8800,N_8322,N_8375);
or U8801 (N_8801,N_8185,N_8159);
or U8802 (N_8802,N_8029,N_8343);
nand U8803 (N_8803,N_8187,N_8498);
xnor U8804 (N_8804,N_8303,N_8070);
or U8805 (N_8805,N_8284,N_8071);
nor U8806 (N_8806,N_8430,N_8389);
or U8807 (N_8807,N_8305,N_8473);
xor U8808 (N_8808,N_8343,N_8371);
nand U8809 (N_8809,N_8447,N_8153);
and U8810 (N_8810,N_8427,N_8050);
and U8811 (N_8811,N_8082,N_8366);
and U8812 (N_8812,N_8323,N_8302);
and U8813 (N_8813,N_8089,N_8424);
or U8814 (N_8814,N_8191,N_8390);
nand U8815 (N_8815,N_8379,N_8424);
nor U8816 (N_8816,N_8381,N_8430);
nand U8817 (N_8817,N_8022,N_8442);
nand U8818 (N_8818,N_8013,N_8059);
nand U8819 (N_8819,N_8399,N_8321);
xnor U8820 (N_8820,N_8112,N_8147);
or U8821 (N_8821,N_8422,N_8114);
nor U8822 (N_8822,N_8281,N_8286);
xor U8823 (N_8823,N_8328,N_8114);
and U8824 (N_8824,N_8468,N_8211);
nand U8825 (N_8825,N_8078,N_8005);
nor U8826 (N_8826,N_8424,N_8284);
nor U8827 (N_8827,N_8234,N_8273);
or U8828 (N_8828,N_8106,N_8165);
nand U8829 (N_8829,N_8413,N_8054);
or U8830 (N_8830,N_8263,N_8143);
xnor U8831 (N_8831,N_8481,N_8198);
nand U8832 (N_8832,N_8252,N_8457);
and U8833 (N_8833,N_8008,N_8159);
nand U8834 (N_8834,N_8313,N_8414);
xnor U8835 (N_8835,N_8296,N_8172);
nor U8836 (N_8836,N_8262,N_8176);
or U8837 (N_8837,N_8443,N_8238);
and U8838 (N_8838,N_8200,N_8378);
nand U8839 (N_8839,N_8156,N_8360);
nor U8840 (N_8840,N_8071,N_8005);
xor U8841 (N_8841,N_8004,N_8134);
nand U8842 (N_8842,N_8087,N_8124);
and U8843 (N_8843,N_8409,N_8222);
nand U8844 (N_8844,N_8464,N_8440);
or U8845 (N_8845,N_8185,N_8383);
and U8846 (N_8846,N_8419,N_8398);
nand U8847 (N_8847,N_8271,N_8406);
nor U8848 (N_8848,N_8185,N_8270);
nor U8849 (N_8849,N_8016,N_8290);
or U8850 (N_8850,N_8281,N_8034);
nand U8851 (N_8851,N_8066,N_8356);
nand U8852 (N_8852,N_8401,N_8225);
xnor U8853 (N_8853,N_8239,N_8112);
and U8854 (N_8854,N_8138,N_8115);
nor U8855 (N_8855,N_8159,N_8193);
or U8856 (N_8856,N_8006,N_8472);
nand U8857 (N_8857,N_8494,N_8482);
nand U8858 (N_8858,N_8224,N_8394);
xnor U8859 (N_8859,N_8193,N_8467);
nand U8860 (N_8860,N_8409,N_8244);
nand U8861 (N_8861,N_8491,N_8313);
nor U8862 (N_8862,N_8326,N_8129);
xnor U8863 (N_8863,N_8166,N_8049);
nand U8864 (N_8864,N_8158,N_8228);
nor U8865 (N_8865,N_8417,N_8214);
and U8866 (N_8866,N_8255,N_8470);
nand U8867 (N_8867,N_8481,N_8001);
or U8868 (N_8868,N_8028,N_8460);
nand U8869 (N_8869,N_8410,N_8100);
nor U8870 (N_8870,N_8276,N_8020);
or U8871 (N_8871,N_8102,N_8227);
and U8872 (N_8872,N_8481,N_8183);
nor U8873 (N_8873,N_8076,N_8142);
nand U8874 (N_8874,N_8144,N_8179);
nor U8875 (N_8875,N_8469,N_8239);
or U8876 (N_8876,N_8035,N_8380);
xnor U8877 (N_8877,N_8434,N_8193);
nand U8878 (N_8878,N_8309,N_8010);
nand U8879 (N_8879,N_8492,N_8485);
or U8880 (N_8880,N_8216,N_8246);
xor U8881 (N_8881,N_8448,N_8000);
and U8882 (N_8882,N_8032,N_8231);
xor U8883 (N_8883,N_8491,N_8319);
nor U8884 (N_8884,N_8091,N_8462);
and U8885 (N_8885,N_8457,N_8134);
and U8886 (N_8886,N_8279,N_8116);
and U8887 (N_8887,N_8268,N_8032);
nor U8888 (N_8888,N_8183,N_8339);
nand U8889 (N_8889,N_8150,N_8035);
nor U8890 (N_8890,N_8224,N_8411);
nand U8891 (N_8891,N_8004,N_8080);
xor U8892 (N_8892,N_8067,N_8189);
and U8893 (N_8893,N_8444,N_8227);
or U8894 (N_8894,N_8167,N_8438);
nor U8895 (N_8895,N_8065,N_8329);
xor U8896 (N_8896,N_8209,N_8095);
nand U8897 (N_8897,N_8275,N_8359);
nor U8898 (N_8898,N_8029,N_8287);
and U8899 (N_8899,N_8464,N_8043);
and U8900 (N_8900,N_8070,N_8467);
and U8901 (N_8901,N_8310,N_8152);
or U8902 (N_8902,N_8223,N_8203);
xor U8903 (N_8903,N_8423,N_8346);
or U8904 (N_8904,N_8206,N_8355);
and U8905 (N_8905,N_8457,N_8378);
nand U8906 (N_8906,N_8495,N_8002);
nor U8907 (N_8907,N_8092,N_8235);
and U8908 (N_8908,N_8249,N_8190);
and U8909 (N_8909,N_8043,N_8093);
or U8910 (N_8910,N_8019,N_8405);
xnor U8911 (N_8911,N_8460,N_8370);
nor U8912 (N_8912,N_8084,N_8203);
nor U8913 (N_8913,N_8388,N_8210);
or U8914 (N_8914,N_8132,N_8303);
nand U8915 (N_8915,N_8070,N_8202);
nor U8916 (N_8916,N_8061,N_8365);
xnor U8917 (N_8917,N_8016,N_8098);
or U8918 (N_8918,N_8112,N_8028);
or U8919 (N_8919,N_8319,N_8238);
and U8920 (N_8920,N_8363,N_8016);
xnor U8921 (N_8921,N_8207,N_8290);
or U8922 (N_8922,N_8249,N_8301);
and U8923 (N_8923,N_8387,N_8186);
xnor U8924 (N_8924,N_8351,N_8107);
xnor U8925 (N_8925,N_8413,N_8169);
or U8926 (N_8926,N_8108,N_8259);
nand U8927 (N_8927,N_8442,N_8461);
xnor U8928 (N_8928,N_8206,N_8041);
nor U8929 (N_8929,N_8316,N_8374);
nand U8930 (N_8930,N_8490,N_8498);
xor U8931 (N_8931,N_8272,N_8090);
nor U8932 (N_8932,N_8026,N_8345);
and U8933 (N_8933,N_8418,N_8437);
xnor U8934 (N_8934,N_8089,N_8120);
nand U8935 (N_8935,N_8117,N_8011);
and U8936 (N_8936,N_8006,N_8133);
xnor U8937 (N_8937,N_8037,N_8210);
nand U8938 (N_8938,N_8367,N_8041);
xnor U8939 (N_8939,N_8254,N_8273);
nor U8940 (N_8940,N_8099,N_8275);
nor U8941 (N_8941,N_8160,N_8267);
xor U8942 (N_8942,N_8207,N_8089);
and U8943 (N_8943,N_8171,N_8241);
and U8944 (N_8944,N_8304,N_8293);
nand U8945 (N_8945,N_8459,N_8144);
xnor U8946 (N_8946,N_8321,N_8173);
or U8947 (N_8947,N_8035,N_8288);
and U8948 (N_8948,N_8250,N_8433);
and U8949 (N_8949,N_8219,N_8063);
xor U8950 (N_8950,N_8211,N_8022);
xor U8951 (N_8951,N_8471,N_8148);
and U8952 (N_8952,N_8187,N_8226);
nor U8953 (N_8953,N_8457,N_8300);
nor U8954 (N_8954,N_8124,N_8137);
or U8955 (N_8955,N_8094,N_8228);
nor U8956 (N_8956,N_8037,N_8111);
or U8957 (N_8957,N_8232,N_8452);
and U8958 (N_8958,N_8398,N_8431);
nor U8959 (N_8959,N_8489,N_8425);
and U8960 (N_8960,N_8270,N_8404);
and U8961 (N_8961,N_8304,N_8069);
nand U8962 (N_8962,N_8239,N_8332);
and U8963 (N_8963,N_8495,N_8462);
or U8964 (N_8964,N_8395,N_8125);
nand U8965 (N_8965,N_8484,N_8343);
or U8966 (N_8966,N_8002,N_8485);
or U8967 (N_8967,N_8212,N_8349);
or U8968 (N_8968,N_8376,N_8028);
or U8969 (N_8969,N_8425,N_8453);
nor U8970 (N_8970,N_8316,N_8425);
nor U8971 (N_8971,N_8364,N_8089);
xnor U8972 (N_8972,N_8012,N_8281);
and U8973 (N_8973,N_8017,N_8327);
nand U8974 (N_8974,N_8310,N_8259);
nand U8975 (N_8975,N_8112,N_8285);
nand U8976 (N_8976,N_8292,N_8106);
nor U8977 (N_8977,N_8357,N_8381);
xnor U8978 (N_8978,N_8395,N_8086);
and U8979 (N_8979,N_8039,N_8081);
and U8980 (N_8980,N_8292,N_8193);
nor U8981 (N_8981,N_8066,N_8014);
xor U8982 (N_8982,N_8346,N_8124);
nor U8983 (N_8983,N_8450,N_8055);
xor U8984 (N_8984,N_8229,N_8305);
and U8985 (N_8985,N_8033,N_8423);
xnor U8986 (N_8986,N_8022,N_8011);
or U8987 (N_8987,N_8205,N_8337);
and U8988 (N_8988,N_8276,N_8319);
and U8989 (N_8989,N_8179,N_8479);
or U8990 (N_8990,N_8414,N_8050);
nor U8991 (N_8991,N_8167,N_8305);
nor U8992 (N_8992,N_8412,N_8438);
nor U8993 (N_8993,N_8024,N_8337);
nand U8994 (N_8994,N_8451,N_8010);
xor U8995 (N_8995,N_8415,N_8121);
and U8996 (N_8996,N_8204,N_8425);
nand U8997 (N_8997,N_8455,N_8022);
nand U8998 (N_8998,N_8198,N_8048);
and U8999 (N_8999,N_8282,N_8119);
and U9000 (N_9000,N_8901,N_8801);
xor U9001 (N_9001,N_8780,N_8894);
and U9002 (N_9002,N_8590,N_8524);
or U9003 (N_9003,N_8976,N_8807);
and U9004 (N_9004,N_8935,N_8567);
and U9005 (N_9005,N_8815,N_8881);
nor U9006 (N_9006,N_8650,N_8861);
xor U9007 (N_9007,N_8790,N_8566);
or U9008 (N_9008,N_8616,N_8765);
nand U9009 (N_9009,N_8946,N_8930);
xnor U9010 (N_9010,N_8809,N_8731);
nor U9011 (N_9011,N_8793,N_8867);
nand U9012 (N_9012,N_8882,N_8820);
and U9013 (N_9013,N_8938,N_8663);
nor U9014 (N_9014,N_8942,N_8971);
xor U9015 (N_9015,N_8680,N_8887);
or U9016 (N_9016,N_8763,N_8506);
and U9017 (N_9017,N_8692,N_8899);
nor U9018 (N_9018,N_8510,N_8501);
and U9019 (N_9019,N_8905,N_8879);
and U9020 (N_9020,N_8522,N_8551);
xnor U9021 (N_9021,N_8963,N_8577);
or U9022 (N_9022,N_8523,N_8778);
and U9023 (N_9023,N_8592,N_8825);
or U9024 (N_9024,N_8803,N_8742);
or U9025 (N_9025,N_8579,N_8621);
nand U9026 (N_9026,N_8540,N_8814);
and U9027 (N_9027,N_8827,N_8953);
xor U9028 (N_9028,N_8569,N_8535);
xor U9029 (N_9029,N_8955,N_8915);
and U9030 (N_9030,N_8728,N_8533);
nand U9031 (N_9031,N_8902,N_8829);
xor U9032 (N_9032,N_8860,N_8549);
xnor U9033 (N_9033,N_8805,N_8896);
nand U9034 (N_9034,N_8545,N_8858);
or U9035 (N_9035,N_8673,N_8676);
nand U9036 (N_9036,N_8672,N_8812);
and U9037 (N_9037,N_8695,N_8679);
and U9038 (N_9038,N_8924,N_8707);
nand U9039 (N_9039,N_8652,N_8844);
nand U9040 (N_9040,N_8677,N_8993);
or U9041 (N_9041,N_8624,N_8697);
or U9042 (N_9042,N_8968,N_8768);
nand U9043 (N_9043,N_8589,N_8872);
or U9044 (N_9044,N_8618,N_8956);
nor U9045 (N_9045,N_8675,N_8594);
or U9046 (N_9046,N_8819,N_8727);
or U9047 (N_9047,N_8880,N_8772);
nand U9048 (N_9048,N_8684,N_8761);
nand U9049 (N_9049,N_8746,N_8563);
and U9050 (N_9050,N_8631,N_8989);
nand U9051 (N_9051,N_8668,N_8611);
and U9052 (N_9052,N_8840,N_8623);
nor U9053 (N_9053,N_8914,N_8713);
nor U9054 (N_9054,N_8913,N_8775);
xnor U9055 (N_9055,N_8599,N_8889);
nand U9056 (N_9056,N_8568,N_8512);
nand U9057 (N_9057,N_8705,N_8646);
and U9058 (N_9058,N_8620,N_8947);
nand U9059 (N_9059,N_8674,N_8565);
xnor U9060 (N_9060,N_8641,N_8527);
nor U9061 (N_9061,N_8700,N_8683);
nand U9062 (N_9062,N_8838,N_8588);
nor U9063 (N_9063,N_8874,N_8559);
nand U9064 (N_9064,N_8714,N_8831);
nand U9065 (N_9065,N_8910,N_8762);
nor U9066 (N_9066,N_8800,N_8606);
nor U9067 (N_9067,N_8550,N_8810);
and U9068 (N_9068,N_8632,N_8521);
nor U9069 (N_9069,N_8647,N_8633);
nand U9070 (N_9070,N_8835,N_8669);
xor U9071 (N_9071,N_8863,N_8767);
nand U9072 (N_9072,N_8597,N_8857);
nor U9073 (N_9073,N_8974,N_8784);
and U9074 (N_9074,N_8954,N_8659);
or U9075 (N_9075,N_8733,N_8515);
xnor U9076 (N_9076,N_8785,N_8824);
xnor U9077 (N_9077,N_8922,N_8529);
and U9078 (N_9078,N_8629,N_8717);
nand U9079 (N_9079,N_8667,N_8759);
nand U9080 (N_9080,N_8917,N_8895);
or U9081 (N_9081,N_8712,N_8797);
nand U9082 (N_9082,N_8747,N_8514);
nand U9083 (N_9083,N_8834,N_8586);
xnor U9084 (N_9084,N_8998,N_8836);
xor U9085 (N_9085,N_8926,N_8817);
and U9086 (N_9086,N_8525,N_8970);
nand U9087 (N_9087,N_8898,N_8859);
nor U9088 (N_9088,N_8711,N_8709);
and U9089 (N_9089,N_8997,N_8919);
and U9090 (N_9090,N_8832,N_8511);
or U9091 (N_9091,N_8945,N_8878);
nor U9092 (N_9092,N_8552,N_8749);
and U9093 (N_9093,N_8718,N_8554);
xnor U9094 (N_9094,N_8702,N_8774);
xnor U9095 (N_9095,N_8601,N_8741);
nor U9096 (N_9096,N_8977,N_8973);
nand U9097 (N_9097,N_8833,N_8873);
and U9098 (N_9098,N_8936,N_8609);
nor U9099 (N_9099,N_8958,N_8724);
nand U9100 (N_9100,N_8622,N_8757);
or U9101 (N_9101,N_8806,N_8986);
nand U9102 (N_9102,N_8939,N_8595);
nand U9103 (N_9103,N_8852,N_8781);
and U9104 (N_9104,N_8870,N_8804);
and U9105 (N_9105,N_8980,N_8990);
and U9106 (N_9106,N_8773,N_8703);
or U9107 (N_9107,N_8580,N_8520);
xor U9108 (N_9108,N_8900,N_8735);
or U9109 (N_9109,N_8690,N_8918);
nand U9110 (N_9110,N_8888,N_8694);
or U9111 (N_9111,N_8605,N_8587);
xnor U9112 (N_9112,N_8604,N_8513);
nand U9113 (N_9113,N_8755,N_8612);
or U9114 (N_9114,N_8754,N_8725);
and U9115 (N_9115,N_8634,N_8992);
or U9116 (N_9116,N_8940,N_8658);
nor U9117 (N_9117,N_8813,N_8642);
nand U9118 (N_9118,N_8734,N_8967);
nand U9119 (N_9119,N_8987,N_8999);
or U9120 (N_9120,N_8644,N_8526);
or U9121 (N_9121,N_8931,N_8584);
or U9122 (N_9122,N_8822,N_8625);
nor U9123 (N_9123,N_8837,N_8903);
nor U9124 (N_9124,N_8950,N_8908);
xnor U9125 (N_9125,N_8541,N_8504);
nor U9126 (N_9126,N_8932,N_8855);
xor U9127 (N_9127,N_8706,N_8869);
or U9128 (N_9128,N_8560,N_8508);
and U9129 (N_9129,N_8710,N_8626);
and U9130 (N_9130,N_8885,N_8897);
nor U9131 (N_9131,N_8651,N_8591);
or U9132 (N_9132,N_8614,N_8635);
xnor U9133 (N_9133,N_8720,N_8505);
and U9134 (N_9134,N_8701,N_8909);
xnor U9135 (N_9135,N_8912,N_8516);
nand U9136 (N_9136,N_8681,N_8722);
or U9137 (N_9137,N_8553,N_8729);
and U9138 (N_9138,N_8818,N_8839);
nand U9139 (N_9139,N_8583,N_8744);
or U9140 (N_9140,N_8911,N_8661);
and U9141 (N_9141,N_8556,N_8868);
nand U9142 (N_9142,N_8688,N_8699);
xnor U9143 (N_9143,N_8730,N_8608);
nor U9144 (N_9144,N_8928,N_8862);
or U9145 (N_9145,N_8978,N_8962);
xnor U9146 (N_9146,N_8920,N_8685);
xnor U9147 (N_9147,N_8794,N_8937);
and U9148 (N_9148,N_8687,N_8600);
nor U9149 (N_9149,N_8983,N_8921);
xnor U9150 (N_9150,N_8751,N_8994);
xor U9151 (N_9151,N_8715,N_8666);
and U9152 (N_9152,N_8846,N_8607);
or U9153 (N_9153,N_8509,N_8648);
xor U9154 (N_9154,N_8984,N_8538);
xnor U9155 (N_9155,N_8670,N_8948);
or U9156 (N_9156,N_8581,N_8788);
nand U9157 (N_9157,N_8830,N_8960);
nor U9158 (N_9158,N_8649,N_8791);
and U9159 (N_9159,N_8573,N_8517);
nand U9160 (N_9160,N_8877,N_8555);
nor U9161 (N_9161,N_8638,N_8544);
or U9162 (N_9162,N_8764,N_8941);
nor U9163 (N_9163,N_8854,N_8528);
xnor U9164 (N_9164,N_8721,N_8795);
xnor U9165 (N_9165,N_8662,N_8548);
or U9166 (N_9166,N_8726,N_8723);
nand U9167 (N_9167,N_8906,N_8850);
or U9168 (N_9168,N_8886,N_8656);
nor U9169 (N_9169,N_8864,N_8578);
nor U9170 (N_9170,N_8637,N_8756);
nor U9171 (N_9171,N_8585,N_8853);
and U9172 (N_9172,N_8923,N_8871);
and U9173 (N_9173,N_8750,N_8570);
nor U9174 (N_9174,N_8891,N_8949);
nor U9175 (N_9175,N_8671,N_8500);
xor U9176 (N_9176,N_8883,N_8865);
nand U9177 (N_9177,N_8654,N_8708);
nand U9178 (N_9178,N_8686,N_8816);
nor U9179 (N_9179,N_8982,N_8849);
xor U9180 (N_9180,N_8736,N_8798);
xnor U9181 (N_9181,N_8503,N_8678);
nor U9182 (N_9182,N_8575,N_8536);
nand U9183 (N_9183,N_8691,N_8653);
or U9184 (N_9184,N_8696,N_8617);
or U9185 (N_9185,N_8952,N_8969);
nand U9186 (N_9186,N_8802,N_8664);
nand U9187 (N_9187,N_8826,N_8636);
nor U9188 (N_9188,N_8934,N_8619);
or U9189 (N_9189,N_8657,N_8907);
nand U9190 (N_9190,N_8739,N_8786);
nor U9191 (N_9191,N_8593,N_8966);
and U9192 (N_9192,N_8776,N_8777);
nand U9193 (N_9193,N_8539,N_8975);
or U9194 (N_9194,N_8848,N_8890);
and U9195 (N_9195,N_8602,N_8760);
xnor U9196 (N_9196,N_8655,N_8665);
xnor U9197 (N_9197,N_8979,N_8689);
nor U9198 (N_9198,N_8972,N_8787);
nor U9199 (N_9199,N_8719,N_8643);
and U9200 (N_9200,N_8640,N_8933);
xor U9201 (N_9201,N_8660,N_8847);
xor U9202 (N_9202,N_8738,N_8603);
or U9203 (N_9203,N_8766,N_8995);
nor U9204 (N_9204,N_8758,N_8951);
nand U9205 (N_9205,N_8698,N_8875);
and U9206 (N_9206,N_8502,N_8743);
nand U9207 (N_9207,N_8916,N_8682);
xor U9208 (N_9208,N_8530,N_8630);
xor U9209 (N_9209,N_8799,N_8925);
nand U9210 (N_9210,N_8811,N_8964);
nor U9211 (N_9211,N_8792,N_8856);
and U9212 (N_9212,N_8789,N_8534);
nand U9213 (N_9213,N_8531,N_8927);
or U9214 (N_9214,N_8537,N_8866);
and U9215 (N_9215,N_8843,N_8543);
and U9216 (N_9216,N_8753,N_8740);
nor U9217 (N_9217,N_8845,N_8828);
and U9218 (N_9218,N_8904,N_8532);
nand U9219 (N_9219,N_8893,N_8991);
xor U9220 (N_9220,N_8821,N_8598);
xor U9221 (N_9221,N_8518,N_8929);
or U9222 (N_9222,N_8716,N_8752);
nand U9223 (N_9223,N_8613,N_8745);
nand U9224 (N_9224,N_8985,N_8769);
nor U9225 (N_9225,N_8693,N_8639);
or U9226 (N_9226,N_8610,N_8996);
or U9227 (N_9227,N_8562,N_8576);
or U9228 (N_9228,N_8704,N_8546);
or U9229 (N_9229,N_8732,N_8771);
or U9230 (N_9230,N_8558,N_8782);
and U9231 (N_9231,N_8574,N_8582);
and U9232 (N_9232,N_8957,N_8823);
nor U9233 (N_9233,N_8988,N_8961);
or U9234 (N_9234,N_8572,N_8851);
xor U9235 (N_9235,N_8628,N_8507);
xor U9236 (N_9236,N_8943,N_8876);
xnor U9237 (N_9237,N_8944,N_8615);
and U9238 (N_9238,N_8571,N_8884);
or U9239 (N_9239,N_8892,N_8770);
or U9240 (N_9240,N_8965,N_8557);
or U9241 (N_9241,N_8779,N_8737);
nor U9242 (N_9242,N_8542,N_8808);
nor U9243 (N_9243,N_8981,N_8547);
or U9244 (N_9244,N_8596,N_8842);
xor U9245 (N_9245,N_8748,N_8959);
xnor U9246 (N_9246,N_8564,N_8561);
xnor U9247 (N_9247,N_8783,N_8627);
xnor U9248 (N_9248,N_8519,N_8796);
nand U9249 (N_9249,N_8645,N_8841);
nand U9250 (N_9250,N_8701,N_8798);
or U9251 (N_9251,N_8911,N_8626);
and U9252 (N_9252,N_8765,N_8656);
and U9253 (N_9253,N_8902,N_8952);
and U9254 (N_9254,N_8558,N_8549);
and U9255 (N_9255,N_8589,N_8795);
nand U9256 (N_9256,N_8682,N_8997);
or U9257 (N_9257,N_8944,N_8735);
or U9258 (N_9258,N_8759,N_8780);
and U9259 (N_9259,N_8670,N_8672);
nor U9260 (N_9260,N_8580,N_8747);
and U9261 (N_9261,N_8775,N_8929);
xnor U9262 (N_9262,N_8754,N_8916);
or U9263 (N_9263,N_8912,N_8674);
nor U9264 (N_9264,N_8845,N_8614);
nor U9265 (N_9265,N_8915,N_8699);
or U9266 (N_9266,N_8822,N_8558);
nand U9267 (N_9267,N_8981,N_8991);
xnor U9268 (N_9268,N_8582,N_8567);
or U9269 (N_9269,N_8736,N_8952);
nor U9270 (N_9270,N_8980,N_8637);
nor U9271 (N_9271,N_8652,N_8557);
nor U9272 (N_9272,N_8887,N_8512);
and U9273 (N_9273,N_8551,N_8990);
or U9274 (N_9274,N_8661,N_8528);
nand U9275 (N_9275,N_8658,N_8539);
nand U9276 (N_9276,N_8577,N_8844);
nor U9277 (N_9277,N_8994,N_8520);
or U9278 (N_9278,N_8984,N_8880);
xnor U9279 (N_9279,N_8939,N_8558);
nor U9280 (N_9280,N_8804,N_8893);
xnor U9281 (N_9281,N_8638,N_8629);
and U9282 (N_9282,N_8896,N_8826);
nand U9283 (N_9283,N_8688,N_8531);
and U9284 (N_9284,N_8588,N_8604);
nor U9285 (N_9285,N_8578,N_8776);
and U9286 (N_9286,N_8593,N_8812);
nor U9287 (N_9287,N_8790,N_8828);
nor U9288 (N_9288,N_8581,N_8881);
nand U9289 (N_9289,N_8848,N_8714);
xor U9290 (N_9290,N_8548,N_8671);
and U9291 (N_9291,N_8612,N_8724);
nand U9292 (N_9292,N_8534,N_8877);
or U9293 (N_9293,N_8648,N_8877);
nand U9294 (N_9294,N_8864,N_8869);
and U9295 (N_9295,N_8652,N_8841);
nor U9296 (N_9296,N_8689,N_8632);
nand U9297 (N_9297,N_8897,N_8551);
nor U9298 (N_9298,N_8671,N_8549);
nand U9299 (N_9299,N_8923,N_8866);
nand U9300 (N_9300,N_8645,N_8684);
nor U9301 (N_9301,N_8712,N_8571);
and U9302 (N_9302,N_8512,N_8934);
xnor U9303 (N_9303,N_8966,N_8651);
and U9304 (N_9304,N_8825,N_8703);
nand U9305 (N_9305,N_8905,N_8950);
xor U9306 (N_9306,N_8606,N_8743);
nand U9307 (N_9307,N_8819,N_8766);
nor U9308 (N_9308,N_8597,N_8629);
xnor U9309 (N_9309,N_8562,N_8652);
nand U9310 (N_9310,N_8783,N_8531);
nor U9311 (N_9311,N_8906,N_8641);
and U9312 (N_9312,N_8911,N_8865);
nand U9313 (N_9313,N_8995,N_8779);
nor U9314 (N_9314,N_8528,N_8783);
and U9315 (N_9315,N_8671,N_8923);
nand U9316 (N_9316,N_8757,N_8682);
and U9317 (N_9317,N_8625,N_8821);
or U9318 (N_9318,N_8538,N_8762);
or U9319 (N_9319,N_8740,N_8700);
nand U9320 (N_9320,N_8701,N_8523);
xnor U9321 (N_9321,N_8537,N_8541);
or U9322 (N_9322,N_8643,N_8562);
or U9323 (N_9323,N_8705,N_8600);
xor U9324 (N_9324,N_8594,N_8632);
nor U9325 (N_9325,N_8832,N_8733);
xnor U9326 (N_9326,N_8948,N_8506);
nor U9327 (N_9327,N_8947,N_8522);
nor U9328 (N_9328,N_8773,N_8866);
or U9329 (N_9329,N_8565,N_8563);
or U9330 (N_9330,N_8781,N_8806);
and U9331 (N_9331,N_8920,N_8679);
nor U9332 (N_9332,N_8690,N_8604);
xor U9333 (N_9333,N_8505,N_8696);
and U9334 (N_9334,N_8800,N_8969);
nor U9335 (N_9335,N_8613,N_8650);
or U9336 (N_9336,N_8968,N_8920);
nor U9337 (N_9337,N_8972,N_8733);
or U9338 (N_9338,N_8975,N_8957);
or U9339 (N_9339,N_8949,N_8548);
and U9340 (N_9340,N_8522,N_8797);
or U9341 (N_9341,N_8657,N_8837);
or U9342 (N_9342,N_8794,N_8679);
and U9343 (N_9343,N_8523,N_8615);
nand U9344 (N_9344,N_8836,N_8588);
and U9345 (N_9345,N_8861,N_8511);
or U9346 (N_9346,N_8983,N_8667);
and U9347 (N_9347,N_8544,N_8891);
and U9348 (N_9348,N_8703,N_8610);
and U9349 (N_9349,N_8603,N_8531);
nand U9350 (N_9350,N_8951,N_8566);
nand U9351 (N_9351,N_8564,N_8792);
and U9352 (N_9352,N_8697,N_8625);
nor U9353 (N_9353,N_8621,N_8924);
and U9354 (N_9354,N_8603,N_8949);
nor U9355 (N_9355,N_8763,N_8963);
nand U9356 (N_9356,N_8525,N_8543);
xor U9357 (N_9357,N_8932,N_8810);
and U9358 (N_9358,N_8587,N_8814);
nand U9359 (N_9359,N_8550,N_8933);
nor U9360 (N_9360,N_8896,N_8880);
or U9361 (N_9361,N_8967,N_8563);
xnor U9362 (N_9362,N_8959,N_8571);
or U9363 (N_9363,N_8812,N_8580);
xor U9364 (N_9364,N_8699,N_8558);
and U9365 (N_9365,N_8620,N_8805);
and U9366 (N_9366,N_8686,N_8571);
nand U9367 (N_9367,N_8884,N_8763);
nand U9368 (N_9368,N_8786,N_8820);
or U9369 (N_9369,N_8942,N_8730);
xnor U9370 (N_9370,N_8734,N_8588);
nor U9371 (N_9371,N_8959,N_8538);
nand U9372 (N_9372,N_8806,N_8938);
nor U9373 (N_9373,N_8732,N_8634);
and U9374 (N_9374,N_8908,N_8797);
nand U9375 (N_9375,N_8695,N_8703);
and U9376 (N_9376,N_8855,N_8725);
and U9377 (N_9377,N_8754,N_8649);
nand U9378 (N_9378,N_8772,N_8621);
and U9379 (N_9379,N_8848,N_8878);
nor U9380 (N_9380,N_8833,N_8543);
nor U9381 (N_9381,N_8713,N_8773);
or U9382 (N_9382,N_8587,N_8656);
and U9383 (N_9383,N_8776,N_8510);
and U9384 (N_9384,N_8688,N_8973);
nor U9385 (N_9385,N_8921,N_8512);
or U9386 (N_9386,N_8881,N_8637);
or U9387 (N_9387,N_8672,N_8865);
nand U9388 (N_9388,N_8658,N_8504);
nor U9389 (N_9389,N_8511,N_8608);
xnor U9390 (N_9390,N_8701,N_8969);
xnor U9391 (N_9391,N_8991,N_8754);
nor U9392 (N_9392,N_8546,N_8913);
nor U9393 (N_9393,N_8671,N_8704);
or U9394 (N_9394,N_8530,N_8992);
or U9395 (N_9395,N_8822,N_8954);
or U9396 (N_9396,N_8653,N_8789);
and U9397 (N_9397,N_8806,N_8675);
nand U9398 (N_9398,N_8811,N_8777);
and U9399 (N_9399,N_8708,N_8805);
or U9400 (N_9400,N_8533,N_8727);
or U9401 (N_9401,N_8887,N_8563);
and U9402 (N_9402,N_8967,N_8625);
nand U9403 (N_9403,N_8782,N_8792);
or U9404 (N_9404,N_8989,N_8697);
and U9405 (N_9405,N_8543,N_8954);
xor U9406 (N_9406,N_8849,N_8978);
and U9407 (N_9407,N_8850,N_8901);
nand U9408 (N_9408,N_8780,N_8576);
and U9409 (N_9409,N_8937,N_8528);
nor U9410 (N_9410,N_8969,N_8767);
xnor U9411 (N_9411,N_8553,N_8680);
nor U9412 (N_9412,N_8667,N_8705);
and U9413 (N_9413,N_8991,N_8647);
xnor U9414 (N_9414,N_8776,N_8546);
nor U9415 (N_9415,N_8705,N_8887);
nand U9416 (N_9416,N_8828,N_8987);
nor U9417 (N_9417,N_8711,N_8736);
or U9418 (N_9418,N_8574,N_8809);
nand U9419 (N_9419,N_8954,N_8948);
xor U9420 (N_9420,N_8926,N_8707);
and U9421 (N_9421,N_8822,N_8903);
or U9422 (N_9422,N_8506,N_8634);
nor U9423 (N_9423,N_8838,N_8931);
xnor U9424 (N_9424,N_8666,N_8943);
and U9425 (N_9425,N_8671,N_8895);
nor U9426 (N_9426,N_8555,N_8904);
xor U9427 (N_9427,N_8718,N_8923);
or U9428 (N_9428,N_8802,N_8792);
nor U9429 (N_9429,N_8680,N_8672);
nor U9430 (N_9430,N_8525,N_8504);
xnor U9431 (N_9431,N_8521,N_8643);
or U9432 (N_9432,N_8973,N_8689);
nand U9433 (N_9433,N_8730,N_8733);
or U9434 (N_9434,N_8947,N_8610);
nand U9435 (N_9435,N_8782,N_8902);
nand U9436 (N_9436,N_8688,N_8749);
xnor U9437 (N_9437,N_8550,N_8610);
nand U9438 (N_9438,N_8889,N_8757);
and U9439 (N_9439,N_8870,N_8915);
nor U9440 (N_9440,N_8784,N_8555);
and U9441 (N_9441,N_8559,N_8716);
nand U9442 (N_9442,N_8998,N_8921);
nand U9443 (N_9443,N_8924,N_8677);
and U9444 (N_9444,N_8597,N_8736);
xnor U9445 (N_9445,N_8653,N_8595);
xnor U9446 (N_9446,N_8665,N_8690);
xor U9447 (N_9447,N_8778,N_8952);
or U9448 (N_9448,N_8897,N_8846);
nor U9449 (N_9449,N_8780,N_8767);
and U9450 (N_9450,N_8802,N_8832);
nand U9451 (N_9451,N_8825,N_8754);
or U9452 (N_9452,N_8689,N_8980);
nand U9453 (N_9453,N_8729,N_8735);
nand U9454 (N_9454,N_8805,N_8946);
nand U9455 (N_9455,N_8898,N_8860);
nand U9456 (N_9456,N_8910,N_8505);
and U9457 (N_9457,N_8770,N_8611);
xor U9458 (N_9458,N_8620,N_8576);
nand U9459 (N_9459,N_8684,N_8870);
and U9460 (N_9460,N_8869,N_8975);
nor U9461 (N_9461,N_8532,N_8718);
xnor U9462 (N_9462,N_8939,N_8589);
nand U9463 (N_9463,N_8818,N_8719);
or U9464 (N_9464,N_8903,N_8919);
nand U9465 (N_9465,N_8507,N_8983);
nand U9466 (N_9466,N_8768,N_8678);
and U9467 (N_9467,N_8797,N_8762);
nand U9468 (N_9468,N_8506,N_8841);
or U9469 (N_9469,N_8994,N_8555);
xnor U9470 (N_9470,N_8888,N_8785);
and U9471 (N_9471,N_8758,N_8766);
xor U9472 (N_9472,N_8953,N_8965);
xor U9473 (N_9473,N_8818,N_8848);
or U9474 (N_9474,N_8652,N_8866);
nand U9475 (N_9475,N_8621,N_8944);
nor U9476 (N_9476,N_8825,N_8724);
and U9477 (N_9477,N_8737,N_8823);
xnor U9478 (N_9478,N_8761,N_8780);
xnor U9479 (N_9479,N_8895,N_8619);
nand U9480 (N_9480,N_8991,N_8531);
or U9481 (N_9481,N_8809,N_8694);
and U9482 (N_9482,N_8924,N_8865);
nor U9483 (N_9483,N_8649,N_8773);
nand U9484 (N_9484,N_8665,N_8629);
nand U9485 (N_9485,N_8919,N_8651);
or U9486 (N_9486,N_8749,N_8830);
xor U9487 (N_9487,N_8528,N_8799);
nor U9488 (N_9488,N_8899,N_8837);
nand U9489 (N_9489,N_8947,N_8597);
nand U9490 (N_9490,N_8991,N_8968);
nand U9491 (N_9491,N_8984,N_8684);
nor U9492 (N_9492,N_8888,N_8817);
or U9493 (N_9493,N_8628,N_8885);
xnor U9494 (N_9494,N_8740,N_8737);
nor U9495 (N_9495,N_8999,N_8504);
nand U9496 (N_9496,N_8882,N_8530);
xor U9497 (N_9497,N_8856,N_8836);
and U9498 (N_9498,N_8824,N_8772);
and U9499 (N_9499,N_8699,N_8686);
nand U9500 (N_9500,N_9472,N_9354);
xnor U9501 (N_9501,N_9140,N_9183);
xor U9502 (N_9502,N_9407,N_9361);
xnor U9503 (N_9503,N_9335,N_9185);
xnor U9504 (N_9504,N_9018,N_9269);
xnor U9505 (N_9505,N_9163,N_9282);
nor U9506 (N_9506,N_9108,N_9436);
xor U9507 (N_9507,N_9062,N_9315);
and U9508 (N_9508,N_9481,N_9423);
nand U9509 (N_9509,N_9458,N_9128);
nor U9510 (N_9510,N_9428,N_9124);
xor U9511 (N_9511,N_9205,N_9162);
and U9512 (N_9512,N_9337,N_9118);
and U9513 (N_9513,N_9331,N_9422);
and U9514 (N_9514,N_9122,N_9478);
or U9515 (N_9515,N_9115,N_9365);
or U9516 (N_9516,N_9297,N_9158);
nor U9517 (N_9517,N_9306,N_9184);
or U9518 (N_9518,N_9217,N_9203);
nand U9519 (N_9519,N_9208,N_9479);
nand U9520 (N_9520,N_9041,N_9287);
or U9521 (N_9521,N_9311,N_9492);
xnor U9522 (N_9522,N_9491,N_9357);
and U9523 (N_9523,N_9447,N_9055);
or U9524 (N_9524,N_9415,N_9264);
nand U9525 (N_9525,N_9267,N_9125);
or U9526 (N_9526,N_9091,N_9419);
nor U9527 (N_9527,N_9343,N_9072);
and U9528 (N_9528,N_9196,N_9249);
nand U9529 (N_9529,N_9393,N_9098);
nand U9530 (N_9530,N_9236,N_9172);
or U9531 (N_9531,N_9084,N_9291);
or U9532 (N_9532,N_9056,N_9440);
nor U9533 (N_9533,N_9023,N_9453);
nand U9534 (N_9534,N_9401,N_9188);
or U9535 (N_9535,N_9304,N_9350);
nor U9536 (N_9536,N_9252,N_9151);
xor U9537 (N_9537,N_9160,N_9024);
nand U9538 (N_9538,N_9459,N_9089);
xor U9539 (N_9539,N_9338,N_9054);
or U9540 (N_9540,N_9347,N_9079);
and U9541 (N_9541,N_9011,N_9190);
and U9542 (N_9542,N_9004,N_9366);
nand U9543 (N_9543,N_9460,N_9199);
or U9544 (N_9544,N_9068,N_9212);
nor U9545 (N_9545,N_9139,N_9327);
xnor U9546 (N_9546,N_9058,N_9138);
or U9547 (N_9547,N_9180,N_9229);
and U9548 (N_9548,N_9421,N_9144);
nand U9549 (N_9549,N_9495,N_9257);
xor U9550 (N_9550,N_9164,N_9157);
nand U9551 (N_9551,N_9120,N_9074);
and U9552 (N_9552,N_9279,N_9238);
and U9553 (N_9553,N_9080,N_9483);
nor U9554 (N_9554,N_9107,N_9227);
nor U9555 (N_9555,N_9454,N_9109);
nand U9556 (N_9556,N_9466,N_9182);
and U9557 (N_9557,N_9087,N_9211);
nand U9558 (N_9558,N_9461,N_9441);
and U9559 (N_9559,N_9251,N_9165);
xnor U9560 (N_9560,N_9284,N_9016);
and U9561 (N_9561,N_9134,N_9475);
nand U9562 (N_9562,N_9009,N_9137);
xnor U9563 (N_9563,N_9187,N_9029);
and U9564 (N_9564,N_9406,N_9194);
xor U9565 (N_9565,N_9235,N_9006);
or U9566 (N_9566,N_9470,N_9399);
nand U9567 (N_9567,N_9223,N_9039);
nand U9568 (N_9568,N_9070,N_9376);
or U9569 (N_9569,N_9310,N_9169);
and U9570 (N_9570,N_9324,N_9156);
nand U9571 (N_9571,N_9312,N_9012);
xnor U9572 (N_9572,N_9330,N_9100);
nor U9573 (N_9573,N_9232,N_9026);
nor U9574 (N_9574,N_9474,N_9341);
nand U9575 (N_9575,N_9209,N_9290);
and U9576 (N_9576,N_9382,N_9416);
nor U9577 (N_9577,N_9445,N_9123);
xor U9578 (N_9578,N_9020,N_9285);
xor U9579 (N_9579,N_9061,N_9408);
xor U9580 (N_9580,N_9277,N_9028);
or U9581 (N_9581,N_9412,N_9239);
xor U9582 (N_9582,N_9225,N_9276);
or U9583 (N_9583,N_9069,N_9051);
and U9584 (N_9584,N_9387,N_9222);
or U9585 (N_9585,N_9414,N_9334);
nand U9586 (N_9586,N_9336,N_9093);
and U9587 (N_9587,N_9030,N_9083);
or U9588 (N_9588,N_9342,N_9218);
nand U9589 (N_9589,N_9048,N_9221);
nand U9590 (N_9590,N_9186,N_9497);
xnor U9591 (N_9591,N_9281,N_9404);
nor U9592 (N_9592,N_9106,N_9463);
nand U9593 (N_9593,N_9457,N_9411);
nor U9594 (N_9594,N_9246,N_9219);
nand U9595 (N_9595,N_9313,N_9424);
nand U9596 (N_9596,N_9325,N_9273);
and U9597 (N_9597,N_9166,N_9136);
nor U9598 (N_9598,N_9121,N_9110);
nor U9599 (N_9599,N_9161,N_9326);
or U9600 (N_9600,N_9231,N_9202);
or U9601 (N_9601,N_9052,N_9170);
or U9602 (N_9602,N_9234,N_9059);
nand U9603 (N_9603,N_9145,N_9237);
or U9604 (N_9604,N_9038,N_9473);
nor U9605 (N_9605,N_9374,N_9254);
nand U9606 (N_9606,N_9022,N_9034);
or U9607 (N_9607,N_9097,N_9067);
nand U9608 (N_9608,N_9035,N_9405);
xnor U9609 (N_9609,N_9258,N_9216);
xor U9610 (N_9610,N_9308,N_9198);
nor U9611 (N_9611,N_9245,N_9292);
xor U9612 (N_9612,N_9081,N_9450);
nand U9613 (N_9613,N_9005,N_9270);
nand U9614 (N_9614,N_9451,N_9490);
xor U9615 (N_9615,N_9485,N_9425);
nor U9616 (N_9616,N_9014,N_9213);
xnor U9617 (N_9617,N_9323,N_9309);
nand U9618 (N_9618,N_9439,N_9119);
xor U9619 (N_9619,N_9426,N_9349);
or U9620 (N_9620,N_9402,N_9126);
nor U9621 (N_9621,N_9046,N_9367);
and U9622 (N_9622,N_9266,N_9105);
nand U9623 (N_9623,N_9111,N_9021);
and U9624 (N_9624,N_9220,N_9319);
and U9625 (N_9625,N_9400,N_9263);
xnor U9626 (N_9626,N_9103,N_9380);
and U9627 (N_9627,N_9177,N_9200);
xnor U9628 (N_9628,N_9036,N_9362);
nor U9629 (N_9629,N_9274,N_9044);
nand U9630 (N_9630,N_9131,N_9075);
nand U9631 (N_9631,N_9228,N_9013);
xnor U9632 (N_9632,N_9372,N_9389);
and U9633 (N_9633,N_9314,N_9339);
or U9634 (N_9634,N_9379,N_9168);
nor U9635 (N_9635,N_9000,N_9477);
and U9636 (N_9636,N_9493,N_9003);
or U9637 (N_9637,N_9214,N_9037);
xnor U9638 (N_9638,N_9390,N_9435);
xnor U9639 (N_9639,N_9275,N_9296);
and U9640 (N_9640,N_9049,N_9242);
nor U9641 (N_9641,N_9096,N_9010);
or U9642 (N_9642,N_9375,N_9063);
xnor U9643 (N_9643,N_9329,N_9053);
or U9644 (N_9644,N_9300,N_9019);
and U9645 (N_9645,N_9127,N_9189);
or U9646 (N_9646,N_9363,N_9398);
xor U9647 (N_9647,N_9429,N_9193);
nand U9648 (N_9648,N_9159,N_9448);
xor U9649 (N_9649,N_9360,N_9344);
nand U9650 (N_9650,N_9465,N_9065);
or U9651 (N_9651,N_9496,N_9386);
xor U9652 (N_9652,N_9057,N_9153);
or U9653 (N_9653,N_9307,N_9204);
or U9654 (N_9654,N_9371,N_9452);
nand U9655 (N_9655,N_9455,N_9112);
nand U9656 (N_9656,N_9295,N_9333);
nand U9657 (N_9657,N_9432,N_9077);
and U9658 (N_9658,N_9101,N_9095);
or U9659 (N_9659,N_9265,N_9409);
or U9660 (N_9660,N_9345,N_9176);
or U9661 (N_9661,N_9207,N_9262);
nand U9662 (N_9662,N_9352,N_9288);
and U9663 (N_9663,N_9253,N_9280);
xor U9664 (N_9664,N_9073,N_9002);
or U9665 (N_9665,N_9394,N_9179);
or U9666 (N_9666,N_9033,N_9464);
and U9667 (N_9667,N_9129,N_9142);
nand U9668 (N_9668,N_9130,N_9484);
and U9669 (N_9669,N_9316,N_9351);
xnor U9670 (N_9670,N_9149,N_9171);
nor U9671 (N_9671,N_9355,N_9418);
nor U9672 (N_9672,N_9260,N_9403);
and U9673 (N_9673,N_9240,N_9480);
nand U9674 (N_9674,N_9317,N_9173);
nor U9675 (N_9675,N_9494,N_9303);
nand U9676 (N_9676,N_9498,N_9410);
nand U9677 (N_9677,N_9045,N_9085);
nand U9678 (N_9678,N_9241,N_9174);
or U9679 (N_9679,N_9431,N_9082);
nand U9680 (N_9680,N_9175,N_9353);
and U9681 (N_9681,N_9146,N_9047);
nor U9682 (N_9682,N_9417,N_9181);
or U9683 (N_9683,N_9104,N_9446);
nand U9684 (N_9684,N_9116,N_9373);
and U9685 (N_9685,N_9286,N_9150);
or U9686 (N_9686,N_9434,N_9391);
xnor U9687 (N_9687,N_9243,N_9283);
or U9688 (N_9688,N_9442,N_9340);
nor U9689 (N_9689,N_9356,N_9358);
nand U9690 (N_9690,N_9261,N_9301);
and U9691 (N_9691,N_9449,N_9396);
xnor U9692 (N_9692,N_9259,N_9268);
or U9693 (N_9693,N_9064,N_9433);
and U9694 (N_9694,N_9167,N_9178);
xnor U9695 (N_9695,N_9395,N_9226);
and U9696 (N_9696,N_9094,N_9247);
nor U9697 (N_9697,N_9364,N_9192);
and U9698 (N_9698,N_9377,N_9348);
or U9699 (N_9699,N_9388,N_9430);
or U9700 (N_9700,N_9215,N_9099);
or U9701 (N_9701,N_9076,N_9031);
xor U9702 (N_9702,N_9294,N_9032);
xnor U9703 (N_9703,N_9201,N_9488);
nand U9704 (N_9704,N_9328,N_9420);
and U9705 (N_9705,N_9233,N_9332);
and U9706 (N_9706,N_9487,N_9385);
and U9707 (N_9707,N_9413,N_9381);
or U9708 (N_9708,N_9092,N_9113);
or U9709 (N_9709,N_9248,N_9117);
or U9710 (N_9710,N_9133,N_9397);
and U9711 (N_9711,N_9469,N_9499);
nand U9712 (N_9712,N_9148,N_9255);
or U9713 (N_9713,N_9132,N_9078);
nand U9714 (N_9714,N_9467,N_9147);
nor U9715 (N_9715,N_9086,N_9210);
or U9716 (N_9716,N_9256,N_9486);
xnor U9717 (N_9717,N_9152,N_9154);
nor U9718 (N_9718,N_9289,N_9001);
xor U9719 (N_9719,N_9071,N_9456);
nor U9720 (N_9720,N_9191,N_9244);
and U9721 (N_9721,N_9427,N_9368);
and U9722 (N_9722,N_9050,N_9299);
nand U9723 (N_9723,N_9155,N_9066);
and U9724 (N_9724,N_9017,N_9250);
nor U9725 (N_9725,N_9383,N_9322);
or U9726 (N_9726,N_9040,N_9043);
nor U9727 (N_9727,N_9090,N_9025);
or U9728 (N_9728,N_9271,N_9359);
nand U9729 (N_9729,N_9489,N_9114);
nor U9730 (N_9730,N_9278,N_9008);
and U9731 (N_9731,N_9007,N_9320);
xor U9732 (N_9732,N_9370,N_9443);
nand U9733 (N_9733,N_9088,N_9369);
xnor U9734 (N_9734,N_9471,N_9135);
nand U9735 (N_9735,N_9392,N_9141);
xnor U9736 (N_9736,N_9224,N_9384);
nand U9737 (N_9737,N_9378,N_9143);
xnor U9738 (N_9738,N_9197,N_9318);
or U9739 (N_9739,N_9042,N_9195);
and U9740 (N_9740,N_9437,N_9102);
or U9741 (N_9741,N_9305,N_9302);
and U9742 (N_9742,N_9027,N_9298);
nor U9743 (N_9743,N_9015,N_9230);
nor U9744 (N_9744,N_9272,N_9462);
or U9745 (N_9745,N_9444,N_9476);
or U9746 (N_9746,N_9468,N_9482);
nand U9747 (N_9747,N_9321,N_9346);
nor U9748 (N_9748,N_9293,N_9206);
nor U9749 (N_9749,N_9438,N_9060);
nand U9750 (N_9750,N_9126,N_9305);
or U9751 (N_9751,N_9399,N_9398);
xnor U9752 (N_9752,N_9095,N_9302);
and U9753 (N_9753,N_9082,N_9492);
nor U9754 (N_9754,N_9186,N_9160);
nor U9755 (N_9755,N_9230,N_9308);
and U9756 (N_9756,N_9157,N_9317);
and U9757 (N_9757,N_9258,N_9205);
nor U9758 (N_9758,N_9402,N_9207);
nand U9759 (N_9759,N_9433,N_9283);
nand U9760 (N_9760,N_9111,N_9053);
and U9761 (N_9761,N_9485,N_9052);
xor U9762 (N_9762,N_9212,N_9190);
and U9763 (N_9763,N_9343,N_9227);
and U9764 (N_9764,N_9266,N_9447);
and U9765 (N_9765,N_9249,N_9442);
nand U9766 (N_9766,N_9166,N_9098);
nand U9767 (N_9767,N_9449,N_9045);
or U9768 (N_9768,N_9283,N_9203);
or U9769 (N_9769,N_9054,N_9052);
or U9770 (N_9770,N_9042,N_9046);
nor U9771 (N_9771,N_9077,N_9208);
or U9772 (N_9772,N_9395,N_9422);
or U9773 (N_9773,N_9191,N_9219);
nor U9774 (N_9774,N_9373,N_9263);
and U9775 (N_9775,N_9171,N_9320);
xnor U9776 (N_9776,N_9310,N_9225);
or U9777 (N_9777,N_9181,N_9088);
or U9778 (N_9778,N_9151,N_9306);
nor U9779 (N_9779,N_9262,N_9368);
nor U9780 (N_9780,N_9272,N_9407);
xnor U9781 (N_9781,N_9325,N_9164);
and U9782 (N_9782,N_9272,N_9032);
nor U9783 (N_9783,N_9493,N_9296);
and U9784 (N_9784,N_9042,N_9376);
and U9785 (N_9785,N_9491,N_9184);
nand U9786 (N_9786,N_9476,N_9379);
or U9787 (N_9787,N_9229,N_9070);
or U9788 (N_9788,N_9334,N_9061);
or U9789 (N_9789,N_9493,N_9103);
nand U9790 (N_9790,N_9327,N_9071);
and U9791 (N_9791,N_9309,N_9199);
or U9792 (N_9792,N_9109,N_9363);
nor U9793 (N_9793,N_9149,N_9331);
nor U9794 (N_9794,N_9299,N_9021);
nor U9795 (N_9795,N_9083,N_9368);
and U9796 (N_9796,N_9424,N_9194);
nand U9797 (N_9797,N_9480,N_9076);
xor U9798 (N_9798,N_9090,N_9265);
xnor U9799 (N_9799,N_9014,N_9269);
xor U9800 (N_9800,N_9045,N_9261);
nor U9801 (N_9801,N_9041,N_9263);
xnor U9802 (N_9802,N_9255,N_9418);
and U9803 (N_9803,N_9234,N_9490);
nand U9804 (N_9804,N_9142,N_9271);
or U9805 (N_9805,N_9388,N_9203);
or U9806 (N_9806,N_9364,N_9022);
or U9807 (N_9807,N_9087,N_9489);
and U9808 (N_9808,N_9438,N_9471);
and U9809 (N_9809,N_9435,N_9363);
and U9810 (N_9810,N_9285,N_9327);
nand U9811 (N_9811,N_9087,N_9377);
or U9812 (N_9812,N_9331,N_9275);
xnor U9813 (N_9813,N_9187,N_9201);
xor U9814 (N_9814,N_9085,N_9103);
or U9815 (N_9815,N_9251,N_9499);
xor U9816 (N_9816,N_9011,N_9081);
and U9817 (N_9817,N_9006,N_9114);
xor U9818 (N_9818,N_9136,N_9005);
xnor U9819 (N_9819,N_9477,N_9308);
and U9820 (N_9820,N_9014,N_9152);
nand U9821 (N_9821,N_9032,N_9249);
nand U9822 (N_9822,N_9415,N_9178);
nor U9823 (N_9823,N_9477,N_9492);
xnor U9824 (N_9824,N_9111,N_9499);
xor U9825 (N_9825,N_9403,N_9096);
xnor U9826 (N_9826,N_9032,N_9022);
and U9827 (N_9827,N_9079,N_9145);
xor U9828 (N_9828,N_9394,N_9312);
xor U9829 (N_9829,N_9372,N_9126);
nand U9830 (N_9830,N_9100,N_9068);
or U9831 (N_9831,N_9492,N_9042);
or U9832 (N_9832,N_9466,N_9443);
nand U9833 (N_9833,N_9188,N_9005);
and U9834 (N_9834,N_9129,N_9423);
xnor U9835 (N_9835,N_9286,N_9330);
nor U9836 (N_9836,N_9032,N_9111);
and U9837 (N_9837,N_9142,N_9401);
and U9838 (N_9838,N_9290,N_9475);
and U9839 (N_9839,N_9240,N_9098);
xnor U9840 (N_9840,N_9041,N_9144);
nor U9841 (N_9841,N_9363,N_9336);
nor U9842 (N_9842,N_9006,N_9381);
or U9843 (N_9843,N_9270,N_9011);
xnor U9844 (N_9844,N_9024,N_9293);
or U9845 (N_9845,N_9367,N_9126);
nor U9846 (N_9846,N_9267,N_9132);
or U9847 (N_9847,N_9488,N_9292);
and U9848 (N_9848,N_9344,N_9182);
xor U9849 (N_9849,N_9437,N_9237);
xnor U9850 (N_9850,N_9047,N_9448);
xnor U9851 (N_9851,N_9339,N_9183);
and U9852 (N_9852,N_9336,N_9276);
nand U9853 (N_9853,N_9041,N_9457);
nand U9854 (N_9854,N_9060,N_9018);
or U9855 (N_9855,N_9496,N_9134);
nand U9856 (N_9856,N_9259,N_9234);
xnor U9857 (N_9857,N_9278,N_9305);
nand U9858 (N_9858,N_9137,N_9120);
and U9859 (N_9859,N_9437,N_9188);
nand U9860 (N_9860,N_9052,N_9432);
nor U9861 (N_9861,N_9094,N_9290);
xnor U9862 (N_9862,N_9086,N_9091);
and U9863 (N_9863,N_9345,N_9210);
and U9864 (N_9864,N_9243,N_9435);
nor U9865 (N_9865,N_9300,N_9198);
nor U9866 (N_9866,N_9114,N_9026);
or U9867 (N_9867,N_9404,N_9164);
or U9868 (N_9868,N_9249,N_9014);
nor U9869 (N_9869,N_9401,N_9208);
nand U9870 (N_9870,N_9376,N_9445);
or U9871 (N_9871,N_9176,N_9186);
and U9872 (N_9872,N_9490,N_9001);
xor U9873 (N_9873,N_9465,N_9194);
and U9874 (N_9874,N_9190,N_9299);
nand U9875 (N_9875,N_9233,N_9367);
or U9876 (N_9876,N_9266,N_9421);
nor U9877 (N_9877,N_9370,N_9315);
xnor U9878 (N_9878,N_9180,N_9491);
or U9879 (N_9879,N_9328,N_9194);
and U9880 (N_9880,N_9163,N_9269);
or U9881 (N_9881,N_9114,N_9337);
xor U9882 (N_9882,N_9406,N_9297);
nor U9883 (N_9883,N_9145,N_9117);
or U9884 (N_9884,N_9300,N_9183);
and U9885 (N_9885,N_9166,N_9388);
or U9886 (N_9886,N_9224,N_9342);
nand U9887 (N_9887,N_9100,N_9026);
or U9888 (N_9888,N_9489,N_9486);
xor U9889 (N_9889,N_9368,N_9389);
and U9890 (N_9890,N_9339,N_9373);
and U9891 (N_9891,N_9179,N_9429);
nor U9892 (N_9892,N_9184,N_9136);
or U9893 (N_9893,N_9448,N_9328);
or U9894 (N_9894,N_9360,N_9402);
nor U9895 (N_9895,N_9055,N_9228);
xnor U9896 (N_9896,N_9240,N_9278);
and U9897 (N_9897,N_9131,N_9300);
nor U9898 (N_9898,N_9445,N_9213);
or U9899 (N_9899,N_9301,N_9472);
xnor U9900 (N_9900,N_9182,N_9009);
and U9901 (N_9901,N_9062,N_9308);
nand U9902 (N_9902,N_9334,N_9289);
nor U9903 (N_9903,N_9135,N_9305);
or U9904 (N_9904,N_9310,N_9453);
and U9905 (N_9905,N_9001,N_9333);
or U9906 (N_9906,N_9314,N_9289);
and U9907 (N_9907,N_9147,N_9476);
nand U9908 (N_9908,N_9442,N_9418);
nand U9909 (N_9909,N_9168,N_9267);
xnor U9910 (N_9910,N_9109,N_9239);
and U9911 (N_9911,N_9151,N_9115);
and U9912 (N_9912,N_9462,N_9136);
and U9913 (N_9913,N_9008,N_9193);
and U9914 (N_9914,N_9463,N_9229);
nor U9915 (N_9915,N_9272,N_9244);
or U9916 (N_9916,N_9390,N_9303);
xnor U9917 (N_9917,N_9277,N_9266);
nor U9918 (N_9918,N_9229,N_9414);
nor U9919 (N_9919,N_9065,N_9143);
nand U9920 (N_9920,N_9104,N_9139);
xor U9921 (N_9921,N_9314,N_9198);
xnor U9922 (N_9922,N_9210,N_9336);
nor U9923 (N_9923,N_9441,N_9155);
nand U9924 (N_9924,N_9132,N_9273);
xor U9925 (N_9925,N_9058,N_9086);
nor U9926 (N_9926,N_9311,N_9370);
or U9927 (N_9927,N_9355,N_9459);
nor U9928 (N_9928,N_9168,N_9061);
or U9929 (N_9929,N_9233,N_9006);
nand U9930 (N_9930,N_9397,N_9059);
nor U9931 (N_9931,N_9271,N_9235);
or U9932 (N_9932,N_9354,N_9416);
or U9933 (N_9933,N_9403,N_9064);
and U9934 (N_9934,N_9444,N_9019);
or U9935 (N_9935,N_9251,N_9034);
xnor U9936 (N_9936,N_9308,N_9073);
nor U9937 (N_9937,N_9057,N_9469);
nand U9938 (N_9938,N_9159,N_9105);
nand U9939 (N_9939,N_9353,N_9452);
or U9940 (N_9940,N_9058,N_9440);
nor U9941 (N_9941,N_9025,N_9220);
or U9942 (N_9942,N_9351,N_9289);
xnor U9943 (N_9943,N_9094,N_9019);
nand U9944 (N_9944,N_9168,N_9396);
or U9945 (N_9945,N_9146,N_9019);
nand U9946 (N_9946,N_9202,N_9335);
xnor U9947 (N_9947,N_9231,N_9263);
nor U9948 (N_9948,N_9172,N_9178);
xnor U9949 (N_9949,N_9045,N_9330);
xnor U9950 (N_9950,N_9485,N_9165);
or U9951 (N_9951,N_9172,N_9125);
and U9952 (N_9952,N_9059,N_9187);
or U9953 (N_9953,N_9491,N_9452);
xor U9954 (N_9954,N_9113,N_9214);
nand U9955 (N_9955,N_9351,N_9056);
xor U9956 (N_9956,N_9241,N_9086);
and U9957 (N_9957,N_9418,N_9317);
nor U9958 (N_9958,N_9423,N_9240);
nand U9959 (N_9959,N_9461,N_9380);
or U9960 (N_9960,N_9080,N_9355);
nand U9961 (N_9961,N_9460,N_9261);
or U9962 (N_9962,N_9098,N_9193);
xor U9963 (N_9963,N_9070,N_9402);
xnor U9964 (N_9964,N_9011,N_9198);
nand U9965 (N_9965,N_9251,N_9493);
xnor U9966 (N_9966,N_9479,N_9294);
and U9967 (N_9967,N_9169,N_9290);
and U9968 (N_9968,N_9251,N_9355);
or U9969 (N_9969,N_9235,N_9224);
and U9970 (N_9970,N_9396,N_9375);
or U9971 (N_9971,N_9118,N_9479);
nor U9972 (N_9972,N_9261,N_9305);
or U9973 (N_9973,N_9462,N_9268);
xor U9974 (N_9974,N_9043,N_9011);
nor U9975 (N_9975,N_9179,N_9280);
and U9976 (N_9976,N_9146,N_9052);
nor U9977 (N_9977,N_9492,N_9257);
nand U9978 (N_9978,N_9133,N_9130);
xor U9979 (N_9979,N_9325,N_9490);
and U9980 (N_9980,N_9018,N_9354);
or U9981 (N_9981,N_9499,N_9358);
or U9982 (N_9982,N_9027,N_9316);
xnor U9983 (N_9983,N_9306,N_9371);
nor U9984 (N_9984,N_9384,N_9470);
and U9985 (N_9985,N_9009,N_9387);
nand U9986 (N_9986,N_9490,N_9294);
nand U9987 (N_9987,N_9384,N_9014);
or U9988 (N_9988,N_9254,N_9152);
and U9989 (N_9989,N_9278,N_9033);
nand U9990 (N_9990,N_9207,N_9355);
nand U9991 (N_9991,N_9407,N_9493);
nand U9992 (N_9992,N_9121,N_9294);
nor U9993 (N_9993,N_9298,N_9163);
nor U9994 (N_9994,N_9283,N_9489);
or U9995 (N_9995,N_9285,N_9239);
nand U9996 (N_9996,N_9105,N_9033);
or U9997 (N_9997,N_9208,N_9187);
and U9998 (N_9998,N_9093,N_9394);
nand U9999 (N_9999,N_9139,N_9179);
nor U10000 (N_10000,N_9681,N_9834);
nand U10001 (N_10001,N_9801,N_9537);
xnor U10002 (N_10002,N_9778,N_9968);
and U10003 (N_10003,N_9880,N_9536);
or U10004 (N_10004,N_9823,N_9898);
nor U10005 (N_10005,N_9572,N_9566);
nor U10006 (N_10006,N_9752,N_9630);
nand U10007 (N_10007,N_9580,N_9985);
and U10008 (N_10008,N_9816,N_9557);
or U10009 (N_10009,N_9613,N_9797);
nor U10010 (N_10010,N_9606,N_9984);
nand U10011 (N_10011,N_9550,N_9881);
and U10012 (N_10012,N_9977,N_9709);
xnor U10013 (N_10013,N_9730,N_9517);
nor U10014 (N_10014,N_9887,N_9590);
xnor U10015 (N_10015,N_9689,N_9657);
or U10016 (N_10016,N_9745,N_9819);
xnor U10017 (N_10017,N_9850,N_9784);
or U10018 (N_10018,N_9629,N_9561);
or U10019 (N_10019,N_9610,N_9775);
nor U10020 (N_10020,N_9812,N_9978);
or U10021 (N_10021,N_9736,N_9967);
nor U10022 (N_10022,N_9651,N_9997);
nor U10023 (N_10023,N_9665,N_9937);
or U10024 (N_10024,N_9548,N_9739);
nand U10025 (N_10025,N_9760,N_9858);
and U10026 (N_10026,N_9905,N_9699);
xor U10027 (N_10027,N_9746,N_9735);
nand U10028 (N_10028,N_9722,N_9632);
or U10029 (N_10029,N_9565,N_9799);
nand U10030 (N_10030,N_9608,N_9941);
and U10031 (N_10031,N_9779,N_9747);
nor U10032 (N_10032,N_9900,N_9913);
xnor U10033 (N_10033,N_9914,N_9811);
nand U10034 (N_10034,N_9586,N_9936);
xnor U10035 (N_10035,N_9790,N_9966);
xor U10036 (N_10036,N_9999,N_9687);
and U10037 (N_10037,N_9970,N_9923);
nor U10038 (N_10038,N_9636,N_9675);
nor U10039 (N_10039,N_9964,N_9943);
nor U10040 (N_10040,N_9912,N_9695);
xor U10041 (N_10041,N_9756,N_9932);
or U10042 (N_10042,N_9893,N_9869);
xnor U10043 (N_10043,N_9983,N_9719);
or U10044 (N_10044,N_9568,N_9539);
nand U10045 (N_10045,N_9653,N_9728);
nand U10046 (N_10046,N_9680,N_9960);
or U10047 (N_10047,N_9770,N_9963);
nor U10048 (N_10048,N_9826,N_9975);
nor U10049 (N_10049,N_9830,N_9721);
or U10050 (N_10050,N_9712,N_9979);
or U10051 (N_10051,N_9875,N_9810);
and U10052 (N_10052,N_9922,N_9871);
and U10053 (N_10053,N_9600,N_9659);
nor U10054 (N_10054,N_9969,N_9777);
nor U10055 (N_10055,N_9592,N_9530);
nand U10056 (N_10056,N_9639,N_9944);
nor U10057 (N_10057,N_9835,N_9940);
xor U10058 (N_10058,N_9621,N_9718);
or U10059 (N_10059,N_9611,N_9771);
xor U10060 (N_10060,N_9702,N_9883);
or U10061 (N_10061,N_9895,N_9618);
nand U10062 (N_10062,N_9872,N_9848);
nor U10063 (N_10063,N_9583,N_9748);
xor U10064 (N_10064,N_9844,N_9828);
and U10065 (N_10065,N_9879,N_9800);
nand U10066 (N_10066,N_9540,N_9825);
nor U10067 (N_10067,N_9522,N_9786);
xor U10068 (N_10068,N_9925,N_9740);
xor U10069 (N_10069,N_9824,N_9598);
or U10070 (N_10070,N_9504,N_9501);
nor U10071 (N_10071,N_9649,N_9711);
xnor U10072 (N_10072,N_9663,N_9954);
nor U10073 (N_10073,N_9605,N_9994);
nor U10074 (N_10074,N_9715,N_9688);
nor U10075 (N_10075,N_9671,N_9965);
or U10076 (N_10076,N_9862,N_9924);
nand U10077 (N_10077,N_9757,N_9725);
xor U10078 (N_10078,N_9918,N_9512);
nand U10079 (N_10079,N_9755,N_9807);
nor U10080 (N_10080,N_9677,N_9714);
nor U10081 (N_10081,N_9578,N_9956);
xor U10082 (N_10082,N_9597,N_9759);
or U10083 (N_10083,N_9669,N_9981);
or U10084 (N_10084,N_9909,N_9768);
or U10085 (N_10085,N_9603,N_9973);
nor U10086 (N_10086,N_9931,N_9792);
nor U10087 (N_10087,N_9762,N_9676);
nand U10088 (N_10088,N_9958,N_9554);
and U10089 (N_10089,N_9556,N_9518);
and U10090 (N_10090,N_9662,N_9926);
and U10091 (N_10091,N_9541,N_9713);
and U10092 (N_10092,N_9577,N_9827);
nor U10093 (N_10093,N_9789,N_9515);
xor U10094 (N_10094,N_9935,N_9587);
and U10095 (N_10095,N_9749,N_9591);
xnor U10096 (N_10096,N_9614,N_9953);
nand U10097 (N_10097,N_9776,N_9545);
or U10098 (N_10098,N_9737,N_9859);
or U10099 (N_10099,N_9694,N_9903);
nor U10100 (N_10100,N_9708,N_9511);
and U10101 (N_10101,N_9831,N_9683);
nand U10102 (N_10102,N_9576,N_9938);
nor U10103 (N_10103,N_9849,N_9724);
xor U10104 (N_10104,N_9729,N_9650);
nand U10105 (N_10105,N_9635,N_9891);
nor U10106 (N_10106,N_9503,N_9527);
and U10107 (N_10107,N_9641,N_9990);
xnor U10108 (N_10108,N_9804,N_9692);
xnor U10109 (N_10109,N_9531,N_9809);
or U10110 (N_10110,N_9581,N_9678);
xor U10111 (N_10111,N_9652,N_9854);
nand U10112 (N_10112,N_9877,N_9894);
nor U10113 (N_10113,N_9866,N_9627);
and U10114 (N_10114,N_9500,N_9582);
xor U10115 (N_10115,N_9674,N_9667);
xnor U10116 (N_10116,N_9682,N_9948);
or U10117 (N_10117,N_9817,N_9876);
nand U10118 (N_10118,N_9584,N_9589);
and U10119 (N_10119,N_9787,N_9904);
nand U10120 (N_10120,N_9951,N_9882);
xor U10121 (N_10121,N_9506,N_9813);
nor U10122 (N_10122,N_9716,N_9705);
nor U10123 (N_10123,N_9933,N_9796);
xor U10124 (N_10124,N_9622,N_9783);
and U10125 (N_10125,N_9696,N_9782);
or U10126 (N_10126,N_9625,N_9982);
nor U10127 (N_10127,N_9899,N_9788);
nand U10128 (N_10128,N_9562,N_9832);
nand U10129 (N_10129,N_9766,N_9575);
xnor U10130 (N_10130,N_9555,N_9971);
nor U10131 (N_10131,N_9806,N_9794);
and U10132 (N_10132,N_9889,N_9957);
and U10133 (N_10133,N_9602,N_9656);
nor U10134 (N_10134,N_9642,N_9845);
xor U10135 (N_10135,N_9732,N_9731);
nand U10136 (N_10136,N_9528,N_9570);
or U10137 (N_10137,N_9523,N_9774);
xor U10138 (N_10138,N_9726,N_9685);
nand U10139 (N_10139,N_9679,N_9623);
nand U10140 (N_10140,N_9761,N_9911);
nor U10141 (N_10141,N_9664,N_9612);
or U10142 (N_10142,N_9772,N_9573);
xnor U10143 (N_10143,N_9640,N_9851);
nor U10144 (N_10144,N_9703,N_9673);
and U10145 (N_10145,N_9995,N_9805);
and U10146 (N_10146,N_9626,N_9553);
nor U10147 (N_10147,N_9560,N_9508);
or U10148 (N_10148,N_9836,N_9874);
xor U10149 (N_10149,N_9633,N_9993);
or U10150 (N_10150,N_9947,N_9764);
nor U10151 (N_10151,N_9628,N_9765);
nand U10152 (N_10152,N_9526,N_9961);
or U10153 (N_10153,N_9617,N_9750);
or U10154 (N_10154,N_9559,N_9886);
and U10155 (N_10155,N_9547,N_9535);
nor U10156 (N_10156,N_9707,N_9596);
nand U10157 (N_10157,N_9896,N_9795);
xor U10158 (N_10158,N_9833,N_9873);
and U10159 (N_10159,N_9704,N_9502);
or U10160 (N_10160,N_9793,N_9920);
xnor U10161 (N_10161,N_9509,N_9595);
or U10162 (N_10162,N_9564,N_9906);
xor U10163 (N_10163,N_9910,N_9571);
nand U10164 (N_10164,N_9525,N_9668);
nor U10165 (N_10165,N_9723,N_9563);
nand U10166 (N_10166,N_9945,N_9615);
or U10167 (N_10167,N_9654,N_9686);
xor U10168 (N_10168,N_9690,N_9754);
nor U10169 (N_10169,N_9601,N_9646);
xor U10170 (N_10170,N_9520,N_9700);
or U10171 (N_10171,N_9986,N_9638);
nand U10172 (N_10172,N_9829,N_9791);
nor U10173 (N_10173,N_9885,N_9802);
nand U10174 (N_10174,N_9594,N_9767);
and U10175 (N_10175,N_9842,N_9857);
or U10176 (N_10176,N_9631,N_9989);
xor U10177 (N_10177,N_9542,N_9852);
and U10178 (N_10178,N_9820,N_9660);
nor U10179 (N_10179,N_9734,N_9930);
or U10180 (N_10180,N_9785,N_9666);
or U10181 (N_10181,N_9670,N_9655);
or U10182 (N_10182,N_9908,N_9843);
and U10183 (N_10183,N_9697,N_9552);
nor U10184 (N_10184,N_9607,N_9534);
xnor U10185 (N_10185,N_9822,N_9996);
xnor U10186 (N_10186,N_9706,N_9864);
and U10187 (N_10187,N_9658,N_9741);
or U10188 (N_10188,N_9865,N_9928);
or U10189 (N_10189,N_9916,N_9616);
xor U10190 (N_10190,N_9609,N_9878);
xnor U10191 (N_10191,N_9643,N_9840);
or U10192 (N_10192,N_9962,N_9888);
xnor U10193 (N_10193,N_9604,N_9645);
nor U10194 (N_10194,N_9856,N_9516);
and U10195 (N_10195,N_9543,N_9942);
xor U10196 (N_10196,N_9815,N_9972);
xnor U10197 (N_10197,N_9620,N_9934);
nor U10198 (N_10198,N_9949,N_9853);
or U10199 (N_10199,N_9892,N_9647);
nor U10200 (N_10200,N_9567,N_9959);
xnor U10201 (N_10201,N_9599,N_9780);
xnor U10202 (N_10202,N_9952,N_9546);
nor U10203 (N_10203,N_9579,N_9974);
and U10204 (N_10204,N_9644,N_9855);
nor U10205 (N_10205,N_9698,N_9870);
nand U10206 (N_10206,N_9538,N_9763);
xor U10207 (N_10207,N_9861,N_9738);
nor U10208 (N_10208,N_9846,N_9585);
and U10209 (N_10209,N_9505,N_9569);
and U10210 (N_10210,N_9991,N_9514);
nor U10211 (N_10211,N_9648,N_9742);
or U10212 (N_10212,N_9841,N_9867);
nand U10213 (N_10213,N_9574,N_9838);
nand U10214 (N_10214,N_9532,N_9558);
nand U10215 (N_10215,N_9691,N_9684);
nand U10216 (N_10216,N_9847,N_9510);
nand U10217 (N_10217,N_9549,N_9744);
nor U10218 (N_10218,N_9929,N_9693);
and U10219 (N_10219,N_9917,N_9727);
xnor U10220 (N_10220,N_9839,N_9837);
xor U10221 (N_10221,N_9907,N_9619);
and U10222 (N_10222,N_9818,N_9733);
and U10223 (N_10223,N_9533,N_9743);
nand U10224 (N_10224,N_9634,N_9998);
nand U10225 (N_10225,N_9890,N_9939);
nor U10226 (N_10226,N_9988,N_9927);
and U10227 (N_10227,N_9751,N_9521);
nor U10228 (N_10228,N_9593,N_9808);
nand U10229 (N_10229,N_9980,N_9717);
xnor U10230 (N_10230,N_9798,N_9915);
or U10231 (N_10231,N_9507,N_9519);
nor U10232 (N_10232,N_9637,N_9868);
xor U10233 (N_10233,N_9919,N_9987);
and U10234 (N_10234,N_9946,N_9624);
nor U10235 (N_10235,N_9544,N_9955);
xnor U10236 (N_10236,N_9551,N_9769);
nand U10237 (N_10237,N_9588,N_9803);
xor U10238 (N_10238,N_9950,N_9524);
xnor U10239 (N_10239,N_9921,N_9897);
nor U10240 (N_10240,N_9720,N_9902);
nand U10241 (N_10241,N_9758,N_9513);
nor U10242 (N_10242,N_9672,N_9821);
and U10243 (N_10243,N_9773,N_9884);
and U10244 (N_10244,N_9863,N_9992);
and U10245 (N_10245,N_9753,N_9781);
nand U10246 (N_10246,N_9860,N_9661);
xnor U10247 (N_10247,N_9976,N_9814);
and U10248 (N_10248,N_9701,N_9710);
or U10249 (N_10249,N_9529,N_9901);
and U10250 (N_10250,N_9619,N_9994);
or U10251 (N_10251,N_9733,N_9952);
and U10252 (N_10252,N_9755,N_9927);
nor U10253 (N_10253,N_9940,N_9503);
xor U10254 (N_10254,N_9715,N_9905);
nand U10255 (N_10255,N_9876,N_9843);
xor U10256 (N_10256,N_9982,N_9802);
or U10257 (N_10257,N_9823,N_9869);
and U10258 (N_10258,N_9624,N_9724);
nor U10259 (N_10259,N_9925,N_9708);
nand U10260 (N_10260,N_9535,N_9585);
nor U10261 (N_10261,N_9604,N_9606);
xor U10262 (N_10262,N_9752,N_9679);
or U10263 (N_10263,N_9718,N_9781);
nand U10264 (N_10264,N_9604,N_9924);
or U10265 (N_10265,N_9902,N_9528);
xor U10266 (N_10266,N_9503,N_9750);
and U10267 (N_10267,N_9644,N_9965);
nand U10268 (N_10268,N_9910,N_9631);
nor U10269 (N_10269,N_9786,N_9960);
nand U10270 (N_10270,N_9580,N_9715);
xnor U10271 (N_10271,N_9689,N_9515);
nor U10272 (N_10272,N_9702,N_9832);
or U10273 (N_10273,N_9845,N_9736);
and U10274 (N_10274,N_9693,N_9859);
nor U10275 (N_10275,N_9602,N_9565);
xor U10276 (N_10276,N_9793,N_9513);
nand U10277 (N_10277,N_9517,N_9962);
or U10278 (N_10278,N_9990,N_9589);
xor U10279 (N_10279,N_9724,N_9948);
xor U10280 (N_10280,N_9643,N_9705);
and U10281 (N_10281,N_9803,N_9686);
and U10282 (N_10282,N_9679,N_9902);
nor U10283 (N_10283,N_9830,N_9781);
nor U10284 (N_10284,N_9807,N_9922);
nor U10285 (N_10285,N_9640,N_9669);
or U10286 (N_10286,N_9953,N_9722);
nor U10287 (N_10287,N_9974,N_9955);
nand U10288 (N_10288,N_9982,N_9697);
nand U10289 (N_10289,N_9623,N_9601);
nor U10290 (N_10290,N_9910,N_9672);
nor U10291 (N_10291,N_9577,N_9712);
nand U10292 (N_10292,N_9807,N_9952);
xor U10293 (N_10293,N_9659,N_9806);
or U10294 (N_10294,N_9743,N_9549);
xnor U10295 (N_10295,N_9675,N_9825);
and U10296 (N_10296,N_9816,N_9616);
nor U10297 (N_10297,N_9844,N_9651);
nand U10298 (N_10298,N_9714,N_9957);
nand U10299 (N_10299,N_9913,N_9644);
nor U10300 (N_10300,N_9914,N_9595);
or U10301 (N_10301,N_9670,N_9755);
and U10302 (N_10302,N_9646,N_9719);
nand U10303 (N_10303,N_9772,N_9950);
nand U10304 (N_10304,N_9703,N_9686);
xor U10305 (N_10305,N_9731,N_9985);
and U10306 (N_10306,N_9758,N_9908);
and U10307 (N_10307,N_9665,N_9734);
or U10308 (N_10308,N_9956,N_9624);
nor U10309 (N_10309,N_9598,N_9989);
nor U10310 (N_10310,N_9908,N_9996);
nand U10311 (N_10311,N_9573,N_9614);
nand U10312 (N_10312,N_9551,N_9820);
or U10313 (N_10313,N_9547,N_9971);
nor U10314 (N_10314,N_9523,N_9527);
or U10315 (N_10315,N_9796,N_9770);
and U10316 (N_10316,N_9700,N_9697);
xnor U10317 (N_10317,N_9728,N_9720);
and U10318 (N_10318,N_9617,N_9964);
xnor U10319 (N_10319,N_9516,N_9653);
xor U10320 (N_10320,N_9601,N_9678);
nor U10321 (N_10321,N_9528,N_9685);
and U10322 (N_10322,N_9946,N_9880);
or U10323 (N_10323,N_9591,N_9594);
xnor U10324 (N_10324,N_9813,N_9673);
nand U10325 (N_10325,N_9915,N_9574);
xnor U10326 (N_10326,N_9656,N_9784);
nor U10327 (N_10327,N_9851,N_9639);
nor U10328 (N_10328,N_9536,N_9682);
nor U10329 (N_10329,N_9605,N_9988);
nand U10330 (N_10330,N_9981,N_9663);
and U10331 (N_10331,N_9701,N_9938);
xor U10332 (N_10332,N_9740,N_9526);
and U10333 (N_10333,N_9841,N_9585);
and U10334 (N_10334,N_9735,N_9933);
nor U10335 (N_10335,N_9926,N_9871);
or U10336 (N_10336,N_9971,N_9970);
and U10337 (N_10337,N_9551,N_9667);
xnor U10338 (N_10338,N_9500,N_9583);
nand U10339 (N_10339,N_9826,N_9981);
nand U10340 (N_10340,N_9586,N_9822);
nor U10341 (N_10341,N_9755,N_9548);
and U10342 (N_10342,N_9647,N_9705);
and U10343 (N_10343,N_9676,N_9736);
and U10344 (N_10344,N_9604,N_9667);
nor U10345 (N_10345,N_9676,N_9761);
nor U10346 (N_10346,N_9894,N_9566);
or U10347 (N_10347,N_9507,N_9783);
or U10348 (N_10348,N_9636,N_9663);
xnor U10349 (N_10349,N_9823,N_9640);
and U10350 (N_10350,N_9796,N_9552);
and U10351 (N_10351,N_9666,N_9826);
nor U10352 (N_10352,N_9717,N_9978);
and U10353 (N_10353,N_9829,N_9766);
nand U10354 (N_10354,N_9868,N_9804);
xor U10355 (N_10355,N_9816,N_9857);
nand U10356 (N_10356,N_9597,N_9571);
and U10357 (N_10357,N_9702,N_9849);
nand U10358 (N_10358,N_9960,N_9530);
nand U10359 (N_10359,N_9610,N_9914);
nand U10360 (N_10360,N_9521,N_9624);
or U10361 (N_10361,N_9990,N_9860);
xnor U10362 (N_10362,N_9551,N_9992);
xor U10363 (N_10363,N_9597,N_9732);
xor U10364 (N_10364,N_9929,N_9875);
and U10365 (N_10365,N_9723,N_9586);
nor U10366 (N_10366,N_9871,N_9894);
nor U10367 (N_10367,N_9518,N_9625);
and U10368 (N_10368,N_9977,N_9545);
xor U10369 (N_10369,N_9870,N_9543);
nor U10370 (N_10370,N_9951,N_9582);
and U10371 (N_10371,N_9956,N_9601);
nor U10372 (N_10372,N_9519,N_9644);
xnor U10373 (N_10373,N_9530,N_9928);
and U10374 (N_10374,N_9758,N_9723);
or U10375 (N_10375,N_9792,N_9759);
xor U10376 (N_10376,N_9793,N_9932);
nor U10377 (N_10377,N_9952,N_9746);
nand U10378 (N_10378,N_9501,N_9616);
and U10379 (N_10379,N_9557,N_9715);
nor U10380 (N_10380,N_9893,N_9664);
xnor U10381 (N_10381,N_9993,N_9674);
and U10382 (N_10382,N_9898,N_9524);
nor U10383 (N_10383,N_9902,N_9736);
xor U10384 (N_10384,N_9846,N_9734);
and U10385 (N_10385,N_9990,N_9861);
or U10386 (N_10386,N_9981,N_9681);
nand U10387 (N_10387,N_9765,N_9599);
nor U10388 (N_10388,N_9645,N_9989);
or U10389 (N_10389,N_9591,N_9590);
xnor U10390 (N_10390,N_9864,N_9645);
xor U10391 (N_10391,N_9871,N_9735);
or U10392 (N_10392,N_9951,N_9812);
or U10393 (N_10393,N_9897,N_9977);
nor U10394 (N_10394,N_9678,N_9862);
nand U10395 (N_10395,N_9641,N_9657);
nor U10396 (N_10396,N_9619,N_9978);
xnor U10397 (N_10397,N_9605,N_9970);
xnor U10398 (N_10398,N_9851,N_9895);
nand U10399 (N_10399,N_9607,N_9869);
xnor U10400 (N_10400,N_9964,N_9759);
xnor U10401 (N_10401,N_9892,N_9740);
or U10402 (N_10402,N_9860,N_9961);
or U10403 (N_10403,N_9781,N_9687);
nor U10404 (N_10404,N_9724,N_9601);
or U10405 (N_10405,N_9736,N_9662);
and U10406 (N_10406,N_9876,N_9607);
or U10407 (N_10407,N_9713,N_9837);
or U10408 (N_10408,N_9546,N_9593);
nor U10409 (N_10409,N_9800,N_9978);
nor U10410 (N_10410,N_9736,N_9846);
and U10411 (N_10411,N_9905,N_9798);
nand U10412 (N_10412,N_9607,N_9655);
or U10413 (N_10413,N_9994,N_9855);
or U10414 (N_10414,N_9824,N_9544);
xnor U10415 (N_10415,N_9838,N_9841);
xor U10416 (N_10416,N_9728,N_9673);
and U10417 (N_10417,N_9587,N_9657);
or U10418 (N_10418,N_9838,N_9804);
xor U10419 (N_10419,N_9611,N_9543);
and U10420 (N_10420,N_9573,N_9881);
or U10421 (N_10421,N_9978,N_9605);
nor U10422 (N_10422,N_9699,N_9912);
or U10423 (N_10423,N_9863,N_9712);
xnor U10424 (N_10424,N_9810,N_9860);
xnor U10425 (N_10425,N_9762,N_9669);
nand U10426 (N_10426,N_9650,N_9576);
xnor U10427 (N_10427,N_9515,N_9942);
nor U10428 (N_10428,N_9818,N_9829);
or U10429 (N_10429,N_9508,N_9991);
nor U10430 (N_10430,N_9845,N_9556);
and U10431 (N_10431,N_9726,N_9542);
xnor U10432 (N_10432,N_9626,N_9682);
nand U10433 (N_10433,N_9898,N_9533);
nor U10434 (N_10434,N_9835,N_9661);
and U10435 (N_10435,N_9727,N_9946);
nor U10436 (N_10436,N_9809,N_9796);
or U10437 (N_10437,N_9815,N_9604);
xnor U10438 (N_10438,N_9987,N_9969);
and U10439 (N_10439,N_9873,N_9527);
nor U10440 (N_10440,N_9721,N_9824);
xnor U10441 (N_10441,N_9532,N_9654);
xor U10442 (N_10442,N_9851,N_9524);
xnor U10443 (N_10443,N_9899,N_9739);
nor U10444 (N_10444,N_9719,N_9554);
xnor U10445 (N_10445,N_9768,N_9743);
nor U10446 (N_10446,N_9646,N_9721);
or U10447 (N_10447,N_9999,N_9875);
or U10448 (N_10448,N_9633,N_9893);
xor U10449 (N_10449,N_9746,N_9507);
nand U10450 (N_10450,N_9860,N_9687);
xor U10451 (N_10451,N_9987,N_9932);
nand U10452 (N_10452,N_9647,N_9570);
nand U10453 (N_10453,N_9537,N_9996);
nand U10454 (N_10454,N_9608,N_9518);
xnor U10455 (N_10455,N_9863,N_9911);
xor U10456 (N_10456,N_9976,N_9842);
or U10457 (N_10457,N_9758,N_9690);
xor U10458 (N_10458,N_9759,N_9967);
nor U10459 (N_10459,N_9979,N_9869);
nand U10460 (N_10460,N_9511,N_9594);
nor U10461 (N_10461,N_9698,N_9801);
nor U10462 (N_10462,N_9672,N_9542);
xor U10463 (N_10463,N_9732,N_9793);
nand U10464 (N_10464,N_9770,N_9697);
xnor U10465 (N_10465,N_9809,N_9790);
nand U10466 (N_10466,N_9776,N_9587);
or U10467 (N_10467,N_9841,N_9624);
xor U10468 (N_10468,N_9807,N_9769);
or U10469 (N_10469,N_9897,N_9876);
nand U10470 (N_10470,N_9830,N_9591);
or U10471 (N_10471,N_9901,N_9625);
nor U10472 (N_10472,N_9780,N_9579);
xor U10473 (N_10473,N_9968,N_9800);
nand U10474 (N_10474,N_9965,N_9893);
or U10475 (N_10475,N_9510,N_9771);
nor U10476 (N_10476,N_9993,N_9676);
xnor U10477 (N_10477,N_9630,N_9623);
xnor U10478 (N_10478,N_9818,N_9960);
or U10479 (N_10479,N_9579,N_9696);
and U10480 (N_10480,N_9539,N_9896);
xnor U10481 (N_10481,N_9958,N_9690);
or U10482 (N_10482,N_9583,N_9628);
nor U10483 (N_10483,N_9646,N_9535);
and U10484 (N_10484,N_9599,N_9511);
nand U10485 (N_10485,N_9561,N_9912);
nor U10486 (N_10486,N_9982,N_9668);
nand U10487 (N_10487,N_9902,N_9780);
xor U10488 (N_10488,N_9882,N_9959);
and U10489 (N_10489,N_9755,N_9773);
nor U10490 (N_10490,N_9923,N_9911);
nor U10491 (N_10491,N_9942,N_9828);
nor U10492 (N_10492,N_9798,N_9786);
nand U10493 (N_10493,N_9937,N_9888);
and U10494 (N_10494,N_9651,N_9656);
nand U10495 (N_10495,N_9643,N_9704);
or U10496 (N_10496,N_9856,N_9676);
nor U10497 (N_10497,N_9838,N_9798);
nor U10498 (N_10498,N_9759,N_9687);
and U10499 (N_10499,N_9673,N_9760);
nand U10500 (N_10500,N_10344,N_10106);
or U10501 (N_10501,N_10017,N_10138);
and U10502 (N_10502,N_10490,N_10141);
and U10503 (N_10503,N_10395,N_10198);
xor U10504 (N_10504,N_10264,N_10021);
nor U10505 (N_10505,N_10208,N_10183);
nor U10506 (N_10506,N_10057,N_10329);
nand U10507 (N_10507,N_10045,N_10091);
nor U10508 (N_10508,N_10493,N_10054);
or U10509 (N_10509,N_10014,N_10466);
and U10510 (N_10510,N_10423,N_10210);
nor U10511 (N_10511,N_10366,N_10376);
nor U10512 (N_10512,N_10327,N_10098);
and U10513 (N_10513,N_10131,N_10371);
nand U10514 (N_10514,N_10246,N_10253);
xnor U10515 (N_10515,N_10209,N_10100);
and U10516 (N_10516,N_10486,N_10140);
xnor U10517 (N_10517,N_10002,N_10353);
or U10518 (N_10518,N_10165,N_10034);
nand U10519 (N_10519,N_10185,N_10328);
or U10520 (N_10520,N_10146,N_10375);
xnor U10521 (N_10521,N_10211,N_10278);
xnor U10522 (N_10522,N_10405,N_10319);
and U10523 (N_10523,N_10364,N_10242);
nor U10524 (N_10524,N_10060,N_10063);
xor U10525 (N_10525,N_10385,N_10051);
or U10526 (N_10526,N_10042,N_10425);
nand U10527 (N_10527,N_10429,N_10473);
or U10528 (N_10528,N_10426,N_10194);
nand U10529 (N_10529,N_10201,N_10020);
xor U10530 (N_10530,N_10262,N_10167);
nand U10531 (N_10531,N_10118,N_10450);
or U10532 (N_10532,N_10256,N_10010);
or U10533 (N_10533,N_10396,N_10199);
or U10534 (N_10534,N_10235,N_10024);
xnor U10535 (N_10535,N_10133,N_10424);
nand U10536 (N_10536,N_10357,N_10207);
and U10537 (N_10537,N_10145,N_10267);
nor U10538 (N_10538,N_10221,N_10187);
nand U10539 (N_10539,N_10471,N_10044);
or U10540 (N_10540,N_10276,N_10484);
or U10541 (N_10541,N_10491,N_10005);
nand U10542 (N_10542,N_10186,N_10386);
or U10543 (N_10543,N_10340,N_10402);
nor U10544 (N_10544,N_10022,N_10065);
and U10545 (N_10545,N_10004,N_10108);
xor U10546 (N_10546,N_10325,N_10206);
nand U10547 (N_10547,N_10321,N_10121);
or U10548 (N_10548,N_10290,N_10422);
xor U10549 (N_10549,N_10409,N_10309);
xor U10550 (N_10550,N_10317,N_10233);
or U10551 (N_10551,N_10069,N_10388);
or U10552 (N_10552,N_10492,N_10369);
nand U10553 (N_10553,N_10417,N_10461);
and U10554 (N_10554,N_10124,N_10299);
or U10555 (N_10555,N_10096,N_10303);
nand U10556 (N_10556,N_10048,N_10348);
nor U10557 (N_10557,N_10190,N_10270);
nand U10558 (N_10558,N_10012,N_10377);
or U10559 (N_10559,N_10197,N_10305);
and U10560 (N_10560,N_10127,N_10240);
or U10561 (N_10561,N_10286,N_10237);
xnor U10562 (N_10562,N_10238,N_10283);
nand U10563 (N_10563,N_10463,N_10056);
nor U10564 (N_10564,N_10431,N_10081);
nor U10565 (N_10565,N_10322,N_10093);
and U10566 (N_10566,N_10026,N_10367);
and U10567 (N_10567,N_10115,N_10273);
nand U10568 (N_10568,N_10482,N_10153);
xor U10569 (N_10569,N_10159,N_10119);
and U10570 (N_10570,N_10293,N_10488);
or U10571 (N_10571,N_10403,N_10339);
xor U10572 (N_10572,N_10252,N_10176);
or U10573 (N_10573,N_10180,N_10025);
nand U10574 (N_10574,N_10363,N_10448);
nand U10575 (N_10575,N_10228,N_10084);
and U10576 (N_10576,N_10204,N_10362);
xor U10577 (N_10577,N_10112,N_10430);
or U10578 (N_10578,N_10464,N_10092);
nor U10579 (N_10579,N_10037,N_10090);
and U10580 (N_10580,N_10035,N_10487);
and U10581 (N_10581,N_10458,N_10314);
or U10582 (N_10582,N_10134,N_10408);
nand U10583 (N_10583,N_10465,N_10156);
nand U10584 (N_10584,N_10105,N_10343);
xnor U10585 (N_10585,N_10421,N_10263);
nand U10586 (N_10586,N_10415,N_10177);
nor U10587 (N_10587,N_10076,N_10323);
xor U10588 (N_10588,N_10447,N_10496);
nor U10589 (N_10589,N_10498,N_10128);
or U10590 (N_10590,N_10383,N_10439);
nand U10591 (N_10591,N_10453,N_10370);
xnor U10592 (N_10592,N_10341,N_10088);
nor U10593 (N_10593,N_10116,N_10077);
xnor U10594 (N_10594,N_10297,N_10427);
xnor U10595 (N_10595,N_10070,N_10315);
xor U10596 (N_10596,N_10481,N_10301);
xor U10597 (N_10597,N_10231,N_10387);
nor U10598 (N_10598,N_10311,N_10279);
xor U10599 (N_10599,N_10347,N_10298);
nor U10600 (N_10600,N_10178,N_10324);
nor U10601 (N_10601,N_10248,N_10239);
nor U10602 (N_10602,N_10470,N_10372);
and U10603 (N_10603,N_10030,N_10226);
xnor U10604 (N_10604,N_10359,N_10313);
or U10605 (N_10605,N_10288,N_10399);
and U10606 (N_10606,N_10277,N_10354);
nor U10607 (N_10607,N_10023,N_10457);
or U10608 (N_10608,N_10038,N_10438);
xor U10609 (N_10609,N_10175,N_10280);
xnor U10610 (N_10610,N_10113,N_10310);
xor U10611 (N_10611,N_10222,N_10203);
nand U10612 (N_10612,N_10123,N_10161);
nor U10613 (N_10613,N_10166,N_10214);
or U10614 (N_10614,N_10043,N_10342);
or U10615 (N_10615,N_10467,N_10179);
or U10616 (N_10616,N_10384,N_10182);
xor U10617 (N_10617,N_10346,N_10250);
nand U10618 (N_10618,N_10041,N_10160);
and U10619 (N_10619,N_10188,N_10304);
or U10620 (N_10620,N_10483,N_10072);
nand U10621 (N_10621,N_10468,N_10040);
and U10622 (N_10622,N_10073,N_10068);
or U10623 (N_10623,N_10085,N_10373);
and U10624 (N_10624,N_10169,N_10011);
and U10625 (N_10625,N_10232,N_10079);
and U10626 (N_10626,N_10397,N_10401);
xnor U10627 (N_10627,N_10260,N_10476);
and U10628 (N_10628,N_10337,N_10196);
nand U10629 (N_10629,N_10082,N_10016);
nand U10630 (N_10630,N_10087,N_10053);
xor U10631 (N_10631,N_10406,N_10202);
nand U10632 (N_10632,N_10110,N_10215);
nand U10633 (N_10633,N_10007,N_10061);
xor U10634 (N_10634,N_10331,N_10219);
and U10635 (N_10635,N_10358,N_10174);
or U10636 (N_10636,N_10360,N_10410);
nand U10637 (N_10637,N_10257,N_10200);
xor U10638 (N_10638,N_10195,N_10157);
and U10639 (N_10639,N_10454,N_10411);
xor U10640 (N_10640,N_10381,N_10052);
and U10641 (N_10641,N_10152,N_10352);
and U10642 (N_10642,N_10398,N_10058);
nand U10643 (N_10643,N_10216,N_10374);
nor U10644 (N_10644,N_10055,N_10125);
nand U10645 (N_10645,N_10265,N_10379);
nand U10646 (N_10646,N_10338,N_10300);
xnor U10647 (N_10647,N_10400,N_10320);
nand U10648 (N_10648,N_10436,N_10130);
nand U10649 (N_10649,N_10050,N_10001);
nor U10650 (N_10650,N_10318,N_10129);
nor U10651 (N_10651,N_10143,N_10142);
nor U10652 (N_10652,N_10191,N_10258);
nand U10653 (N_10653,N_10170,N_10220);
and U10654 (N_10654,N_10393,N_10064);
xnor U10655 (N_10655,N_10472,N_10149);
or U10656 (N_10656,N_10217,N_10158);
nor U10657 (N_10657,N_10066,N_10378);
and U10658 (N_10658,N_10028,N_10489);
nor U10659 (N_10659,N_10245,N_10459);
and U10660 (N_10660,N_10111,N_10412);
xnor U10661 (N_10661,N_10099,N_10441);
or U10662 (N_10662,N_10418,N_10289);
nor U10663 (N_10663,N_10150,N_10102);
nand U10664 (N_10664,N_10462,N_10469);
and U10665 (N_10665,N_10281,N_10485);
nor U10666 (N_10666,N_10274,N_10224);
nand U10667 (N_10667,N_10032,N_10046);
nand U10668 (N_10668,N_10306,N_10189);
xor U10669 (N_10669,N_10446,N_10122);
xnor U10670 (N_10670,N_10181,N_10332);
nor U10671 (N_10671,N_10452,N_10365);
nand U10672 (N_10672,N_10047,N_10137);
or U10673 (N_10673,N_10101,N_10266);
xnor U10674 (N_10674,N_10184,N_10368);
xnor U10675 (N_10675,N_10009,N_10247);
xor U10676 (N_10676,N_10413,N_10497);
or U10677 (N_10677,N_10480,N_10404);
nand U10678 (N_10678,N_10031,N_10036);
and U10679 (N_10679,N_10243,N_10033);
nand U10680 (N_10680,N_10162,N_10294);
nor U10681 (N_10681,N_10495,N_10390);
or U10682 (N_10682,N_10229,N_10269);
nand U10683 (N_10683,N_10335,N_10168);
nor U10684 (N_10684,N_10435,N_10312);
nor U10685 (N_10685,N_10336,N_10259);
or U10686 (N_10686,N_10205,N_10382);
nor U10687 (N_10687,N_10356,N_10451);
xor U10688 (N_10688,N_10027,N_10287);
xnor U10689 (N_10689,N_10475,N_10499);
or U10690 (N_10690,N_10330,N_10249);
nor U10691 (N_10691,N_10416,N_10104);
xor U10692 (N_10692,N_10097,N_10244);
nor U10693 (N_10693,N_10478,N_10477);
or U10694 (N_10694,N_10443,N_10282);
or U10695 (N_10695,N_10271,N_10013);
or U10696 (N_10696,N_10349,N_10455);
nor U10697 (N_10697,N_10275,N_10172);
nor U10698 (N_10698,N_10261,N_10444);
and U10699 (N_10699,N_10049,N_10139);
or U10700 (N_10700,N_10193,N_10227);
and U10701 (N_10701,N_10285,N_10018);
nand U10702 (N_10702,N_10456,N_10272);
nand U10703 (N_10703,N_10414,N_10291);
nand U10704 (N_10704,N_10241,N_10086);
or U10705 (N_10705,N_10000,N_10223);
nand U10706 (N_10706,N_10155,N_10136);
nor U10707 (N_10707,N_10039,N_10292);
or U10708 (N_10708,N_10059,N_10420);
xor U10709 (N_10709,N_10135,N_10302);
nand U10710 (N_10710,N_10334,N_10164);
or U10711 (N_10711,N_10019,N_10144);
nand U10712 (N_10712,N_10015,N_10008);
nand U10713 (N_10713,N_10163,N_10440);
xor U10714 (N_10714,N_10460,N_10428);
and U10715 (N_10715,N_10062,N_10089);
and U10716 (N_10716,N_10437,N_10361);
and U10717 (N_10717,N_10080,N_10445);
or U10718 (N_10718,N_10254,N_10003);
nand U10719 (N_10719,N_10107,N_10350);
or U10720 (N_10720,N_10434,N_10132);
xnor U10721 (N_10721,N_10255,N_10442);
nor U10722 (N_10722,N_10268,N_10029);
or U10723 (N_10723,N_10151,N_10078);
nand U10724 (N_10724,N_10074,N_10083);
nor U10725 (N_10725,N_10114,N_10433);
and U10726 (N_10726,N_10213,N_10474);
xor U10727 (N_10727,N_10192,N_10380);
nand U10728 (N_10728,N_10126,N_10345);
or U10729 (N_10729,N_10148,N_10351);
and U10730 (N_10730,N_10284,N_10391);
nor U10731 (N_10731,N_10308,N_10154);
nor U10732 (N_10732,N_10394,N_10071);
or U10733 (N_10733,N_10171,N_10449);
xnor U10734 (N_10734,N_10479,N_10389);
or U10735 (N_10735,N_10307,N_10173);
nor U10736 (N_10736,N_10006,N_10296);
and U10737 (N_10737,N_10117,N_10432);
or U10738 (N_10738,N_10419,N_10316);
xor U10739 (N_10739,N_10230,N_10212);
or U10740 (N_10740,N_10095,N_10120);
and U10741 (N_10741,N_10109,N_10094);
xnor U10742 (N_10742,N_10234,N_10147);
or U10743 (N_10743,N_10251,N_10407);
nand U10744 (N_10744,N_10225,N_10075);
or U10745 (N_10745,N_10218,N_10355);
or U10746 (N_10746,N_10236,N_10326);
and U10747 (N_10747,N_10295,N_10103);
or U10748 (N_10748,N_10494,N_10333);
nand U10749 (N_10749,N_10067,N_10392);
or U10750 (N_10750,N_10387,N_10278);
nor U10751 (N_10751,N_10165,N_10424);
or U10752 (N_10752,N_10132,N_10049);
and U10753 (N_10753,N_10058,N_10424);
nor U10754 (N_10754,N_10182,N_10208);
and U10755 (N_10755,N_10272,N_10005);
or U10756 (N_10756,N_10270,N_10244);
or U10757 (N_10757,N_10011,N_10475);
nand U10758 (N_10758,N_10493,N_10405);
nor U10759 (N_10759,N_10481,N_10254);
xnor U10760 (N_10760,N_10182,N_10030);
or U10761 (N_10761,N_10144,N_10016);
nor U10762 (N_10762,N_10362,N_10167);
and U10763 (N_10763,N_10420,N_10020);
xnor U10764 (N_10764,N_10242,N_10133);
nand U10765 (N_10765,N_10439,N_10450);
nor U10766 (N_10766,N_10272,N_10187);
and U10767 (N_10767,N_10037,N_10438);
and U10768 (N_10768,N_10043,N_10223);
or U10769 (N_10769,N_10287,N_10234);
nor U10770 (N_10770,N_10072,N_10161);
nor U10771 (N_10771,N_10091,N_10489);
xor U10772 (N_10772,N_10387,N_10025);
xor U10773 (N_10773,N_10368,N_10185);
nand U10774 (N_10774,N_10120,N_10078);
or U10775 (N_10775,N_10273,N_10141);
and U10776 (N_10776,N_10430,N_10069);
nand U10777 (N_10777,N_10354,N_10210);
xor U10778 (N_10778,N_10045,N_10150);
xnor U10779 (N_10779,N_10095,N_10252);
nand U10780 (N_10780,N_10387,N_10044);
nor U10781 (N_10781,N_10158,N_10336);
xor U10782 (N_10782,N_10456,N_10233);
xnor U10783 (N_10783,N_10160,N_10179);
nor U10784 (N_10784,N_10191,N_10007);
or U10785 (N_10785,N_10292,N_10470);
nor U10786 (N_10786,N_10000,N_10272);
nor U10787 (N_10787,N_10037,N_10077);
nor U10788 (N_10788,N_10072,N_10420);
or U10789 (N_10789,N_10396,N_10248);
nor U10790 (N_10790,N_10054,N_10287);
nor U10791 (N_10791,N_10261,N_10091);
xnor U10792 (N_10792,N_10494,N_10392);
or U10793 (N_10793,N_10416,N_10165);
and U10794 (N_10794,N_10233,N_10226);
nor U10795 (N_10795,N_10493,N_10477);
nor U10796 (N_10796,N_10091,N_10352);
or U10797 (N_10797,N_10313,N_10133);
and U10798 (N_10798,N_10337,N_10262);
nor U10799 (N_10799,N_10125,N_10057);
nor U10800 (N_10800,N_10227,N_10390);
and U10801 (N_10801,N_10459,N_10417);
and U10802 (N_10802,N_10222,N_10193);
nand U10803 (N_10803,N_10467,N_10437);
or U10804 (N_10804,N_10383,N_10316);
and U10805 (N_10805,N_10433,N_10237);
xor U10806 (N_10806,N_10386,N_10280);
nand U10807 (N_10807,N_10332,N_10178);
or U10808 (N_10808,N_10333,N_10116);
nand U10809 (N_10809,N_10344,N_10088);
or U10810 (N_10810,N_10356,N_10029);
xnor U10811 (N_10811,N_10236,N_10162);
xnor U10812 (N_10812,N_10114,N_10401);
nor U10813 (N_10813,N_10064,N_10276);
nor U10814 (N_10814,N_10112,N_10154);
xor U10815 (N_10815,N_10039,N_10309);
or U10816 (N_10816,N_10161,N_10281);
nand U10817 (N_10817,N_10401,N_10480);
nor U10818 (N_10818,N_10218,N_10114);
nor U10819 (N_10819,N_10015,N_10394);
or U10820 (N_10820,N_10374,N_10272);
or U10821 (N_10821,N_10345,N_10010);
or U10822 (N_10822,N_10293,N_10034);
or U10823 (N_10823,N_10392,N_10309);
and U10824 (N_10824,N_10436,N_10429);
and U10825 (N_10825,N_10232,N_10093);
and U10826 (N_10826,N_10416,N_10273);
xnor U10827 (N_10827,N_10300,N_10484);
nand U10828 (N_10828,N_10401,N_10015);
nor U10829 (N_10829,N_10137,N_10195);
nor U10830 (N_10830,N_10069,N_10088);
or U10831 (N_10831,N_10091,N_10389);
nand U10832 (N_10832,N_10188,N_10296);
or U10833 (N_10833,N_10226,N_10496);
and U10834 (N_10834,N_10372,N_10024);
or U10835 (N_10835,N_10106,N_10460);
and U10836 (N_10836,N_10116,N_10063);
nor U10837 (N_10837,N_10138,N_10246);
xor U10838 (N_10838,N_10440,N_10380);
or U10839 (N_10839,N_10217,N_10344);
and U10840 (N_10840,N_10421,N_10428);
nand U10841 (N_10841,N_10172,N_10150);
nor U10842 (N_10842,N_10060,N_10483);
nor U10843 (N_10843,N_10073,N_10076);
nand U10844 (N_10844,N_10199,N_10090);
and U10845 (N_10845,N_10337,N_10447);
nand U10846 (N_10846,N_10384,N_10451);
xnor U10847 (N_10847,N_10359,N_10064);
nand U10848 (N_10848,N_10344,N_10182);
and U10849 (N_10849,N_10176,N_10397);
nor U10850 (N_10850,N_10341,N_10245);
or U10851 (N_10851,N_10414,N_10373);
or U10852 (N_10852,N_10310,N_10060);
and U10853 (N_10853,N_10403,N_10472);
and U10854 (N_10854,N_10360,N_10002);
or U10855 (N_10855,N_10124,N_10148);
nor U10856 (N_10856,N_10443,N_10303);
xnor U10857 (N_10857,N_10187,N_10420);
nor U10858 (N_10858,N_10415,N_10154);
and U10859 (N_10859,N_10424,N_10157);
xor U10860 (N_10860,N_10285,N_10082);
or U10861 (N_10861,N_10018,N_10267);
or U10862 (N_10862,N_10487,N_10183);
xnor U10863 (N_10863,N_10030,N_10082);
xor U10864 (N_10864,N_10084,N_10257);
xnor U10865 (N_10865,N_10083,N_10238);
xor U10866 (N_10866,N_10309,N_10412);
xnor U10867 (N_10867,N_10385,N_10121);
or U10868 (N_10868,N_10356,N_10312);
nand U10869 (N_10869,N_10394,N_10471);
xnor U10870 (N_10870,N_10372,N_10195);
nor U10871 (N_10871,N_10216,N_10167);
or U10872 (N_10872,N_10069,N_10145);
or U10873 (N_10873,N_10363,N_10452);
or U10874 (N_10874,N_10265,N_10331);
nor U10875 (N_10875,N_10137,N_10135);
xnor U10876 (N_10876,N_10076,N_10365);
nand U10877 (N_10877,N_10158,N_10259);
nor U10878 (N_10878,N_10172,N_10299);
nand U10879 (N_10879,N_10366,N_10060);
xnor U10880 (N_10880,N_10453,N_10361);
xnor U10881 (N_10881,N_10084,N_10087);
or U10882 (N_10882,N_10309,N_10099);
nor U10883 (N_10883,N_10162,N_10128);
or U10884 (N_10884,N_10358,N_10253);
xor U10885 (N_10885,N_10425,N_10330);
nand U10886 (N_10886,N_10309,N_10224);
or U10887 (N_10887,N_10238,N_10126);
nor U10888 (N_10888,N_10413,N_10011);
xnor U10889 (N_10889,N_10126,N_10013);
nor U10890 (N_10890,N_10341,N_10167);
or U10891 (N_10891,N_10224,N_10153);
nand U10892 (N_10892,N_10084,N_10369);
nand U10893 (N_10893,N_10449,N_10003);
and U10894 (N_10894,N_10222,N_10173);
nor U10895 (N_10895,N_10493,N_10184);
nand U10896 (N_10896,N_10482,N_10263);
or U10897 (N_10897,N_10430,N_10332);
nand U10898 (N_10898,N_10270,N_10383);
and U10899 (N_10899,N_10499,N_10102);
xnor U10900 (N_10900,N_10055,N_10462);
nor U10901 (N_10901,N_10058,N_10149);
and U10902 (N_10902,N_10201,N_10132);
and U10903 (N_10903,N_10404,N_10368);
nand U10904 (N_10904,N_10237,N_10456);
or U10905 (N_10905,N_10361,N_10117);
nand U10906 (N_10906,N_10348,N_10085);
and U10907 (N_10907,N_10222,N_10429);
xnor U10908 (N_10908,N_10143,N_10091);
or U10909 (N_10909,N_10139,N_10375);
nand U10910 (N_10910,N_10070,N_10250);
nand U10911 (N_10911,N_10208,N_10318);
and U10912 (N_10912,N_10080,N_10102);
nor U10913 (N_10913,N_10189,N_10266);
and U10914 (N_10914,N_10214,N_10446);
and U10915 (N_10915,N_10073,N_10256);
or U10916 (N_10916,N_10350,N_10230);
xor U10917 (N_10917,N_10222,N_10440);
xnor U10918 (N_10918,N_10273,N_10285);
xor U10919 (N_10919,N_10108,N_10213);
or U10920 (N_10920,N_10320,N_10009);
nor U10921 (N_10921,N_10432,N_10007);
nor U10922 (N_10922,N_10414,N_10429);
nor U10923 (N_10923,N_10063,N_10049);
nor U10924 (N_10924,N_10015,N_10217);
nand U10925 (N_10925,N_10016,N_10359);
nand U10926 (N_10926,N_10168,N_10306);
or U10927 (N_10927,N_10358,N_10444);
xor U10928 (N_10928,N_10430,N_10150);
xnor U10929 (N_10929,N_10042,N_10095);
nor U10930 (N_10930,N_10467,N_10001);
nor U10931 (N_10931,N_10491,N_10169);
nand U10932 (N_10932,N_10387,N_10385);
or U10933 (N_10933,N_10289,N_10147);
nor U10934 (N_10934,N_10035,N_10042);
nor U10935 (N_10935,N_10216,N_10484);
nand U10936 (N_10936,N_10411,N_10146);
nor U10937 (N_10937,N_10433,N_10472);
xnor U10938 (N_10938,N_10023,N_10304);
xnor U10939 (N_10939,N_10274,N_10415);
or U10940 (N_10940,N_10428,N_10366);
nand U10941 (N_10941,N_10162,N_10374);
and U10942 (N_10942,N_10006,N_10037);
nor U10943 (N_10943,N_10394,N_10365);
or U10944 (N_10944,N_10438,N_10252);
xor U10945 (N_10945,N_10323,N_10054);
nor U10946 (N_10946,N_10037,N_10132);
or U10947 (N_10947,N_10409,N_10049);
or U10948 (N_10948,N_10379,N_10145);
xor U10949 (N_10949,N_10364,N_10245);
or U10950 (N_10950,N_10290,N_10129);
xnor U10951 (N_10951,N_10327,N_10052);
nor U10952 (N_10952,N_10101,N_10334);
or U10953 (N_10953,N_10038,N_10182);
nor U10954 (N_10954,N_10165,N_10472);
and U10955 (N_10955,N_10128,N_10013);
xnor U10956 (N_10956,N_10264,N_10427);
or U10957 (N_10957,N_10073,N_10286);
and U10958 (N_10958,N_10443,N_10022);
nor U10959 (N_10959,N_10019,N_10487);
nand U10960 (N_10960,N_10114,N_10021);
or U10961 (N_10961,N_10142,N_10152);
nor U10962 (N_10962,N_10373,N_10474);
or U10963 (N_10963,N_10225,N_10221);
nor U10964 (N_10964,N_10264,N_10117);
nand U10965 (N_10965,N_10242,N_10225);
or U10966 (N_10966,N_10420,N_10243);
or U10967 (N_10967,N_10420,N_10192);
nor U10968 (N_10968,N_10086,N_10476);
or U10969 (N_10969,N_10008,N_10042);
nor U10970 (N_10970,N_10226,N_10122);
or U10971 (N_10971,N_10026,N_10244);
nand U10972 (N_10972,N_10454,N_10329);
nor U10973 (N_10973,N_10343,N_10317);
nor U10974 (N_10974,N_10259,N_10352);
xnor U10975 (N_10975,N_10051,N_10126);
nand U10976 (N_10976,N_10044,N_10016);
nor U10977 (N_10977,N_10331,N_10277);
and U10978 (N_10978,N_10110,N_10158);
or U10979 (N_10979,N_10296,N_10433);
or U10980 (N_10980,N_10054,N_10347);
or U10981 (N_10981,N_10075,N_10083);
nand U10982 (N_10982,N_10215,N_10175);
and U10983 (N_10983,N_10432,N_10489);
and U10984 (N_10984,N_10199,N_10099);
nor U10985 (N_10985,N_10080,N_10408);
and U10986 (N_10986,N_10210,N_10374);
or U10987 (N_10987,N_10216,N_10155);
or U10988 (N_10988,N_10004,N_10486);
or U10989 (N_10989,N_10290,N_10023);
and U10990 (N_10990,N_10015,N_10284);
nand U10991 (N_10991,N_10086,N_10429);
xor U10992 (N_10992,N_10166,N_10365);
or U10993 (N_10993,N_10148,N_10077);
and U10994 (N_10994,N_10272,N_10301);
xor U10995 (N_10995,N_10249,N_10084);
nor U10996 (N_10996,N_10128,N_10404);
and U10997 (N_10997,N_10041,N_10368);
nor U10998 (N_10998,N_10193,N_10241);
or U10999 (N_10999,N_10249,N_10364);
or U11000 (N_11000,N_10598,N_10988);
nor U11001 (N_11001,N_10503,N_10507);
and U11002 (N_11002,N_10792,N_10809);
nor U11003 (N_11003,N_10837,N_10512);
nor U11004 (N_11004,N_10618,N_10818);
nor U11005 (N_11005,N_10690,N_10681);
or U11006 (N_11006,N_10637,N_10955);
nand U11007 (N_11007,N_10509,N_10536);
and U11008 (N_11008,N_10985,N_10606);
or U11009 (N_11009,N_10776,N_10798);
xnor U11010 (N_11010,N_10870,N_10580);
and U11011 (N_11011,N_10656,N_10605);
xor U11012 (N_11012,N_10811,N_10884);
nor U11013 (N_11013,N_10881,N_10930);
nand U11014 (N_11014,N_10890,N_10511);
xor U11015 (N_11015,N_10629,N_10749);
nand U11016 (N_11016,N_10584,N_10938);
nand U11017 (N_11017,N_10953,N_10773);
xnor U11018 (N_11018,N_10970,N_10980);
nand U11019 (N_11019,N_10824,N_10672);
xnor U11020 (N_11020,N_10735,N_10500);
xor U11021 (N_11021,N_10857,N_10942);
and U11022 (N_11022,N_10558,N_10934);
and U11023 (N_11023,N_10704,N_10533);
or U11024 (N_11024,N_10997,N_10582);
xnor U11025 (N_11025,N_10796,N_10520);
nor U11026 (N_11026,N_10995,N_10635);
nand U11027 (N_11027,N_10611,N_10647);
nor U11028 (N_11028,N_10855,N_10543);
nor U11029 (N_11029,N_10803,N_10914);
or U11030 (N_11030,N_10548,N_10686);
and U11031 (N_11031,N_10570,N_10909);
or U11032 (N_11032,N_10717,N_10880);
nor U11033 (N_11033,N_10514,N_10730);
xor U11034 (N_11034,N_10941,N_10994);
or U11035 (N_11035,N_10555,N_10673);
or U11036 (N_11036,N_10604,N_10648);
xor U11037 (N_11037,N_10869,N_10778);
xor U11038 (N_11038,N_10845,N_10940);
or U11039 (N_11039,N_10614,N_10624);
nand U11040 (N_11040,N_10990,N_10891);
and U11041 (N_11041,N_10563,N_10767);
or U11042 (N_11042,N_10682,N_10562);
or U11043 (N_11043,N_10963,N_10725);
or U11044 (N_11044,N_10879,N_10593);
or U11045 (N_11045,N_10554,N_10685);
and U11046 (N_11046,N_10766,N_10783);
or U11047 (N_11047,N_10978,N_10810);
xor U11048 (N_11048,N_10949,N_10616);
nand U11049 (N_11049,N_10713,N_10873);
and U11050 (N_11050,N_10699,N_10758);
nor U11051 (N_11051,N_10784,N_10993);
nand U11052 (N_11052,N_10969,N_10788);
xor U11053 (N_11053,N_10566,N_10760);
or U11054 (N_11054,N_10744,N_10908);
xor U11055 (N_11055,N_10660,N_10862);
and U11056 (N_11056,N_10849,N_10721);
nand U11057 (N_11057,N_10587,N_10762);
or U11058 (N_11058,N_10989,N_10799);
nand U11059 (N_11059,N_10772,N_10828);
nand U11060 (N_11060,N_10984,N_10950);
or U11061 (N_11061,N_10835,N_10751);
nand U11062 (N_11062,N_10755,N_10831);
and U11063 (N_11063,N_10638,N_10865);
xor U11064 (N_11064,N_10759,N_10677);
xor U11065 (N_11065,N_10928,N_10684);
xor U11066 (N_11066,N_10820,N_10797);
nor U11067 (N_11067,N_10781,N_10972);
and U11068 (N_11068,N_10557,N_10607);
nor U11069 (N_11069,N_10898,N_10896);
nand U11070 (N_11070,N_10750,N_10707);
or U11071 (N_11071,N_10851,N_10737);
xnor U11072 (N_11072,N_10723,N_10868);
or U11073 (N_11073,N_10519,N_10692);
xnor U11074 (N_11074,N_10731,N_10626);
and U11075 (N_11075,N_10859,N_10537);
nand U11076 (N_11076,N_10669,N_10631);
and U11077 (N_11077,N_10588,N_10747);
and U11078 (N_11078,N_10510,N_10528);
nand U11079 (N_11079,N_10675,N_10623);
xnor U11080 (N_11080,N_10931,N_10667);
nand U11081 (N_11081,N_10608,N_10874);
nor U11082 (N_11082,N_10829,N_10960);
nand U11083 (N_11083,N_10695,N_10535);
nor U11084 (N_11084,N_10714,N_10912);
nor U11085 (N_11085,N_10551,N_10569);
xnor U11086 (N_11086,N_10559,N_10517);
and U11087 (N_11087,N_10866,N_10863);
xnor U11088 (N_11088,N_10589,N_10697);
nand U11089 (N_11089,N_10753,N_10998);
nand U11090 (N_11090,N_10944,N_10904);
nor U11091 (N_11091,N_10987,N_10933);
xnor U11092 (N_11092,N_10756,N_10687);
nor U11093 (N_11093,N_10703,N_10504);
or U11094 (N_11094,N_10875,N_10644);
nor U11095 (N_11095,N_10550,N_10823);
xnor U11096 (N_11096,N_10668,N_10646);
and U11097 (N_11097,N_10991,N_10757);
and U11098 (N_11098,N_10733,N_10951);
xor U11099 (N_11099,N_10889,N_10954);
nand U11100 (N_11100,N_10903,N_10625);
and U11101 (N_11101,N_10892,N_10728);
or U11102 (N_11102,N_10806,N_10974);
nand U11103 (N_11103,N_10878,N_10741);
or U11104 (N_11104,N_10917,N_10915);
nor U11105 (N_11105,N_10542,N_10545);
or U11106 (N_11106,N_10779,N_10771);
or U11107 (N_11107,N_10708,N_10549);
nand U11108 (N_11108,N_10794,N_10621);
xor U11109 (N_11109,N_10929,N_10547);
or U11110 (N_11110,N_10659,N_10641);
xor U11111 (N_11111,N_10992,N_10975);
or U11112 (N_11112,N_10977,N_10864);
and U11113 (N_11113,N_10576,N_10657);
nor U11114 (N_11114,N_10578,N_10586);
nor U11115 (N_11115,N_10847,N_10948);
nor U11116 (N_11116,N_10508,N_10945);
or U11117 (N_11117,N_10632,N_10680);
xnor U11118 (N_11118,N_10683,N_10833);
nor U11119 (N_11119,N_10743,N_10952);
and U11120 (N_11120,N_10802,N_10665);
nand U11121 (N_11121,N_10722,N_10654);
nand U11122 (N_11122,N_10817,N_10959);
nor U11123 (N_11123,N_10574,N_10622);
or U11124 (N_11124,N_10825,N_10523);
or U11125 (N_11125,N_10612,N_10590);
or U11126 (N_11126,N_10872,N_10782);
nand U11127 (N_11127,N_10719,N_10645);
nand U11128 (N_11128,N_10615,N_10853);
nor U11129 (N_11129,N_10702,N_10516);
nor U11130 (N_11130,N_10765,N_10848);
xor U11131 (N_11131,N_10585,N_10877);
and U11132 (N_11132,N_10513,N_10630);
nor U11133 (N_11133,N_10712,N_10964);
nor U11134 (N_11134,N_10716,N_10663);
or U11135 (N_11135,N_10724,N_10642);
and U11136 (N_11136,N_10601,N_10739);
nand U11137 (N_11137,N_10594,N_10894);
or U11138 (N_11138,N_10981,N_10946);
or U11139 (N_11139,N_10826,N_10775);
and U11140 (N_11140,N_10577,N_10807);
nor U11141 (N_11141,N_10666,N_10812);
and U11142 (N_11142,N_10777,N_10653);
nand U11143 (N_11143,N_10899,N_10501);
nor U11144 (N_11144,N_10958,N_10962);
and U11145 (N_11145,N_10640,N_10842);
nor U11146 (N_11146,N_10764,N_10619);
nand U11147 (N_11147,N_10564,N_10922);
nand U11148 (N_11148,N_10532,N_10652);
nor U11149 (N_11149,N_10661,N_10650);
and U11150 (N_11150,N_10800,N_10814);
or U11151 (N_11151,N_10732,N_10836);
nand U11152 (N_11152,N_10726,N_10957);
or U11153 (N_11153,N_10526,N_10736);
nand U11154 (N_11154,N_10649,N_10738);
xnor U11155 (N_11155,N_10709,N_10936);
and U11156 (N_11156,N_10693,N_10919);
nand U11157 (N_11157,N_10740,N_10698);
xnor U11158 (N_11158,N_10926,N_10943);
xnor U11159 (N_11159,N_10567,N_10575);
xnor U11160 (N_11160,N_10620,N_10846);
nand U11161 (N_11161,N_10540,N_10634);
nand U11162 (N_11162,N_10591,N_10602);
and U11163 (N_11163,N_10924,N_10871);
or U11164 (N_11164,N_10902,N_10805);
or U11165 (N_11165,N_10754,N_10761);
nor U11166 (N_11166,N_10546,N_10808);
xor U11167 (N_11167,N_10861,N_10600);
nand U11168 (N_11168,N_10572,N_10561);
and U11169 (N_11169,N_10844,N_10900);
or U11170 (N_11170,N_10858,N_10920);
nand U11171 (N_11171,N_10789,N_10711);
or U11172 (N_11172,N_10923,N_10748);
or U11173 (N_11173,N_10530,N_10617);
nand U11174 (N_11174,N_10838,N_10529);
nand U11175 (N_11175,N_10583,N_10795);
or U11176 (N_11176,N_10973,N_10860);
and U11177 (N_11177,N_10983,N_10999);
or U11178 (N_11178,N_10552,N_10701);
nand U11179 (N_11179,N_10700,N_10895);
nand U11180 (N_11180,N_10882,N_10639);
and U11181 (N_11181,N_10907,N_10786);
xnor U11182 (N_11182,N_10839,N_10966);
nor U11183 (N_11183,N_10534,N_10843);
and U11184 (N_11184,N_10734,N_10705);
nor U11185 (N_11185,N_10925,N_10876);
xor U11186 (N_11186,N_10888,N_10592);
or U11187 (N_11187,N_10918,N_10935);
and U11188 (N_11188,N_10785,N_10581);
and U11189 (N_11189,N_10671,N_10752);
nand U11190 (N_11190,N_10518,N_10815);
and U11191 (N_11191,N_10763,N_10670);
nand U11192 (N_11192,N_10706,N_10599);
xor U11193 (N_11193,N_10819,N_10961);
nand U11194 (N_11194,N_10885,N_10633);
nand U11195 (N_11195,N_10718,N_10780);
nand U11196 (N_11196,N_10793,N_10976);
or U11197 (N_11197,N_10841,N_10906);
nor U11198 (N_11198,N_10971,N_10813);
nor U11199 (N_11199,N_10636,N_10729);
or U11200 (N_11200,N_10774,N_10541);
or U11201 (N_11201,N_10676,N_10901);
xor U11202 (N_11202,N_10965,N_10502);
xor U11203 (N_11203,N_10627,N_10834);
nand U11204 (N_11204,N_10967,N_10787);
nor U11205 (N_11205,N_10506,N_10610);
nor U11206 (N_11206,N_10694,N_10852);
nand U11207 (N_11207,N_10745,N_10664);
xnor U11208 (N_11208,N_10515,N_10897);
nor U11209 (N_11209,N_10538,N_10553);
xnor U11210 (N_11210,N_10932,N_10968);
and U11211 (N_11211,N_10727,N_10939);
nand U11212 (N_11212,N_10822,N_10790);
or U11213 (N_11213,N_10651,N_10609);
nand U11214 (N_11214,N_10710,N_10883);
and U11215 (N_11215,N_10613,N_10521);
and U11216 (N_11216,N_10571,N_10821);
or U11217 (N_11217,N_10643,N_10544);
xor U11218 (N_11218,N_10688,N_10524);
nand U11219 (N_11219,N_10927,N_10850);
xnor U11220 (N_11220,N_10579,N_10887);
nor U11221 (N_11221,N_10911,N_10505);
or U11222 (N_11222,N_10678,N_10979);
or U11223 (N_11223,N_10662,N_10560);
and U11224 (N_11224,N_10658,N_10691);
nor U11225 (N_11225,N_10522,N_10827);
nor U11226 (N_11226,N_10982,N_10893);
and U11227 (N_11227,N_10573,N_10746);
and U11228 (N_11228,N_10804,N_10867);
or U11229 (N_11229,N_10921,N_10905);
xor U11230 (N_11230,N_10715,N_10816);
xnor U11231 (N_11231,N_10556,N_10596);
xor U11232 (N_11232,N_10769,N_10720);
nand U11233 (N_11233,N_10840,N_10956);
nand U11234 (N_11234,N_10832,N_10996);
nand U11235 (N_11235,N_10655,N_10830);
nor U11236 (N_11236,N_10791,N_10854);
xnor U11237 (N_11237,N_10986,N_10689);
xnor U11238 (N_11238,N_10679,N_10597);
xnor U11239 (N_11239,N_10539,N_10595);
xor U11240 (N_11240,N_10916,N_10674);
and U11241 (N_11241,N_10525,N_10770);
or U11242 (N_11242,N_10603,N_10696);
nand U11243 (N_11243,N_10886,N_10856);
or U11244 (N_11244,N_10531,N_10913);
xor U11245 (N_11245,N_10910,N_10947);
xor U11246 (N_11246,N_10801,N_10768);
nand U11247 (N_11247,N_10527,N_10568);
nor U11248 (N_11248,N_10565,N_10937);
nand U11249 (N_11249,N_10742,N_10628);
xor U11250 (N_11250,N_10756,N_10818);
and U11251 (N_11251,N_10898,N_10654);
or U11252 (N_11252,N_10609,N_10741);
nor U11253 (N_11253,N_10866,N_10509);
xor U11254 (N_11254,N_10968,N_10795);
and U11255 (N_11255,N_10791,N_10804);
and U11256 (N_11256,N_10769,N_10989);
xnor U11257 (N_11257,N_10761,N_10964);
xnor U11258 (N_11258,N_10959,N_10985);
nor U11259 (N_11259,N_10831,N_10810);
nor U11260 (N_11260,N_10626,N_10606);
nand U11261 (N_11261,N_10833,N_10542);
and U11262 (N_11262,N_10527,N_10935);
nand U11263 (N_11263,N_10988,N_10948);
xnor U11264 (N_11264,N_10811,N_10871);
nand U11265 (N_11265,N_10583,N_10969);
nor U11266 (N_11266,N_10667,N_10747);
nand U11267 (N_11267,N_10881,N_10713);
and U11268 (N_11268,N_10557,N_10827);
xor U11269 (N_11269,N_10975,N_10769);
xor U11270 (N_11270,N_10809,N_10540);
nand U11271 (N_11271,N_10955,N_10716);
and U11272 (N_11272,N_10696,N_10740);
nor U11273 (N_11273,N_10734,N_10962);
and U11274 (N_11274,N_10745,N_10917);
or U11275 (N_11275,N_10526,N_10647);
nand U11276 (N_11276,N_10611,N_10991);
nand U11277 (N_11277,N_10709,N_10809);
and U11278 (N_11278,N_10588,N_10928);
and U11279 (N_11279,N_10798,N_10777);
and U11280 (N_11280,N_10572,N_10818);
nand U11281 (N_11281,N_10631,N_10703);
or U11282 (N_11282,N_10855,N_10655);
or U11283 (N_11283,N_10520,N_10981);
nand U11284 (N_11284,N_10707,N_10747);
nor U11285 (N_11285,N_10555,N_10669);
and U11286 (N_11286,N_10926,N_10878);
and U11287 (N_11287,N_10961,N_10893);
xnor U11288 (N_11288,N_10834,N_10552);
or U11289 (N_11289,N_10501,N_10760);
xor U11290 (N_11290,N_10544,N_10648);
xor U11291 (N_11291,N_10544,N_10587);
xnor U11292 (N_11292,N_10517,N_10671);
xnor U11293 (N_11293,N_10625,N_10973);
or U11294 (N_11294,N_10878,N_10698);
nand U11295 (N_11295,N_10934,N_10867);
xnor U11296 (N_11296,N_10794,N_10529);
or U11297 (N_11297,N_10981,N_10765);
nand U11298 (N_11298,N_10884,N_10501);
nor U11299 (N_11299,N_10724,N_10668);
xnor U11300 (N_11300,N_10926,N_10752);
nor U11301 (N_11301,N_10983,N_10755);
nor U11302 (N_11302,N_10526,N_10965);
nand U11303 (N_11303,N_10695,N_10721);
xnor U11304 (N_11304,N_10967,N_10509);
nor U11305 (N_11305,N_10843,N_10509);
and U11306 (N_11306,N_10980,N_10823);
xor U11307 (N_11307,N_10965,N_10621);
xor U11308 (N_11308,N_10699,N_10514);
nand U11309 (N_11309,N_10891,N_10732);
nand U11310 (N_11310,N_10534,N_10755);
nand U11311 (N_11311,N_10992,N_10855);
xor U11312 (N_11312,N_10959,N_10509);
or U11313 (N_11313,N_10954,N_10613);
or U11314 (N_11314,N_10562,N_10834);
nor U11315 (N_11315,N_10728,N_10955);
nand U11316 (N_11316,N_10716,N_10950);
xnor U11317 (N_11317,N_10614,N_10659);
nor U11318 (N_11318,N_10838,N_10667);
xnor U11319 (N_11319,N_10685,N_10649);
xor U11320 (N_11320,N_10547,N_10958);
nand U11321 (N_11321,N_10544,N_10833);
and U11322 (N_11322,N_10843,N_10983);
or U11323 (N_11323,N_10793,N_10896);
nor U11324 (N_11324,N_10725,N_10932);
or U11325 (N_11325,N_10518,N_10917);
and U11326 (N_11326,N_10886,N_10842);
or U11327 (N_11327,N_10563,N_10506);
nand U11328 (N_11328,N_10556,N_10839);
or U11329 (N_11329,N_10527,N_10584);
xnor U11330 (N_11330,N_10773,N_10948);
xor U11331 (N_11331,N_10610,N_10518);
or U11332 (N_11332,N_10935,N_10817);
nand U11333 (N_11333,N_10545,N_10871);
or U11334 (N_11334,N_10727,N_10643);
nor U11335 (N_11335,N_10798,N_10588);
xor U11336 (N_11336,N_10890,N_10744);
and U11337 (N_11337,N_10703,N_10849);
nand U11338 (N_11338,N_10896,N_10967);
nor U11339 (N_11339,N_10937,N_10735);
or U11340 (N_11340,N_10535,N_10648);
xor U11341 (N_11341,N_10870,N_10827);
xnor U11342 (N_11342,N_10983,N_10846);
or U11343 (N_11343,N_10906,N_10726);
or U11344 (N_11344,N_10754,N_10543);
xor U11345 (N_11345,N_10804,N_10596);
xnor U11346 (N_11346,N_10575,N_10627);
nand U11347 (N_11347,N_10534,N_10612);
nand U11348 (N_11348,N_10573,N_10786);
and U11349 (N_11349,N_10767,N_10540);
and U11350 (N_11350,N_10961,N_10706);
or U11351 (N_11351,N_10962,N_10856);
nand U11352 (N_11352,N_10533,N_10904);
nand U11353 (N_11353,N_10882,N_10953);
nand U11354 (N_11354,N_10728,N_10983);
and U11355 (N_11355,N_10981,N_10766);
xor U11356 (N_11356,N_10913,N_10979);
nand U11357 (N_11357,N_10860,N_10632);
and U11358 (N_11358,N_10593,N_10602);
nand U11359 (N_11359,N_10575,N_10775);
and U11360 (N_11360,N_10746,N_10523);
xnor U11361 (N_11361,N_10645,N_10750);
or U11362 (N_11362,N_10579,N_10967);
nand U11363 (N_11363,N_10547,N_10953);
xor U11364 (N_11364,N_10723,N_10604);
nand U11365 (N_11365,N_10972,N_10531);
and U11366 (N_11366,N_10599,N_10646);
and U11367 (N_11367,N_10720,N_10995);
or U11368 (N_11368,N_10813,N_10729);
nor U11369 (N_11369,N_10929,N_10876);
nand U11370 (N_11370,N_10779,N_10737);
xnor U11371 (N_11371,N_10596,N_10866);
or U11372 (N_11372,N_10807,N_10920);
nand U11373 (N_11373,N_10762,N_10636);
nand U11374 (N_11374,N_10906,N_10778);
or U11375 (N_11375,N_10819,N_10986);
and U11376 (N_11376,N_10891,N_10996);
and U11377 (N_11377,N_10741,N_10771);
and U11378 (N_11378,N_10813,N_10975);
or U11379 (N_11379,N_10930,N_10750);
nor U11380 (N_11380,N_10703,N_10651);
and U11381 (N_11381,N_10674,N_10779);
xor U11382 (N_11382,N_10535,N_10761);
or U11383 (N_11383,N_10518,N_10572);
xnor U11384 (N_11384,N_10874,N_10971);
nand U11385 (N_11385,N_10728,N_10740);
nor U11386 (N_11386,N_10537,N_10684);
nand U11387 (N_11387,N_10671,N_10787);
or U11388 (N_11388,N_10812,N_10938);
nand U11389 (N_11389,N_10938,N_10866);
nand U11390 (N_11390,N_10640,N_10785);
xor U11391 (N_11391,N_10849,N_10658);
nor U11392 (N_11392,N_10506,N_10720);
nand U11393 (N_11393,N_10587,N_10928);
nand U11394 (N_11394,N_10703,N_10888);
nor U11395 (N_11395,N_10780,N_10919);
and U11396 (N_11396,N_10680,N_10721);
xor U11397 (N_11397,N_10550,N_10618);
nor U11398 (N_11398,N_10898,N_10548);
nand U11399 (N_11399,N_10949,N_10914);
nor U11400 (N_11400,N_10935,N_10858);
nand U11401 (N_11401,N_10631,N_10561);
and U11402 (N_11402,N_10861,N_10529);
and U11403 (N_11403,N_10645,N_10632);
and U11404 (N_11404,N_10786,N_10828);
or U11405 (N_11405,N_10648,N_10731);
and U11406 (N_11406,N_10599,N_10532);
or U11407 (N_11407,N_10818,N_10669);
or U11408 (N_11408,N_10665,N_10624);
nand U11409 (N_11409,N_10682,N_10645);
nand U11410 (N_11410,N_10619,N_10759);
or U11411 (N_11411,N_10967,N_10552);
nor U11412 (N_11412,N_10699,N_10584);
and U11413 (N_11413,N_10953,N_10609);
or U11414 (N_11414,N_10610,N_10597);
or U11415 (N_11415,N_10965,N_10755);
nand U11416 (N_11416,N_10761,N_10675);
nand U11417 (N_11417,N_10650,N_10993);
or U11418 (N_11418,N_10670,N_10510);
or U11419 (N_11419,N_10722,N_10950);
nor U11420 (N_11420,N_10733,N_10711);
and U11421 (N_11421,N_10771,N_10542);
nand U11422 (N_11422,N_10900,N_10705);
xnor U11423 (N_11423,N_10601,N_10880);
nand U11424 (N_11424,N_10554,N_10640);
and U11425 (N_11425,N_10604,N_10607);
nor U11426 (N_11426,N_10638,N_10974);
xnor U11427 (N_11427,N_10983,N_10848);
nor U11428 (N_11428,N_10943,N_10770);
nor U11429 (N_11429,N_10913,N_10522);
nand U11430 (N_11430,N_10881,N_10515);
nor U11431 (N_11431,N_10901,N_10823);
or U11432 (N_11432,N_10696,N_10791);
nand U11433 (N_11433,N_10540,N_10661);
or U11434 (N_11434,N_10546,N_10538);
nor U11435 (N_11435,N_10609,N_10779);
xnor U11436 (N_11436,N_10922,N_10593);
or U11437 (N_11437,N_10910,N_10733);
and U11438 (N_11438,N_10679,N_10937);
and U11439 (N_11439,N_10531,N_10506);
and U11440 (N_11440,N_10773,N_10889);
or U11441 (N_11441,N_10949,N_10718);
nand U11442 (N_11442,N_10759,N_10966);
and U11443 (N_11443,N_10959,N_10801);
xnor U11444 (N_11444,N_10834,N_10851);
nor U11445 (N_11445,N_10839,N_10892);
xor U11446 (N_11446,N_10527,N_10704);
nor U11447 (N_11447,N_10590,N_10693);
nand U11448 (N_11448,N_10696,N_10525);
nor U11449 (N_11449,N_10615,N_10871);
xnor U11450 (N_11450,N_10594,N_10995);
or U11451 (N_11451,N_10912,N_10664);
nand U11452 (N_11452,N_10853,N_10860);
xor U11453 (N_11453,N_10560,N_10779);
nor U11454 (N_11454,N_10678,N_10628);
and U11455 (N_11455,N_10816,N_10736);
or U11456 (N_11456,N_10654,N_10577);
or U11457 (N_11457,N_10845,N_10526);
nor U11458 (N_11458,N_10712,N_10860);
or U11459 (N_11459,N_10629,N_10911);
or U11460 (N_11460,N_10850,N_10996);
and U11461 (N_11461,N_10566,N_10691);
nor U11462 (N_11462,N_10686,N_10719);
and U11463 (N_11463,N_10830,N_10523);
or U11464 (N_11464,N_10754,N_10863);
nand U11465 (N_11465,N_10690,N_10583);
xnor U11466 (N_11466,N_10839,N_10749);
and U11467 (N_11467,N_10534,N_10625);
nor U11468 (N_11468,N_10662,N_10882);
nand U11469 (N_11469,N_10694,N_10756);
and U11470 (N_11470,N_10634,N_10654);
nand U11471 (N_11471,N_10944,N_10658);
or U11472 (N_11472,N_10636,N_10864);
or U11473 (N_11473,N_10946,N_10979);
xor U11474 (N_11474,N_10752,N_10916);
or U11475 (N_11475,N_10645,N_10986);
or U11476 (N_11476,N_10691,N_10734);
nor U11477 (N_11477,N_10583,N_10764);
xnor U11478 (N_11478,N_10965,N_10619);
or U11479 (N_11479,N_10735,N_10972);
xnor U11480 (N_11480,N_10761,N_10993);
nor U11481 (N_11481,N_10794,N_10604);
nor U11482 (N_11482,N_10832,N_10602);
nand U11483 (N_11483,N_10900,N_10969);
or U11484 (N_11484,N_10778,N_10855);
nand U11485 (N_11485,N_10552,N_10920);
nand U11486 (N_11486,N_10605,N_10815);
nand U11487 (N_11487,N_10901,N_10995);
xnor U11488 (N_11488,N_10703,N_10570);
xnor U11489 (N_11489,N_10811,N_10594);
nand U11490 (N_11490,N_10564,N_10730);
or U11491 (N_11491,N_10902,N_10663);
nor U11492 (N_11492,N_10824,N_10835);
nand U11493 (N_11493,N_10872,N_10529);
or U11494 (N_11494,N_10602,N_10907);
and U11495 (N_11495,N_10611,N_10629);
nand U11496 (N_11496,N_10892,N_10874);
nor U11497 (N_11497,N_10503,N_10617);
nand U11498 (N_11498,N_10942,N_10898);
nand U11499 (N_11499,N_10566,N_10579);
nor U11500 (N_11500,N_11378,N_11022);
xor U11501 (N_11501,N_11205,N_11414);
nand U11502 (N_11502,N_11028,N_11270);
and U11503 (N_11503,N_11395,N_11450);
or U11504 (N_11504,N_11273,N_11260);
or U11505 (N_11505,N_11377,N_11372);
nand U11506 (N_11506,N_11451,N_11193);
and U11507 (N_11507,N_11335,N_11298);
nor U11508 (N_11508,N_11245,N_11485);
and U11509 (N_11509,N_11488,N_11139);
and U11510 (N_11510,N_11177,N_11452);
nand U11511 (N_11511,N_11444,N_11064);
xor U11512 (N_11512,N_11490,N_11351);
nand U11513 (N_11513,N_11122,N_11363);
or U11514 (N_11514,N_11459,N_11478);
or U11515 (N_11515,N_11076,N_11436);
xor U11516 (N_11516,N_11465,N_11180);
nand U11517 (N_11517,N_11396,N_11247);
nor U11518 (N_11518,N_11191,N_11067);
nor U11519 (N_11519,N_11101,N_11498);
and U11520 (N_11520,N_11116,N_11188);
nand U11521 (N_11521,N_11388,N_11127);
nand U11522 (N_11522,N_11142,N_11013);
xnor U11523 (N_11523,N_11220,N_11329);
nand U11524 (N_11524,N_11364,N_11054);
nor U11525 (N_11525,N_11340,N_11232);
or U11526 (N_11526,N_11401,N_11128);
nand U11527 (N_11527,N_11472,N_11442);
or U11528 (N_11528,N_11063,N_11283);
xnor U11529 (N_11529,N_11005,N_11321);
or U11530 (N_11530,N_11182,N_11299);
and U11531 (N_11531,N_11155,N_11084);
nand U11532 (N_11532,N_11447,N_11429);
nand U11533 (N_11533,N_11079,N_11412);
nor U11534 (N_11534,N_11337,N_11333);
nor U11535 (N_11535,N_11322,N_11303);
or U11536 (N_11536,N_11201,N_11249);
xor U11537 (N_11537,N_11132,N_11227);
or U11538 (N_11538,N_11104,N_11124);
and U11539 (N_11539,N_11456,N_11475);
nand U11540 (N_11540,N_11400,N_11460);
and U11541 (N_11541,N_11496,N_11292);
xnor U11542 (N_11542,N_11417,N_11163);
nor U11543 (N_11543,N_11256,N_11103);
nand U11544 (N_11544,N_11240,N_11257);
or U11545 (N_11545,N_11106,N_11462);
or U11546 (N_11546,N_11243,N_11194);
nor U11547 (N_11547,N_11092,N_11165);
and U11548 (N_11548,N_11466,N_11373);
xnor U11549 (N_11549,N_11031,N_11074);
xnor U11550 (N_11550,N_11131,N_11175);
and U11551 (N_11551,N_11278,N_11289);
nor U11552 (N_11552,N_11046,N_11050);
or U11553 (N_11553,N_11150,N_11157);
and U11554 (N_11554,N_11187,N_11294);
and U11555 (N_11555,N_11037,N_11441);
or U11556 (N_11556,N_11072,N_11136);
nand U11557 (N_11557,N_11241,N_11130);
or U11558 (N_11558,N_11371,N_11204);
and U11559 (N_11559,N_11448,N_11085);
and U11560 (N_11560,N_11374,N_11407);
nor U11561 (N_11561,N_11184,N_11439);
nor U11562 (N_11562,N_11423,N_11110);
and U11563 (N_11563,N_11481,N_11231);
nor U11564 (N_11564,N_11087,N_11471);
and U11565 (N_11565,N_11406,N_11222);
or U11566 (N_11566,N_11196,N_11387);
nor U11567 (N_11567,N_11168,N_11261);
nand U11568 (N_11568,N_11107,N_11347);
or U11569 (N_11569,N_11015,N_11237);
and U11570 (N_11570,N_11176,N_11129);
or U11571 (N_11571,N_11493,N_11334);
and U11572 (N_11572,N_11148,N_11234);
xor U11573 (N_11573,N_11034,N_11318);
nand U11574 (N_11574,N_11319,N_11411);
nor U11575 (N_11575,N_11291,N_11145);
nand U11576 (N_11576,N_11235,N_11152);
nand U11577 (N_11577,N_11223,N_11408);
nor U11578 (N_11578,N_11437,N_11086);
and U11579 (N_11579,N_11265,N_11454);
xnor U11580 (N_11580,N_11469,N_11003);
nand U11581 (N_11581,N_11305,N_11147);
nor U11582 (N_11582,N_11065,N_11166);
xnor U11583 (N_11583,N_11370,N_11416);
and U11584 (N_11584,N_11263,N_11413);
and U11585 (N_11585,N_11095,N_11361);
nand U11586 (N_11586,N_11380,N_11255);
or U11587 (N_11587,N_11440,N_11006);
nand U11588 (N_11588,N_11049,N_11008);
nor U11589 (N_11589,N_11487,N_11228);
and U11590 (N_11590,N_11403,N_11153);
xnor U11591 (N_11591,N_11059,N_11082);
xor U11592 (N_11592,N_11474,N_11113);
and U11593 (N_11593,N_11126,N_11286);
xnor U11594 (N_11594,N_11424,N_11057);
or U11595 (N_11595,N_11258,N_11202);
nor U11596 (N_11596,N_11445,N_11069);
xnor U11597 (N_11597,N_11355,N_11285);
or U11598 (N_11598,N_11405,N_11356);
xor U11599 (N_11599,N_11125,N_11239);
or U11600 (N_11600,N_11016,N_11038);
xnor U11601 (N_11601,N_11495,N_11393);
or U11602 (N_11602,N_11123,N_11404);
or U11603 (N_11603,N_11042,N_11078);
or U11604 (N_11604,N_11271,N_11089);
nand U11605 (N_11605,N_11217,N_11409);
xnor U11606 (N_11606,N_11183,N_11173);
or U11607 (N_11607,N_11272,N_11419);
nor U11608 (N_11608,N_11111,N_11207);
nand U11609 (N_11609,N_11225,N_11169);
nor U11610 (N_11610,N_11149,N_11345);
and U11611 (N_11611,N_11219,N_11327);
nor U11612 (N_11612,N_11362,N_11433);
or U11613 (N_11613,N_11002,N_11181);
xnor U11614 (N_11614,N_11199,N_11040);
and U11615 (N_11615,N_11309,N_11427);
and U11616 (N_11616,N_11117,N_11200);
or U11617 (N_11617,N_11338,N_11310);
or U11618 (N_11618,N_11317,N_11203);
nand U11619 (N_11619,N_11159,N_11178);
xnor U11620 (N_11620,N_11097,N_11246);
or U11621 (N_11621,N_11375,N_11218);
nand U11622 (N_11622,N_11236,N_11140);
nand U11623 (N_11623,N_11422,N_11012);
nand U11624 (N_11624,N_11009,N_11489);
or U11625 (N_11625,N_11281,N_11379);
nand U11626 (N_11626,N_11053,N_11385);
or U11627 (N_11627,N_11052,N_11021);
or U11628 (N_11628,N_11386,N_11011);
nor U11629 (N_11629,N_11277,N_11392);
nor U11630 (N_11630,N_11342,N_11398);
nand U11631 (N_11631,N_11114,N_11047);
nand U11632 (N_11632,N_11287,N_11151);
nor U11633 (N_11633,N_11029,N_11135);
xor U11634 (N_11634,N_11036,N_11343);
xnor U11635 (N_11635,N_11266,N_11100);
nor U11636 (N_11636,N_11426,N_11238);
nor U11637 (N_11637,N_11352,N_11119);
nand U11638 (N_11638,N_11192,N_11244);
and U11639 (N_11639,N_11384,N_11492);
xor U11640 (N_11640,N_11458,N_11430);
nand U11641 (N_11641,N_11102,N_11360);
nand U11642 (N_11642,N_11081,N_11455);
and U11643 (N_11643,N_11250,N_11453);
or U11644 (N_11644,N_11051,N_11144);
nor U11645 (N_11645,N_11376,N_11120);
nor U11646 (N_11646,N_11214,N_11105);
nor U11647 (N_11647,N_11499,N_11216);
or U11648 (N_11648,N_11328,N_11172);
and U11649 (N_11649,N_11279,N_11083);
xnor U11650 (N_11650,N_11369,N_11160);
xnor U11651 (N_11651,N_11033,N_11354);
nor U11652 (N_11652,N_11267,N_11336);
and U11653 (N_11653,N_11174,N_11094);
nor U11654 (N_11654,N_11491,N_11170);
nand U11655 (N_11655,N_11295,N_11007);
nand U11656 (N_11656,N_11262,N_11366);
xnor U11657 (N_11657,N_11195,N_11023);
nor U11658 (N_11658,N_11099,N_11320);
nor U11659 (N_11659,N_11325,N_11230);
and U11660 (N_11660,N_11397,N_11402);
or U11661 (N_11661,N_11061,N_11133);
xnor U11662 (N_11662,N_11324,N_11368);
nor U11663 (N_11663,N_11323,N_11226);
nor U11664 (N_11664,N_11461,N_11476);
or U11665 (N_11665,N_11004,N_11014);
and U11666 (N_11666,N_11020,N_11483);
and U11667 (N_11667,N_11457,N_11293);
nand U11668 (N_11668,N_11330,N_11350);
or U11669 (N_11669,N_11039,N_11041);
nor U11670 (N_11670,N_11365,N_11269);
nand U11671 (N_11671,N_11066,N_11058);
nor U11672 (N_11672,N_11391,N_11121);
and U11673 (N_11673,N_11399,N_11000);
nor U11674 (N_11674,N_11443,N_11449);
xnor U11675 (N_11675,N_11045,N_11274);
nor U11676 (N_11676,N_11068,N_11096);
nand U11677 (N_11677,N_11486,N_11302);
nor U11678 (N_11678,N_11154,N_11221);
nor U11679 (N_11679,N_11035,N_11118);
nand U11680 (N_11680,N_11332,N_11307);
and U11681 (N_11681,N_11311,N_11143);
nand U11682 (N_11682,N_11410,N_11482);
or U11683 (N_11683,N_11316,N_11186);
or U11684 (N_11684,N_11389,N_11315);
nand U11685 (N_11685,N_11190,N_11115);
nor U11686 (N_11686,N_11428,N_11314);
and U11687 (N_11687,N_11357,N_11434);
nor U11688 (N_11688,N_11473,N_11060);
nand U11689 (N_11689,N_11027,N_11189);
and U11690 (N_11690,N_11141,N_11259);
xor U11691 (N_11691,N_11358,N_11432);
nor U11692 (N_11692,N_11167,N_11497);
nor U11693 (N_11693,N_11044,N_11206);
nand U11694 (N_11694,N_11349,N_11224);
or U11695 (N_11695,N_11019,N_11229);
xor U11696 (N_11696,N_11251,N_11137);
nor U11697 (N_11697,N_11339,N_11138);
or U11698 (N_11698,N_11344,N_11326);
nor U11699 (N_11699,N_11017,N_11026);
or U11700 (N_11700,N_11030,N_11435);
nand U11701 (N_11701,N_11070,N_11276);
nand U11702 (N_11702,N_11197,N_11264);
nor U11703 (N_11703,N_11112,N_11468);
xnor U11704 (N_11704,N_11282,N_11073);
nor U11705 (N_11705,N_11179,N_11248);
xor U11706 (N_11706,N_11394,N_11080);
nand U11707 (N_11707,N_11098,N_11341);
nor U11708 (N_11708,N_11438,N_11348);
xnor U11709 (N_11709,N_11484,N_11018);
xor U11710 (N_11710,N_11093,N_11109);
or U11711 (N_11711,N_11024,N_11209);
xor U11712 (N_11712,N_11390,N_11381);
xnor U11713 (N_11713,N_11463,N_11383);
or U11714 (N_11714,N_11171,N_11043);
xnor U11715 (N_11715,N_11161,N_11331);
nor U11716 (N_11716,N_11075,N_11090);
or U11717 (N_11717,N_11480,N_11284);
and U11718 (N_11718,N_11467,N_11425);
nand U11719 (N_11719,N_11048,N_11359);
or U11720 (N_11720,N_11268,N_11242);
xor U11721 (N_11721,N_11306,N_11208);
nand U11722 (N_11722,N_11494,N_11477);
or U11723 (N_11723,N_11062,N_11290);
nor U11724 (N_11724,N_11108,N_11211);
and U11725 (N_11725,N_11156,N_11312);
and U11726 (N_11726,N_11446,N_11353);
nand U11727 (N_11727,N_11297,N_11252);
or U11728 (N_11728,N_11308,N_11313);
or U11729 (N_11729,N_11091,N_11146);
nand U11730 (N_11730,N_11056,N_11134);
nand U11731 (N_11731,N_11032,N_11215);
and U11732 (N_11732,N_11479,N_11280);
or U11733 (N_11733,N_11288,N_11010);
nand U11734 (N_11734,N_11421,N_11420);
nor U11735 (N_11735,N_11071,N_11382);
nor U11736 (N_11736,N_11164,N_11088);
or U11737 (N_11737,N_11346,N_11254);
nor U11738 (N_11738,N_11233,N_11213);
xnor U11739 (N_11739,N_11055,N_11212);
or U11740 (N_11740,N_11077,N_11415);
and U11741 (N_11741,N_11464,N_11162);
nor U11742 (N_11742,N_11301,N_11210);
nand U11743 (N_11743,N_11304,N_11253);
and U11744 (N_11744,N_11001,N_11025);
or U11745 (N_11745,N_11185,N_11158);
xor U11746 (N_11746,N_11367,N_11300);
nor U11747 (N_11747,N_11198,N_11470);
or U11748 (N_11748,N_11296,N_11418);
and U11749 (N_11749,N_11431,N_11275);
nand U11750 (N_11750,N_11119,N_11383);
nor U11751 (N_11751,N_11422,N_11148);
and U11752 (N_11752,N_11408,N_11196);
or U11753 (N_11753,N_11468,N_11060);
and U11754 (N_11754,N_11124,N_11384);
nand U11755 (N_11755,N_11449,N_11059);
xnor U11756 (N_11756,N_11076,N_11366);
nor U11757 (N_11757,N_11365,N_11427);
xor U11758 (N_11758,N_11397,N_11166);
nand U11759 (N_11759,N_11018,N_11373);
or U11760 (N_11760,N_11309,N_11070);
or U11761 (N_11761,N_11378,N_11310);
or U11762 (N_11762,N_11412,N_11366);
nor U11763 (N_11763,N_11180,N_11060);
and U11764 (N_11764,N_11429,N_11093);
nor U11765 (N_11765,N_11005,N_11141);
xor U11766 (N_11766,N_11478,N_11352);
nand U11767 (N_11767,N_11459,N_11258);
nor U11768 (N_11768,N_11047,N_11215);
or U11769 (N_11769,N_11004,N_11110);
nor U11770 (N_11770,N_11406,N_11445);
xnor U11771 (N_11771,N_11408,N_11130);
or U11772 (N_11772,N_11456,N_11025);
or U11773 (N_11773,N_11461,N_11125);
nor U11774 (N_11774,N_11011,N_11003);
or U11775 (N_11775,N_11491,N_11370);
nand U11776 (N_11776,N_11130,N_11058);
xor U11777 (N_11777,N_11028,N_11085);
and U11778 (N_11778,N_11242,N_11125);
nor U11779 (N_11779,N_11421,N_11067);
nand U11780 (N_11780,N_11034,N_11202);
nand U11781 (N_11781,N_11100,N_11080);
nor U11782 (N_11782,N_11012,N_11308);
xor U11783 (N_11783,N_11127,N_11159);
and U11784 (N_11784,N_11494,N_11146);
xor U11785 (N_11785,N_11363,N_11338);
and U11786 (N_11786,N_11015,N_11050);
nor U11787 (N_11787,N_11482,N_11287);
xnor U11788 (N_11788,N_11036,N_11025);
xor U11789 (N_11789,N_11087,N_11314);
xor U11790 (N_11790,N_11492,N_11447);
xor U11791 (N_11791,N_11151,N_11449);
and U11792 (N_11792,N_11021,N_11406);
xor U11793 (N_11793,N_11294,N_11147);
xnor U11794 (N_11794,N_11389,N_11108);
nand U11795 (N_11795,N_11296,N_11129);
and U11796 (N_11796,N_11372,N_11301);
xnor U11797 (N_11797,N_11446,N_11094);
xnor U11798 (N_11798,N_11208,N_11494);
and U11799 (N_11799,N_11058,N_11294);
and U11800 (N_11800,N_11011,N_11457);
nor U11801 (N_11801,N_11375,N_11062);
nor U11802 (N_11802,N_11411,N_11477);
and U11803 (N_11803,N_11104,N_11290);
xor U11804 (N_11804,N_11016,N_11271);
or U11805 (N_11805,N_11289,N_11185);
or U11806 (N_11806,N_11195,N_11132);
and U11807 (N_11807,N_11277,N_11080);
xnor U11808 (N_11808,N_11390,N_11048);
nand U11809 (N_11809,N_11354,N_11491);
xor U11810 (N_11810,N_11386,N_11175);
nand U11811 (N_11811,N_11179,N_11387);
xnor U11812 (N_11812,N_11480,N_11307);
or U11813 (N_11813,N_11021,N_11151);
and U11814 (N_11814,N_11223,N_11390);
and U11815 (N_11815,N_11036,N_11207);
nor U11816 (N_11816,N_11059,N_11300);
or U11817 (N_11817,N_11424,N_11355);
and U11818 (N_11818,N_11489,N_11250);
and U11819 (N_11819,N_11055,N_11149);
xnor U11820 (N_11820,N_11455,N_11129);
nor U11821 (N_11821,N_11174,N_11260);
xnor U11822 (N_11822,N_11186,N_11081);
nand U11823 (N_11823,N_11146,N_11194);
and U11824 (N_11824,N_11283,N_11092);
and U11825 (N_11825,N_11467,N_11274);
nand U11826 (N_11826,N_11416,N_11386);
nand U11827 (N_11827,N_11392,N_11365);
nand U11828 (N_11828,N_11008,N_11248);
or U11829 (N_11829,N_11398,N_11200);
nand U11830 (N_11830,N_11215,N_11204);
or U11831 (N_11831,N_11466,N_11125);
and U11832 (N_11832,N_11312,N_11277);
and U11833 (N_11833,N_11373,N_11383);
or U11834 (N_11834,N_11012,N_11168);
xor U11835 (N_11835,N_11145,N_11347);
or U11836 (N_11836,N_11425,N_11416);
nand U11837 (N_11837,N_11481,N_11445);
and U11838 (N_11838,N_11409,N_11122);
nand U11839 (N_11839,N_11465,N_11423);
or U11840 (N_11840,N_11132,N_11364);
xor U11841 (N_11841,N_11291,N_11283);
xnor U11842 (N_11842,N_11137,N_11362);
xor U11843 (N_11843,N_11263,N_11226);
nor U11844 (N_11844,N_11379,N_11015);
or U11845 (N_11845,N_11251,N_11087);
or U11846 (N_11846,N_11033,N_11308);
nor U11847 (N_11847,N_11408,N_11160);
nand U11848 (N_11848,N_11175,N_11033);
xnor U11849 (N_11849,N_11027,N_11415);
nand U11850 (N_11850,N_11259,N_11064);
or U11851 (N_11851,N_11247,N_11496);
nor U11852 (N_11852,N_11428,N_11480);
and U11853 (N_11853,N_11024,N_11159);
or U11854 (N_11854,N_11496,N_11175);
xor U11855 (N_11855,N_11480,N_11455);
or U11856 (N_11856,N_11395,N_11054);
nand U11857 (N_11857,N_11086,N_11012);
or U11858 (N_11858,N_11064,N_11258);
nand U11859 (N_11859,N_11294,N_11287);
or U11860 (N_11860,N_11299,N_11376);
nand U11861 (N_11861,N_11392,N_11333);
and U11862 (N_11862,N_11243,N_11138);
xor U11863 (N_11863,N_11107,N_11186);
nor U11864 (N_11864,N_11416,N_11360);
xor U11865 (N_11865,N_11485,N_11106);
xor U11866 (N_11866,N_11031,N_11418);
nor U11867 (N_11867,N_11401,N_11383);
nand U11868 (N_11868,N_11246,N_11325);
or U11869 (N_11869,N_11066,N_11327);
nand U11870 (N_11870,N_11233,N_11021);
xnor U11871 (N_11871,N_11025,N_11165);
and U11872 (N_11872,N_11076,N_11305);
xor U11873 (N_11873,N_11101,N_11135);
nand U11874 (N_11874,N_11330,N_11267);
nor U11875 (N_11875,N_11126,N_11203);
nor U11876 (N_11876,N_11480,N_11154);
nand U11877 (N_11877,N_11422,N_11178);
nor U11878 (N_11878,N_11091,N_11003);
or U11879 (N_11879,N_11444,N_11359);
or U11880 (N_11880,N_11333,N_11301);
xnor U11881 (N_11881,N_11279,N_11149);
nand U11882 (N_11882,N_11292,N_11397);
nor U11883 (N_11883,N_11186,N_11434);
nand U11884 (N_11884,N_11332,N_11082);
nand U11885 (N_11885,N_11019,N_11337);
nand U11886 (N_11886,N_11235,N_11069);
or U11887 (N_11887,N_11431,N_11340);
xnor U11888 (N_11888,N_11439,N_11218);
nand U11889 (N_11889,N_11188,N_11135);
xor U11890 (N_11890,N_11384,N_11334);
and U11891 (N_11891,N_11198,N_11365);
nand U11892 (N_11892,N_11277,N_11354);
and U11893 (N_11893,N_11480,N_11412);
nand U11894 (N_11894,N_11296,N_11057);
nor U11895 (N_11895,N_11170,N_11292);
and U11896 (N_11896,N_11468,N_11274);
and U11897 (N_11897,N_11434,N_11177);
nand U11898 (N_11898,N_11490,N_11064);
nand U11899 (N_11899,N_11045,N_11035);
or U11900 (N_11900,N_11214,N_11179);
and U11901 (N_11901,N_11131,N_11031);
and U11902 (N_11902,N_11431,N_11188);
nor U11903 (N_11903,N_11093,N_11069);
xor U11904 (N_11904,N_11005,N_11167);
and U11905 (N_11905,N_11438,N_11473);
nand U11906 (N_11906,N_11395,N_11223);
and U11907 (N_11907,N_11374,N_11441);
xor U11908 (N_11908,N_11364,N_11168);
nor U11909 (N_11909,N_11487,N_11360);
and U11910 (N_11910,N_11191,N_11254);
xor U11911 (N_11911,N_11268,N_11483);
nor U11912 (N_11912,N_11282,N_11348);
xor U11913 (N_11913,N_11152,N_11009);
and U11914 (N_11914,N_11391,N_11202);
xor U11915 (N_11915,N_11418,N_11012);
nand U11916 (N_11916,N_11457,N_11355);
xnor U11917 (N_11917,N_11276,N_11232);
nor U11918 (N_11918,N_11368,N_11421);
and U11919 (N_11919,N_11317,N_11196);
nor U11920 (N_11920,N_11385,N_11007);
nor U11921 (N_11921,N_11272,N_11181);
nand U11922 (N_11922,N_11163,N_11202);
and U11923 (N_11923,N_11104,N_11146);
or U11924 (N_11924,N_11397,N_11168);
or U11925 (N_11925,N_11170,N_11497);
nand U11926 (N_11926,N_11193,N_11072);
and U11927 (N_11927,N_11093,N_11387);
nor U11928 (N_11928,N_11322,N_11422);
xor U11929 (N_11929,N_11451,N_11197);
nand U11930 (N_11930,N_11146,N_11203);
nand U11931 (N_11931,N_11165,N_11480);
or U11932 (N_11932,N_11161,N_11052);
or U11933 (N_11933,N_11200,N_11144);
and U11934 (N_11934,N_11138,N_11470);
or U11935 (N_11935,N_11476,N_11301);
nand U11936 (N_11936,N_11130,N_11013);
xor U11937 (N_11937,N_11051,N_11139);
nand U11938 (N_11938,N_11302,N_11077);
nand U11939 (N_11939,N_11120,N_11388);
nand U11940 (N_11940,N_11148,N_11002);
nor U11941 (N_11941,N_11425,N_11451);
nor U11942 (N_11942,N_11336,N_11090);
xor U11943 (N_11943,N_11374,N_11249);
nor U11944 (N_11944,N_11342,N_11106);
or U11945 (N_11945,N_11261,N_11220);
or U11946 (N_11946,N_11499,N_11106);
nand U11947 (N_11947,N_11085,N_11187);
nand U11948 (N_11948,N_11213,N_11459);
nand U11949 (N_11949,N_11041,N_11174);
or U11950 (N_11950,N_11125,N_11065);
and U11951 (N_11951,N_11440,N_11022);
nand U11952 (N_11952,N_11414,N_11236);
xor U11953 (N_11953,N_11364,N_11176);
xnor U11954 (N_11954,N_11218,N_11067);
and U11955 (N_11955,N_11168,N_11150);
nor U11956 (N_11956,N_11301,N_11027);
and U11957 (N_11957,N_11394,N_11214);
xnor U11958 (N_11958,N_11317,N_11239);
xor U11959 (N_11959,N_11017,N_11152);
nand U11960 (N_11960,N_11318,N_11457);
nor U11961 (N_11961,N_11455,N_11366);
or U11962 (N_11962,N_11368,N_11099);
or U11963 (N_11963,N_11103,N_11324);
or U11964 (N_11964,N_11406,N_11486);
and U11965 (N_11965,N_11086,N_11319);
xnor U11966 (N_11966,N_11135,N_11042);
nor U11967 (N_11967,N_11193,N_11447);
and U11968 (N_11968,N_11348,N_11147);
nor U11969 (N_11969,N_11405,N_11180);
and U11970 (N_11970,N_11083,N_11077);
or U11971 (N_11971,N_11321,N_11044);
and U11972 (N_11972,N_11089,N_11486);
nor U11973 (N_11973,N_11465,N_11260);
or U11974 (N_11974,N_11337,N_11304);
nand U11975 (N_11975,N_11013,N_11201);
nand U11976 (N_11976,N_11043,N_11062);
nand U11977 (N_11977,N_11062,N_11250);
nand U11978 (N_11978,N_11027,N_11010);
nor U11979 (N_11979,N_11271,N_11005);
and U11980 (N_11980,N_11330,N_11102);
nand U11981 (N_11981,N_11233,N_11292);
or U11982 (N_11982,N_11405,N_11053);
nor U11983 (N_11983,N_11237,N_11123);
nand U11984 (N_11984,N_11434,N_11199);
and U11985 (N_11985,N_11056,N_11054);
or U11986 (N_11986,N_11325,N_11475);
nor U11987 (N_11987,N_11310,N_11259);
or U11988 (N_11988,N_11140,N_11052);
and U11989 (N_11989,N_11423,N_11072);
or U11990 (N_11990,N_11125,N_11395);
and U11991 (N_11991,N_11306,N_11043);
xnor U11992 (N_11992,N_11122,N_11432);
or U11993 (N_11993,N_11025,N_11494);
and U11994 (N_11994,N_11222,N_11374);
xnor U11995 (N_11995,N_11332,N_11134);
xor U11996 (N_11996,N_11279,N_11232);
or U11997 (N_11997,N_11134,N_11036);
nand U11998 (N_11998,N_11413,N_11124);
or U11999 (N_11999,N_11350,N_11123);
nor U12000 (N_12000,N_11549,N_11961);
nand U12001 (N_12001,N_11616,N_11563);
nand U12002 (N_12002,N_11707,N_11558);
nor U12003 (N_12003,N_11648,N_11790);
nor U12004 (N_12004,N_11710,N_11685);
nand U12005 (N_12005,N_11939,N_11583);
and U12006 (N_12006,N_11829,N_11721);
or U12007 (N_12007,N_11669,N_11723);
or U12008 (N_12008,N_11573,N_11565);
xnor U12009 (N_12009,N_11856,N_11993);
and U12010 (N_12010,N_11955,N_11525);
and U12011 (N_12011,N_11699,N_11883);
or U12012 (N_12012,N_11854,N_11657);
and U12013 (N_12013,N_11546,N_11950);
and U12014 (N_12014,N_11968,N_11996);
xor U12015 (N_12015,N_11954,N_11914);
xnor U12016 (N_12016,N_11832,N_11841);
xnor U12017 (N_12017,N_11767,N_11755);
nand U12018 (N_12018,N_11526,N_11766);
or U12019 (N_12019,N_11609,N_11527);
or U12020 (N_12020,N_11973,N_11646);
and U12021 (N_12021,N_11948,N_11636);
nand U12022 (N_12022,N_11849,N_11506);
or U12023 (N_12023,N_11888,N_11679);
and U12024 (N_12024,N_11754,N_11663);
xnor U12025 (N_12025,N_11581,N_11629);
nand U12026 (N_12026,N_11960,N_11524);
or U12027 (N_12027,N_11726,N_11643);
or U12028 (N_12028,N_11659,N_11964);
or U12029 (N_12029,N_11789,N_11575);
nor U12030 (N_12030,N_11981,N_11942);
and U12031 (N_12031,N_11979,N_11574);
or U12032 (N_12032,N_11998,N_11514);
or U12033 (N_12033,N_11800,N_11706);
nor U12034 (N_12034,N_11953,N_11803);
or U12035 (N_12035,N_11830,N_11610);
xnor U12036 (N_12036,N_11631,N_11694);
nand U12037 (N_12037,N_11802,N_11984);
and U12038 (N_12038,N_11559,N_11896);
and U12039 (N_12039,N_11768,N_11686);
nor U12040 (N_12040,N_11840,N_11658);
and U12041 (N_12041,N_11744,N_11889);
nand U12042 (N_12042,N_11827,N_11536);
and U12043 (N_12043,N_11639,N_11617);
nor U12044 (N_12044,N_11667,N_11569);
xnor U12045 (N_12045,N_11600,N_11628);
nand U12046 (N_12046,N_11893,N_11831);
nand U12047 (N_12047,N_11518,N_11963);
nor U12048 (N_12048,N_11891,N_11731);
nand U12049 (N_12049,N_11930,N_11861);
nand U12050 (N_12050,N_11995,N_11627);
nor U12051 (N_12051,N_11638,N_11670);
or U12052 (N_12052,N_11588,N_11582);
xnor U12053 (N_12053,N_11622,N_11823);
nor U12054 (N_12054,N_11900,N_11985);
nand U12055 (N_12055,N_11735,N_11912);
xor U12056 (N_12056,N_11999,N_11791);
and U12057 (N_12057,N_11738,N_11796);
and U12058 (N_12058,N_11875,N_11931);
nand U12059 (N_12059,N_11966,N_11668);
nor U12060 (N_12060,N_11647,N_11806);
xor U12061 (N_12061,N_11903,N_11894);
nor U12062 (N_12062,N_11971,N_11556);
and U12063 (N_12063,N_11925,N_11517);
nand U12064 (N_12064,N_11509,N_11906);
nand U12065 (N_12065,N_11613,N_11828);
or U12066 (N_12066,N_11705,N_11808);
nor U12067 (N_12067,N_11879,N_11634);
or U12068 (N_12068,N_11936,N_11701);
or U12069 (N_12069,N_11732,N_11741);
or U12070 (N_12070,N_11562,N_11605);
nand U12071 (N_12071,N_11538,N_11714);
nor U12072 (N_12072,N_11910,N_11580);
nor U12073 (N_12073,N_11994,N_11683);
nor U12074 (N_12074,N_11990,N_11528);
nand U12075 (N_12075,N_11771,N_11779);
nand U12076 (N_12076,N_11774,N_11920);
or U12077 (N_12077,N_11750,N_11834);
nand U12078 (N_12078,N_11867,N_11797);
xnor U12079 (N_12079,N_11807,N_11594);
and U12080 (N_12080,N_11623,N_11678);
nor U12081 (N_12081,N_11899,N_11974);
nor U12082 (N_12082,N_11632,N_11637);
and U12083 (N_12083,N_11544,N_11591);
nand U12084 (N_12084,N_11897,N_11868);
and U12085 (N_12085,N_11795,N_11916);
nor U12086 (N_12086,N_11871,N_11817);
nand U12087 (N_12087,N_11599,N_11652);
and U12088 (N_12088,N_11501,N_11872);
nand U12089 (N_12089,N_11579,N_11585);
xor U12090 (N_12090,N_11842,N_11703);
or U12091 (N_12091,N_11760,N_11748);
and U12092 (N_12092,N_11641,N_11805);
xnor U12093 (N_12093,N_11598,N_11568);
xnor U12094 (N_12094,N_11590,N_11650);
nand U12095 (N_12095,N_11855,N_11870);
nand U12096 (N_12096,N_11813,N_11727);
and U12097 (N_12097,N_11933,N_11552);
nand U12098 (N_12098,N_11662,N_11940);
or U12099 (N_12099,N_11988,N_11725);
nor U12100 (N_12100,N_11844,N_11786);
and U12101 (N_12101,N_11740,N_11548);
xnor U12102 (N_12102,N_11826,N_11711);
and U12103 (N_12103,N_11708,N_11895);
nor U12104 (N_12104,N_11747,N_11520);
nand U12105 (N_12105,N_11851,N_11787);
and U12106 (N_12106,N_11737,N_11991);
and U12107 (N_12107,N_11783,N_11713);
xor U12108 (N_12108,N_11927,N_11530);
or U12109 (N_12109,N_11722,N_11926);
and U12110 (N_12110,N_11957,N_11773);
and U12111 (N_12111,N_11908,N_11655);
or U12112 (N_12112,N_11507,N_11976);
or U12113 (N_12113,N_11719,N_11642);
or U12114 (N_12114,N_11845,N_11715);
and U12115 (N_12115,N_11540,N_11775);
nor U12116 (N_12116,N_11918,N_11688);
nor U12117 (N_12117,N_11572,N_11929);
xor U12118 (N_12118,N_11718,N_11566);
or U12119 (N_12119,N_11794,N_11664);
and U12120 (N_12120,N_11809,N_11630);
and U12121 (N_12121,N_11839,N_11736);
or U12122 (N_12122,N_11874,N_11547);
xor U12123 (N_12123,N_11983,N_11850);
and U12124 (N_12124,N_11923,N_11989);
and U12125 (N_12125,N_11537,N_11612);
nand U12126 (N_12126,N_11919,N_11550);
xnor U12127 (N_12127,N_11947,N_11611);
or U12128 (N_12128,N_11969,N_11941);
nor U12129 (N_12129,N_11877,N_11656);
and U12130 (N_12130,N_11607,N_11762);
xor U12131 (N_12131,N_11586,N_11784);
nand U12132 (N_12132,N_11788,N_11907);
xor U12133 (N_12133,N_11557,N_11804);
nand U12134 (N_12134,N_11970,N_11621);
nor U12135 (N_12135,N_11858,N_11700);
xor U12136 (N_12136,N_11626,N_11661);
nand U12137 (N_12137,N_11570,N_11502);
or U12138 (N_12138,N_11618,N_11846);
nand U12139 (N_12139,N_11752,N_11690);
nand U12140 (N_12140,N_11676,N_11578);
or U12141 (N_12141,N_11510,N_11902);
nand U12142 (N_12142,N_11682,N_11560);
and U12143 (N_12143,N_11982,N_11772);
and U12144 (N_12144,N_11959,N_11620);
nor U12145 (N_12145,N_11958,N_11597);
xnor U12146 (N_12146,N_11887,N_11943);
and U12147 (N_12147,N_11977,N_11869);
and U12148 (N_12148,N_11848,N_11539);
and U12149 (N_12149,N_11666,N_11965);
xor U12150 (N_12150,N_11697,N_11522);
and U12151 (N_12151,N_11757,N_11519);
nor U12152 (N_12152,N_11833,N_11730);
xnor U12153 (N_12153,N_11535,N_11733);
or U12154 (N_12154,N_11820,N_11674);
or U12155 (N_12155,N_11975,N_11531);
and U12156 (N_12156,N_11751,N_11533);
or U12157 (N_12157,N_11904,N_11500);
or U12158 (N_12158,N_11951,N_11884);
and U12159 (N_12159,N_11799,N_11793);
xnor U12160 (N_12160,N_11952,N_11724);
or U12161 (N_12161,N_11753,N_11821);
nor U12162 (N_12162,N_11614,N_11709);
or U12163 (N_12163,N_11944,N_11625);
and U12164 (N_12164,N_11689,N_11759);
xor U12165 (N_12165,N_11997,N_11921);
nor U12166 (N_12166,N_11935,N_11693);
nor U12167 (N_12167,N_11601,N_11635);
xnor U12168 (N_12168,N_11967,N_11515);
or U12169 (N_12169,N_11822,N_11672);
or U12170 (N_12170,N_11847,N_11913);
xnor U12171 (N_12171,N_11778,N_11764);
and U12172 (N_12172,N_11541,N_11956);
nor U12173 (N_12173,N_11843,N_11878);
xor U12174 (N_12174,N_11838,N_11862);
nor U12175 (N_12175,N_11645,N_11593);
xnor U12176 (N_12176,N_11742,N_11521);
xnor U12177 (N_12177,N_11649,N_11513);
xnor U12178 (N_12178,N_11729,N_11567);
and U12179 (N_12179,N_11619,N_11587);
and U12180 (N_12180,N_11825,N_11886);
or U12181 (N_12181,N_11924,N_11746);
and U12182 (N_12182,N_11835,N_11633);
or U12183 (N_12183,N_11863,N_11584);
or U12184 (N_12184,N_11534,N_11545);
nor U12185 (N_12185,N_11511,N_11695);
nand U12186 (N_12186,N_11798,N_11712);
or U12187 (N_12187,N_11812,N_11553);
nand U12188 (N_12188,N_11922,N_11592);
and U12189 (N_12189,N_11720,N_11523);
xnor U12190 (N_12190,N_11882,N_11651);
and U12191 (N_12191,N_11728,N_11819);
xnor U12192 (N_12192,N_11743,N_11564);
nand U12193 (N_12193,N_11980,N_11785);
nor U12194 (N_12194,N_11665,N_11691);
or U12195 (N_12195,N_11640,N_11576);
and U12196 (N_12196,N_11692,N_11529);
nand U12197 (N_12197,N_11769,N_11684);
nor U12198 (N_12198,N_11836,N_11765);
nand U12199 (N_12199,N_11716,N_11704);
nor U12200 (N_12200,N_11905,N_11532);
and U12201 (N_12201,N_11503,N_11859);
xor U12202 (N_12202,N_11880,N_11873);
nand U12203 (N_12203,N_11675,N_11780);
and U12204 (N_12204,N_11987,N_11654);
nor U12205 (N_12205,N_11946,N_11653);
and U12206 (N_12206,N_11595,N_11673);
nor U12207 (N_12207,N_11660,N_11949);
or U12208 (N_12208,N_11677,N_11776);
nand U12209 (N_12209,N_11561,N_11758);
and U12210 (N_12210,N_11671,N_11551);
nand U12211 (N_12211,N_11938,N_11763);
and U12212 (N_12212,N_11978,N_11554);
xor U12213 (N_12213,N_11745,N_11749);
nor U12214 (N_12214,N_11892,N_11898);
nand U12215 (N_12215,N_11865,N_11603);
xnor U12216 (N_12216,N_11698,N_11508);
or U12217 (N_12217,N_11624,N_11986);
and U12218 (N_12218,N_11577,N_11687);
nand U12219 (N_12219,N_11937,N_11680);
and U12220 (N_12220,N_11909,N_11860);
xnor U12221 (N_12221,N_11885,N_11818);
nor U12222 (N_12222,N_11571,N_11702);
xor U12223 (N_12223,N_11604,N_11696);
nor U12224 (N_12224,N_11901,N_11615);
nor U12225 (N_12225,N_11837,N_11857);
nand U12226 (N_12226,N_11644,N_11516);
and U12227 (N_12227,N_11934,N_11717);
nor U12228 (N_12228,N_11890,N_11917);
or U12229 (N_12229,N_11852,N_11734);
xnor U12230 (N_12230,N_11816,N_11543);
and U12231 (N_12231,N_11815,N_11866);
and U12232 (N_12232,N_11810,N_11915);
xor U12233 (N_12233,N_11824,N_11876);
or U12234 (N_12234,N_11811,N_11555);
xnor U12235 (N_12235,N_11512,N_11608);
nand U12236 (N_12236,N_11739,N_11881);
nand U12237 (N_12237,N_11589,N_11756);
and U12238 (N_12238,N_11761,N_11853);
nor U12239 (N_12239,N_11781,N_11864);
xnor U12240 (N_12240,N_11928,N_11606);
and U12241 (N_12241,N_11770,N_11596);
nand U12242 (N_12242,N_11911,N_11542);
nand U12243 (N_12243,N_11945,N_11932);
nand U12244 (N_12244,N_11814,N_11504);
nand U12245 (N_12245,N_11505,N_11962);
xnor U12246 (N_12246,N_11681,N_11992);
and U12247 (N_12247,N_11792,N_11801);
or U12248 (N_12248,N_11972,N_11602);
nand U12249 (N_12249,N_11782,N_11777);
and U12250 (N_12250,N_11816,N_11931);
or U12251 (N_12251,N_11709,N_11704);
nand U12252 (N_12252,N_11502,N_11671);
xor U12253 (N_12253,N_11570,N_11690);
nor U12254 (N_12254,N_11938,N_11954);
and U12255 (N_12255,N_11814,N_11940);
xor U12256 (N_12256,N_11915,N_11512);
nand U12257 (N_12257,N_11610,N_11626);
and U12258 (N_12258,N_11722,N_11607);
or U12259 (N_12259,N_11855,N_11979);
nor U12260 (N_12260,N_11575,N_11724);
and U12261 (N_12261,N_11946,N_11521);
and U12262 (N_12262,N_11540,N_11617);
and U12263 (N_12263,N_11999,N_11526);
nor U12264 (N_12264,N_11953,N_11849);
or U12265 (N_12265,N_11966,N_11728);
nand U12266 (N_12266,N_11826,N_11861);
and U12267 (N_12267,N_11624,N_11633);
nor U12268 (N_12268,N_11526,N_11543);
nand U12269 (N_12269,N_11826,N_11886);
nand U12270 (N_12270,N_11573,N_11586);
nor U12271 (N_12271,N_11897,N_11569);
and U12272 (N_12272,N_11707,N_11695);
nand U12273 (N_12273,N_11994,N_11702);
xor U12274 (N_12274,N_11631,N_11638);
and U12275 (N_12275,N_11586,N_11550);
and U12276 (N_12276,N_11635,N_11803);
or U12277 (N_12277,N_11879,N_11655);
or U12278 (N_12278,N_11877,N_11989);
and U12279 (N_12279,N_11579,N_11613);
and U12280 (N_12280,N_11750,N_11699);
and U12281 (N_12281,N_11730,N_11639);
nand U12282 (N_12282,N_11994,N_11849);
nand U12283 (N_12283,N_11939,N_11515);
xor U12284 (N_12284,N_11960,N_11933);
nand U12285 (N_12285,N_11537,N_11954);
or U12286 (N_12286,N_11538,N_11652);
xor U12287 (N_12287,N_11724,N_11859);
xnor U12288 (N_12288,N_11584,N_11779);
xor U12289 (N_12289,N_11681,N_11603);
or U12290 (N_12290,N_11925,N_11694);
nor U12291 (N_12291,N_11745,N_11799);
xnor U12292 (N_12292,N_11515,N_11738);
or U12293 (N_12293,N_11950,N_11715);
nor U12294 (N_12294,N_11873,N_11805);
and U12295 (N_12295,N_11935,N_11960);
xnor U12296 (N_12296,N_11687,N_11791);
nor U12297 (N_12297,N_11982,N_11606);
xnor U12298 (N_12298,N_11837,N_11560);
or U12299 (N_12299,N_11644,N_11840);
and U12300 (N_12300,N_11569,N_11528);
nand U12301 (N_12301,N_11565,N_11589);
and U12302 (N_12302,N_11820,N_11675);
nand U12303 (N_12303,N_11751,N_11986);
xor U12304 (N_12304,N_11522,N_11520);
xnor U12305 (N_12305,N_11931,N_11708);
xnor U12306 (N_12306,N_11615,N_11697);
xor U12307 (N_12307,N_11741,N_11593);
nand U12308 (N_12308,N_11912,N_11524);
nor U12309 (N_12309,N_11924,N_11986);
xnor U12310 (N_12310,N_11970,N_11683);
or U12311 (N_12311,N_11901,N_11696);
xor U12312 (N_12312,N_11540,N_11743);
nor U12313 (N_12313,N_11906,N_11770);
xnor U12314 (N_12314,N_11558,N_11912);
or U12315 (N_12315,N_11926,N_11831);
nand U12316 (N_12316,N_11797,N_11970);
xor U12317 (N_12317,N_11767,N_11857);
or U12318 (N_12318,N_11870,N_11726);
and U12319 (N_12319,N_11655,N_11705);
and U12320 (N_12320,N_11997,N_11875);
or U12321 (N_12321,N_11691,N_11704);
and U12322 (N_12322,N_11581,N_11729);
nand U12323 (N_12323,N_11872,N_11954);
nor U12324 (N_12324,N_11868,N_11731);
or U12325 (N_12325,N_11856,N_11758);
nand U12326 (N_12326,N_11675,N_11524);
nor U12327 (N_12327,N_11986,N_11885);
and U12328 (N_12328,N_11997,N_11594);
and U12329 (N_12329,N_11809,N_11880);
xnor U12330 (N_12330,N_11620,N_11755);
or U12331 (N_12331,N_11717,N_11677);
nand U12332 (N_12332,N_11759,N_11900);
xor U12333 (N_12333,N_11907,N_11523);
nand U12334 (N_12334,N_11970,N_11542);
xor U12335 (N_12335,N_11785,N_11745);
and U12336 (N_12336,N_11747,N_11754);
nand U12337 (N_12337,N_11905,N_11949);
nand U12338 (N_12338,N_11611,N_11992);
xor U12339 (N_12339,N_11793,N_11774);
nand U12340 (N_12340,N_11873,N_11794);
and U12341 (N_12341,N_11648,N_11607);
nand U12342 (N_12342,N_11860,N_11882);
nor U12343 (N_12343,N_11952,N_11629);
and U12344 (N_12344,N_11833,N_11688);
nand U12345 (N_12345,N_11810,N_11943);
nand U12346 (N_12346,N_11707,N_11619);
or U12347 (N_12347,N_11731,N_11583);
xnor U12348 (N_12348,N_11765,N_11802);
or U12349 (N_12349,N_11653,N_11985);
and U12350 (N_12350,N_11760,N_11596);
or U12351 (N_12351,N_11872,N_11870);
nand U12352 (N_12352,N_11871,N_11922);
xnor U12353 (N_12353,N_11817,N_11628);
and U12354 (N_12354,N_11793,N_11948);
or U12355 (N_12355,N_11864,N_11734);
nor U12356 (N_12356,N_11535,N_11826);
nand U12357 (N_12357,N_11645,N_11870);
nand U12358 (N_12358,N_11501,N_11757);
or U12359 (N_12359,N_11861,N_11530);
or U12360 (N_12360,N_11537,N_11586);
and U12361 (N_12361,N_11639,N_11747);
and U12362 (N_12362,N_11945,N_11637);
and U12363 (N_12363,N_11797,N_11790);
nor U12364 (N_12364,N_11637,N_11819);
xnor U12365 (N_12365,N_11962,N_11960);
or U12366 (N_12366,N_11850,N_11696);
xor U12367 (N_12367,N_11772,N_11754);
or U12368 (N_12368,N_11663,N_11522);
and U12369 (N_12369,N_11854,N_11669);
nor U12370 (N_12370,N_11529,N_11555);
nand U12371 (N_12371,N_11929,N_11765);
xor U12372 (N_12372,N_11611,N_11678);
or U12373 (N_12373,N_11642,N_11654);
xor U12374 (N_12374,N_11583,N_11610);
and U12375 (N_12375,N_11731,N_11636);
or U12376 (N_12376,N_11529,N_11864);
nand U12377 (N_12377,N_11824,N_11968);
nor U12378 (N_12378,N_11758,N_11936);
or U12379 (N_12379,N_11974,N_11838);
xnor U12380 (N_12380,N_11975,N_11764);
or U12381 (N_12381,N_11993,N_11750);
xor U12382 (N_12382,N_11572,N_11577);
xor U12383 (N_12383,N_11713,N_11551);
or U12384 (N_12384,N_11834,N_11589);
or U12385 (N_12385,N_11862,N_11721);
nand U12386 (N_12386,N_11907,N_11980);
nand U12387 (N_12387,N_11808,N_11842);
nand U12388 (N_12388,N_11740,N_11946);
nand U12389 (N_12389,N_11683,N_11641);
nand U12390 (N_12390,N_11665,N_11792);
and U12391 (N_12391,N_11814,N_11991);
nand U12392 (N_12392,N_11710,N_11766);
nand U12393 (N_12393,N_11761,N_11601);
or U12394 (N_12394,N_11993,N_11824);
and U12395 (N_12395,N_11588,N_11868);
and U12396 (N_12396,N_11892,N_11961);
nor U12397 (N_12397,N_11973,N_11931);
xnor U12398 (N_12398,N_11993,N_11746);
nor U12399 (N_12399,N_11963,N_11573);
xor U12400 (N_12400,N_11788,N_11844);
nor U12401 (N_12401,N_11906,N_11568);
xor U12402 (N_12402,N_11696,N_11739);
nor U12403 (N_12403,N_11913,N_11824);
nand U12404 (N_12404,N_11996,N_11875);
and U12405 (N_12405,N_11791,N_11974);
xor U12406 (N_12406,N_11753,N_11882);
and U12407 (N_12407,N_11769,N_11532);
nor U12408 (N_12408,N_11916,N_11965);
xor U12409 (N_12409,N_11847,N_11524);
nor U12410 (N_12410,N_11928,N_11867);
and U12411 (N_12411,N_11900,N_11556);
nor U12412 (N_12412,N_11929,N_11850);
nand U12413 (N_12413,N_11500,N_11529);
xnor U12414 (N_12414,N_11787,N_11693);
nand U12415 (N_12415,N_11972,N_11509);
xnor U12416 (N_12416,N_11902,N_11587);
or U12417 (N_12417,N_11833,N_11799);
nor U12418 (N_12418,N_11770,N_11798);
xor U12419 (N_12419,N_11509,N_11886);
and U12420 (N_12420,N_11978,N_11733);
and U12421 (N_12421,N_11604,N_11551);
xor U12422 (N_12422,N_11974,N_11703);
nand U12423 (N_12423,N_11714,N_11670);
xnor U12424 (N_12424,N_11898,N_11758);
nor U12425 (N_12425,N_11709,N_11848);
or U12426 (N_12426,N_11933,N_11628);
nor U12427 (N_12427,N_11594,N_11906);
or U12428 (N_12428,N_11750,N_11758);
and U12429 (N_12429,N_11644,N_11592);
nand U12430 (N_12430,N_11546,N_11832);
and U12431 (N_12431,N_11560,N_11828);
and U12432 (N_12432,N_11785,N_11859);
nor U12433 (N_12433,N_11851,N_11885);
and U12434 (N_12434,N_11831,N_11761);
and U12435 (N_12435,N_11928,N_11706);
and U12436 (N_12436,N_11787,N_11732);
xor U12437 (N_12437,N_11908,N_11510);
or U12438 (N_12438,N_11800,N_11645);
xnor U12439 (N_12439,N_11734,N_11924);
nor U12440 (N_12440,N_11739,N_11779);
and U12441 (N_12441,N_11849,N_11724);
nand U12442 (N_12442,N_11699,N_11763);
xor U12443 (N_12443,N_11987,N_11538);
xnor U12444 (N_12444,N_11973,N_11771);
and U12445 (N_12445,N_11527,N_11734);
nor U12446 (N_12446,N_11874,N_11625);
and U12447 (N_12447,N_11805,N_11781);
xnor U12448 (N_12448,N_11909,N_11653);
nand U12449 (N_12449,N_11790,N_11781);
nor U12450 (N_12450,N_11534,N_11526);
or U12451 (N_12451,N_11869,N_11563);
nand U12452 (N_12452,N_11863,N_11872);
nor U12453 (N_12453,N_11645,N_11669);
nand U12454 (N_12454,N_11519,N_11916);
xor U12455 (N_12455,N_11619,N_11940);
nand U12456 (N_12456,N_11710,N_11585);
xnor U12457 (N_12457,N_11737,N_11990);
or U12458 (N_12458,N_11917,N_11941);
nor U12459 (N_12459,N_11965,N_11737);
or U12460 (N_12460,N_11614,N_11560);
nand U12461 (N_12461,N_11797,N_11505);
nor U12462 (N_12462,N_11701,N_11571);
xnor U12463 (N_12463,N_11741,N_11802);
nand U12464 (N_12464,N_11625,N_11865);
and U12465 (N_12465,N_11626,N_11739);
xor U12466 (N_12466,N_11974,N_11767);
nor U12467 (N_12467,N_11817,N_11759);
and U12468 (N_12468,N_11954,N_11897);
nand U12469 (N_12469,N_11544,N_11903);
and U12470 (N_12470,N_11514,N_11755);
and U12471 (N_12471,N_11866,N_11980);
xor U12472 (N_12472,N_11746,N_11957);
nor U12473 (N_12473,N_11913,N_11712);
or U12474 (N_12474,N_11668,N_11557);
xnor U12475 (N_12475,N_11767,N_11854);
nand U12476 (N_12476,N_11723,N_11893);
or U12477 (N_12477,N_11901,N_11865);
xnor U12478 (N_12478,N_11889,N_11996);
nor U12479 (N_12479,N_11795,N_11726);
xnor U12480 (N_12480,N_11679,N_11939);
and U12481 (N_12481,N_11772,N_11966);
and U12482 (N_12482,N_11950,N_11897);
nor U12483 (N_12483,N_11829,N_11743);
and U12484 (N_12484,N_11714,N_11645);
nor U12485 (N_12485,N_11786,N_11600);
or U12486 (N_12486,N_11751,N_11823);
xnor U12487 (N_12487,N_11983,N_11999);
nor U12488 (N_12488,N_11515,N_11944);
xnor U12489 (N_12489,N_11995,N_11743);
or U12490 (N_12490,N_11552,N_11877);
nand U12491 (N_12491,N_11954,N_11946);
and U12492 (N_12492,N_11882,N_11503);
nand U12493 (N_12493,N_11866,N_11623);
and U12494 (N_12494,N_11800,N_11610);
xnor U12495 (N_12495,N_11867,N_11677);
and U12496 (N_12496,N_11755,N_11686);
nand U12497 (N_12497,N_11578,N_11856);
or U12498 (N_12498,N_11823,N_11598);
nand U12499 (N_12499,N_11903,N_11857);
nor U12500 (N_12500,N_12135,N_12172);
and U12501 (N_12501,N_12428,N_12370);
nor U12502 (N_12502,N_12312,N_12401);
xnor U12503 (N_12503,N_12026,N_12450);
xnor U12504 (N_12504,N_12284,N_12002);
xnor U12505 (N_12505,N_12111,N_12231);
nand U12506 (N_12506,N_12466,N_12241);
nand U12507 (N_12507,N_12394,N_12039);
nor U12508 (N_12508,N_12001,N_12009);
xnor U12509 (N_12509,N_12119,N_12485);
nand U12510 (N_12510,N_12107,N_12341);
nand U12511 (N_12511,N_12057,N_12388);
and U12512 (N_12512,N_12049,N_12131);
xor U12513 (N_12513,N_12353,N_12071);
nor U12514 (N_12514,N_12165,N_12088);
nor U12515 (N_12515,N_12294,N_12102);
or U12516 (N_12516,N_12117,N_12140);
nand U12517 (N_12517,N_12464,N_12174);
and U12518 (N_12518,N_12025,N_12058);
and U12519 (N_12519,N_12348,N_12308);
and U12520 (N_12520,N_12461,N_12151);
nor U12521 (N_12521,N_12304,N_12458);
nor U12522 (N_12522,N_12323,N_12068);
or U12523 (N_12523,N_12300,N_12113);
or U12524 (N_12524,N_12031,N_12277);
and U12525 (N_12525,N_12351,N_12380);
nor U12526 (N_12526,N_12330,N_12175);
or U12527 (N_12527,N_12305,N_12374);
nor U12528 (N_12528,N_12115,N_12448);
and U12529 (N_12529,N_12099,N_12093);
and U12530 (N_12530,N_12298,N_12095);
nand U12531 (N_12531,N_12391,N_12038);
xnor U12532 (N_12532,N_12494,N_12293);
xor U12533 (N_12533,N_12084,N_12322);
xnor U12534 (N_12534,N_12121,N_12120);
and U12535 (N_12535,N_12456,N_12110);
nand U12536 (N_12536,N_12015,N_12340);
nor U12537 (N_12537,N_12460,N_12367);
or U12538 (N_12538,N_12359,N_12048);
and U12539 (N_12539,N_12287,N_12496);
or U12540 (N_12540,N_12027,N_12018);
xor U12541 (N_12541,N_12422,N_12385);
nor U12542 (N_12542,N_12372,N_12378);
nor U12543 (N_12543,N_12389,N_12316);
and U12544 (N_12544,N_12130,N_12282);
xnor U12545 (N_12545,N_12265,N_12419);
nor U12546 (N_12546,N_12166,N_12347);
and U12547 (N_12547,N_12288,N_12339);
nor U12548 (N_12548,N_12257,N_12143);
nand U12549 (N_12549,N_12318,N_12008);
or U12550 (N_12550,N_12133,N_12278);
or U12551 (N_12551,N_12263,N_12290);
nor U12552 (N_12552,N_12200,N_12204);
and U12553 (N_12553,N_12486,N_12234);
and U12554 (N_12554,N_12237,N_12346);
xnor U12555 (N_12555,N_12499,N_12045);
nor U12556 (N_12556,N_12315,N_12210);
xor U12557 (N_12557,N_12427,N_12202);
xnor U12558 (N_12558,N_12451,N_12495);
nand U12559 (N_12559,N_12307,N_12404);
or U12560 (N_12560,N_12064,N_12381);
xnor U12561 (N_12561,N_12044,N_12283);
xor U12562 (N_12562,N_12016,N_12443);
and U12563 (N_12563,N_12157,N_12452);
nand U12564 (N_12564,N_12345,N_12075);
xnor U12565 (N_12565,N_12144,N_12435);
nand U12566 (N_12566,N_12050,N_12148);
nor U12567 (N_12567,N_12269,N_12441);
and U12568 (N_12568,N_12261,N_12053);
nand U12569 (N_12569,N_12332,N_12418);
or U12570 (N_12570,N_12080,N_12276);
or U12571 (N_12571,N_12396,N_12386);
nand U12572 (N_12572,N_12147,N_12361);
and U12573 (N_12573,N_12303,N_12226);
or U12574 (N_12574,N_12336,N_12470);
and U12575 (N_12575,N_12349,N_12221);
nor U12576 (N_12576,N_12214,N_12463);
and U12577 (N_12577,N_12056,N_12465);
xor U12578 (N_12578,N_12258,N_12420);
and U12579 (N_12579,N_12264,N_12247);
and U12580 (N_12580,N_12407,N_12434);
xor U12581 (N_12581,N_12393,N_12207);
and U12582 (N_12582,N_12397,N_12061);
nand U12583 (N_12583,N_12155,N_12362);
nor U12584 (N_12584,N_12091,N_12171);
or U12585 (N_12585,N_12487,N_12227);
nor U12586 (N_12586,N_12392,N_12311);
and U12587 (N_12587,N_12037,N_12299);
or U12588 (N_12588,N_12125,N_12090);
nand U12589 (N_12589,N_12302,N_12357);
and U12590 (N_12590,N_12182,N_12124);
and U12591 (N_12591,N_12096,N_12161);
xor U12592 (N_12592,N_12270,N_12471);
and U12593 (N_12593,N_12051,N_12245);
or U12594 (N_12594,N_12235,N_12371);
and U12595 (N_12595,N_12403,N_12179);
or U12596 (N_12596,N_12178,N_12167);
nand U12597 (N_12597,N_12216,N_12104);
nor U12598 (N_12598,N_12097,N_12063);
and U12599 (N_12599,N_12498,N_12424);
or U12600 (N_12600,N_12156,N_12036);
and U12601 (N_12601,N_12432,N_12255);
or U12602 (N_12602,N_12368,N_12366);
nor U12603 (N_12603,N_12350,N_12275);
nand U12604 (N_12604,N_12077,N_12272);
or U12605 (N_12605,N_12190,N_12203);
or U12606 (N_12606,N_12342,N_12395);
nand U12607 (N_12607,N_12154,N_12076);
nor U12608 (N_12608,N_12289,N_12415);
xnor U12609 (N_12609,N_12473,N_12006);
xnor U12610 (N_12610,N_12239,N_12320);
or U12611 (N_12611,N_12236,N_12297);
nand U12612 (N_12612,N_12209,N_12028);
nor U12613 (N_12613,N_12136,N_12042);
nand U12614 (N_12614,N_12313,N_12319);
and U12615 (N_12615,N_12122,N_12399);
and U12616 (N_12616,N_12326,N_12032);
or U12617 (N_12617,N_12047,N_12205);
nand U12618 (N_12618,N_12138,N_12081);
and U12619 (N_12619,N_12023,N_12431);
and U12620 (N_12620,N_12052,N_12497);
nor U12621 (N_12621,N_12029,N_12333);
nor U12622 (N_12622,N_12079,N_12334);
and U12623 (N_12623,N_12177,N_12163);
xor U12624 (N_12624,N_12112,N_12426);
or U12625 (N_12625,N_12256,N_12437);
or U12626 (N_12626,N_12478,N_12453);
xor U12627 (N_12627,N_12267,N_12343);
and U12628 (N_12628,N_12149,N_12365);
nor U12629 (N_12629,N_12108,N_12373);
and U12630 (N_12630,N_12408,N_12011);
xnor U12631 (N_12631,N_12176,N_12129);
nand U12632 (N_12632,N_12109,N_12195);
nand U12633 (N_12633,N_12309,N_12014);
nor U12634 (N_12634,N_12295,N_12150);
nand U12635 (N_12635,N_12457,N_12273);
nor U12636 (N_12636,N_12271,N_12410);
or U12637 (N_12637,N_12220,N_12477);
and U12638 (N_12638,N_12335,N_12480);
or U12639 (N_12639,N_12445,N_12442);
and U12640 (N_12640,N_12159,N_12067);
xor U12641 (N_12641,N_12358,N_12327);
and U12642 (N_12642,N_12429,N_12082);
nor U12643 (N_12643,N_12484,N_12035);
and U12644 (N_12644,N_12065,N_12022);
or U12645 (N_12645,N_12017,N_12232);
xnor U12646 (N_12646,N_12387,N_12253);
nor U12647 (N_12647,N_12436,N_12199);
nand U12648 (N_12648,N_12225,N_12352);
nand U12649 (N_12649,N_12010,N_12060);
nor U12650 (N_12650,N_12364,N_12041);
xor U12651 (N_12651,N_12127,N_12406);
and U12652 (N_12652,N_12325,N_12173);
and U12653 (N_12653,N_12416,N_12005);
or U12654 (N_12654,N_12337,N_12375);
nand U12655 (N_12655,N_12012,N_12242);
xnor U12656 (N_12656,N_12310,N_12033);
nor U12657 (N_12657,N_12398,N_12417);
or U12658 (N_12658,N_12493,N_12123);
nand U12659 (N_12659,N_12369,N_12142);
and U12660 (N_12660,N_12212,N_12376);
and U12661 (N_12661,N_12462,N_12070);
or U12662 (N_12662,N_12101,N_12145);
xor U12663 (N_12663,N_12098,N_12191);
nand U12664 (N_12664,N_12438,N_12043);
or U12665 (N_12665,N_12279,N_12400);
xnor U12666 (N_12666,N_12222,N_12092);
nand U12667 (N_12667,N_12083,N_12383);
or U12668 (N_12668,N_12296,N_12197);
or U12669 (N_12669,N_12160,N_12479);
and U12670 (N_12670,N_12411,N_12338);
nor U12671 (N_12671,N_12162,N_12089);
and U12672 (N_12672,N_12004,N_12238);
and U12673 (N_12673,N_12446,N_12188);
and U12674 (N_12674,N_12317,N_12003);
xnor U12675 (N_12675,N_12158,N_12331);
or U12676 (N_12676,N_12344,N_12449);
nor U12677 (N_12677,N_12066,N_12246);
nor U12678 (N_12678,N_12180,N_12377);
and U12679 (N_12679,N_12306,N_12013);
xor U12680 (N_12680,N_12094,N_12414);
nor U12681 (N_12681,N_12467,N_12324);
nand U12682 (N_12682,N_12329,N_12228);
or U12683 (N_12683,N_12072,N_12314);
or U12684 (N_12684,N_12440,N_12421);
nor U12685 (N_12685,N_12244,N_12137);
or U12686 (N_12686,N_12168,N_12430);
xnor U12687 (N_12687,N_12116,N_12134);
nor U12688 (N_12688,N_12229,N_12074);
nor U12689 (N_12689,N_12413,N_12285);
and U12690 (N_12690,N_12185,N_12217);
or U12691 (N_12691,N_12034,N_12062);
nor U12692 (N_12692,N_12233,N_12251);
nor U12693 (N_12693,N_12024,N_12046);
xnor U12694 (N_12694,N_12249,N_12186);
or U12695 (N_12695,N_12482,N_12274);
and U12696 (N_12696,N_12382,N_12280);
nor U12697 (N_12697,N_12248,N_12196);
and U12698 (N_12698,N_12439,N_12447);
nand U12699 (N_12699,N_12489,N_12030);
or U12700 (N_12700,N_12146,N_12481);
nor U12701 (N_12701,N_12132,N_12189);
and U12702 (N_12702,N_12240,N_12183);
and U12703 (N_12703,N_12118,N_12286);
nand U12704 (N_12704,N_12390,N_12198);
or U12705 (N_12705,N_12301,N_12328);
nand U12706 (N_12706,N_12476,N_12219);
and U12707 (N_12707,N_12184,N_12468);
and U12708 (N_12708,N_12490,N_12218);
nand U12709 (N_12709,N_12250,N_12360);
nand U12710 (N_12710,N_12356,N_12412);
nand U12711 (N_12711,N_12019,N_12433);
nand U12712 (N_12712,N_12259,N_12187);
nor U12713 (N_12713,N_12201,N_12223);
and U12714 (N_12714,N_12262,N_12106);
nand U12715 (N_12715,N_12254,N_12105);
nor U12716 (N_12716,N_12100,N_12152);
nor U12717 (N_12717,N_12169,N_12455);
nor U12718 (N_12718,N_12069,N_12073);
xor U12719 (N_12719,N_12488,N_12192);
xor U12720 (N_12720,N_12164,N_12086);
or U12721 (N_12721,N_12139,N_12475);
or U12722 (N_12722,N_12054,N_12021);
xor U12723 (N_12723,N_12085,N_12128);
nor U12724 (N_12724,N_12252,N_12078);
nand U12725 (N_12725,N_12483,N_12492);
nand U12726 (N_12726,N_12230,N_12211);
xor U12727 (N_12727,N_12194,N_12141);
or U12728 (N_12728,N_12103,N_12291);
xor U12729 (N_12729,N_12206,N_12409);
nand U12730 (N_12730,N_12170,N_12292);
nand U12731 (N_12731,N_12243,N_12469);
or U12732 (N_12732,N_12423,N_12384);
nand U12733 (N_12733,N_12425,N_12268);
nand U12734 (N_12734,N_12321,N_12355);
and U12735 (N_12735,N_12153,N_12354);
nand U12736 (N_12736,N_12454,N_12266);
or U12737 (N_12737,N_12059,N_12193);
nand U12738 (N_12738,N_12007,N_12224);
nor U12739 (N_12739,N_12020,N_12281);
and U12740 (N_12740,N_12213,N_12114);
and U12741 (N_12741,N_12087,N_12126);
xnor U12742 (N_12742,N_12459,N_12405);
nand U12743 (N_12743,N_12472,N_12363);
xor U12744 (N_12744,N_12402,N_12379);
and U12745 (N_12745,N_12040,N_12055);
or U12746 (N_12746,N_12215,N_12181);
or U12747 (N_12747,N_12208,N_12491);
xor U12748 (N_12748,N_12000,N_12474);
and U12749 (N_12749,N_12260,N_12444);
nand U12750 (N_12750,N_12019,N_12202);
xnor U12751 (N_12751,N_12239,N_12203);
nor U12752 (N_12752,N_12444,N_12109);
xnor U12753 (N_12753,N_12024,N_12010);
xor U12754 (N_12754,N_12127,N_12303);
or U12755 (N_12755,N_12111,N_12130);
nor U12756 (N_12756,N_12123,N_12079);
xnor U12757 (N_12757,N_12216,N_12211);
and U12758 (N_12758,N_12155,N_12111);
xor U12759 (N_12759,N_12383,N_12325);
nor U12760 (N_12760,N_12255,N_12402);
or U12761 (N_12761,N_12437,N_12231);
and U12762 (N_12762,N_12083,N_12390);
and U12763 (N_12763,N_12473,N_12210);
and U12764 (N_12764,N_12038,N_12268);
or U12765 (N_12765,N_12366,N_12104);
nand U12766 (N_12766,N_12249,N_12110);
xnor U12767 (N_12767,N_12211,N_12026);
and U12768 (N_12768,N_12108,N_12183);
and U12769 (N_12769,N_12072,N_12081);
nand U12770 (N_12770,N_12002,N_12277);
and U12771 (N_12771,N_12224,N_12137);
nor U12772 (N_12772,N_12198,N_12042);
nand U12773 (N_12773,N_12312,N_12335);
nor U12774 (N_12774,N_12474,N_12232);
or U12775 (N_12775,N_12042,N_12163);
nand U12776 (N_12776,N_12249,N_12424);
xor U12777 (N_12777,N_12129,N_12021);
or U12778 (N_12778,N_12093,N_12163);
and U12779 (N_12779,N_12394,N_12327);
nor U12780 (N_12780,N_12119,N_12332);
xor U12781 (N_12781,N_12095,N_12017);
nand U12782 (N_12782,N_12409,N_12373);
nand U12783 (N_12783,N_12477,N_12359);
nor U12784 (N_12784,N_12197,N_12248);
nor U12785 (N_12785,N_12219,N_12253);
xnor U12786 (N_12786,N_12065,N_12124);
xor U12787 (N_12787,N_12206,N_12184);
xor U12788 (N_12788,N_12329,N_12144);
or U12789 (N_12789,N_12208,N_12277);
and U12790 (N_12790,N_12347,N_12308);
or U12791 (N_12791,N_12464,N_12210);
nand U12792 (N_12792,N_12292,N_12028);
nand U12793 (N_12793,N_12448,N_12091);
xnor U12794 (N_12794,N_12110,N_12177);
or U12795 (N_12795,N_12305,N_12114);
or U12796 (N_12796,N_12198,N_12441);
nor U12797 (N_12797,N_12102,N_12458);
xnor U12798 (N_12798,N_12028,N_12036);
or U12799 (N_12799,N_12444,N_12197);
and U12800 (N_12800,N_12027,N_12133);
nand U12801 (N_12801,N_12043,N_12279);
nand U12802 (N_12802,N_12001,N_12486);
nand U12803 (N_12803,N_12409,N_12401);
and U12804 (N_12804,N_12046,N_12097);
nor U12805 (N_12805,N_12363,N_12138);
or U12806 (N_12806,N_12056,N_12390);
or U12807 (N_12807,N_12212,N_12404);
nor U12808 (N_12808,N_12168,N_12024);
nand U12809 (N_12809,N_12418,N_12152);
nor U12810 (N_12810,N_12017,N_12051);
xnor U12811 (N_12811,N_12344,N_12159);
nand U12812 (N_12812,N_12103,N_12050);
or U12813 (N_12813,N_12145,N_12236);
nand U12814 (N_12814,N_12020,N_12189);
nor U12815 (N_12815,N_12027,N_12175);
xnor U12816 (N_12816,N_12421,N_12024);
or U12817 (N_12817,N_12293,N_12136);
nand U12818 (N_12818,N_12082,N_12116);
and U12819 (N_12819,N_12292,N_12490);
and U12820 (N_12820,N_12290,N_12205);
or U12821 (N_12821,N_12455,N_12353);
nand U12822 (N_12822,N_12113,N_12047);
and U12823 (N_12823,N_12079,N_12357);
xnor U12824 (N_12824,N_12156,N_12204);
nor U12825 (N_12825,N_12093,N_12208);
or U12826 (N_12826,N_12238,N_12181);
and U12827 (N_12827,N_12055,N_12212);
nor U12828 (N_12828,N_12299,N_12357);
and U12829 (N_12829,N_12258,N_12282);
nor U12830 (N_12830,N_12160,N_12013);
and U12831 (N_12831,N_12235,N_12003);
or U12832 (N_12832,N_12132,N_12376);
nor U12833 (N_12833,N_12061,N_12417);
xor U12834 (N_12834,N_12036,N_12187);
nor U12835 (N_12835,N_12052,N_12026);
or U12836 (N_12836,N_12308,N_12215);
xnor U12837 (N_12837,N_12303,N_12126);
xnor U12838 (N_12838,N_12303,N_12441);
nor U12839 (N_12839,N_12001,N_12152);
nand U12840 (N_12840,N_12223,N_12342);
and U12841 (N_12841,N_12328,N_12363);
and U12842 (N_12842,N_12387,N_12498);
and U12843 (N_12843,N_12163,N_12002);
and U12844 (N_12844,N_12422,N_12298);
or U12845 (N_12845,N_12110,N_12347);
xnor U12846 (N_12846,N_12491,N_12129);
xnor U12847 (N_12847,N_12091,N_12321);
or U12848 (N_12848,N_12245,N_12072);
and U12849 (N_12849,N_12040,N_12453);
or U12850 (N_12850,N_12435,N_12082);
nor U12851 (N_12851,N_12165,N_12143);
nor U12852 (N_12852,N_12353,N_12299);
nor U12853 (N_12853,N_12476,N_12099);
nand U12854 (N_12854,N_12319,N_12253);
and U12855 (N_12855,N_12082,N_12482);
nor U12856 (N_12856,N_12079,N_12064);
or U12857 (N_12857,N_12025,N_12117);
and U12858 (N_12858,N_12329,N_12421);
xnor U12859 (N_12859,N_12005,N_12177);
nand U12860 (N_12860,N_12218,N_12092);
xnor U12861 (N_12861,N_12136,N_12459);
xor U12862 (N_12862,N_12286,N_12476);
nor U12863 (N_12863,N_12427,N_12121);
or U12864 (N_12864,N_12421,N_12059);
xnor U12865 (N_12865,N_12403,N_12212);
xnor U12866 (N_12866,N_12363,N_12265);
or U12867 (N_12867,N_12039,N_12396);
and U12868 (N_12868,N_12456,N_12050);
xnor U12869 (N_12869,N_12034,N_12043);
or U12870 (N_12870,N_12253,N_12336);
nand U12871 (N_12871,N_12028,N_12326);
nor U12872 (N_12872,N_12008,N_12387);
nor U12873 (N_12873,N_12444,N_12023);
or U12874 (N_12874,N_12250,N_12374);
nand U12875 (N_12875,N_12214,N_12241);
xor U12876 (N_12876,N_12120,N_12493);
nor U12877 (N_12877,N_12428,N_12349);
nor U12878 (N_12878,N_12426,N_12051);
nor U12879 (N_12879,N_12265,N_12311);
xnor U12880 (N_12880,N_12078,N_12283);
and U12881 (N_12881,N_12402,N_12364);
or U12882 (N_12882,N_12404,N_12349);
nand U12883 (N_12883,N_12426,N_12291);
xnor U12884 (N_12884,N_12210,N_12441);
or U12885 (N_12885,N_12029,N_12048);
xor U12886 (N_12886,N_12174,N_12293);
nor U12887 (N_12887,N_12469,N_12016);
and U12888 (N_12888,N_12358,N_12303);
or U12889 (N_12889,N_12195,N_12435);
and U12890 (N_12890,N_12352,N_12054);
xnor U12891 (N_12891,N_12476,N_12073);
nand U12892 (N_12892,N_12396,N_12414);
or U12893 (N_12893,N_12103,N_12095);
xnor U12894 (N_12894,N_12409,N_12140);
or U12895 (N_12895,N_12029,N_12045);
nand U12896 (N_12896,N_12056,N_12290);
and U12897 (N_12897,N_12323,N_12368);
and U12898 (N_12898,N_12453,N_12329);
xnor U12899 (N_12899,N_12070,N_12330);
nand U12900 (N_12900,N_12103,N_12420);
xnor U12901 (N_12901,N_12153,N_12213);
xnor U12902 (N_12902,N_12295,N_12297);
and U12903 (N_12903,N_12096,N_12081);
or U12904 (N_12904,N_12031,N_12102);
and U12905 (N_12905,N_12154,N_12242);
nor U12906 (N_12906,N_12260,N_12198);
or U12907 (N_12907,N_12040,N_12203);
nor U12908 (N_12908,N_12295,N_12144);
xnor U12909 (N_12909,N_12469,N_12295);
and U12910 (N_12910,N_12308,N_12275);
or U12911 (N_12911,N_12373,N_12016);
xnor U12912 (N_12912,N_12019,N_12203);
nor U12913 (N_12913,N_12179,N_12117);
or U12914 (N_12914,N_12472,N_12063);
and U12915 (N_12915,N_12357,N_12050);
and U12916 (N_12916,N_12177,N_12087);
and U12917 (N_12917,N_12459,N_12217);
nor U12918 (N_12918,N_12174,N_12428);
and U12919 (N_12919,N_12091,N_12326);
nand U12920 (N_12920,N_12320,N_12058);
and U12921 (N_12921,N_12025,N_12101);
or U12922 (N_12922,N_12097,N_12472);
and U12923 (N_12923,N_12455,N_12178);
or U12924 (N_12924,N_12441,N_12176);
xnor U12925 (N_12925,N_12078,N_12383);
and U12926 (N_12926,N_12243,N_12293);
and U12927 (N_12927,N_12188,N_12314);
or U12928 (N_12928,N_12405,N_12061);
nand U12929 (N_12929,N_12132,N_12342);
xnor U12930 (N_12930,N_12442,N_12247);
xnor U12931 (N_12931,N_12024,N_12382);
and U12932 (N_12932,N_12353,N_12392);
and U12933 (N_12933,N_12392,N_12265);
and U12934 (N_12934,N_12408,N_12062);
nand U12935 (N_12935,N_12363,N_12113);
or U12936 (N_12936,N_12457,N_12128);
or U12937 (N_12937,N_12277,N_12150);
nor U12938 (N_12938,N_12214,N_12125);
nor U12939 (N_12939,N_12290,N_12456);
and U12940 (N_12940,N_12055,N_12464);
or U12941 (N_12941,N_12299,N_12111);
nand U12942 (N_12942,N_12251,N_12299);
xor U12943 (N_12943,N_12198,N_12299);
nand U12944 (N_12944,N_12385,N_12453);
and U12945 (N_12945,N_12101,N_12060);
nand U12946 (N_12946,N_12357,N_12392);
and U12947 (N_12947,N_12104,N_12413);
nor U12948 (N_12948,N_12235,N_12447);
nor U12949 (N_12949,N_12181,N_12397);
or U12950 (N_12950,N_12100,N_12146);
or U12951 (N_12951,N_12034,N_12351);
xor U12952 (N_12952,N_12439,N_12321);
or U12953 (N_12953,N_12356,N_12328);
and U12954 (N_12954,N_12003,N_12035);
nor U12955 (N_12955,N_12184,N_12081);
or U12956 (N_12956,N_12254,N_12033);
and U12957 (N_12957,N_12460,N_12075);
nor U12958 (N_12958,N_12181,N_12322);
nor U12959 (N_12959,N_12288,N_12107);
nor U12960 (N_12960,N_12060,N_12221);
or U12961 (N_12961,N_12350,N_12117);
xor U12962 (N_12962,N_12287,N_12477);
nor U12963 (N_12963,N_12060,N_12471);
nand U12964 (N_12964,N_12408,N_12252);
and U12965 (N_12965,N_12370,N_12254);
xor U12966 (N_12966,N_12073,N_12482);
xnor U12967 (N_12967,N_12414,N_12047);
and U12968 (N_12968,N_12255,N_12034);
and U12969 (N_12969,N_12412,N_12383);
nand U12970 (N_12970,N_12222,N_12133);
and U12971 (N_12971,N_12221,N_12097);
nand U12972 (N_12972,N_12391,N_12404);
xnor U12973 (N_12973,N_12360,N_12107);
xnor U12974 (N_12974,N_12027,N_12287);
and U12975 (N_12975,N_12406,N_12382);
nor U12976 (N_12976,N_12136,N_12059);
nand U12977 (N_12977,N_12476,N_12194);
or U12978 (N_12978,N_12020,N_12015);
and U12979 (N_12979,N_12203,N_12467);
or U12980 (N_12980,N_12379,N_12109);
nor U12981 (N_12981,N_12312,N_12147);
nand U12982 (N_12982,N_12257,N_12408);
nor U12983 (N_12983,N_12346,N_12160);
xor U12984 (N_12984,N_12366,N_12336);
xor U12985 (N_12985,N_12003,N_12196);
or U12986 (N_12986,N_12116,N_12251);
and U12987 (N_12987,N_12337,N_12013);
and U12988 (N_12988,N_12142,N_12015);
nor U12989 (N_12989,N_12362,N_12043);
xor U12990 (N_12990,N_12000,N_12222);
and U12991 (N_12991,N_12427,N_12298);
nor U12992 (N_12992,N_12250,N_12279);
nand U12993 (N_12993,N_12295,N_12420);
nor U12994 (N_12994,N_12470,N_12179);
nand U12995 (N_12995,N_12427,N_12291);
nand U12996 (N_12996,N_12330,N_12415);
or U12997 (N_12997,N_12101,N_12268);
nand U12998 (N_12998,N_12257,N_12305);
xor U12999 (N_12999,N_12298,N_12223);
xnor U13000 (N_13000,N_12957,N_12817);
nor U13001 (N_13001,N_12677,N_12571);
nor U13002 (N_13002,N_12714,N_12829);
and U13003 (N_13003,N_12919,N_12818);
nand U13004 (N_13004,N_12551,N_12899);
or U13005 (N_13005,N_12972,N_12687);
nor U13006 (N_13006,N_12888,N_12519);
xor U13007 (N_13007,N_12999,N_12596);
xor U13008 (N_13008,N_12708,N_12757);
or U13009 (N_13009,N_12780,N_12942);
nand U13010 (N_13010,N_12807,N_12769);
and U13011 (N_13011,N_12800,N_12644);
or U13012 (N_13012,N_12837,N_12946);
nand U13013 (N_13013,N_12742,N_12938);
nor U13014 (N_13014,N_12896,N_12789);
or U13015 (N_13015,N_12977,N_12993);
nand U13016 (N_13016,N_12759,N_12808);
nor U13017 (N_13017,N_12795,N_12569);
nor U13018 (N_13018,N_12730,N_12512);
and U13019 (N_13019,N_12636,N_12924);
nand U13020 (N_13020,N_12657,N_12563);
and U13021 (N_13021,N_12768,N_12621);
nand U13022 (N_13022,N_12593,N_12735);
or U13023 (N_13023,N_12516,N_12874);
xnor U13024 (N_13024,N_12839,N_12589);
nand U13025 (N_13025,N_12989,N_12565);
xnor U13026 (N_13026,N_12860,N_12517);
nor U13027 (N_13027,N_12573,N_12727);
xnor U13028 (N_13028,N_12965,N_12941);
and U13029 (N_13029,N_12664,N_12642);
xor U13030 (N_13030,N_12908,N_12509);
nand U13031 (N_13031,N_12980,N_12988);
nand U13032 (N_13032,N_12926,N_12884);
nand U13033 (N_13033,N_12683,N_12674);
nor U13034 (N_13034,N_12766,N_12917);
xnor U13035 (N_13035,N_12658,N_12929);
xnor U13036 (N_13036,N_12685,N_12895);
and U13037 (N_13037,N_12557,N_12877);
nor U13038 (N_13038,N_12579,N_12982);
nand U13039 (N_13039,N_12580,N_12893);
nand U13040 (N_13040,N_12543,N_12947);
or U13041 (N_13041,N_12653,N_12562);
xnor U13042 (N_13042,N_12521,N_12691);
xor U13043 (N_13043,N_12602,N_12690);
nor U13044 (N_13044,N_12564,N_12639);
xor U13045 (N_13045,N_12904,N_12663);
and U13046 (N_13046,N_12552,N_12640);
nor U13047 (N_13047,N_12676,N_12985);
and U13048 (N_13048,N_12886,N_12614);
nand U13049 (N_13049,N_12587,N_12963);
xnor U13050 (N_13050,N_12554,N_12654);
nor U13051 (N_13051,N_12525,N_12921);
nand U13052 (N_13052,N_12722,N_12936);
nor U13053 (N_13053,N_12756,N_12558);
and U13054 (N_13054,N_12968,N_12918);
or U13055 (N_13055,N_12843,N_12538);
or U13056 (N_13056,N_12611,N_12616);
nor U13057 (N_13057,N_12869,N_12828);
nor U13058 (N_13058,N_12831,N_12816);
xor U13059 (N_13059,N_12739,N_12827);
nand U13060 (N_13060,N_12976,N_12594);
and U13061 (N_13061,N_12885,N_12528);
and U13062 (N_13062,N_12995,N_12514);
xnor U13063 (N_13063,N_12699,N_12850);
and U13064 (N_13064,N_12502,N_12631);
nor U13065 (N_13065,N_12555,N_12851);
or U13066 (N_13066,N_12841,N_12669);
nor U13067 (N_13067,N_12923,N_12864);
and U13068 (N_13068,N_12994,N_12794);
nor U13069 (N_13069,N_12620,N_12842);
xnor U13070 (N_13070,N_12720,N_12612);
nor U13071 (N_13071,N_12629,N_12617);
nor U13072 (N_13072,N_12544,N_12732);
nand U13073 (N_13073,N_12651,N_12873);
and U13074 (N_13074,N_12530,N_12858);
nor U13075 (N_13075,N_12849,N_12799);
xor U13076 (N_13076,N_12624,N_12753);
nand U13077 (N_13077,N_12656,N_12898);
nand U13078 (N_13078,N_12761,N_12608);
and U13079 (N_13079,N_12572,N_12513);
nand U13080 (N_13080,N_12578,N_12511);
or U13081 (N_13081,N_12504,N_12583);
or U13082 (N_13082,N_12660,N_12711);
or U13083 (N_13083,N_12894,N_12848);
and U13084 (N_13084,N_12574,N_12678);
nor U13085 (N_13085,N_12609,N_12992);
nor U13086 (N_13086,N_12772,N_12830);
and U13087 (N_13087,N_12782,N_12906);
xor U13088 (N_13088,N_12506,N_12943);
and U13089 (N_13089,N_12760,N_12679);
and U13090 (N_13090,N_12803,N_12997);
xnor U13091 (N_13091,N_12695,N_12747);
nor U13092 (N_13092,N_12500,N_12966);
xor U13093 (N_13093,N_12623,N_12710);
and U13094 (N_13094,N_12672,N_12702);
nand U13095 (N_13095,N_12582,N_12954);
nand U13096 (N_13096,N_12836,N_12840);
nand U13097 (N_13097,N_12556,N_12802);
or U13098 (N_13098,N_12713,N_12726);
or U13099 (N_13099,N_12689,N_12868);
and U13100 (N_13100,N_12812,N_12969);
nor U13101 (N_13101,N_12878,N_12667);
and U13102 (N_13102,N_12650,N_12854);
or U13103 (N_13103,N_12834,N_12698);
xor U13104 (N_13104,N_12939,N_12570);
nor U13105 (N_13105,N_12591,N_12974);
or U13106 (N_13106,N_12529,N_12527);
or U13107 (N_13107,N_12984,N_12568);
nand U13108 (N_13108,N_12887,N_12673);
xor U13109 (N_13109,N_12890,N_12978);
nor U13110 (N_13110,N_12870,N_12838);
and U13111 (N_13111,N_12703,N_12659);
and U13112 (N_13112,N_12522,N_12964);
nor U13113 (N_13113,N_12607,N_12927);
nand U13114 (N_13114,N_12649,N_12585);
nand U13115 (N_13115,N_12910,N_12945);
xnor U13116 (N_13116,N_12603,N_12606);
or U13117 (N_13117,N_12814,N_12889);
or U13118 (N_13118,N_12619,N_12736);
nand U13119 (N_13119,N_12692,N_12809);
nor U13120 (N_13120,N_12643,N_12542);
xor U13121 (N_13121,N_12961,N_12820);
or U13122 (N_13122,N_12520,N_12787);
xor U13123 (N_13123,N_12539,N_12930);
xor U13124 (N_13124,N_12973,N_12902);
and U13125 (N_13125,N_12645,N_12721);
nand U13126 (N_13126,N_12741,N_12916);
xnor U13127 (N_13127,N_12531,N_12833);
nor U13128 (N_13128,N_12953,N_12971);
or U13129 (N_13129,N_12566,N_12666);
nand U13130 (N_13130,N_12990,N_12680);
nand U13131 (N_13131,N_12626,N_12777);
xor U13132 (N_13132,N_12706,N_12536);
or U13133 (N_13133,N_12765,N_12610);
nor U13134 (N_13134,N_12955,N_12781);
and U13135 (N_13135,N_12712,N_12754);
xor U13136 (N_13136,N_12588,N_12738);
nor U13137 (N_13137,N_12892,N_12745);
nand U13138 (N_13138,N_12832,N_12670);
nor U13139 (N_13139,N_12905,N_12724);
or U13140 (N_13140,N_12646,N_12567);
nor U13141 (N_13141,N_12637,N_12790);
nor U13142 (N_13142,N_12665,N_12604);
or U13143 (N_13143,N_12779,N_12792);
xor U13144 (N_13144,N_12857,N_12684);
nand U13145 (N_13145,N_12524,N_12935);
or U13146 (N_13146,N_12897,N_12737);
nor U13147 (N_13147,N_12881,N_12875);
xor U13148 (N_13148,N_12682,N_12694);
xnor U13149 (N_13149,N_12863,N_12847);
nand U13150 (N_13150,N_12882,N_12605);
nand U13151 (N_13151,N_12796,N_12959);
xor U13152 (N_13152,N_12776,N_12852);
xor U13153 (N_13153,N_12937,N_12534);
nor U13154 (N_13154,N_12715,N_12821);
and U13155 (N_13155,N_12758,N_12773);
nor U13156 (N_13156,N_12576,N_12883);
nor U13157 (N_13157,N_12647,N_12783);
or U13158 (N_13158,N_12791,N_12835);
or U13159 (N_13159,N_12950,N_12951);
and U13160 (N_13160,N_12987,N_12744);
and U13161 (N_13161,N_12805,N_12763);
nand U13162 (N_13162,N_12846,N_12668);
or U13163 (N_13163,N_12810,N_12503);
xnor U13164 (N_13164,N_12901,N_12662);
nand U13165 (N_13165,N_12770,N_12598);
and U13166 (N_13166,N_12584,N_12734);
xnor U13167 (N_13167,N_12547,N_12633);
nand U13168 (N_13168,N_12824,N_12933);
nor U13169 (N_13169,N_12535,N_12934);
or U13170 (N_13170,N_12618,N_12751);
and U13171 (N_13171,N_12537,N_12853);
nand U13172 (N_13172,N_12798,N_12775);
nand U13173 (N_13173,N_12731,N_12625);
and U13174 (N_13174,N_12746,N_12526);
nand U13175 (N_13175,N_12597,N_12733);
nor U13176 (N_13176,N_12728,N_12911);
and U13177 (N_13177,N_12778,N_12743);
nand U13178 (N_13178,N_12634,N_12806);
or U13179 (N_13179,N_12872,N_12804);
xor U13180 (N_13180,N_12983,N_12518);
xor U13181 (N_13181,N_12697,N_12581);
xnor U13182 (N_13182,N_12940,N_12590);
and U13183 (N_13183,N_12635,N_12866);
nand U13184 (N_13184,N_12823,N_12671);
nand U13185 (N_13185,N_12546,N_12915);
xnor U13186 (N_13186,N_12786,N_12948);
xor U13187 (N_13187,N_12891,N_12627);
nand U13188 (N_13188,N_12856,N_12719);
xnor U13189 (N_13189,N_12913,N_12767);
nor U13190 (N_13190,N_12541,N_12648);
nand U13191 (N_13191,N_12880,N_12845);
nor U13192 (N_13192,N_12559,N_12723);
nor U13193 (N_13193,N_12652,N_12819);
nor U13194 (N_13194,N_12920,N_12975);
and U13195 (N_13195,N_12788,N_12928);
and U13196 (N_13196,N_12601,N_12986);
nor U13197 (N_13197,N_12784,N_12979);
nor U13198 (N_13198,N_12962,N_12599);
nor U13199 (N_13199,N_12996,N_12914);
or U13200 (N_13200,N_12879,N_12825);
nand U13201 (N_13201,N_12813,N_12586);
xnor U13202 (N_13202,N_12553,N_12793);
nor U13203 (N_13203,N_12903,N_12970);
xor U13204 (N_13204,N_12909,N_12709);
xnor U13205 (N_13205,N_12630,N_12764);
nor U13206 (N_13206,N_12797,N_12859);
or U13207 (N_13207,N_12922,N_12661);
or U13208 (N_13208,N_12704,N_12912);
nand U13209 (N_13209,N_12755,N_12540);
nand U13210 (N_13210,N_12718,N_12628);
or U13211 (N_13211,N_12801,N_12615);
or U13212 (N_13212,N_12729,N_12508);
nand U13213 (N_13213,N_12811,N_12998);
and U13214 (N_13214,N_12956,N_12549);
or U13215 (N_13215,N_12705,N_12944);
xnor U13216 (N_13216,N_12952,N_12641);
or U13217 (N_13217,N_12774,N_12688);
nor U13218 (N_13218,N_12991,N_12981);
and U13219 (N_13219,N_12510,N_12696);
xor U13220 (N_13220,N_12862,N_12876);
xnor U13221 (N_13221,N_12958,N_12577);
and U13222 (N_13222,N_12561,N_12750);
and U13223 (N_13223,N_12844,N_12675);
nor U13224 (N_13224,N_12967,N_12907);
and U13225 (N_13225,N_12622,N_12523);
nand U13226 (N_13226,N_12545,N_12826);
and U13227 (N_13227,N_12740,N_12638);
and U13228 (N_13228,N_12717,N_12900);
and U13229 (N_13229,N_12632,N_12865);
and U13230 (N_13230,N_12505,N_12861);
nor U13231 (N_13231,N_12501,N_12871);
xnor U13232 (N_13232,N_12707,N_12532);
and U13233 (N_13233,N_12949,N_12960);
or U13234 (N_13234,N_12681,N_12613);
and U13235 (N_13235,N_12771,N_12533);
or U13236 (N_13236,N_12855,N_12701);
and U13237 (N_13237,N_12592,N_12507);
and U13238 (N_13238,N_12815,N_12550);
xnor U13239 (N_13239,N_12575,N_12867);
or U13240 (N_13240,N_12925,N_12749);
and U13241 (N_13241,N_12700,N_12560);
and U13242 (N_13242,N_12932,N_12600);
nor U13243 (N_13243,N_12693,N_12548);
nand U13244 (N_13244,N_12931,N_12752);
xnor U13245 (N_13245,N_12595,N_12822);
xnor U13246 (N_13246,N_12655,N_12716);
or U13247 (N_13247,N_12785,N_12748);
nand U13248 (N_13248,N_12725,N_12762);
nand U13249 (N_13249,N_12515,N_12686);
nor U13250 (N_13250,N_12987,N_12686);
xnor U13251 (N_13251,N_12519,N_12920);
or U13252 (N_13252,N_12937,N_12511);
nand U13253 (N_13253,N_12978,N_12581);
nand U13254 (N_13254,N_12812,N_12799);
or U13255 (N_13255,N_12759,N_12650);
nor U13256 (N_13256,N_12674,N_12775);
and U13257 (N_13257,N_12924,N_12631);
nand U13258 (N_13258,N_12697,N_12968);
xnor U13259 (N_13259,N_12978,N_12660);
xor U13260 (N_13260,N_12539,N_12927);
xor U13261 (N_13261,N_12898,N_12690);
nand U13262 (N_13262,N_12916,N_12610);
and U13263 (N_13263,N_12526,N_12521);
and U13264 (N_13264,N_12648,N_12640);
xnor U13265 (N_13265,N_12671,N_12887);
or U13266 (N_13266,N_12845,N_12964);
nand U13267 (N_13267,N_12503,N_12562);
or U13268 (N_13268,N_12578,N_12781);
or U13269 (N_13269,N_12933,N_12978);
or U13270 (N_13270,N_12969,N_12803);
and U13271 (N_13271,N_12739,N_12578);
and U13272 (N_13272,N_12886,N_12956);
xnor U13273 (N_13273,N_12613,N_12710);
xnor U13274 (N_13274,N_12815,N_12638);
nand U13275 (N_13275,N_12743,N_12985);
and U13276 (N_13276,N_12718,N_12968);
or U13277 (N_13277,N_12859,N_12647);
nor U13278 (N_13278,N_12540,N_12567);
and U13279 (N_13279,N_12968,N_12554);
and U13280 (N_13280,N_12720,N_12706);
nor U13281 (N_13281,N_12891,N_12779);
xnor U13282 (N_13282,N_12664,N_12674);
xor U13283 (N_13283,N_12914,N_12753);
and U13284 (N_13284,N_12608,N_12799);
nor U13285 (N_13285,N_12749,N_12640);
or U13286 (N_13286,N_12964,N_12769);
xor U13287 (N_13287,N_12515,N_12991);
or U13288 (N_13288,N_12698,N_12551);
nand U13289 (N_13289,N_12515,N_12649);
and U13290 (N_13290,N_12518,N_12733);
and U13291 (N_13291,N_12623,N_12544);
or U13292 (N_13292,N_12931,N_12946);
nor U13293 (N_13293,N_12936,N_12918);
nor U13294 (N_13294,N_12959,N_12560);
or U13295 (N_13295,N_12758,N_12529);
nand U13296 (N_13296,N_12602,N_12932);
xnor U13297 (N_13297,N_12824,N_12696);
xor U13298 (N_13298,N_12641,N_12528);
or U13299 (N_13299,N_12811,N_12766);
or U13300 (N_13300,N_12948,N_12686);
xor U13301 (N_13301,N_12520,N_12681);
nor U13302 (N_13302,N_12815,N_12819);
and U13303 (N_13303,N_12851,N_12500);
or U13304 (N_13304,N_12599,N_12800);
nor U13305 (N_13305,N_12802,N_12775);
and U13306 (N_13306,N_12950,N_12765);
and U13307 (N_13307,N_12555,N_12689);
xor U13308 (N_13308,N_12863,N_12533);
nand U13309 (N_13309,N_12928,N_12938);
or U13310 (N_13310,N_12675,N_12997);
xor U13311 (N_13311,N_12592,N_12541);
or U13312 (N_13312,N_12587,N_12529);
xnor U13313 (N_13313,N_12739,N_12708);
and U13314 (N_13314,N_12558,N_12912);
and U13315 (N_13315,N_12631,N_12524);
or U13316 (N_13316,N_12905,N_12670);
nand U13317 (N_13317,N_12625,N_12634);
or U13318 (N_13318,N_12557,N_12906);
nor U13319 (N_13319,N_12914,N_12965);
and U13320 (N_13320,N_12705,N_12801);
and U13321 (N_13321,N_12682,N_12632);
and U13322 (N_13322,N_12761,N_12780);
nand U13323 (N_13323,N_12622,N_12911);
and U13324 (N_13324,N_12702,N_12817);
nor U13325 (N_13325,N_12700,N_12751);
xor U13326 (N_13326,N_12785,N_12792);
nor U13327 (N_13327,N_12721,N_12699);
or U13328 (N_13328,N_12849,N_12705);
nor U13329 (N_13329,N_12915,N_12561);
nand U13330 (N_13330,N_12657,N_12783);
nor U13331 (N_13331,N_12562,N_12516);
xnor U13332 (N_13332,N_12644,N_12659);
nor U13333 (N_13333,N_12773,N_12830);
and U13334 (N_13334,N_12985,N_12751);
or U13335 (N_13335,N_12555,N_12926);
and U13336 (N_13336,N_12851,N_12798);
xnor U13337 (N_13337,N_12711,N_12777);
nor U13338 (N_13338,N_12983,N_12768);
xnor U13339 (N_13339,N_12562,N_12538);
nand U13340 (N_13340,N_12808,N_12878);
xnor U13341 (N_13341,N_12905,N_12749);
and U13342 (N_13342,N_12903,N_12583);
or U13343 (N_13343,N_12820,N_12552);
nor U13344 (N_13344,N_12881,N_12882);
or U13345 (N_13345,N_12795,N_12530);
nand U13346 (N_13346,N_12822,N_12588);
nand U13347 (N_13347,N_12680,N_12575);
xnor U13348 (N_13348,N_12912,N_12823);
and U13349 (N_13349,N_12734,N_12986);
nand U13350 (N_13350,N_12614,N_12812);
or U13351 (N_13351,N_12637,N_12639);
or U13352 (N_13352,N_12814,N_12711);
and U13353 (N_13353,N_12785,N_12931);
xor U13354 (N_13354,N_12728,N_12723);
nand U13355 (N_13355,N_12950,N_12838);
xor U13356 (N_13356,N_12977,N_12753);
xor U13357 (N_13357,N_12652,N_12937);
and U13358 (N_13358,N_12874,N_12974);
nor U13359 (N_13359,N_12757,N_12649);
nor U13360 (N_13360,N_12612,N_12988);
nand U13361 (N_13361,N_12523,N_12926);
xnor U13362 (N_13362,N_12825,N_12587);
nand U13363 (N_13363,N_12833,N_12674);
xor U13364 (N_13364,N_12767,N_12791);
and U13365 (N_13365,N_12530,N_12583);
xor U13366 (N_13366,N_12883,N_12586);
xnor U13367 (N_13367,N_12643,N_12780);
or U13368 (N_13368,N_12798,N_12888);
nand U13369 (N_13369,N_12564,N_12953);
xor U13370 (N_13370,N_12967,N_12925);
or U13371 (N_13371,N_12612,N_12710);
nand U13372 (N_13372,N_12539,N_12592);
xor U13373 (N_13373,N_12557,N_12814);
and U13374 (N_13374,N_12542,N_12902);
nand U13375 (N_13375,N_12879,N_12672);
nand U13376 (N_13376,N_12841,N_12730);
xnor U13377 (N_13377,N_12946,N_12648);
nor U13378 (N_13378,N_12667,N_12856);
nor U13379 (N_13379,N_12578,N_12783);
and U13380 (N_13380,N_12761,N_12692);
xnor U13381 (N_13381,N_12506,N_12912);
nand U13382 (N_13382,N_12690,N_12529);
nand U13383 (N_13383,N_12577,N_12857);
and U13384 (N_13384,N_12851,N_12896);
nor U13385 (N_13385,N_12951,N_12869);
nand U13386 (N_13386,N_12785,N_12949);
or U13387 (N_13387,N_12669,N_12671);
nand U13388 (N_13388,N_12768,N_12545);
and U13389 (N_13389,N_12521,N_12972);
or U13390 (N_13390,N_12520,N_12940);
nand U13391 (N_13391,N_12682,N_12731);
nor U13392 (N_13392,N_12637,N_12992);
nand U13393 (N_13393,N_12721,N_12584);
nand U13394 (N_13394,N_12822,N_12680);
nand U13395 (N_13395,N_12670,N_12922);
nand U13396 (N_13396,N_12948,N_12516);
nor U13397 (N_13397,N_12743,N_12995);
nor U13398 (N_13398,N_12764,N_12911);
nor U13399 (N_13399,N_12845,N_12730);
xor U13400 (N_13400,N_12907,N_12771);
xnor U13401 (N_13401,N_12783,N_12557);
nor U13402 (N_13402,N_12665,N_12872);
nor U13403 (N_13403,N_12581,N_12896);
xnor U13404 (N_13404,N_12707,N_12686);
or U13405 (N_13405,N_12596,N_12716);
xnor U13406 (N_13406,N_12582,N_12936);
xor U13407 (N_13407,N_12857,N_12591);
and U13408 (N_13408,N_12871,N_12543);
or U13409 (N_13409,N_12568,N_12580);
xnor U13410 (N_13410,N_12648,N_12815);
nand U13411 (N_13411,N_12752,N_12626);
and U13412 (N_13412,N_12675,N_12673);
or U13413 (N_13413,N_12980,N_12733);
or U13414 (N_13414,N_12608,N_12886);
and U13415 (N_13415,N_12752,N_12637);
and U13416 (N_13416,N_12616,N_12631);
or U13417 (N_13417,N_12786,N_12811);
xnor U13418 (N_13418,N_12623,N_12597);
nand U13419 (N_13419,N_12904,N_12867);
nor U13420 (N_13420,N_12752,N_12689);
nor U13421 (N_13421,N_12508,N_12863);
nor U13422 (N_13422,N_12971,N_12717);
nor U13423 (N_13423,N_12520,N_12992);
nor U13424 (N_13424,N_12932,N_12755);
or U13425 (N_13425,N_12679,N_12697);
nor U13426 (N_13426,N_12900,N_12658);
xor U13427 (N_13427,N_12585,N_12535);
and U13428 (N_13428,N_12818,N_12701);
xor U13429 (N_13429,N_12982,N_12585);
xor U13430 (N_13430,N_12666,N_12976);
nor U13431 (N_13431,N_12873,N_12614);
nor U13432 (N_13432,N_12733,N_12756);
xor U13433 (N_13433,N_12805,N_12519);
xnor U13434 (N_13434,N_12691,N_12815);
and U13435 (N_13435,N_12825,N_12924);
and U13436 (N_13436,N_12675,N_12904);
and U13437 (N_13437,N_12969,N_12839);
nor U13438 (N_13438,N_12882,N_12760);
or U13439 (N_13439,N_12966,N_12761);
nor U13440 (N_13440,N_12648,N_12713);
or U13441 (N_13441,N_12634,N_12525);
or U13442 (N_13442,N_12624,N_12519);
or U13443 (N_13443,N_12540,N_12526);
nand U13444 (N_13444,N_12537,N_12655);
or U13445 (N_13445,N_12978,N_12965);
or U13446 (N_13446,N_12695,N_12791);
nand U13447 (N_13447,N_12986,N_12702);
nor U13448 (N_13448,N_12900,N_12835);
or U13449 (N_13449,N_12585,N_12794);
xnor U13450 (N_13450,N_12843,N_12814);
nand U13451 (N_13451,N_12599,N_12897);
xnor U13452 (N_13452,N_12921,N_12635);
or U13453 (N_13453,N_12733,N_12662);
nor U13454 (N_13454,N_12584,N_12595);
or U13455 (N_13455,N_12509,N_12610);
xor U13456 (N_13456,N_12926,N_12562);
nand U13457 (N_13457,N_12737,N_12872);
and U13458 (N_13458,N_12937,N_12692);
nand U13459 (N_13459,N_12775,N_12730);
nor U13460 (N_13460,N_12793,N_12695);
and U13461 (N_13461,N_12869,N_12557);
or U13462 (N_13462,N_12637,N_12837);
nor U13463 (N_13463,N_12631,N_12966);
and U13464 (N_13464,N_12742,N_12645);
nand U13465 (N_13465,N_12807,N_12797);
xor U13466 (N_13466,N_12757,N_12828);
xnor U13467 (N_13467,N_12600,N_12746);
xor U13468 (N_13468,N_12936,N_12585);
nor U13469 (N_13469,N_12659,N_12820);
xor U13470 (N_13470,N_12798,N_12774);
or U13471 (N_13471,N_12508,N_12603);
and U13472 (N_13472,N_12694,N_12787);
xor U13473 (N_13473,N_12803,N_12942);
nand U13474 (N_13474,N_12891,N_12887);
nand U13475 (N_13475,N_12970,N_12586);
or U13476 (N_13476,N_12827,N_12922);
nor U13477 (N_13477,N_12938,N_12501);
xor U13478 (N_13478,N_12613,N_12628);
nor U13479 (N_13479,N_12524,N_12605);
xnor U13480 (N_13480,N_12743,N_12939);
or U13481 (N_13481,N_12658,N_12760);
or U13482 (N_13482,N_12910,N_12712);
xnor U13483 (N_13483,N_12520,N_12718);
nor U13484 (N_13484,N_12611,N_12917);
nor U13485 (N_13485,N_12614,N_12849);
and U13486 (N_13486,N_12596,N_12626);
xor U13487 (N_13487,N_12670,N_12954);
nor U13488 (N_13488,N_12915,N_12726);
or U13489 (N_13489,N_12895,N_12543);
nand U13490 (N_13490,N_12533,N_12811);
xor U13491 (N_13491,N_12844,N_12649);
nor U13492 (N_13492,N_12982,N_12976);
and U13493 (N_13493,N_12966,N_12948);
and U13494 (N_13494,N_12722,N_12619);
or U13495 (N_13495,N_12926,N_12724);
and U13496 (N_13496,N_12932,N_12746);
nand U13497 (N_13497,N_12965,N_12899);
xor U13498 (N_13498,N_12710,N_12518);
nand U13499 (N_13499,N_12754,N_12583);
nor U13500 (N_13500,N_13048,N_13068);
xnor U13501 (N_13501,N_13066,N_13255);
xnor U13502 (N_13502,N_13455,N_13220);
or U13503 (N_13503,N_13184,N_13069);
nor U13504 (N_13504,N_13326,N_13350);
nand U13505 (N_13505,N_13451,N_13264);
xnor U13506 (N_13506,N_13034,N_13221);
nor U13507 (N_13507,N_13022,N_13115);
or U13508 (N_13508,N_13174,N_13027);
xor U13509 (N_13509,N_13037,N_13071);
or U13510 (N_13510,N_13269,N_13017);
and U13511 (N_13511,N_13003,N_13143);
nand U13512 (N_13512,N_13147,N_13236);
and U13513 (N_13513,N_13279,N_13043);
nor U13514 (N_13514,N_13086,N_13189);
or U13515 (N_13515,N_13408,N_13010);
and U13516 (N_13516,N_13134,N_13401);
nor U13517 (N_13517,N_13302,N_13435);
and U13518 (N_13518,N_13132,N_13493);
and U13519 (N_13519,N_13073,N_13310);
nand U13520 (N_13520,N_13213,N_13433);
nand U13521 (N_13521,N_13355,N_13489);
and U13522 (N_13522,N_13207,N_13397);
or U13523 (N_13523,N_13060,N_13178);
and U13524 (N_13524,N_13338,N_13212);
and U13525 (N_13525,N_13271,N_13137);
nor U13526 (N_13526,N_13230,N_13026);
nor U13527 (N_13527,N_13331,N_13488);
nor U13528 (N_13528,N_13272,N_13280);
nor U13529 (N_13529,N_13064,N_13361);
nand U13530 (N_13530,N_13124,N_13434);
nand U13531 (N_13531,N_13468,N_13226);
or U13532 (N_13532,N_13033,N_13393);
nand U13533 (N_13533,N_13395,N_13238);
or U13534 (N_13534,N_13363,N_13260);
nor U13535 (N_13535,N_13047,N_13299);
or U13536 (N_13536,N_13389,N_13459);
or U13537 (N_13537,N_13157,N_13456);
xnor U13538 (N_13538,N_13254,N_13411);
or U13539 (N_13539,N_13258,N_13002);
nor U13540 (N_13540,N_13369,N_13289);
xor U13541 (N_13541,N_13076,N_13441);
and U13542 (N_13542,N_13392,N_13407);
or U13543 (N_13543,N_13123,N_13497);
and U13544 (N_13544,N_13443,N_13371);
nor U13545 (N_13545,N_13245,N_13243);
nor U13546 (N_13546,N_13130,N_13466);
or U13547 (N_13547,N_13422,N_13428);
nor U13548 (N_13548,N_13463,N_13417);
or U13549 (N_13549,N_13112,N_13253);
nor U13550 (N_13550,N_13045,N_13172);
and U13551 (N_13551,N_13372,N_13335);
xor U13552 (N_13552,N_13241,N_13276);
and U13553 (N_13553,N_13259,N_13457);
nor U13554 (N_13554,N_13256,N_13185);
and U13555 (N_13555,N_13458,N_13445);
and U13556 (N_13556,N_13117,N_13050);
nand U13557 (N_13557,N_13474,N_13227);
xor U13558 (N_13558,N_13291,N_13467);
or U13559 (N_13559,N_13019,N_13431);
or U13560 (N_13560,N_13074,N_13345);
nor U13561 (N_13561,N_13438,N_13413);
or U13562 (N_13562,N_13290,N_13181);
xor U13563 (N_13563,N_13358,N_13439);
nor U13564 (N_13564,N_13078,N_13054);
nor U13565 (N_13565,N_13469,N_13183);
nor U13566 (N_13566,N_13107,N_13442);
and U13567 (N_13567,N_13266,N_13426);
nor U13568 (N_13568,N_13315,N_13347);
or U13569 (N_13569,N_13378,N_13138);
xor U13570 (N_13570,N_13316,N_13101);
and U13571 (N_13571,N_13484,N_13400);
nor U13572 (N_13572,N_13496,N_13150);
or U13573 (N_13573,N_13287,N_13175);
nor U13574 (N_13574,N_13306,N_13399);
xor U13575 (N_13575,N_13224,N_13121);
xor U13576 (N_13576,N_13294,N_13268);
nand U13577 (N_13577,N_13228,N_13454);
xnor U13578 (N_13578,N_13041,N_13270);
or U13579 (N_13579,N_13232,N_13148);
nand U13580 (N_13580,N_13229,N_13349);
nand U13581 (N_13581,N_13359,N_13402);
and U13582 (N_13582,N_13007,N_13160);
nor U13583 (N_13583,N_13430,N_13028);
xnor U13584 (N_13584,N_13406,N_13379);
nand U13585 (N_13585,N_13244,N_13490);
nand U13586 (N_13586,N_13444,N_13154);
xnor U13587 (N_13587,N_13165,N_13367);
and U13588 (N_13588,N_13014,N_13267);
and U13589 (N_13589,N_13319,N_13095);
xnor U13590 (N_13590,N_13263,N_13472);
or U13591 (N_13591,N_13352,N_13257);
and U13592 (N_13592,N_13199,N_13087);
or U13593 (N_13593,N_13437,N_13161);
and U13594 (N_13594,N_13390,N_13159);
nand U13595 (N_13595,N_13478,N_13204);
nand U13596 (N_13596,N_13385,N_13333);
nand U13597 (N_13597,N_13317,N_13274);
or U13598 (N_13598,N_13099,N_13155);
and U13599 (N_13599,N_13334,N_13125);
xor U13600 (N_13600,N_13169,N_13214);
xor U13601 (N_13601,N_13351,N_13119);
and U13602 (N_13602,N_13176,N_13193);
and U13603 (N_13603,N_13336,N_13133);
and U13604 (N_13604,N_13200,N_13421);
and U13605 (N_13605,N_13035,N_13140);
and U13606 (N_13606,N_13149,N_13360);
and U13607 (N_13607,N_13219,N_13065);
xor U13608 (N_13608,N_13151,N_13348);
and U13609 (N_13609,N_13031,N_13006);
or U13610 (N_13610,N_13203,N_13483);
and U13611 (N_13611,N_13011,N_13072);
nand U13612 (N_13612,N_13144,N_13320);
and U13613 (N_13613,N_13039,N_13303);
xnor U13614 (N_13614,N_13001,N_13201);
or U13615 (N_13615,N_13288,N_13323);
or U13616 (N_13616,N_13215,N_13314);
or U13617 (N_13617,N_13242,N_13362);
xor U13618 (N_13618,N_13479,N_13285);
or U13619 (N_13619,N_13491,N_13225);
and U13620 (N_13620,N_13487,N_13084);
xor U13621 (N_13621,N_13449,N_13322);
and U13622 (N_13622,N_13436,N_13388);
and U13623 (N_13623,N_13180,N_13067);
xnor U13624 (N_13624,N_13195,N_13312);
xor U13625 (N_13625,N_13305,N_13108);
nor U13626 (N_13626,N_13321,N_13246);
nor U13627 (N_13627,N_13146,N_13222);
nor U13628 (N_13628,N_13296,N_13191);
xor U13629 (N_13629,N_13110,N_13208);
and U13630 (N_13630,N_13364,N_13261);
nand U13631 (N_13631,N_13109,N_13168);
xor U13632 (N_13632,N_13082,N_13330);
or U13633 (N_13633,N_13136,N_13218);
nor U13634 (N_13634,N_13300,N_13324);
nand U13635 (N_13635,N_13286,N_13453);
nor U13636 (N_13636,N_13089,N_13036);
nand U13637 (N_13637,N_13403,N_13394);
xnor U13638 (N_13638,N_13366,N_13234);
xnor U13639 (N_13639,N_13091,N_13104);
or U13640 (N_13640,N_13318,N_13063);
nand U13641 (N_13641,N_13171,N_13308);
and U13642 (N_13642,N_13309,N_13432);
nand U13643 (N_13643,N_13052,N_13410);
xnor U13644 (N_13644,N_13032,N_13325);
nand U13645 (N_13645,N_13423,N_13145);
or U13646 (N_13646,N_13081,N_13216);
nand U13647 (N_13647,N_13384,N_13197);
nor U13648 (N_13648,N_13179,N_13008);
and U13649 (N_13649,N_13342,N_13278);
nand U13650 (N_13650,N_13190,N_13000);
nor U13651 (N_13651,N_13495,N_13102);
xor U13652 (N_13652,N_13059,N_13103);
and U13653 (N_13653,N_13141,N_13249);
xor U13654 (N_13654,N_13235,N_13370);
and U13655 (N_13655,N_13482,N_13485);
and U13656 (N_13656,N_13038,N_13339);
or U13657 (N_13657,N_13177,N_13153);
nor U13658 (N_13658,N_13111,N_13452);
nor U13659 (N_13659,N_13049,N_13284);
nor U13660 (N_13660,N_13205,N_13387);
nor U13661 (N_13661,N_13020,N_13128);
nand U13662 (N_13662,N_13327,N_13187);
nor U13663 (N_13663,N_13447,N_13373);
nand U13664 (N_13664,N_13061,N_13462);
xor U13665 (N_13665,N_13446,N_13281);
nor U13666 (N_13666,N_13016,N_13120);
xor U13667 (N_13667,N_13166,N_13062);
and U13668 (N_13668,N_13353,N_13044);
xor U13669 (N_13669,N_13156,N_13404);
xor U13670 (N_13670,N_13346,N_13233);
and U13671 (N_13671,N_13475,N_13420);
or U13672 (N_13672,N_13092,N_13051);
nand U13673 (N_13673,N_13492,N_13237);
nor U13674 (N_13674,N_13470,N_13486);
xor U13675 (N_13675,N_13398,N_13412);
nor U13676 (N_13676,N_13301,N_13298);
or U13677 (N_13677,N_13476,N_13198);
nand U13678 (N_13678,N_13498,N_13055);
nor U13679 (N_13679,N_13409,N_13277);
nand U13680 (N_13680,N_13192,N_13024);
nand U13681 (N_13681,N_13382,N_13098);
and U13682 (N_13682,N_13405,N_13013);
nor U13683 (N_13683,N_13262,N_13365);
nor U13684 (N_13684,N_13004,N_13295);
nand U13685 (N_13685,N_13162,N_13424);
or U13686 (N_13686,N_13465,N_13293);
nand U13687 (N_13687,N_13217,N_13313);
or U13688 (N_13688,N_13391,N_13223);
or U13689 (N_13689,N_13240,N_13377);
and U13690 (N_13690,N_13374,N_13211);
and U13691 (N_13691,N_13005,N_13418);
xor U13692 (N_13692,N_13058,N_13292);
nor U13693 (N_13693,N_13481,N_13196);
and U13694 (N_13694,N_13340,N_13164);
and U13695 (N_13695,N_13070,N_13448);
nor U13696 (N_13696,N_13053,N_13499);
xnor U13697 (N_13697,N_13250,N_13343);
xnor U13698 (N_13698,N_13354,N_13114);
or U13699 (N_13699,N_13015,N_13186);
nand U13700 (N_13700,N_13273,N_13332);
xnor U13701 (N_13701,N_13328,N_13009);
nand U13702 (N_13702,N_13040,N_13473);
nand U13703 (N_13703,N_13158,N_13450);
xnor U13704 (N_13704,N_13085,N_13167);
nor U13705 (N_13705,N_13173,N_13282);
or U13706 (N_13706,N_13056,N_13380);
or U13707 (N_13707,N_13080,N_13297);
or U13708 (N_13708,N_13376,N_13427);
nor U13709 (N_13709,N_13356,N_13021);
nand U13710 (N_13710,N_13093,N_13464);
xnor U13711 (N_13711,N_13097,N_13170);
nor U13712 (N_13712,N_13210,N_13096);
nor U13713 (N_13713,N_13118,N_13419);
or U13714 (N_13714,N_13029,N_13231);
or U13715 (N_13715,N_13357,N_13381);
nand U13716 (N_13716,N_13142,N_13090);
nand U13717 (N_13717,N_13152,N_13163);
and U13718 (N_13718,N_13480,N_13429);
nand U13719 (N_13719,N_13461,N_13075);
and U13720 (N_13720,N_13023,N_13460);
nor U13721 (N_13721,N_13337,N_13283);
and U13722 (N_13722,N_13239,N_13129);
or U13723 (N_13723,N_13341,N_13116);
or U13724 (N_13724,N_13202,N_13018);
nand U13725 (N_13725,N_13127,N_13304);
xnor U13726 (N_13726,N_13025,N_13126);
nor U13727 (N_13727,N_13139,N_13042);
nand U13728 (N_13728,N_13135,N_13386);
nand U13729 (N_13729,N_13106,N_13113);
or U13730 (N_13730,N_13368,N_13105);
nand U13731 (N_13731,N_13307,N_13030);
xnor U13732 (N_13732,N_13209,N_13252);
nor U13733 (N_13733,N_13344,N_13415);
nand U13734 (N_13734,N_13329,N_13077);
nand U13735 (N_13735,N_13416,N_13425);
or U13736 (N_13736,N_13079,N_13057);
xor U13737 (N_13737,N_13046,N_13012);
and U13738 (N_13738,N_13083,N_13206);
or U13739 (N_13739,N_13182,N_13440);
or U13740 (N_13740,N_13383,N_13122);
or U13741 (N_13741,N_13265,N_13251);
nor U13742 (N_13742,N_13471,N_13477);
nand U13743 (N_13743,N_13088,N_13311);
and U13744 (N_13744,N_13375,N_13194);
and U13745 (N_13745,N_13188,N_13494);
xor U13746 (N_13746,N_13131,N_13248);
and U13747 (N_13747,N_13100,N_13247);
nor U13748 (N_13748,N_13396,N_13414);
or U13749 (N_13749,N_13275,N_13094);
or U13750 (N_13750,N_13474,N_13137);
nor U13751 (N_13751,N_13178,N_13308);
nor U13752 (N_13752,N_13186,N_13482);
and U13753 (N_13753,N_13368,N_13299);
or U13754 (N_13754,N_13199,N_13045);
xor U13755 (N_13755,N_13064,N_13109);
or U13756 (N_13756,N_13334,N_13166);
nand U13757 (N_13757,N_13335,N_13223);
xnor U13758 (N_13758,N_13438,N_13381);
nor U13759 (N_13759,N_13160,N_13249);
nand U13760 (N_13760,N_13281,N_13331);
and U13761 (N_13761,N_13103,N_13480);
or U13762 (N_13762,N_13315,N_13460);
and U13763 (N_13763,N_13380,N_13176);
or U13764 (N_13764,N_13420,N_13395);
and U13765 (N_13765,N_13204,N_13282);
or U13766 (N_13766,N_13205,N_13333);
or U13767 (N_13767,N_13089,N_13428);
xnor U13768 (N_13768,N_13092,N_13403);
or U13769 (N_13769,N_13372,N_13348);
and U13770 (N_13770,N_13472,N_13102);
and U13771 (N_13771,N_13461,N_13496);
and U13772 (N_13772,N_13143,N_13215);
and U13773 (N_13773,N_13472,N_13221);
or U13774 (N_13774,N_13410,N_13198);
nor U13775 (N_13775,N_13184,N_13002);
xor U13776 (N_13776,N_13261,N_13146);
and U13777 (N_13777,N_13291,N_13386);
or U13778 (N_13778,N_13277,N_13464);
xor U13779 (N_13779,N_13453,N_13467);
xor U13780 (N_13780,N_13482,N_13466);
xor U13781 (N_13781,N_13462,N_13438);
and U13782 (N_13782,N_13292,N_13033);
xnor U13783 (N_13783,N_13045,N_13083);
nor U13784 (N_13784,N_13267,N_13206);
xnor U13785 (N_13785,N_13484,N_13473);
nand U13786 (N_13786,N_13161,N_13205);
nor U13787 (N_13787,N_13097,N_13062);
and U13788 (N_13788,N_13454,N_13491);
xor U13789 (N_13789,N_13002,N_13019);
and U13790 (N_13790,N_13395,N_13173);
and U13791 (N_13791,N_13047,N_13157);
nor U13792 (N_13792,N_13403,N_13057);
or U13793 (N_13793,N_13188,N_13190);
or U13794 (N_13794,N_13464,N_13039);
nor U13795 (N_13795,N_13229,N_13233);
and U13796 (N_13796,N_13041,N_13426);
nand U13797 (N_13797,N_13314,N_13179);
xor U13798 (N_13798,N_13083,N_13376);
xnor U13799 (N_13799,N_13430,N_13367);
nand U13800 (N_13800,N_13113,N_13361);
nor U13801 (N_13801,N_13248,N_13421);
and U13802 (N_13802,N_13080,N_13226);
nand U13803 (N_13803,N_13443,N_13126);
nor U13804 (N_13804,N_13437,N_13306);
nor U13805 (N_13805,N_13320,N_13457);
and U13806 (N_13806,N_13316,N_13392);
nor U13807 (N_13807,N_13186,N_13101);
nand U13808 (N_13808,N_13328,N_13373);
xnor U13809 (N_13809,N_13359,N_13386);
or U13810 (N_13810,N_13493,N_13106);
or U13811 (N_13811,N_13098,N_13057);
or U13812 (N_13812,N_13452,N_13189);
and U13813 (N_13813,N_13086,N_13382);
nand U13814 (N_13814,N_13047,N_13409);
xor U13815 (N_13815,N_13151,N_13261);
and U13816 (N_13816,N_13435,N_13415);
and U13817 (N_13817,N_13440,N_13326);
or U13818 (N_13818,N_13182,N_13281);
and U13819 (N_13819,N_13165,N_13310);
nor U13820 (N_13820,N_13270,N_13057);
nand U13821 (N_13821,N_13353,N_13485);
and U13822 (N_13822,N_13153,N_13170);
nor U13823 (N_13823,N_13145,N_13195);
or U13824 (N_13824,N_13379,N_13121);
xnor U13825 (N_13825,N_13394,N_13253);
nand U13826 (N_13826,N_13368,N_13041);
nand U13827 (N_13827,N_13369,N_13254);
and U13828 (N_13828,N_13495,N_13219);
or U13829 (N_13829,N_13443,N_13343);
or U13830 (N_13830,N_13422,N_13153);
xnor U13831 (N_13831,N_13314,N_13035);
or U13832 (N_13832,N_13231,N_13276);
xor U13833 (N_13833,N_13255,N_13083);
nor U13834 (N_13834,N_13073,N_13148);
xor U13835 (N_13835,N_13357,N_13276);
nand U13836 (N_13836,N_13391,N_13064);
xnor U13837 (N_13837,N_13432,N_13043);
and U13838 (N_13838,N_13067,N_13301);
xnor U13839 (N_13839,N_13436,N_13000);
xnor U13840 (N_13840,N_13245,N_13201);
xor U13841 (N_13841,N_13055,N_13107);
xnor U13842 (N_13842,N_13190,N_13370);
xnor U13843 (N_13843,N_13061,N_13384);
and U13844 (N_13844,N_13095,N_13216);
or U13845 (N_13845,N_13312,N_13115);
and U13846 (N_13846,N_13465,N_13287);
and U13847 (N_13847,N_13254,N_13013);
or U13848 (N_13848,N_13402,N_13484);
or U13849 (N_13849,N_13358,N_13256);
nand U13850 (N_13850,N_13491,N_13330);
nand U13851 (N_13851,N_13276,N_13461);
nand U13852 (N_13852,N_13293,N_13444);
nand U13853 (N_13853,N_13055,N_13172);
xnor U13854 (N_13854,N_13495,N_13316);
xnor U13855 (N_13855,N_13156,N_13137);
nor U13856 (N_13856,N_13072,N_13205);
nand U13857 (N_13857,N_13093,N_13363);
nor U13858 (N_13858,N_13422,N_13304);
nor U13859 (N_13859,N_13328,N_13023);
xnor U13860 (N_13860,N_13364,N_13321);
nand U13861 (N_13861,N_13154,N_13424);
or U13862 (N_13862,N_13107,N_13236);
or U13863 (N_13863,N_13361,N_13173);
nand U13864 (N_13864,N_13327,N_13110);
or U13865 (N_13865,N_13057,N_13160);
nor U13866 (N_13866,N_13115,N_13098);
xnor U13867 (N_13867,N_13173,N_13000);
and U13868 (N_13868,N_13170,N_13403);
nand U13869 (N_13869,N_13423,N_13036);
and U13870 (N_13870,N_13179,N_13273);
nand U13871 (N_13871,N_13398,N_13194);
and U13872 (N_13872,N_13236,N_13496);
nor U13873 (N_13873,N_13444,N_13417);
nor U13874 (N_13874,N_13143,N_13427);
and U13875 (N_13875,N_13216,N_13467);
xor U13876 (N_13876,N_13002,N_13398);
or U13877 (N_13877,N_13337,N_13082);
and U13878 (N_13878,N_13110,N_13242);
nor U13879 (N_13879,N_13248,N_13182);
nor U13880 (N_13880,N_13458,N_13431);
nor U13881 (N_13881,N_13397,N_13392);
or U13882 (N_13882,N_13471,N_13038);
xor U13883 (N_13883,N_13493,N_13139);
or U13884 (N_13884,N_13401,N_13079);
xor U13885 (N_13885,N_13245,N_13480);
nand U13886 (N_13886,N_13050,N_13054);
nand U13887 (N_13887,N_13077,N_13042);
nand U13888 (N_13888,N_13119,N_13266);
xor U13889 (N_13889,N_13224,N_13249);
nor U13890 (N_13890,N_13307,N_13177);
xor U13891 (N_13891,N_13403,N_13277);
and U13892 (N_13892,N_13446,N_13111);
and U13893 (N_13893,N_13474,N_13494);
nor U13894 (N_13894,N_13340,N_13126);
xor U13895 (N_13895,N_13365,N_13323);
and U13896 (N_13896,N_13455,N_13225);
nor U13897 (N_13897,N_13398,N_13162);
and U13898 (N_13898,N_13375,N_13186);
or U13899 (N_13899,N_13409,N_13188);
xnor U13900 (N_13900,N_13097,N_13066);
nand U13901 (N_13901,N_13306,N_13370);
xor U13902 (N_13902,N_13071,N_13413);
xnor U13903 (N_13903,N_13213,N_13360);
nor U13904 (N_13904,N_13353,N_13351);
nand U13905 (N_13905,N_13144,N_13045);
xnor U13906 (N_13906,N_13218,N_13454);
and U13907 (N_13907,N_13492,N_13497);
or U13908 (N_13908,N_13408,N_13327);
nand U13909 (N_13909,N_13242,N_13248);
nor U13910 (N_13910,N_13201,N_13293);
nand U13911 (N_13911,N_13372,N_13179);
nand U13912 (N_13912,N_13493,N_13137);
xnor U13913 (N_13913,N_13331,N_13387);
or U13914 (N_13914,N_13114,N_13325);
or U13915 (N_13915,N_13483,N_13012);
nor U13916 (N_13916,N_13096,N_13310);
xor U13917 (N_13917,N_13247,N_13091);
xnor U13918 (N_13918,N_13416,N_13005);
and U13919 (N_13919,N_13369,N_13132);
xnor U13920 (N_13920,N_13125,N_13008);
xnor U13921 (N_13921,N_13454,N_13088);
xor U13922 (N_13922,N_13119,N_13254);
nand U13923 (N_13923,N_13487,N_13178);
and U13924 (N_13924,N_13057,N_13320);
nand U13925 (N_13925,N_13468,N_13027);
nor U13926 (N_13926,N_13474,N_13163);
or U13927 (N_13927,N_13046,N_13197);
xor U13928 (N_13928,N_13201,N_13479);
nand U13929 (N_13929,N_13005,N_13079);
or U13930 (N_13930,N_13071,N_13399);
xor U13931 (N_13931,N_13422,N_13030);
or U13932 (N_13932,N_13155,N_13068);
nor U13933 (N_13933,N_13129,N_13375);
and U13934 (N_13934,N_13443,N_13175);
nor U13935 (N_13935,N_13130,N_13252);
and U13936 (N_13936,N_13334,N_13344);
or U13937 (N_13937,N_13000,N_13326);
xnor U13938 (N_13938,N_13005,N_13469);
nand U13939 (N_13939,N_13428,N_13490);
and U13940 (N_13940,N_13074,N_13087);
nand U13941 (N_13941,N_13104,N_13258);
nor U13942 (N_13942,N_13414,N_13196);
nor U13943 (N_13943,N_13239,N_13098);
nor U13944 (N_13944,N_13441,N_13387);
xnor U13945 (N_13945,N_13229,N_13139);
nand U13946 (N_13946,N_13089,N_13279);
and U13947 (N_13947,N_13360,N_13162);
nand U13948 (N_13948,N_13067,N_13147);
xnor U13949 (N_13949,N_13216,N_13003);
and U13950 (N_13950,N_13248,N_13037);
nand U13951 (N_13951,N_13141,N_13313);
xor U13952 (N_13952,N_13250,N_13446);
nor U13953 (N_13953,N_13292,N_13201);
and U13954 (N_13954,N_13026,N_13267);
nor U13955 (N_13955,N_13351,N_13386);
nor U13956 (N_13956,N_13493,N_13101);
xnor U13957 (N_13957,N_13140,N_13064);
and U13958 (N_13958,N_13385,N_13142);
or U13959 (N_13959,N_13260,N_13048);
nand U13960 (N_13960,N_13498,N_13011);
nor U13961 (N_13961,N_13068,N_13489);
xnor U13962 (N_13962,N_13242,N_13062);
or U13963 (N_13963,N_13419,N_13051);
nor U13964 (N_13964,N_13320,N_13394);
nand U13965 (N_13965,N_13026,N_13228);
xnor U13966 (N_13966,N_13173,N_13188);
xor U13967 (N_13967,N_13291,N_13040);
xnor U13968 (N_13968,N_13433,N_13043);
nand U13969 (N_13969,N_13048,N_13429);
xor U13970 (N_13970,N_13315,N_13351);
xor U13971 (N_13971,N_13191,N_13203);
xor U13972 (N_13972,N_13495,N_13413);
xnor U13973 (N_13973,N_13268,N_13229);
and U13974 (N_13974,N_13409,N_13211);
nor U13975 (N_13975,N_13209,N_13373);
or U13976 (N_13976,N_13095,N_13224);
xnor U13977 (N_13977,N_13042,N_13105);
or U13978 (N_13978,N_13283,N_13049);
and U13979 (N_13979,N_13222,N_13046);
nor U13980 (N_13980,N_13476,N_13098);
xor U13981 (N_13981,N_13196,N_13292);
or U13982 (N_13982,N_13465,N_13103);
nand U13983 (N_13983,N_13148,N_13300);
or U13984 (N_13984,N_13386,N_13199);
xor U13985 (N_13985,N_13331,N_13332);
nand U13986 (N_13986,N_13210,N_13438);
and U13987 (N_13987,N_13221,N_13450);
or U13988 (N_13988,N_13007,N_13464);
or U13989 (N_13989,N_13059,N_13460);
nor U13990 (N_13990,N_13158,N_13044);
or U13991 (N_13991,N_13305,N_13005);
or U13992 (N_13992,N_13240,N_13054);
and U13993 (N_13993,N_13370,N_13025);
nor U13994 (N_13994,N_13285,N_13001);
or U13995 (N_13995,N_13020,N_13357);
xor U13996 (N_13996,N_13243,N_13452);
xor U13997 (N_13997,N_13020,N_13102);
nand U13998 (N_13998,N_13002,N_13353);
xor U13999 (N_13999,N_13341,N_13347);
nand U14000 (N_14000,N_13805,N_13702);
or U14001 (N_14001,N_13985,N_13789);
xnor U14002 (N_14002,N_13699,N_13882);
nor U14003 (N_14003,N_13550,N_13849);
or U14004 (N_14004,N_13724,N_13636);
nand U14005 (N_14005,N_13774,N_13828);
or U14006 (N_14006,N_13915,N_13810);
and U14007 (N_14007,N_13771,N_13895);
xor U14008 (N_14008,N_13677,N_13742);
nand U14009 (N_14009,N_13638,N_13876);
or U14010 (N_14010,N_13541,N_13544);
or U14011 (N_14011,N_13713,N_13917);
or U14012 (N_14012,N_13987,N_13512);
and U14013 (N_14013,N_13770,N_13662);
or U14014 (N_14014,N_13559,N_13634);
and U14015 (N_14015,N_13884,N_13606);
nand U14016 (N_14016,N_13936,N_13905);
nand U14017 (N_14017,N_13990,N_13957);
xor U14018 (N_14018,N_13986,N_13668);
or U14019 (N_14019,N_13598,N_13618);
xor U14020 (N_14020,N_13546,N_13747);
or U14021 (N_14021,N_13871,N_13931);
nor U14022 (N_14022,N_13651,N_13703);
nand U14023 (N_14023,N_13503,N_13996);
or U14024 (N_14024,N_13570,N_13603);
nand U14025 (N_14025,N_13942,N_13573);
nand U14026 (N_14026,N_13553,N_13617);
and U14027 (N_14027,N_13966,N_13943);
xnor U14028 (N_14028,N_13718,N_13687);
or U14029 (N_14029,N_13625,N_13822);
or U14030 (N_14030,N_13645,N_13960);
nor U14031 (N_14031,N_13949,N_13739);
xor U14032 (N_14032,N_13781,N_13650);
and U14033 (N_14033,N_13814,N_13519);
or U14034 (N_14034,N_13953,N_13902);
or U14035 (N_14035,N_13743,N_13759);
nand U14036 (N_14036,N_13552,N_13580);
xor U14037 (N_14037,N_13528,N_13578);
and U14038 (N_14038,N_13673,N_13794);
or U14039 (N_14039,N_13818,N_13850);
nor U14040 (N_14040,N_13809,N_13660);
and U14041 (N_14041,N_13562,N_13571);
nand U14042 (N_14042,N_13928,N_13522);
nand U14043 (N_14043,N_13654,N_13549);
nand U14044 (N_14044,N_13916,N_13803);
or U14045 (N_14045,N_13568,N_13577);
nand U14046 (N_14046,N_13776,N_13726);
xor U14047 (N_14047,N_13565,N_13854);
and U14048 (N_14048,N_13873,N_13678);
nand U14049 (N_14049,N_13847,N_13741);
and U14050 (N_14050,N_13526,N_13560);
and U14051 (N_14051,N_13710,N_13593);
nor U14052 (N_14052,N_13735,N_13971);
nand U14053 (N_14053,N_13633,N_13995);
or U14054 (N_14054,N_13518,N_13655);
nor U14055 (N_14055,N_13981,N_13683);
nor U14056 (N_14056,N_13701,N_13613);
nand U14057 (N_14057,N_13779,N_13764);
nand U14058 (N_14058,N_13563,N_13551);
nand U14059 (N_14059,N_13845,N_13797);
or U14060 (N_14060,N_13524,N_13783);
nand U14061 (N_14061,N_13740,N_13903);
nand U14062 (N_14062,N_13900,N_13988);
and U14063 (N_14063,N_13510,N_13534);
and U14064 (N_14064,N_13558,N_13842);
xnor U14065 (N_14065,N_13700,N_13939);
and U14066 (N_14066,N_13892,N_13937);
nor U14067 (N_14067,N_13540,N_13689);
or U14068 (N_14068,N_13501,N_13904);
nor U14069 (N_14069,N_13935,N_13542);
and U14070 (N_14070,N_13836,N_13821);
or U14071 (N_14071,N_13817,N_13858);
nor U14072 (N_14072,N_13827,N_13946);
and U14073 (N_14073,N_13793,N_13929);
nand U14074 (N_14074,N_13707,N_13736);
xor U14075 (N_14075,N_13686,N_13863);
nor U14076 (N_14076,N_13629,N_13586);
xnor U14077 (N_14077,N_13567,N_13899);
nand U14078 (N_14078,N_13866,N_13778);
or U14079 (N_14079,N_13667,N_13944);
or U14080 (N_14080,N_13891,N_13865);
or U14081 (N_14081,N_13690,N_13877);
nor U14082 (N_14082,N_13688,N_13808);
or U14083 (N_14083,N_13835,N_13509);
or U14084 (N_14084,N_13912,N_13649);
or U14085 (N_14085,N_13628,N_13555);
and U14086 (N_14086,N_13584,N_13833);
and U14087 (N_14087,N_13993,N_13983);
nor U14088 (N_14088,N_13804,N_13772);
nor U14089 (N_14089,N_13529,N_13978);
nor U14090 (N_14090,N_13914,N_13614);
or U14091 (N_14091,N_13973,N_13640);
or U14092 (N_14092,N_13753,N_13830);
or U14093 (N_14093,N_13525,N_13901);
or U14094 (N_14094,N_13922,N_13685);
and U14095 (N_14095,N_13511,N_13965);
nor U14096 (N_14096,N_13658,N_13661);
nand U14097 (N_14097,N_13870,N_13984);
nor U14098 (N_14098,N_13893,N_13920);
and U14099 (N_14099,N_13588,N_13581);
nand U14100 (N_14100,N_13720,N_13768);
xor U14101 (N_14101,N_13664,N_13755);
nor U14102 (N_14102,N_13924,N_13644);
nand U14103 (N_14103,N_13513,N_13750);
nor U14104 (N_14104,N_13692,N_13769);
xor U14105 (N_14105,N_13947,N_13765);
nand U14106 (N_14106,N_13890,N_13958);
or U14107 (N_14107,N_13516,N_13592);
or U14108 (N_14108,N_13932,N_13705);
xnor U14109 (N_14109,N_13982,N_13575);
xnor U14110 (N_14110,N_13777,N_13906);
and U14111 (N_14111,N_13583,N_13801);
or U14112 (N_14112,N_13715,N_13611);
nor U14113 (N_14113,N_13642,N_13725);
xor U14114 (N_14114,N_13786,N_13886);
or U14115 (N_14115,N_13693,N_13961);
xnor U14116 (N_14116,N_13798,N_13762);
or U14117 (N_14117,N_13969,N_13998);
nand U14118 (N_14118,N_13732,N_13523);
or U14119 (N_14119,N_13788,N_13885);
xnor U14120 (N_14120,N_13896,N_13970);
nor U14121 (N_14121,N_13761,N_13517);
xor U14122 (N_14122,N_13663,N_13545);
and U14123 (N_14123,N_13599,N_13941);
nand U14124 (N_14124,N_13864,N_13635);
and U14125 (N_14125,N_13959,N_13691);
nand U14126 (N_14126,N_13955,N_13566);
nor U14127 (N_14127,N_13733,N_13731);
xor U14128 (N_14128,N_13579,N_13682);
or U14129 (N_14129,N_13576,N_13813);
or U14130 (N_14130,N_13975,N_13952);
nor U14131 (N_14131,N_13859,N_13780);
xor U14132 (N_14132,N_13760,N_13652);
nand U14133 (N_14133,N_13766,N_13727);
nand U14134 (N_14134,N_13659,N_13819);
nand U14135 (N_14135,N_13704,N_13923);
nand U14136 (N_14136,N_13556,N_13956);
or U14137 (N_14137,N_13734,N_13737);
or U14138 (N_14138,N_13802,N_13716);
xnor U14139 (N_14139,N_13840,N_13875);
or U14140 (N_14140,N_13888,N_13601);
nor U14141 (N_14141,N_13841,N_13697);
or U14142 (N_14142,N_13880,N_13530);
nor U14143 (N_14143,N_13874,N_13527);
and U14144 (N_14144,N_13608,N_13600);
nor U14145 (N_14145,N_13826,N_13717);
xor U14146 (N_14146,N_13561,N_13878);
or U14147 (N_14147,N_13962,N_13824);
xnor U14148 (N_14148,N_13612,N_13626);
xnor U14149 (N_14149,N_13506,N_13621);
nand U14150 (N_14150,N_13911,N_13837);
nand U14151 (N_14151,N_13666,N_13507);
nand U14152 (N_14152,N_13537,N_13548);
nor U14153 (N_14153,N_13746,N_13674);
nand U14154 (N_14154,N_13994,N_13728);
or U14155 (N_14155,N_13532,N_13933);
or U14156 (N_14156,N_13812,N_13538);
nand U14157 (N_14157,N_13856,N_13616);
and U14158 (N_14158,N_13589,N_13968);
xor U14159 (N_14159,N_13590,N_13839);
nand U14160 (N_14160,N_13637,N_13773);
nand U14161 (N_14161,N_13572,N_13502);
nand U14162 (N_14162,N_13615,N_13868);
and U14163 (N_14163,N_13574,N_13521);
or U14164 (N_14164,N_13547,N_13730);
nor U14165 (N_14165,N_13684,N_13763);
nor U14166 (N_14166,N_13790,N_13921);
xor U14167 (N_14167,N_13582,N_13853);
xor U14168 (N_14168,N_13602,N_13992);
nor U14169 (N_14169,N_13520,N_13536);
xnor U14170 (N_14170,N_13627,N_13696);
and U14171 (N_14171,N_13676,N_13963);
xnor U14172 (N_14172,N_13775,N_13844);
xor U14173 (N_14173,N_13846,N_13816);
xor U14174 (N_14174,N_13729,N_13980);
or U14175 (N_14175,N_13539,N_13967);
and U14176 (N_14176,N_13504,N_13829);
or U14177 (N_14177,N_13531,N_13622);
xor U14178 (N_14178,N_13694,N_13639);
and U14179 (N_14179,N_13977,N_13754);
or U14180 (N_14180,N_13631,N_13909);
or U14181 (N_14181,N_13670,N_13831);
xnor U14182 (N_14182,N_13989,N_13533);
or U14183 (N_14183,N_13653,N_13721);
nor U14184 (N_14184,N_13596,N_13641);
and U14185 (N_14185,N_13569,N_13834);
and U14186 (N_14186,N_13825,N_13881);
or U14187 (N_14187,N_13894,N_13712);
or U14188 (N_14188,N_13974,N_13945);
and U14189 (N_14189,N_13680,N_13934);
xor U14190 (N_14190,N_13860,N_13948);
nor U14191 (N_14191,N_13869,N_13508);
nand U14192 (N_14192,N_13647,N_13999);
xor U14193 (N_14193,N_13913,N_13938);
nand U14194 (N_14194,N_13723,N_13972);
nor U14195 (N_14195,N_13706,N_13708);
xor U14196 (N_14196,N_13861,N_13675);
or U14197 (N_14197,N_13505,N_13657);
and U14198 (N_14198,N_13709,N_13609);
or U14199 (N_14199,N_13791,N_13695);
or U14200 (N_14200,N_13832,N_13738);
and U14201 (N_14201,N_13823,N_13862);
nand U14202 (N_14202,N_13807,N_13564);
nor U14203 (N_14203,N_13879,N_13554);
nand U14204 (N_14204,N_13951,N_13785);
nor U14205 (N_14205,N_13620,N_13744);
nor U14206 (N_14206,N_13648,N_13630);
nor U14207 (N_14207,N_13806,N_13979);
xnor U14208 (N_14208,N_13587,N_13787);
or U14209 (N_14209,N_13792,N_13665);
nor U14210 (N_14210,N_13883,N_13997);
and U14211 (N_14211,N_13681,N_13848);
nor U14212 (N_14212,N_13619,N_13607);
xnor U14213 (N_14213,N_13926,N_13752);
nand U14214 (N_14214,N_13643,N_13595);
xor U14215 (N_14215,N_13597,N_13679);
and U14216 (N_14216,N_13669,N_13910);
or U14217 (N_14217,N_13711,N_13820);
and U14218 (N_14218,N_13954,N_13889);
nor U14219 (N_14219,N_13795,N_13605);
and U14220 (N_14220,N_13857,N_13991);
nand U14221 (N_14221,N_13714,N_13918);
and U14222 (N_14222,N_13722,N_13623);
nand U14223 (N_14223,N_13782,N_13800);
nand U14224 (N_14224,N_13796,N_13799);
and U14225 (N_14225,N_13515,N_13610);
nand U14226 (N_14226,N_13557,N_13745);
nand U14227 (N_14227,N_13543,N_13767);
and U14228 (N_14228,N_13940,N_13964);
or U14229 (N_14229,N_13591,N_13927);
or U14230 (N_14230,N_13872,N_13851);
nor U14231 (N_14231,N_13585,N_13758);
nor U14232 (N_14232,N_13908,N_13887);
and U14233 (N_14233,N_13535,N_13656);
or U14234 (N_14234,N_13930,N_13843);
nor U14235 (N_14235,N_13698,N_13852);
nor U14236 (N_14236,N_13514,N_13751);
xor U14237 (N_14237,N_13907,N_13719);
nand U14238 (N_14238,N_13925,N_13898);
or U14239 (N_14239,N_13976,N_13784);
nand U14240 (N_14240,N_13756,N_13855);
nor U14241 (N_14241,N_13672,N_13624);
nand U14242 (N_14242,N_13594,N_13500);
and U14243 (N_14243,N_13811,N_13671);
and U14244 (N_14244,N_13867,N_13604);
and U14245 (N_14245,N_13646,N_13632);
nor U14246 (N_14246,N_13919,N_13748);
or U14247 (N_14247,N_13757,N_13815);
nand U14248 (N_14248,N_13950,N_13897);
or U14249 (N_14249,N_13838,N_13749);
or U14250 (N_14250,N_13569,N_13822);
nand U14251 (N_14251,N_13638,N_13580);
nor U14252 (N_14252,N_13980,N_13705);
xor U14253 (N_14253,N_13677,N_13684);
nand U14254 (N_14254,N_13944,N_13999);
or U14255 (N_14255,N_13596,N_13947);
xor U14256 (N_14256,N_13729,N_13551);
nor U14257 (N_14257,N_13748,N_13639);
xor U14258 (N_14258,N_13751,N_13998);
or U14259 (N_14259,N_13861,N_13896);
nand U14260 (N_14260,N_13572,N_13970);
nor U14261 (N_14261,N_13747,N_13983);
and U14262 (N_14262,N_13833,N_13859);
or U14263 (N_14263,N_13615,N_13698);
xor U14264 (N_14264,N_13516,N_13827);
and U14265 (N_14265,N_13974,N_13709);
or U14266 (N_14266,N_13804,N_13562);
or U14267 (N_14267,N_13528,N_13997);
nand U14268 (N_14268,N_13754,N_13614);
xnor U14269 (N_14269,N_13805,N_13718);
xnor U14270 (N_14270,N_13966,N_13880);
xor U14271 (N_14271,N_13964,N_13523);
and U14272 (N_14272,N_13613,N_13580);
nor U14273 (N_14273,N_13915,N_13899);
nor U14274 (N_14274,N_13910,N_13555);
nor U14275 (N_14275,N_13864,N_13512);
xor U14276 (N_14276,N_13784,N_13768);
nor U14277 (N_14277,N_13504,N_13987);
or U14278 (N_14278,N_13680,N_13809);
xnor U14279 (N_14279,N_13607,N_13946);
xnor U14280 (N_14280,N_13537,N_13747);
nor U14281 (N_14281,N_13904,N_13893);
nor U14282 (N_14282,N_13978,N_13714);
and U14283 (N_14283,N_13906,N_13862);
xnor U14284 (N_14284,N_13768,N_13806);
nor U14285 (N_14285,N_13859,N_13762);
xor U14286 (N_14286,N_13922,N_13738);
nand U14287 (N_14287,N_13592,N_13637);
or U14288 (N_14288,N_13946,N_13748);
xnor U14289 (N_14289,N_13879,N_13944);
or U14290 (N_14290,N_13692,N_13857);
xor U14291 (N_14291,N_13571,N_13530);
nand U14292 (N_14292,N_13803,N_13567);
nand U14293 (N_14293,N_13819,N_13590);
xor U14294 (N_14294,N_13745,N_13555);
and U14295 (N_14295,N_13550,N_13739);
or U14296 (N_14296,N_13967,N_13861);
and U14297 (N_14297,N_13552,N_13550);
nand U14298 (N_14298,N_13776,N_13960);
or U14299 (N_14299,N_13669,N_13872);
xor U14300 (N_14300,N_13618,N_13557);
xnor U14301 (N_14301,N_13718,N_13583);
nor U14302 (N_14302,N_13620,N_13678);
and U14303 (N_14303,N_13658,N_13706);
xor U14304 (N_14304,N_13693,N_13598);
xor U14305 (N_14305,N_13645,N_13543);
and U14306 (N_14306,N_13835,N_13686);
and U14307 (N_14307,N_13692,N_13811);
nand U14308 (N_14308,N_13724,N_13589);
nor U14309 (N_14309,N_13933,N_13577);
xor U14310 (N_14310,N_13550,N_13664);
or U14311 (N_14311,N_13590,N_13688);
nand U14312 (N_14312,N_13943,N_13577);
or U14313 (N_14313,N_13987,N_13768);
xnor U14314 (N_14314,N_13779,N_13909);
nor U14315 (N_14315,N_13727,N_13608);
nor U14316 (N_14316,N_13529,N_13783);
xor U14317 (N_14317,N_13993,N_13919);
xnor U14318 (N_14318,N_13960,N_13500);
xor U14319 (N_14319,N_13655,N_13502);
and U14320 (N_14320,N_13681,N_13980);
and U14321 (N_14321,N_13969,N_13939);
nand U14322 (N_14322,N_13671,N_13623);
nor U14323 (N_14323,N_13889,N_13818);
or U14324 (N_14324,N_13983,N_13666);
xor U14325 (N_14325,N_13824,N_13818);
nor U14326 (N_14326,N_13942,N_13655);
nand U14327 (N_14327,N_13906,N_13640);
and U14328 (N_14328,N_13526,N_13730);
nand U14329 (N_14329,N_13766,N_13780);
and U14330 (N_14330,N_13881,N_13791);
xnor U14331 (N_14331,N_13559,N_13524);
nand U14332 (N_14332,N_13626,N_13773);
and U14333 (N_14333,N_13629,N_13808);
nor U14334 (N_14334,N_13691,N_13606);
nor U14335 (N_14335,N_13748,N_13961);
and U14336 (N_14336,N_13967,N_13786);
or U14337 (N_14337,N_13553,N_13871);
and U14338 (N_14338,N_13513,N_13781);
nand U14339 (N_14339,N_13819,N_13806);
and U14340 (N_14340,N_13606,N_13790);
nand U14341 (N_14341,N_13975,N_13742);
or U14342 (N_14342,N_13744,N_13730);
and U14343 (N_14343,N_13509,N_13741);
or U14344 (N_14344,N_13883,N_13794);
nand U14345 (N_14345,N_13504,N_13996);
and U14346 (N_14346,N_13839,N_13738);
or U14347 (N_14347,N_13965,N_13723);
nand U14348 (N_14348,N_13661,N_13926);
or U14349 (N_14349,N_13849,N_13622);
nor U14350 (N_14350,N_13517,N_13804);
nor U14351 (N_14351,N_13535,N_13863);
nor U14352 (N_14352,N_13810,N_13858);
xor U14353 (N_14353,N_13695,N_13768);
or U14354 (N_14354,N_13768,N_13598);
or U14355 (N_14355,N_13776,N_13607);
nor U14356 (N_14356,N_13789,N_13617);
xnor U14357 (N_14357,N_13795,N_13862);
and U14358 (N_14358,N_13540,N_13515);
xnor U14359 (N_14359,N_13640,N_13704);
xor U14360 (N_14360,N_13604,N_13575);
nand U14361 (N_14361,N_13860,N_13573);
nand U14362 (N_14362,N_13914,N_13541);
nand U14363 (N_14363,N_13863,N_13752);
and U14364 (N_14364,N_13661,N_13590);
xnor U14365 (N_14365,N_13989,N_13555);
or U14366 (N_14366,N_13653,N_13611);
xor U14367 (N_14367,N_13745,N_13775);
and U14368 (N_14368,N_13805,N_13672);
or U14369 (N_14369,N_13945,N_13814);
nand U14370 (N_14370,N_13717,N_13899);
and U14371 (N_14371,N_13691,N_13707);
or U14372 (N_14372,N_13890,N_13620);
nand U14373 (N_14373,N_13757,N_13586);
nor U14374 (N_14374,N_13740,N_13861);
nor U14375 (N_14375,N_13979,N_13699);
and U14376 (N_14376,N_13909,N_13813);
or U14377 (N_14377,N_13658,N_13594);
xor U14378 (N_14378,N_13751,N_13582);
or U14379 (N_14379,N_13955,N_13614);
and U14380 (N_14380,N_13648,N_13639);
or U14381 (N_14381,N_13526,N_13712);
or U14382 (N_14382,N_13822,N_13753);
xnor U14383 (N_14383,N_13702,N_13687);
nor U14384 (N_14384,N_13874,N_13566);
or U14385 (N_14385,N_13641,N_13605);
and U14386 (N_14386,N_13820,N_13537);
nand U14387 (N_14387,N_13789,N_13566);
xnor U14388 (N_14388,N_13746,N_13781);
nand U14389 (N_14389,N_13823,N_13776);
and U14390 (N_14390,N_13943,N_13881);
or U14391 (N_14391,N_13690,N_13810);
nand U14392 (N_14392,N_13876,N_13556);
xnor U14393 (N_14393,N_13531,N_13913);
or U14394 (N_14394,N_13915,N_13652);
nor U14395 (N_14395,N_13830,N_13605);
or U14396 (N_14396,N_13732,N_13728);
xor U14397 (N_14397,N_13657,N_13788);
xnor U14398 (N_14398,N_13868,N_13669);
and U14399 (N_14399,N_13996,N_13742);
nor U14400 (N_14400,N_13532,N_13835);
xor U14401 (N_14401,N_13788,N_13945);
xnor U14402 (N_14402,N_13808,N_13880);
xnor U14403 (N_14403,N_13644,N_13916);
or U14404 (N_14404,N_13684,N_13690);
xor U14405 (N_14405,N_13721,N_13740);
or U14406 (N_14406,N_13929,N_13914);
nor U14407 (N_14407,N_13871,N_13998);
nor U14408 (N_14408,N_13515,N_13781);
nand U14409 (N_14409,N_13808,N_13664);
nor U14410 (N_14410,N_13838,N_13768);
or U14411 (N_14411,N_13950,N_13748);
nand U14412 (N_14412,N_13557,N_13865);
or U14413 (N_14413,N_13519,N_13664);
or U14414 (N_14414,N_13602,N_13609);
nor U14415 (N_14415,N_13873,N_13631);
nor U14416 (N_14416,N_13634,N_13851);
nor U14417 (N_14417,N_13604,N_13985);
nor U14418 (N_14418,N_13622,N_13736);
xnor U14419 (N_14419,N_13756,N_13670);
or U14420 (N_14420,N_13949,N_13639);
or U14421 (N_14421,N_13655,N_13951);
xor U14422 (N_14422,N_13864,N_13996);
and U14423 (N_14423,N_13594,N_13543);
or U14424 (N_14424,N_13507,N_13910);
xor U14425 (N_14425,N_13807,N_13621);
and U14426 (N_14426,N_13808,N_13697);
and U14427 (N_14427,N_13736,N_13625);
or U14428 (N_14428,N_13990,N_13656);
xnor U14429 (N_14429,N_13609,N_13630);
or U14430 (N_14430,N_13966,N_13535);
or U14431 (N_14431,N_13853,N_13891);
nor U14432 (N_14432,N_13570,N_13577);
nor U14433 (N_14433,N_13887,N_13847);
nor U14434 (N_14434,N_13809,N_13614);
nor U14435 (N_14435,N_13709,N_13662);
or U14436 (N_14436,N_13913,N_13866);
nand U14437 (N_14437,N_13758,N_13685);
or U14438 (N_14438,N_13856,N_13764);
xor U14439 (N_14439,N_13569,N_13515);
and U14440 (N_14440,N_13670,N_13570);
nand U14441 (N_14441,N_13757,N_13827);
or U14442 (N_14442,N_13712,N_13686);
or U14443 (N_14443,N_13814,N_13535);
nor U14444 (N_14444,N_13847,N_13918);
and U14445 (N_14445,N_13780,N_13998);
nand U14446 (N_14446,N_13816,N_13940);
or U14447 (N_14447,N_13778,N_13661);
nor U14448 (N_14448,N_13743,N_13894);
xnor U14449 (N_14449,N_13713,N_13778);
xnor U14450 (N_14450,N_13923,N_13547);
xnor U14451 (N_14451,N_13509,N_13903);
nand U14452 (N_14452,N_13896,N_13691);
xnor U14453 (N_14453,N_13762,N_13865);
xnor U14454 (N_14454,N_13776,N_13517);
xor U14455 (N_14455,N_13527,N_13906);
nor U14456 (N_14456,N_13578,N_13915);
nand U14457 (N_14457,N_13680,N_13669);
and U14458 (N_14458,N_13580,N_13870);
and U14459 (N_14459,N_13790,N_13788);
nand U14460 (N_14460,N_13765,N_13899);
or U14461 (N_14461,N_13512,N_13911);
xnor U14462 (N_14462,N_13920,N_13766);
nand U14463 (N_14463,N_13539,N_13986);
nor U14464 (N_14464,N_13676,N_13703);
or U14465 (N_14465,N_13620,N_13907);
or U14466 (N_14466,N_13773,N_13912);
nor U14467 (N_14467,N_13673,N_13785);
nand U14468 (N_14468,N_13521,N_13525);
and U14469 (N_14469,N_13718,N_13606);
and U14470 (N_14470,N_13726,N_13624);
or U14471 (N_14471,N_13808,N_13626);
or U14472 (N_14472,N_13973,N_13607);
or U14473 (N_14473,N_13756,N_13982);
xnor U14474 (N_14474,N_13758,N_13951);
nand U14475 (N_14475,N_13599,N_13769);
nand U14476 (N_14476,N_13991,N_13717);
nand U14477 (N_14477,N_13615,N_13827);
nand U14478 (N_14478,N_13923,N_13994);
or U14479 (N_14479,N_13688,N_13700);
nand U14480 (N_14480,N_13623,N_13959);
and U14481 (N_14481,N_13682,N_13506);
nor U14482 (N_14482,N_13695,N_13574);
or U14483 (N_14483,N_13574,N_13697);
and U14484 (N_14484,N_13753,N_13858);
nand U14485 (N_14485,N_13718,N_13535);
nor U14486 (N_14486,N_13611,N_13809);
nand U14487 (N_14487,N_13771,N_13858);
or U14488 (N_14488,N_13520,N_13818);
nand U14489 (N_14489,N_13795,N_13896);
or U14490 (N_14490,N_13666,N_13695);
nand U14491 (N_14491,N_13636,N_13625);
or U14492 (N_14492,N_13668,N_13875);
nor U14493 (N_14493,N_13991,N_13515);
or U14494 (N_14494,N_13934,N_13781);
or U14495 (N_14495,N_13590,N_13630);
xnor U14496 (N_14496,N_13939,N_13611);
or U14497 (N_14497,N_13581,N_13718);
and U14498 (N_14498,N_13634,N_13947);
xnor U14499 (N_14499,N_13615,N_13897);
and U14500 (N_14500,N_14079,N_14345);
or U14501 (N_14501,N_14357,N_14091);
xor U14502 (N_14502,N_14065,N_14273);
xor U14503 (N_14503,N_14329,N_14041);
or U14504 (N_14504,N_14184,N_14212);
or U14505 (N_14505,N_14386,N_14439);
and U14506 (N_14506,N_14189,N_14276);
nand U14507 (N_14507,N_14385,N_14005);
and U14508 (N_14508,N_14169,N_14370);
nand U14509 (N_14509,N_14034,N_14121);
nand U14510 (N_14510,N_14375,N_14368);
or U14511 (N_14511,N_14373,N_14445);
or U14512 (N_14512,N_14266,N_14479);
or U14513 (N_14513,N_14304,N_14076);
xor U14514 (N_14514,N_14424,N_14402);
nor U14515 (N_14515,N_14269,N_14149);
nand U14516 (N_14516,N_14097,N_14294);
nand U14517 (N_14517,N_14448,N_14259);
nor U14518 (N_14518,N_14205,N_14408);
xor U14519 (N_14519,N_14497,N_14422);
and U14520 (N_14520,N_14431,N_14392);
and U14521 (N_14521,N_14100,N_14252);
or U14522 (N_14522,N_14157,N_14261);
nor U14523 (N_14523,N_14440,N_14143);
nand U14524 (N_14524,N_14124,N_14101);
xnor U14525 (N_14525,N_14173,N_14028);
nor U14526 (N_14526,N_14344,N_14475);
or U14527 (N_14527,N_14008,N_14183);
and U14528 (N_14528,N_14415,N_14038);
and U14529 (N_14529,N_14468,N_14281);
nand U14530 (N_14530,N_14372,N_14116);
xor U14531 (N_14531,N_14350,N_14308);
or U14532 (N_14532,N_14061,N_14299);
or U14533 (N_14533,N_14068,N_14496);
nand U14534 (N_14534,N_14327,N_14443);
xor U14535 (N_14535,N_14428,N_14177);
nand U14536 (N_14536,N_14401,N_14070);
nand U14537 (N_14537,N_14360,N_14221);
and U14538 (N_14538,N_14409,N_14336);
nand U14539 (N_14539,N_14247,N_14449);
nor U14540 (N_14540,N_14255,N_14384);
and U14541 (N_14541,N_14403,N_14090);
or U14542 (N_14542,N_14251,N_14238);
xor U14543 (N_14543,N_14035,N_14233);
nor U14544 (N_14544,N_14249,N_14208);
or U14545 (N_14545,N_14355,N_14139);
nor U14546 (N_14546,N_14193,N_14310);
xnor U14547 (N_14547,N_14311,N_14120);
and U14548 (N_14548,N_14314,N_14258);
nor U14549 (N_14549,N_14426,N_14285);
and U14550 (N_14550,N_14330,N_14434);
nand U14551 (N_14551,N_14067,N_14146);
or U14552 (N_14552,N_14486,N_14024);
nor U14553 (N_14553,N_14234,N_14026);
xnor U14554 (N_14554,N_14471,N_14107);
xor U14555 (N_14555,N_14007,N_14018);
nor U14556 (N_14556,N_14337,N_14248);
nor U14557 (N_14557,N_14203,N_14232);
xor U14558 (N_14558,N_14181,N_14225);
nand U14559 (N_14559,N_14331,N_14270);
or U14560 (N_14560,N_14192,N_14213);
xnor U14561 (N_14561,N_14338,N_14323);
nand U14562 (N_14562,N_14462,N_14396);
or U14563 (N_14563,N_14222,N_14312);
xnor U14564 (N_14564,N_14334,N_14482);
or U14565 (N_14565,N_14194,N_14489);
xnor U14566 (N_14566,N_14123,N_14084);
nand U14567 (N_14567,N_14349,N_14347);
or U14568 (N_14568,N_14226,N_14006);
or U14569 (N_14569,N_14122,N_14031);
or U14570 (N_14570,N_14379,N_14180);
or U14571 (N_14571,N_14195,N_14071);
xor U14572 (N_14572,N_14039,N_14051);
nor U14573 (N_14573,N_14140,N_14464);
and U14574 (N_14574,N_14303,N_14019);
nand U14575 (N_14575,N_14348,N_14346);
nor U14576 (N_14576,N_14211,N_14240);
nor U14577 (N_14577,N_14050,N_14250);
xnor U14578 (N_14578,N_14014,N_14075);
nand U14579 (N_14579,N_14296,N_14418);
nor U14580 (N_14580,N_14369,N_14376);
nand U14581 (N_14581,N_14004,N_14412);
nor U14582 (N_14582,N_14490,N_14458);
or U14583 (N_14583,N_14371,N_14118);
or U14584 (N_14584,N_14467,N_14282);
xor U14585 (N_14585,N_14245,N_14231);
nand U14586 (N_14586,N_14047,N_14069);
and U14587 (N_14587,N_14275,N_14129);
nand U14588 (N_14588,N_14013,N_14460);
or U14589 (N_14589,N_14318,N_14280);
or U14590 (N_14590,N_14397,N_14387);
or U14591 (N_14591,N_14277,N_14199);
xnor U14592 (N_14592,N_14104,N_14215);
nor U14593 (N_14593,N_14112,N_14382);
nor U14594 (N_14594,N_14147,N_14400);
and U14595 (N_14595,N_14046,N_14263);
and U14596 (N_14596,N_14291,N_14105);
xor U14597 (N_14597,N_14364,N_14484);
or U14598 (N_14598,N_14244,N_14103);
or U14599 (N_14599,N_14354,N_14113);
xnor U14600 (N_14600,N_14176,N_14117);
or U14601 (N_14601,N_14414,N_14151);
and U14602 (N_14602,N_14362,N_14480);
or U14603 (N_14603,N_14134,N_14466);
and U14604 (N_14604,N_14214,N_14292);
and U14605 (N_14605,N_14253,N_14265);
or U14606 (N_14606,N_14229,N_14416);
and U14607 (N_14607,N_14298,N_14186);
xnor U14608 (N_14608,N_14207,N_14301);
nand U14609 (N_14609,N_14174,N_14145);
nor U14610 (N_14610,N_14469,N_14052);
or U14611 (N_14611,N_14324,N_14491);
or U14612 (N_14612,N_14492,N_14011);
nand U14613 (N_14613,N_14352,N_14405);
nand U14614 (N_14614,N_14335,N_14436);
and U14615 (N_14615,N_14109,N_14210);
nor U14616 (N_14616,N_14135,N_14411);
xor U14617 (N_14617,N_14343,N_14435);
nand U14618 (N_14618,N_14056,N_14243);
or U14619 (N_14619,N_14054,N_14461);
and U14620 (N_14620,N_14452,N_14172);
xor U14621 (N_14621,N_14137,N_14419);
xor U14622 (N_14622,N_14246,N_14165);
nor U14623 (N_14623,N_14074,N_14099);
nand U14624 (N_14624,N_14081,N_14022);
xnor U14625 (N_14625,N_14154,N_14020);
nor U14626 (N_14626,N_14111,N_14055);
nor U14627 (N_14627,N_14478,N_14179);
xor U14628 (N_14628,N_14239,N_14260);
nor U14629 (N_14629,N_14297,N_14170);
xnor U14630 (N_14630,N_14150,N_14086);
or U14631 (N_14631,N_14293,N_14367);
and U14632 (N_14632,N_14358,N_14340);
nand U14633 (N_14633,N_14009,N_14159);
nor U14634 (N_14634,N_14487,N_14224);
or U14635 (N_14635,N_14279,N_14141);
nor U14636 (N_14636,N_14380,N_14420);
xor U14637 (N_14637,N_14217,N_14156);
or U14638 (N_14638,N_14305,N_14102);
nor U14639 (N_14639,N_14309,N_14027);
or U14640 (N_14640,N_14295,N_14393);
xnor U14641 (N_14641,N_14437,N_14288);
nor U14642 (N_14642,N_14030,N_14197);
or U14643 (N_14643,N_14465,N_14187);
and U14644 (N_14644,N_14073,N_14433);
and U14645 (N_14645,N_14237,N_14062);
and U14646 (N_14646,N_14040,N_14058);
nor U14647 (N_14647,N_14206,N_14404);
and U14648 (N_14648,N_14398,N_14453);
nor U14649 (N_14649,N_14495,N_14201);
and U14650 (N_14650,N_14220,N_14307);
or U14651 (N_14651,N_14322,N_14254);
nor U14652 (N_14652,N_14289,N_14493);
xnor U14653 (N_14653,N_14060,N_14332);
or U14654 (N_14654,N_14430,N_14447);
and U14655 (N_14655,N_14094,N_14096);
nor U14656 (N_14656,N_14032,N_14417);
xnor U14657 (N_14657,N_14044,N_14078);
nand U14658 (N_14658,N_14407,N_14363);
or U14659 (N_14659,N_14029,N_14053);
and U14660 (N_14660,N_14286,N_14164);
nor U14661 (N_14661,N_14168,N_14499);
nor U14662 (N_14662,N_14390,N_14163);
xor U14663 (N_14663,N_14048,N_14389);
nand U14664 (N_14664,N_14115,N_14283);
and U14665 (N_14665,N_14142,N_14425);
or U14666 (N_14666,N_14125,N_14128);
or U14667 (N_14667,N_14450,N_14321);
and U14668 (N_14668,N_14162,N_14167);
and U14669 (N_14669,N_14442,N_14356);
and U14670 (N_14670,N_14325,N_14138);
xor U14671 (N_14671,N_14016,N_14476);
nand U14672 (N_14672,N_14175,N_14278);
or U14673 (N_14673,N_14021,N_14095);
and U14674 (N_14674,N_14316,N_14036);
nor U14675 (N_14675,N_14042,N_14130);
nor U14676 (N_14676,N_14342,N_14003);
or U14677 (N_14677,N_14341,N_14395);
and U14678 (N_14678,N_14178,N_14066);
and U14679 (N_14679,N_14488,N_14015);
nor U14680 (N_14680,N_14223,N_14427);
nor U14681 (N_14681,N_14001,N_14087);
or U14682 (N_14682,N_14083,N_14339);
nand U14683 (N_14683,N_14080,N_14191);
or U14684 (N_14684,N_14454,N_14085);
nor U14685 (N_14685,N_14271,N_14377);
nor U14686 (N_14686,N_14494,N_14235);
nor U14687 (N_14687,N_14064,N_14136);
and U14688 (N_14688,N_14126,N_14119);
and U14689 (N_14689,N_14381,N_14002);
nand U14690 (N_14690,N_14012,N_14483);
xnor U14691 (N_14691,N_14158,N_14353);
nand U14692 (N_14692,N_14365,N_14256);
nor U14693 (N_14693,N_14399,N_14209);
xnor U14694 (N_14694,N_14394,N_14262);
nand U14695 (N_14695,N_14045,N_14098);
and U14696 (N_14696,N_14110,N_14171);
and U14697 (N_14697,N_14463,N_14182);
nand U14698 (N_14698,N_14459,N_14216);
xor U14699 (N_14699,N_14300,N_14063);
nor U14700 (N_14700,N_14093,N_14188);
nor U14701 (N_14701,N_14236,N_14328);
or U14702 (N_14702,N_14023,N_14284);
nand U14703 (N_14703,N_14410,N_14132);
nor U14704 (N_14704,N_14290,N_14114);
or U14705 (N_14705,N_14272,N_14152);
and U14706 (N_14706,N_14092,N_14444);
nor U14707 (N_14707,N_14366,N_14025);
nor U14708 (N_14708,N_14326,N_14196);
nand U14709 (N_14709,N_14049,N_14148);
and U14710 (N_14710,N_14333,N_14474);
and U14711 (N_14711,N_14155,N_14082);
or U14712 (N_14712,N_14413,N_14185);
or U14713 (N_14713,N_14160,N_14219);
xor U14714 (N_14714,N_14077,N_14153);
and U14715 (N_14715,N_14438,N_14313);
xor U14716 (N_14716,N_14485,N_14059);
xor U14717 (N_14717,N_14268,N_14472);
xnor U14718 (N_14718,N_14274,N_14383);
xnor U14719 (N_14719,N_14161,N_14423);
or U14720 (N_14720,N_14287,N_14455);
and U14721 (N_14721,N_14432,N_14361);
nand U14722 (N_14722,N_14198,N_14230);
xnor U14723 (N_14723,N_14317,N_14106);
and U14724 (N_14724,N_14320,N_14391);
and U14725 (N_14725,N_14374,N_14441);
xnor U14726 (N_14726,N_14010,N_14200);
xnor U14727 (N_14727,N_14241,N_14264);
nor U14728 (N_14728,N_14481,N_14088);
or U14729 (N_14729,N_14457,N_14218);
or U14730 (N_14730,N_14227,N_14406);
or U14731 (N_14731,N_14033,N_14477);
and U14732 (N_14732,N_14127,N_14319);
and U14733 (N_14733,N_14267,N_14302);
and U14734 (N_14734,N_14421,N_14228);
xor U14735 (N_14735,N_14131,N_14257);
or U14736 (N_14736,N_14470,N_14359);
xnor U14737 (N_14737,N_14315,N_14473);
nor U14738 (N_14738,N_14089,N_14429);
or U14739 (N_14739,N_14351,N_14242);
xor U14740 (N_14740,N_14451,N_14388);
nor U14741 (N_14741,N_14072,N_14108);
or U14742 (N_14742,N_14202,N_14306);
or U14743 (N_14743,N_14498,N_14017);
nor U14744 (N_14744,N_14378,N_14190);
and U14745 (N_14745,N_14456,N_14000);
and U14746 (N_14746,N_14144,N_14204);
and U14747 (N_14747,N_14037,N_14057);
nor U14748 (N_14748,N_14446,N_14043);
nand U14749 (N_14749,N_14166,N_14133);
and U14750 (N_14750,N_14069,N_14018);
nand U14751 (N_14751,N_14491,N_14252);
or U14752 (N_14752,N_14362,N_14292);
or U14753 (N_14753,N_14331,N_14282);
nand U14754 (N_14754,N_14381,N_14213);
and U14755 (N_14755,N_14107,N_14371);
xnor U14756 (N_14756,N_14120,N_14177);
nor U14757 (N_14757,N_14234,N_14314);
and U14758 (N_14758,N_14412,N_14126);
nor U14759 (N_14759,N_14350,N_14341);
or U14760 (N_14760,N_14060,N_14443);
and U14761 (N_14761,N_14329,N_14240);
nor U14762 (N_14762,N_14388,N_14239);
or U14763 (N_14763,N_14015,N_14033);
xor U14764 (N_14764,N_14425,N_14024);
nor U14765 (N_14765,N_14115,N_14434);
or U14766 (N_14766,N_14033,N_14014);
nor U14767 (N_14767,N_14296,N_14398);
and U14768 (N_14768,N_14108,N_14149);
and U14769 (N_14769,N_14293,N_14227);
nor U14770 (N_14770,N_14215,N_14416);
xor U14771 (N_14771,N_14012,N_14352);
nand U14772 (N_14772,N_14226,N_14263);
and U14773 (N_14773,N_14324,N_14287);
xor U14774 (N_14774,N_14048,N_14234);
nor U14775 (N_14775,N_14486,N_14028);
and U14776 (N_14776,N_14260,N_14499);
nand U14777 (N_14777,N_14385,N_14376);
nor U14778 (N_14778,N_14384,N_14358);
or U14779 (N_14779,N_14313,N_14101);
or U14780 (N_14780,N_14030,N_14329);
or U14781 (N_14781,N_14450,N_14460);
nor U14782 (N_14782,N_14471,N_14159);
and U14783 (N_14783,N_14083,N_14480);
or U14784 (N_14784,N_14278,N_14242);
or U14785 (N_14785,N_14469,N_14263);
or U14786 (N_14786,N_14229,N_14110);
and U14787 (N_14787,N_14119,N_14090);
xnor U14788 (N_14788,N_14075,N_14095);
nor U14789 (N_14789,N_14110,N_14054);
xor U14790 (N_14790,N_14150,N_14055);
and U14791 (N_14791,N_14215,N_14227);
nand U14792 (N_14792,N_14072,N_14384);
nand U14793 (N_14793,N_14097,N_14241);
and U14794 (N_14794,N_14094,N_14078);
or U14795 (N_14795,N_14347,N_14397);
xor U14796 (N_14796,N_14301,N_14032);
or U14797 (N_14797,N_14431,N_14095);
nor U14798 (N_14798,N_14157,N_14326);
nor U14799 (N_14799,N_14467,N_14026);
or U14800 (N_14800,N_14069,N_14089);
nand U14801 (N_14801,N_14217,N_14189);
nand U14802 (N_14802,N_14167,N_14338);
and U14803 (N_14803,N_14052,N_14032);
or U14804 (N_14804,N_14397,N_14301);
xor U14805 (N_14805,N_14201,N_14086);
xor U14806 (N_14806,N_14042,N_14251);
xor U14807 (N_14807,N_14063,N_14485);
xnor U14808 (N_14808,N_14195,N_14048);
and U14809 (N_14809,N_14400,N_14431);
xor U14810 (N_14810,N_14361,N_14393);
nor U14811 (N_14811,N_14171,N_14166);
and U14812 (N_14812,N_14445,N_14282);
nand U14813 (N_14813,N_14366,N_14428);
xor U14814 (N_14814,N_14383,N_14060);
nand U14815 (N_14815,N_14314,N_14385);
xor U14816 (N_14816,N_14034,N_14215);
and U14817 (N_14817,N_14254,N_14412);
nand U14818 (N_14818,N_14175,N_14363);
nor U14819 (N_14819,N_14176,N_14087);
xor U14820 (N_14820,N_14313,N_14331);
or U14821 (N_14821,N_14215,N_14263);
or U14822 (N_14822,N_14291,N_14186);
and U14823 (N_14823,N_14199,N_14036);
nor U14824 (N_14824,N_14436,N_14367);
or U14825 (N_14825,N_14398,N_14215);
xor U14826 (N_14826,N_14372,N_14461);
nor U14827 (N_14827,N_14456,N_14088);
or U14828 (N_14828,N_14022,N_14489);
and U14829 (N_14829,N_14022,N_14030);
and U14830 (N_14830,N_14359,N_14032);
nor U14831 (N_14831,N_14332,N_14035);
nor U14832 (N_14832,N_14402,N_14151);
and U14833 (N_14833,N_14478,N_14390);
nor U14834 (N_14834,N_14289,N_14229);
or U14835 (N_14835,N_14214,N_14188);
or U14836 (N_14836,N_14266,N_14079);
nor U14837 (N_14837,N_14082,N_14012);
nand U14838 (N_14838,N_14279,N_14448);
nand U14839 (N_14839,N_14053,N_14185);
xor U14840 (N_14840,N_14163,N_14067);
nand U14841 (N_14841,N_14210,N_14040);
and U14842 (N_14842,N_14015,N_14394);
nand U14843 (N_14843,N_14384,N_14264);
xor U14844 (N_14844,N_14394,N_14364);
and U14845 (N_14845,N_14247,N_14237);
or U14846 (N_14846,N_14362,N_14185);
nor U14847 (N_14847,N_14495,N_14052);
or U14848 (N_14848,N_14112,N_14087);
nor U14849 (N_14849,N_14125,N_14272);
nand U14850 (N_14850,N_14123,N_14343);
nor U14851 (N_14851,N_14263,N_14284);
nand U14852 (N_14852,N_14463,N_14303);
nand U14853 (N_14853,N_14247,N_14332);
nand U14854 (N_14854,N_14485,N_14453);
nand U14855 (N_14855,N_14444,N_14183);
xnor U14856 (N_14856,N_14019,N_14120);
xnor U14857 (N_14857,N_14243,N_14393);
nand U14858 (N_14858,N_14138,N_14071);
or U14859 (N_14859,N_14061,N_14020);
xor U14860 (N_14860,N_14280,N_14121);
nor U14861 (N_14861,N_14402,N_14265);
nand U14862 (N_14862,N_14325,N_14248);
nand U14863 (N_14863,N_14025,N_14172);
xnor U14864 (N_14864,N_14348,N_14224);
xor U14865 (N_14865,N_14302,N_14301);
and U14866 (N_14866,N_14408,N_14469);
nand U14867 (N_14867,N_14431,N_14417);
or U14868 (N_14868,N_14079,N_14263);
nand U14869 (N_14869,N_14093,N_14340);
nor U14870 (N_14870,N_14211,N_14356);
xor U14871 (N_14871,N_14174,N_14451);
or U14872 (N_14872,N_14076,N_14443);
and U14873 (N_14873,N_14232,N_14451);
or U14874 (N_14874,N_14041,N_14160);
nand U14875 (N_14875,N_14488,N_14443);
or U14876 (N_14876,N_14373,N_14186);
or U14877 (N_14877,N_14160,N_14088);
nor U14878 (N_14878,N_14316,N_14371);
nand U14879 (N_14879,N_14295,N_14150);
xor U14880 (N_14880,N_14218,N_14319);
and U14881 (N_14881,N_14264,N_14125);
and U14882 (N_14882,N_14182,N_14111);
nand U14883 (N_14883,N_14471,N_14280);
or U14884 (N_14884,N_14403,N_14389);
nor U14885 (N_14885,N_14074,N_14220);
nand U14886 (N_14886,N_14473,N_14312);
xnor U14887 (N_14887,N_14180,N_14012);
and U14888 (N_14888,N_14017,N_14274);
xor U14889 (N_14889,N_14082,N_14329);
or U14890 (N_14890,N_14431,N_14068);
xnor U14891 (N_14891,N_14361,N_14312);
and U14892 (N_14892,N_14258,N_14174);
nand U14893 (N_14893,N_14145,N_14052);
and U14894 (N_14894,N_14452,N_14336);
and U14895 (N_14895,N_14356,N_14129);
nand U14896 (N_14896,N_14187,N_14395);
xor U14897 (N_14897,N_14261,N_14322);
nor U14898 (N_14898,N_14014,N_14202);
nand U14899 (N_14899,N_14089,N_14078);
nor U14900 (N_14900,N_14403,N_14313);
and U14901 (N_14901,N_14346,N_14184);
nand U14902 (N_14902,N_14384,N_14348);
nor U14903 (N_14903,N_14139,N_14352);
and U14904 (N_14904,N_14428,N_14400);
and U14905 (N_14905,N_14440,N_14199);
and U14906 (N_14906,N_14049,N_14344);
and U14907 (N_14907,N_14118,N_14250);
xor U14908 (N_14908,N_14141,N_14271);
nor U14909 (N_14909,N_14480,N_14004);
xnor U14910 (N_14910,N_14346,N_14391);
and U14911 (N_14911,N_14446,N_14112);
nor U14912 (N_14912,N_14400,N_14090);
nor U14913 (N_14913,N_14276,N_14351);
or U14914 (N_14914,N_14269,N_14448);
or U14915 (N_14915,N_14000,N_14200);
or U14916 (N_14916,N_14144,N_14003);
and U14917 (N_14917,N_14484,N_14226);
or U14918 (N_14918,N_14354,N_14044);
xor U14919 (N_14919,N_14136,N_14340);
or U14920 (N_14920,N_14029,N_14412);
and U14921 (N_14921,N_14116,N_14213);
and U14922 (N_14922,N_14491,N_14301);
xnor U14923 (N_14923,N_14360,N_14331);
nor U14924 (N_14924,N_14217,N_14059);
nand U14925 (N_14925,N_14024,N_14357);
nor U14926 (N_14926,N_14412,N_14231);
nor U14927 (N_14927,N_14409,N_14234);
xor U14928 (N_14928,N_14196,N_14261);
xor U14929 (N_14929,N_14302,N_14177);
xor U14930 (N_14930,N_14458,N_14351);
or U14931 (N_14931,N_14325,N_14408);
or U14932 (N_14932,N_14411,N_14086);
xnor U14933 (N_14933,N_14441,N_14467);
nor U14934 (N_14934,N_14130,N_14107);
or U14935 (N_14935,N_14209,N_14032);
nand U14936 (N_14936,N_14027,N_14433);
and U14937 (N_14937,N_14434,N_14273);
nand U14938 (N_14938,N_14455,N_14251);
nand U14939 (N_14939,N_14182,N_14246);
and U14940 (N_14940,N_14208,N_14079);
xor U14941 (N_14941,N_14443,N_14314);
xor U14942 (N_14942,N_14188,N_14025);
xor U14943 (N_14943,N_14154,N_14109);
or U14944 (N_14944,N_14495,N_14221);
nor U14945 (N_14945,N_14065,N_14449);
nand U14946 (N_14946,N_14102,N_14382);
and U14947 (N_14947,N_14354,N_14170);
or U14948 (N_14948,N_14175,N_14344);
nand U14949 (N_14949,N_14032,N_14358);
and U14950 (N_14950,N_14300,N_14466);
nor U14951 (N_14951,N_14338,N_14109);
and U14952 (N_14952,N_14210,N_14276);
xor U14953 (N_14953,N_14471,N_14000);
or U14954 (N_14954,N_14288,N_14249);
or U14955 (N_14955,N_14140,N_14331);
xnor U14956 (N_14956,N_14475,N_14339);
xor U14957 (N_14957,N_14153,N_14230);
or U14958 (N_14958,N_14132,N_14113);
and U14959 (N_14959,N_14057,N_14424);
or U14960 (N_14960,N_14002,N_14444);
nor U14961 (N_14961,N_14174,N_14161);
nand U14962 (N_14962,N_14023,N_14153);
nand U14963 (N_14963,N_14445,N_14355);
nor U14964 (N_14964,N_14392,N_14436);
xnor U14965 (N_14965,N_14235,N_14253);
nor U14966 (N_14966,N_14313,N_14489);
xnor U14967 (N_14967,N_14189,N_14431);
or U14968 (N_14968,N_14153,N_14253);
nand U14969 (N_14969,N_14195,N_14279);
xor U14970 (N_14970,N_14221,N_14303);
nand U14971 (N_14971,N_14425,N_14058);
or U14972 (N_14972,N_14330,N_14294);
xnor U14973 (N_14973,N_14104,N_14266);
and U14974 (N_14974,N_14094,N_14114);
or U14975 (N_14975,N_14181,N_14404);
and U14976 (N_14976,N_14161,N_14487);
or U14977 (N_14977,N_14275,N_14037);
nand U14978 (N_14978,N_14430,N_14100);
and U14979 (N_14979,N_14460,N_14092);
nand U14980 (N_14980,N_14412,N_14272);
and U14981 (N_14981,N_14166,N_14296);
xnor U14982 (N_14982,N_14315,N_14110);
and U14983 (N_14983,N_14233,N_14316);
or U14984 (N_14984,N_14121,N_14064);
or U14985 (N_14985,N_14020,N_14419);
nor U14986 (N_14986,N_14187,N_14009);
nand U14987 (N_14987,N_14079,N_14284);
nor U14988 (N_14988,N_14097,N_14380);
xnor U14989 (N_14989,N_14180,N_14429);
nand U14990 (N_14990,N_14204,N_14141);
nand U14991 (N_14991,N_14242,N_14133);
or U14992 (N_14992,N_14248,N_14153);
nand U14993 (N_14993,N_14014,N_14424);
and U14994 (N_14994,N_14155,N_14363);
or U14995 (N_14995,N_14048,N_14295);
xor U14996 (N_14996,N_14329,N_14465);
or U14997 (N_14997,N_14489,N_14347);
or U14998 (N_14998,N_14345,N_14191);
xnor U14999 (N_14999,N_14126,N_14118);
xor U15000 (N_15000,N_14552,N_14870);
xor U15001 (N_15001,N_14561,N_14808);
or U15002 (N_15002,N_14921,N_14633);
nor U15003 (N_15003,N_14780,N_14971);
and U15004 (N_15004,N_14629,N_14816);
nand U15005 (N_15005,N_14817,N_14862);
nor U15006 (N_15006,N_14990,N_14518);
nor U15007 (N_15007,N_14650,N_14635);
xnor U15008 (N_15008,N_14915,N_14621);
nand U15009 (N_15009,N_14589,N_14864);
and U15010 (N_15010,N_14595,N_14715);
or U15011 (N_15011,N_14669,N_14770);
xor U15012 (N_15012,N_14695,N_14824);
and U15013 (N_15013,N_14940,N_14722);
nand U15014 (N_15014,N_14582,N_14922);
xor U15015 (N_15015,N_14632,N_14592);
or U15016 (N_15016,N_14784,N_14769);
xor U15017 (N_15017,N_14840,N_14532);
xor U15018 (N_15018,N_14531,N_14679);
or U15019 (N_15019,N_14564,N_14775);
nand U15020 (N_15020,N_14934,N_14622);
nand U15021 (N_15021,N_14642,N_14545);
xnor U15022 (N_15022,N_14952,N_14661);
and U15023 (N_15023,N_14819,N_14603);
nor U15024 (N_15024,N_14999,N_14609);
or U15025 (N_15025,N_14709,N_14513);
or U15026 (N_15026,N_14820,N_14988);
nand U15027 (N_15027,N_14643,N_14904);
and U15028 (N_15028,N_14735,N_14969);
xnor U15029 (N_15029,N_14853,N_14975);
nand U15030 (N_15030,N_14526,N_14730);
and U15031 (N_15031,N_14749,N_14795);
or U15032 (N_15032,N_14884,N_14678);
and U15033 (N_15033,N_14941,N_14638);
and U15034 (N_15034,N_14521,N_14671);
nand U15035 (N_15035,N_14828,N_14747);
nor U15036 (N_15036,N_14551,N_14560);
nor U15037 (N_15037,N_14689,N_14558);
or U15038 (N_15038,N_14666,N_14570);
xor U15039 (N_15039,N_14742,N_14578);
and U15040 (N_15040,N_14524,N_14982);
xnor U15041 (N_15041,N_14811,N_14583);
and U15042 (N_15042,N_14752,N_14852);
and U15043 (N_15043,N_14557,N_14625);
and U15044 (N_15044,N_14882,N_14841);
nand U15045 (N_15045,N_14830,N_14738);
or U15046 (N_15046,N_14670,N_14994);
nand U15047 (N_15047,N_14832,N_14731);
nor U15048 (N_15048,N_14980,N_14979);
nor U15049 (N_15049,N_14891,N_14702);
xnor U15050 (N_15050,N_14781,N_14692);
and U15051 (N_15051,N_14662,N_14674);
and U15052 (N_15052,N_14908,N_14753);
and U15053 (N_15053,N_14759,N_14973);
or U15054 (N_15054,N_14863,N_14829);
nor U15055 (N_15055,N_14879,N_14706);
xor U15056 (N_15056,N_14909,N_14700);
nand U15057 (N_15057,N_14542,N_14726);
or U15058 (N_15058,N_14655,N_14618);
nand U15059 (N_15059,N_14627,N_14528);
nand U15060 (N_15060,N_14651,N_14646);
nand U15061 (N_15061,N_14758,N_14736);
nor U15062 (N_15062,N_14815,N_14810);
nor U15063 (N_15063,N_14794,N_14797);
nand U15064 (N_15064,N_14506,N_14932);
and U15065 (N_15065,N_14918,N_14774);
nand U15066 (N_15066,N_14858,N_14911);
xor U15067 (N_15067,N_14929,N_14639);
or U15068 (N_15068,N_14563,N_14630);
nor U15069 (N_15069,N_14511,N_14572);
or U15070 (N_15070,N_14983,N_14641);
nor U15071 (N_15071,N_14591,N_14588);
xnor U15072 (N_15072,N_14649,N_14772);
xnor U15073 (N_15073,N_14555,N_14871);
and U15074 (N_15074,N_14665,N_14924);
nand U15075 (N_15075,N_14914,N_14765);
and U15076 (N_15076,N_14615,N_14687);
and U15077 (N_15077,N_14574,N_14672);
or U15078 (N_15078,N_14837,N_14806);
and U15079 (N_15079,N_14944,N_14556);
nand U15080 (N_15080,N_14910,N_14834);
and U15081 (N_15081,N_14523,N_14690);
and U15082 (N_15082,N_14698,N_14799);
and U15083 (N_15083,N_14947,N_14903);
and U15084 (N_15084,N_14779,N_14613);
xor U15085 (N_15085,N_14680,N_14843);
nand U15086 (N_15086,N_14798,N_14538);
nor U15087 (N_15087,N_14928,N_14548);
nand U15088 (N_15088,N_14842,N_14939);
or U15089 (N_15089,N_14833,N_14920);
nand U15090 (N_15090,N_14991,N_14516);
xor U15091 (N_15091,N_14529,N_14510);
and U15092 (N_15092,N_14598,N_14734);
and U15093 (N_15093,N_14575,N_14675);
xor U15094 (N_15094,N_14601,N_14916);
or U15095 (N_15095,N_14989,N_14577);
xnor U15096 (N_15096,N_14549,N_14886);
nor U15097 (N_15097,N_14746,N_14992);
nand U15098 (N_15098,N_14697,N_14860);
nor U15099 (N_15099,N_14619,N_14724);
and U15100 (N_15100,N_14898,N_14894);
or U15101 (N_15101,N_14846,N_14663);
and U15102 (N_15102,N_14569,N_14550);
nand U15103 (N_15103,N_14546,N_14567);
nand U15104 (N_15104,N_14984,N_14501);
or U15105 (N_15105,N_14527,N_14782);
xnor U15106 (N_15106,N_14831,N_14517);
xnor U15107 (N_15107,N_14701,N_14590);
nor U15108 (N_15108,N_14660,N_14648);
xnor U15109 (N_15109,N_14606,N_14838);
or U15110 (N_15110,N_14685,N_14554);
xor U15111 (N_15111,N_14525,N_14713);
xnor U15112 (N_15112,N_14901,N_14976);
or U15113 (N_15113,N_14792,N_14540);
and U15114 (N_15114,N_14503,N_14966);
nor U15115 (N_15115,N_14616,N_14508);
or U15116 (N_15116,N_14926,N_14818);
or U15117 (N_15117,N_14751,N_14956);
nand U15118 (N_15118,N_14773,N_14998);
or U15119 (N_15119,N_14803,N_14868);
or U15120 (N_15120,N_14520,N_14541);
and U15121 (N_15121,N_14607,N_14800);
and U15122 (N_15122,N_14981,N_14694);
xnor U15123 (N_15123,N_14801,N_14535);
and U15124 (N_15124,N_14987,N_14938);
xnor U15125 (N_15125,N_14509,N_14696);
xnor U15126 (N_15126,N_14710,N_14919);
xnor U15127 (N_15127,N_14720,N_14767);
nor U15128 (N_15128,N_14530,N_14923);
and U15129 (N_15129,N_14711,N_14614);
and U15130 (N_15130,N_14637,N_14608);
or U15131 (N_15131,N_14899,N_14744);
nor U15132 (N_15132,N_14741,N_14644);
or U15133 (N_15133,N_14883,N_14761);
nand U15134 (N_15134,N_14950,N_14723);
xor U15135 (N_15135,N_14836,N_14628);
nor U15136 (N_15136,N_14626,N_14539);
xor U15137 (N_15137,N_14740,N_14597);
and U15138 (N_15138,N_14851,N_14902);
and U15139 (N_15139,N_14705,N_14768);
or U15140 (N_15140,N_14721,N_14805);
nor U15141 (N_15141,N_14568,N_14640);
xor U15142 (N_15142,N_14714,N_14931);
and U15143 (N_15143,N_14707,N_14855);
and U15144 (N_15144,N_14887,N_14906);
nand U15145 (N_15145,N_14986,N_14913);
and U15146 (N_15146,N_14712,N_14757);
nand U15147 (N_15147,N_14536,N_14907);
nor U15148 (N_15148,N_14996,N_14877);
xor U15149 (N_15149,N_14659,N_14876);
and U15150 (N_15150,N_14872,N_14958);
and U15151 (N_15151,N_14771,N_14847);
nor U15152 (N_15152,N_14576,N_14504);
and U15153 (N_15153,N_14636,N_14543);
nor U15154 (N_15154,N_14878,N_14968);
xor U15155 (N_15155,N_14850,N_14859);
nand U15156 (N_15156,N_14955,N_14587);
and U15157 (N_15157,N_14844,N_14892);
and U15158 (N_15158,N_14813,N_14943);
and U15159 (N_15159,N_14612,N_14776);
nand U15160 (N_15160,N_14566,N_14942);
and U15161 (N_15161,N_14867,N_14949);
or U15162 (N_15162,N_14562,N_14600);
nand U15163 (N_15163,N_14848,N_14573);
nand U15164 (N_15164,N_14533,N_14936);
nand U15165 (N_15165,N_14762,N_14873);
or U15166 (N_15166,N_14764,N_14869);
and U15167 (N_15167,N_14703,N_14977);
nor U15168 (N_15168,N_14547,N_14875);
xnor U15169 (N_15169,N_14748,N_14500);
nand U15170 (N_15170,N_14959,N_14604);
or U15171 (N_15171,N_14676,N_14725);
xnor U15172 (N_15172,N_14645,N_14683);
and U15173 (N_15173,N_14951,N_14664);
nand U15174 (N_15174,N_14945,N_14893);
and U15175 (N_15175,N_14890,N_14974);
or U15176 (N_15176,N_14963,N_14565);
or U15177 (N_15177,N_14845,N_14766);
nor U15178 (N_15178,N_14737,N_14579);
or U15179 (N_15179,N_14656,N_14825);
nor U15180 (N_15180,N_14881,N_14804);
nand U15181 (N_15181,N_14760,N_14927);
or U15182 (N_15182,N_14787,N_14512);
or U15183 (N_15183,N_14681,N_14677);
or U15184 (N_15184,N_14623,N_14967);
xnor U15185 (N_15185,N_14610,N_14791);
xor U15186 (N_15186,N_14571,N_14553);
or U15187 (N_15187,N_14617,N_14937);
xnor U15188 (N_15188,N_14691,N_14502);
and U15189 (N_15189,N_14580,N_14897);
xnor U15190 (N_15190,N_14653,N_14970);
or U15191 (N_15191,N_14611,N_14957);
xor U15192 (N_15192,N_14585,N_14946);
xor U15193 (N_15193,N_14849,N_14515);
nand U15194 (N_15194,N_14605,N_14785);
or U15195 (N_15195,N_14905,N_14874);
or U15196 (N_15196,N_14704,N_14985);
xor U15197 (N_15197,N_14821,N_14935);
and U15198 (N_15198,N_14708,N_14581);
nand U15199 (N_15199,N_14962,N_14954);
nand U15200 (N_15200,N_14812,N_14802);
nor U15201 (N_15201,N_14647,N_14596);
and U15202 (N_15202,N_14634,N_14688);
nor U15203 (N_15203,N_14719,N_14965);
xnor U15204 (N_15204,N_14827,N_14826);
xnor U15205 (N_15205,N_14786,N_14522);
nor U15206 (N_15206,N_14717,N_14796);
nor U15207 (N_15207,N_14885,N_14745);
xor U15208 (N_15208,N_14658,N_14880);
and U15209 (N_15209,N_14861,N_14788);
and U15210 (N_15210,N_14777,N_14732);
and U15211 (N_15211,N_14978,N_14856);
and U15212 (N_15212,N_14514,N_14537);
xnor U15213 (N_15213,N_14896,N_14716);
nand U15214 (N_15214,N_14822,N_14809);
or U15215 (N_15215,N_14684,N_14602);
and U15216 (N_15216,N_14718,N_14727);
nand U15217 (N_15217,N_14763,N_14507);
nand U15218 (N_15218,N_14972,N_14823);
or U15219 (N_15219,N_14925,N_14739);
xor U15220 (N_15220,N_14593,N_14997);
xnor U15221 (N_15221,N_14756,N_14728);
or U15222 (N_15222,N_14750,N_14505);
and U15223 (N_15223,N_14930,N_14857);
xnor U15224 (N_15224,N_14519,N_14599);
and U15225 (N_15225,N_14854,N_14790);
nor U15226 (N_15226,N_14584,N_14654);
xnor U15227 (N_15227,N_14839,N_14835);
nand U15228 (N_15228,N_14807,N_14995);
xor U15229 (N_15229,N_14961,N_14652);
nor U15230 (N_15230,N_14743,N_14865);
xnor U15231 (N_15231,N_14673,N_14699);
or U15232 (N_15232,N_14912,N_14900);
xor U15233 (N_15233,N_14754,N_14783);
or U15234 (N_15234,N_14729,N_14667);
and U15235 (N_15235,N_14686,N_14814);
nor U15236 (N_15236,N_14933,N_14964);
or U15237 (N_15237,N_14917,N_14544);
and U15238 (N_15238,N_14993,N_14755);
or U15239 (N_15239,N_14953,N_14534);
xor U15240 (N_15240,N_14733,N_14620);
or U15241 (N_15241,N_14631,N_14888);
nor U15242 (N_15242,N_14586,N_14624);
or U15243 (N_15243,N_14657,N_14559);
xnor U15244 (N_15244,N_14789,N_14960);
xnor U15245 (N_15245,N_14668,N_14948);
and U15246 (N_15246,N_14778,N_14693);
nor U15247 (N_15247,N_14682,N_14895);
xnor U15248 (N_15248,N_14793,N_14889);
or U15249 (N_15249,N_14594,N_14866);
xnor U15250 (N_15250,N_14598,N_14731);
nor U15251 (N_15251,N_14906,N_14597);
and U15252 (N_15252,N_14818,N_14520);
nor U15253 (N_15253,N_14671,N_14609);
or U15254 (N_15254,N_14998,N_14696);
nor U15255 (N_15255,N_14622,N_14861);
xor U15256 (N_15256,N_14672,N_14547);
or U15257 (N_15257,N_14956,N_14512);
nor U15258 (N_15258,N_14701,N_14504);
xnor U15259 (N_15259,N_14682,N_14645);
nand U15260 (N_15260,N_14846,N_14828);
xnor U15261 (N_15261,N_14556,N_14974);
nand U15262 (N_15262,N_14562,N_14926);
nor U15263 (N_15263,N_14807,N_14588);
or U15264 (N_15264,N_14830,N_14914);
nand U15265 (N_15265,N_14592,N_14528);
nand U15266 (N_15266,N_14586,N_14516);
and U15267 (N_15267,N_14648,N_14632);
xor U15268 (N_15268,N_14800,N_14684);
nor U15269 (N_15269,N_14796,N_14524);
nand U15270 (N_15270,N_14604,N_14700);
and U15271 (N_15271,N_14625,N_14510);
xor U15272 (N_15272,N_14918,N_14715);
or U15273 (N_15273,N_14668,N_14690);
nand U15274 (N_15274,N_14705,N_14760);
and U15275 (N_15275,N_14922,N_14725);
nand U15276 (N_15276,N_14866,N_14880);
nor U15277 (N_15277,N_14592,N_14954);
or U15278 (N_15278,N_14760,N_14969);
nand U15279 (N_15279,N_14543,N_14810);
or U15280 (N_15280,N_14877,N_14995);
nor U15281 (N_15281,N_14771,N_14711);
and U15282 (N_15282,N_14521,N_14937);
and U15283 (N_15283,N_14550,N_14969);
and U15284 (N_15284,N_14638,N_14520);
xnor U15285 (N_15285,N_14790,N_14978);
and U15286 (N_15286,N_14591,N_14688);
nand U15287 (N_15287,N_14664,N_14946);
nor U15288 (N_15288,N_14942,N_14586);
xnor U15289 (N_15289,N_14554,N_14589);
xnor U15290 (N_15290,N_14642,N_14827);
or U15291 (N_15291,N_14823,N_14944);
nor U15292 (N_15292,N_14741,N_14952);
nand U15293 (N_15293,N_14696,N_14957);
nand U15294 (N_15294,N_14962,N_14886);
and U15295 (N_15295,N_14822,N_14777);
and U15296 (N_15296,N_14997,N_14516);
nand U15297 (N_15297,N_14889,N_14799);
and U15298 (N_15298,N_14855,N_14933);
xnor U15299 (N_15299,N_14891,N_14559);
nor U15300 (N_15300,N_14528,N_14536);
nand U15301 (N_15301,N_14737,N_14725);
nand U15302 (N_15302,N_14926,N_14574);
nor U15303 (N_15303,N_14777,N_14983);
and U15304 (N_15304,N_14713,N_14630);
nand U15305 (N_15305,N_14632,N_14988);
xor U15306 (N_15306,N_14596,N_14899);
nor U15307 (N_15307,N_14890,N_14602);
nand U15308 (N_15308,N_14547,N_14553);
or U15309 (N_15309,N_14614,N_14869);
or U15310 (N_15310,N_14694,N_14521);
nor U15311 (N_15311,N_14897,N_14778);
xor U15312 (N_15312,N_14515,N_14727);
nand U15313 (N_15313,N_14913,N_14793);
nor U15314 (N_15314,N_14992,N_14779);
nand U15315 (N_15315,N_14848,N_14541);
xnor U15316 (N_15316,N_14692,N_14646);
or U15317 (N_15317,N_14636,N_14865);
nand U15318 (N_15318,N_14670,N_14818);
nand U15319 (N_15319,N_14659,N_14930);
nor U15320 (N_15320,N_14917,N_14612);
nand U15321 (N_15321,N_14963,N_14952);
or U15322 (N_15322,N_14782,N_14604);
xnor U15323 (N_15323,N_14907,N_14564);
and U15324 (N_15324,N_14875,N_14560);
xor U15325 (N_15325,N_14590,N_14593);
or U15326 (N_15326,N_14556,N_14741);
nand U15327 (N_15327,N_14875,N_14511);
and U15328 (N_15328,N_14783,N_14511);
or U15329 (N_15329,N_14702,N_14719);
xor U15330 (N_15330,N_14998,N_14669);
and U15331 (N_15331,N_14950,N_14617);
or U15332 (N_15332,N_14964,N_14919);
or U15333 (N_15333,N_14773,N_14912);
nor U15334 (N_15334,N_14958,N_14690);
and U15335 (N_15335,N_14967,N_14639);
or U15336 (N_15336,N_14592,N_14999);
and U15337 (N_15337,N_14920,N_14886);
xnor U15338 (N_15338,N_14639,N_14693);
nor U15339 (N_15339,N_14996,N_14828);
and U15340 (N_15340,N_14596,N_14504);
or U15341 (N_15341,N_14841,N_14551);
xnor U15342 (N_15342,N_14825,N_14831);
or U15343 (N_15343,N_14844,N_14829);
and U15344 (N_15344,N_14628,N_14955);
nor U15345 (N_15345,N_14671,N_14685);
nand U15346 (N_15346,N_14590,N_14702);
or U15347 (N_15347,N_14976,N_14910);
xnor U15348 (N_15348,N_14962,N_14937);
or U15349 (N_15349,N_14511,N_14744);
nand U15350 (N_15350,N_14936,N_14647);
nor U15351 (N_15351,N_14593,N_14607);
and U15352 (N_15352,N_14630,N_14788);
xnor U15353 (N_15353,N_14715,N_14773);
or U15354 (N_15354,N_14996,N_14982);
nand U15355 (N_15355,N_14942,N_14965);
nor U15356 (N_15356,N_14933,N_14681);
and U15357 (N_15357,N_14537,N_14937);
and U15358 (N_15358,N_14596,N_14838);
nand U15359 (N_15359,N_14613,N_14923);
and U15360 (N_15360,N_14508,N_14766);
xor U15361 (N_15361,N_14732,N_14505);
nor U15362 (N_15362,N_14700,N_14749);
or U15363 (N_15363,N_14743,N_14698);
xor U15364 (N_15364,N_14621,N_14548);
nand U15365 (N_15365,N_14628,N_14830);
and U15366 (N_15366,N_14966,N_14734);
xnor U15367 (N_15367,N_14936,N_14619);
xor U15368 (N_15368,N_14838,N_14729);
and U15369 (N_15369,N_14623,N_14656);
nand U15370 (N_15370,N_14746,N_14923);
and U15371 (N_15371,N_14666,N_14715);
and U15372 (N_15372,N_14997,N_14896);
or U15373 (N_15373,N_14930,N_14556);
nand U15374 (N_15374,N_14784,N_14634);
nand U15375 (N_15375,N_14976,N_14860);
and U15376 (N_15376,N_14701,N_14822);
nor U15377 (N_15377,N_14955,N_14778);
nor U15378 (N_15378,N_14718,N_14513);
nor U15379 (N_15379,N_14978,N_14624);
and U15380 (N_15380,N_14991,N_14608);
and U15381 (N_15381,N_14623,N_14999);
nand U15382 (N_15382,N_14973,N_14710);
nand U15383 (N_15383,N_14986,N_14577);
and U15384 (N_15384,N_14732,N_14528);
nor U15385 (N_15385,N_14824,N_14606);
xnor U15386 (N_15386,N_14613,N_14616);
nor U15387 (N_15387,N_14759,N_14556);
and U15388 (N_15388,N_14760,N_14813);
xor U15389 (N_15389,N_14746,N_14983);
nand U15390 (N_15390,N_14789,N_14982);
or U15391 (N_15391,N_14975,N_14798);
nand U15392 (N_15392,N_14967,N_14828);
nor U15393 (N_15393,N_14718,N_14555);
nand U15394 (N_15394,N_14719,N_14669);
xnor U15395 (N_15395,N_14712,N_14586);
nor U15396 (N_15396,N_14768,N_14547);
and U15397 (N_15397,N_14662,N_14983);
xnor U15398 (N_15398,N_14718,N_14570);
xor U15399 (N_15399,N_14501,N_14550);
and U15400 (N_15400,N_14914,N_14842);
or U15401 (N_15401,N_14527,N_14661);
nand U15402 (N_15402,N_14942,N_14988);
xnor U15403 (N_15403,N_14765,N_14519);
and U15404 (N_15404,N_14860,N_14862);
nand U15405 (N_15405,N_14954,N_14561);
nor U15406 (N_15406,N_14946,N_14799);
nor U15407 (N_15407,N_14744,N_14560);
and U15408 (N_15408,N_14937,N_14888);
nand U15409 (N_15409,N_14958,N_14657);
xnor U15410 (N_15410,N_14531,N_14870);
or U15411 (N_15411,N_14918,N_14880);
or U15412 (N_15412,N_14644,N_14514);
nor U15413 (N_15413,N_14813,N_14992);
and U15414 (N_15414,N_14847,N_14819);
nand U15415 (N_15415,N_14808,N_14666);
xnor U15416 (N_15416,N_14774,N_14991);
nand U15417 (N_15417,N_14928,N_14612);
or U15418 (N_15418,N_14811,N_14809);
or U15419 (N_15419,N_14689,N_14663);
xnor U15420 (N_15420,N_14959,N_14671);
xnor U15421 (N_15421,N_14992,N_14916);
xor U15422 (N_15422,N_14807,N_14886);
and U15423 (N_15423,N_14702,N_14952);
xor U15424 (N_15424,N_14702,N_14608);
or U15425 (N_15425,N_14894,N_14760);
nor U15426 (N_15426,N_14684,N_14839);
or U15427 (N_15427,N_14807,N_14755);
nor U15428 (N_15428,N_14825,N_14845);
nand U15429 (N_15429,N_14998,N_14906);
nand U15430 (N_15430,N_14935,N_14668);
xnor U15431 (N_15431,N_14768,N_14809);
nor U15432 (N_15432,N_14773,N_14914);
or U15433 (N_15433,N_14531,N_14894);
or U15434 (N_15434,N_14930,N_14886);
xnor U15435 (N_15435,N_14641,N_14902);
xnor U15436 (N_15436,N_14931,N_14909);
and U15437 (N_15437,N_14784,N_14678);
nor U15438 (N_15438,N_14891,N_14651);
or U15439 (N_15439,N_14860,N_14703);
and U15440 (N_15440,N_14780,N_14523);
nand U15441 (N_15441,N_14914,N_14855);
and U15442 (N_15442,N_14527,N_14588);
xor U15443 (N_15443,N_14742,N_14530);
or U15444 (N_15444,N_14512,N_14921);
nand U15445 (N_15445,N_14730,N_14790);
or U15446 (N_15446,N_14523,N_14842);
or U15447 (N_15447,N_14854,N_14571);
nor U15448 (N_15448,N_14821,N_14751);
nor U15449 (N_15449,N_14717,N_14781);
nor U15450 (N_15450,N_14623,N_14678);
and U15451 (N_15451,N_14769,N_14910);
or U15452 (N_15452,N_14832,N_14530);
nand U15453 (N_15453,N_14700,N_14996);
nor U15454 (N_15454,N_14755,N_14756);
and U15455 (N_15455,N_14757,N_14527);
xnor U15456 (N_15456,N_14711,N_14518);
nor U15457 (N_15457,N_14828,N_14954);
or U15458 (N_15458,N_14883,N_14839);
or U15459 (N_15459,N_14668,N_14509);
and U15460 (N_15460,N_14626,N_14805);
xnor U15461 (N_15461,N_14866,N_14823);
xnor U15462 (N_15462,N_14709,N_14631);
and U15463 (N_15463,N_14743,N_14738);
nor U15464 (N_15464,N_14901,N_14528);
xnor U15465 (N_15465,N_14889,N_14975);
or U15466 (N_15466,N_14592,N_14767);
xor U15467 (N_15467,N_14636,N_14525);
xnor U15468 (N_15468,N_14836,N_14573);
xnor U15469 (N_15469,N_14928,N_14567);
or U15470 (N_15470,N_14623,N_14710);
xor U15471 (N_15471,N_14940,N_14659);
or U15472 (N_15472,N_14637,N_14911);
and U15473 (N_15473,N_14653,N_14568);
nor U15474 (N_15474,N_14904,N_14892);
xor U15475 (N_15475,N_14843,N_14658);
nand U15476 (N_15476,N_14916,N_14877);
or U15477 (N_15477,N_14784,N_14670);
nor U15478 (N_15478,N_14627,N_14605);
and U15479 (N_15479,N_14795,N_14971);
nor U15480 (N_15480,N_14947,N_14960);
nand U15481 (N_15481,N_14541,N_14842);
and U15482 (N_15482,N_14633,N_14998);
or U15483 (N_15483,N_14976,N_14940);
xnor U15484 (N_15484,N_14799,N_14834);
or U15485 (N_15485,N_14768,N_14762);
nand U15486 (N_15486,N_14517,N_14525);
and U15487 (N_15487,N_14686,N_14760);
and U15488 (N_15488,N_14712,N_14741);
nor U15489 (N_15489,N_14895,N_14847);
xnor U15490 (N_15490,N_14724,N_14837);
nand U15491 (N_15491,N_14805,N_14564);
xor U15492 (N_15492,N_14998,N_14816);
nor U15493 (N_15493,N_14677,N_14966);
and U15494 (N_15494,N_14680,N_14936);
and U15495 (N_15495,N_14530,N_14584);
xnor U15496 (N_15496,N_14948,N_14703);
nand U15497 (N_15497,N_14635,N_14932);
xnor U15498 (N_15498,N_14941,N_14904);
xnor U15499 (N_15499,N_14561,N_14554);
nand U15500 (N_15500,N_15365,N_15176);
nand U15501 (N_15501,N_15006,N_15455);
xor U15502 (N_15502,N_15045,N_15254);
or U15503 (N_15503,N_15380,N_15408);
or U15504 (N_15504,N_15312,N_15298);
and U15505 (N_15505,N_15160,N_15440);
nor U15506 (N_15506,N_15288,N_15063);
or U15507 (N_15507,N_15232,N_15208);
nand U15508 (N_15508,N_15200,N_15463);
xor U15509 (N_15509,N_15371,N_15084);
nand U15510 (N_15510,N_15235,N_15094);
or U15511 (N_15511,N_15489,N_15282);
xnor U15512 (N_15512,N_15396,N_15334);
and U15513 (N_15513,N_15303,N_15468);
or U15514 (N_15514,N_15086,N_15034);
or U15515 (N_15515,N_15442,N_15384);
and U15516 (N_15516,N_15467,N_15296);
nor U15517 (N_15517,N_15492,N_15243);
nand U15518 (N_15518,N_15238,N_15258);
or U15519 (N_15519,N_15026,N_15197);
xnor U15520 (N_15520,N_15327,N_15198);
and U15521 (N_15521,N_15141,N_15028);
xor U15522 (N_15522,N_15362,N_15255);
nand U15523 (N_15523,N_15432,N_15321);
or U15524 (N_15524,N_15175,N_15343);
nand U15525 (N_15525,N_15316,N_15195);
or U15526 (N_15526,N_15493,N_15484);
or U15527 (N_15527,N_15498,N_15302);
or U15528 (N_15528,N_15406,N_15054);
and U15529 (N_15529,N_15159,N_15415);
or U15530 (N_15530,N_15032,N_15212);
and U15531 (N_15531,N_15482,N_15333);
xor U15532 (N_15532,N_15444,N_15073);
nor U15533 (N_15533,N_15360,N_15130);
or U15534 (N_15534,N_15236,N_15477);
nand U15535 (N_15535,N_15250,N_15299);
nor U15536 (N_15536,N_15107,N_15438);
nor U15537 (N_15537,N_15252,N_15265);
nand U15538 (N_15538,N_15179,N_15125);
or U15539 (N_15539,N_15366,N_15337);
xor U15540 (N_15540,N_15330,N_15344);
and U15541 (N_15541,N_15486,N_15007);
or U15542 (N_15542,N_15354,N_15306);
nand U15543 (N_15543,N_15143,N_15319);
or U15544 (N_15544,N_15294,N_15244);
or U15545 (N_15545,N_15449,N_15429);
and U15546 (N_15546,N_15308,N_15199);
xnor U15547 (N_15547,N_15342,N_15188);
nand U15548 (N_15548,N_15348,N_15328);
and U15549 (N_15549,N_15091,N_15029);
nand U15550 (N_15550,N_15257,N_15012);
nor U15551 (N_15551,N_15315,N_15388);
nor U15552 (N_15552,N_15453,N_15120);
nand U15553 (N_15553,N_15456,N_15099);
nand U15554 (N_15554,N_15185,N_15205);
nor U15555 (N_15555,N_15428,N_15088);
xnor U15556 (N_15556,N_15046,N_15373);
nor U15557 (N_15557,N_15418,N_15065);
or U15558 (N_15558,N_15166,N_15237);
xnor U15559 (N_15559,N_15341,N_15022);
nand U15560 (N_15560,N_15136,N_15082);
or U15561 (N_15561,N_15309,N_15112);
nand U15562 (N_15562,N_15021,N_15289);
nand U15563 (N_15563,N_15119,N_15150);
or U15564 (N_15564,N_15056,N_15370);
or U15565 (N_15565,N_15109,N_15149);
and U15566 (N_15566,N_15496,N_15364);
xnor U15567 (N_15567,N_15009,N_15039);
nor U15568 (N_15568,N_15038,N_15284);
and U15569 (N_15569,N_15431,N_15051);
nor U15570 (N_15570,N_15071,N_15089);
nor U15571 (N_15571,N_15340,N_15245);
nor U15572 (N_15572,N_15399,N_15098);
or U15573 (N_15573,N_15350,N_15052);
nand U15574 (N_15574,N_15481,N_15019);
xnor U15575 (N_15575,N_15323,N_15173);
nand U15576 (N_15576,N_15192,N_15367);
xnor U15577 (N_15577,N_15147,N_15177);
nor U15578 (N_15578,N_15386,N_15471);
or U15579 (N_15579,N_15397,N_15215);
and U15580 (N_15580,N_15387,N_15181);
nand U15581 (N_15581,N_15118,N_15325);
xor U15582 (N_15582,N_15280,N_15152);
nor U15583 (N_15583,N_15078,N_15083);
nor U15584 (N_15584,N_15349,N_15356);
xnor U15585 (N_15585,N_15183,N_15033);
or U15586 (N_15586,N_15283,N_15223);
xnor U15587 (N_15587,N_15194,N_15322);
or U15588 (N_15588,N_15332,N_15115);
and U15589 (N_15589,N_15193,N_15300);
and U15590 (N_15590,N_15172,N_15233);
nand U15591 (N_15591,N_15382,N_15008);
nand U15592 (N_15592,N_15290,N_15357);
nor U15593 (N_15593,N_15097,N_15329);
nor U15594 (N_15594,N_15393,N_15405);
nand U15595 (N_15595,N_15003,N_15184);
nand U15596 (N_15596,N_15494,N_15117);
xor U15597 (N_15597,N_15291,N_15450);
xor U15598 (N_15598,N_15459,N_15355);
nor U15599 (N_15599,N_15155,N_15224);
nor U15600 (N_15600,N_15024,N_15129);
and U15601 (N_15601,N_15466,N_15196);
nor U15602 (N_15602,N_15170,N_15446);
xnor U15603 (N_15603,N_15018,N_15497);
xor U15604 (N_15604,N_15491,N_15042);
nand U15605 (N_15605,N_15061,N_15101);
nor U15606 (N_15606,N_15163,N_15400);
xnor U15607 (N_15607,N_15262,N_15269);
xnor U15608 (N_15608,N_15093,N_15417);
xor U15609 (N_15609,N_15404,N_15326);
and U15610 (N_15610,N_15499,N_15295);
and U15611 (N_15611,N_15377,N_15383);
nor U15612 (N_15612,N_15369,N_15451);
xnor U15613 (N_15613,N_15036,N_15372);
nor U15614 (N_15614,N_15487,N_15234);
or U15615 (N_15615,N_15148,N_15263);
xnor U15616 (N_15616,N_15347,N_15110);
or U15617 (N_15617,N_15128,N_15156);
and U15618 (N_15618,N_15320,N_15058);
and U15619 (N_15619,N_15087,N_15066);
nand U15620 (N_15620,N_15469,N_15273);
and U15621 (N_15621,N_15123,N_15113);
xnor U15622 (N_15622,N_15485,N_15047);
nand U15623 (N_15623,N_15394,N_15488);
and U15624 (N_15624,N_15030,N_15435);
or U15625 (N_15625,N_15075,N_15001);
or U15626 (N_15626,N_15165,N_15264);
and U15627 (N_15627,N_15043,N_15162);
nand U15628 (N_15628,N_15437,N_15187);
xor U15629 (N_15629,N_15070,N_15313);
nor U15630 (N_15630,N_15304,N_15127);
or U15631 (N_15631,N_15293,N_15168);
nor U15632 (N_15632,N_15297,N_15307);
nor U15633 (N_15633,N_15363,N_15274);
nor U15634 (N_15634,N_15324,N_15059);
nand U15635 (N_15635,N_15271,N_15311);
nor U15636 (N_15636,N_15100,N_15207);
and U15637 (N_15637,N_15241,N_15279);
or U15638 (N_15638,N_15014,N_15248);
nand U15639 (N_15639,N_15000,N_15220);
nor U15640 (N_15640,N_15085,N_15102);
or U15641 (N_15641,N_15409,N_15095);
nor U15642 (N_15642,N_15385,N_15005);
nor U15643 (N_15643,N_15457,N_15060);
nand U15644 (N_15644,N_15217,N_15436);
or U15645 (N_15645,N_15473,N_15214);
and U15646 (N_15646,N_15376,N_15253);
nand U15647 (N_15647,N_15227,N_15247);
nor U15648 (N_15648,N_15210,N_15031);
xnor U15649 (N_15649,N_15126,N_15144);
nand U15650 (N_15650,N_15398,N_15275);
nand U15651 (N_15651,N_15465,N_15229);
nor U15652 (N_15652,N_15490,N_15103);
or U15653 (N_15653,N_15260,N_15191);
and U15654 (N_15654,N_15202,N_15057);
nor U15655 (N_15655,N_15401,N_15424);
and U15656 (N_15656,N_15425,N_15226);
nand U15657 (N_15657,N_15483,N_15281);
nand U15658 (N_15658,N_15339,N_15142);
or U15659 (N_15659,N_15010,N_15368);
or U15660 (N_15660,N_15206,N_15246);
nor U15661 (N_15661,N_15211,N_15044);
nand U15662 (N_15662,N_15430,N_15461);
and U15663 (N_15663,N_15164,N_15413);
nand U15664 (N_15664,N_15203,N_15310);
xnor U15665 (N_15665,N_15351,N_15189);
nand U15666 (N_15666,N_15204,N_15104);
nand U15667 (N_15667,N_15261,N_15285);
and U15668 (N_15668,N_15267,N_15423);
nor U15669 (N_15669,N_15331,N_15020);
nor U15670 (N_15670,N_15420,N_15266);
and U15671 (N_15671,N_15472,N_15314);
nor U15672 (N_15672,N_15495,N_15190);
or U15673 (N_15673,N_15427,N_15439);
or U15674 (N_15674,N_15464,N_15378);
xnor U15675 (N_15675,N_15270,N_15055);
or U15676 (N_15676,N_15201,N_15338);
or U15677 (N_15677,N_15256,N_15259);
or U15678 (N_15678,N_15359,N_15422);
nand U15679 (N_15679,N_15135,N_15272);
and U15680 (N_15680,N_15452,N_15230);
nor U15681 (N_15681,N_15414,N_15157);
or U15682 (N_15682,N_15222,N_15301);
nand U15683 (N_15683,N_15426,N_15381);
xor U15684 (N_15684,N_15353,N_15004);
and U15685 (N_15685,N_15447,N_15096);
nor U15686 (N_15686,N_15092,N_15153);
or U15687 (N_15687,N_15268,N_15064);
xnor U15688 (N_15688,N_15434,N_15209);
and U15689 (N_15689,N_15286,N_15124);
nand U15690 (N_15690,N_15395,N_15475);
xor U15691 (N_15691,N_15225,N_15178);
or U15692 (N_15692,N_15167,N_15476);
nand U15693 (N_15693,N_15403,N_15011);
xor U15694 (N_15694,N_15015,N_15221);
nor U15695 (N_15695,N_15076,N_15174);
xor U15696 (N_15696,N_15037,N_15035);
or U15697 (N_15697,N_15421,N_15433);
or U15698 (N_15698,N_15375,N_15448);
xor U15699 (N_15699,N_15002,N_15345);
nand U15700 (N_15700,N_15231,N_15305);
nand U15701 (N_15701,N_15240,N_15049);
xor U15702 (N_15702,N_15138,N_15443);
xnor U15703 (N_15703,N_15287,N_15139);
and U15704 (N_15704,N_15242,N_15121);
and U15705 (N_15705,N_15016,N_15041);
and U15706 (N_15706,N_15480,N_15474);
nand U15707 (N_15707,N_15069,N_15278);
and U15708 (N_15708,N_15122,N_15186);
nor U15709 (N_15709,N_15470,N_15023);
xnor U15710 (N_15710,N_15412,N_15114);
xnor U15711 (N_15711,N_15068,N_15218);
nor U15712 (N_15712,N_15134,N_15392);
xor U15713 (N_15713,N_15140,N_15171);
or U15714 (N_15714,N_15374,N_15137);
and U15715 (N_15715,N_15111,N_15390);
xnor U15716 (N_15716,N_15182,N_15358);
nor U15717 (N_15717,N_15048,N_15458);
and U15718 (N_15718,N_15346,N_15335);
xnor U15719 (N_15719,N_15132,N_15276);
xor U15720 (N_15720,N_15454,N_15151);
nand U15721 (N_15721,N_15361,N_15249);
xor U15722 (N_15722,N_15219,N_15352);
or U15723 (N_15723,N_15062,N_15292);
or U15724 (N_15724,N_15462,N_15213);
nor U15725 (N_15725,N_15116,N_15145);
nand U15726 (N_15726,N_15228,N_15379);
nand U15727 (N_15727,N_15080,N_15146);
nand U15728 (N_15728,N_15251,N_15154);
or U15729 (N_15729,N_15389,N_15239);
nand U15730 (N_15730,N_15318,N_15277);
nor U15731 (N_15731,N_15013,N_15416);
or U15732 (N_15732,N_15441,N_15411);
and U15733 (N_15733,N_15040,N_15391);
and U15734 (N_15734,N_15108,N_15158);
nand U15735 (N_15735,N_15317,N_15407);
or U15736 (N_15736,N_15479,N_15410);
or U15737 (N_15737,N_15081,N_15402);
xnor U15738 (N_15738,N_15131,N_15050);
and U15739 (N_15739,N_15067,N_15027);
and U15740 (N_15740,N_15077,N_15169);
nor U15741 (N_15741,N_15336,N_15106);
nand U15742 (N_15742,N_15105,N_15017);
nor U15743 (N_15743,N_15090,N_15133);
or U15744 (N_15744,N_15161,N_15419);
xnor U15745 (N_15745,N_15460,N_15074);
or U15746 (N_15746,N_15079,N_15025);
nor U15747 (N_15747,N_15445,N_15478);
and U15748 (N_15748,N_15072,N_15180);
or U15749 (N_15749,N_15053,N_15216);
and U15750 (N_15750,N_15051,N_15379);
xnor U15751 (N_15751,N_15243,N_15347);
xnor U15752 (N_15752,N_15375,N_15077);
and U15753 (N_15753,N_15387,N_15381);
xor U15754 (N_15754,N_15357,N_15340);
nor U15755 (N_15755,N_15249,N_15167);
nor U15756 (N_15756,N_15017,N_15429);
xnor U15757 (N_15757,N_15344,N_15053);
xnor U15758 (N_15758,N_15158,N_15272);
nor U15759 (N_15759,N_15495,N_15045);
xnor U15760 (N_15760,N_15293,N_15497);
xor U15761 (N_15761,N_15384,N_15166);
and U15762 (N_15762,N_15304,N_15462);
xnor U15763 (N_15763,N_15026,N_15189);
xnor U15764 (N_15764,N_15084,N_15466);
and U15765 (N_15765,N_15049,N_15009);
xor U15766 (N_15766,N_15171,N_15349);
and U15767 (N_15767,N_15310,N_15489);
nand U15768 (N_15768,N_15003,N_15276);
xor U15769 (N_15769,N_15085,N_15014);
xnor U15770 (N_15770,N_15222,N_15188);
xor U15771 (N_15771,N_15042,N_15200);
nor U15772 (N_15772,N_15070,N_15387);
xnor U15773 (N_15773,N_15364,N_15310);
or U15774 (N_15774,N_15075,N_15276);
or U15775 (N_15775,N_15467,N_15311);
and U15776 (N_15776,N_15351,N_15421);
nand U15777 (N_15777,N_15318,N_15220);
nand U15778 (N_15778,N_15078,N_15284);
xnor U15779 (N_15779,N_15138,N_15477);
nor U15780 (N_15780,N_15073,N_15046);
xnor U15781 (N_15781,N_15274,N_15287);
nor U15782 (N_15782,N_15416,N_15077);
nand U15783 (N_15783,N_15412,N_15310);
and U15784 (N_15784,N_15127,N_15473);
xnor U15785 (N_15785,N_15166,N_15286);
xnor U15786 (N_15786,N_15091,N_15406);
xor U15787 (N_15787,N_15043,N_15312);
and U15788 (N_15788,N_15088,N_15448);
and U15789 (N_15789,N_15354,N_15202);
or U15790 (N_15790,N_15223,N_15146);
or U15791 (N_15791,N_15334,N_15257);
nand U15792 (N_15792,N_15347,N_15194);
nand U15793 (N_15793,N_15263,N_15447);
nand U15794 (N_15794,N_15360,N_15139);
and U15795 (N_15795,N_15229,N_15492);
nor U15796 (N_15796,N_15187,N_15446);
xnor U15797 (N_15797,N_15246,N_15135);
and U15798 (N_15798,N_15280,N_15418);
nand U15799 (N_15799,N_15340,N_15120);
or U15800 (N_15800,N_15097,N_15086);
xnor U15801 (N_15801,N_15431,N_15430);
nor U15802 (N_15802,N_15356,N_15122);
and U15803 (N_15803,N_15258,N_15422);
xnor U15804 (N_15804,N_15241,N_15278);
and U15805 (N_15805,N_15255,N_15470);
or U15806 (N_15806,N_15452,N_15075);
xnor U15807 (N_15807,N_15036,N_15464);
xnor U15808 (N_15808,N_15204,N_15334);
nor U15809 (N_15809,N_15106,N_15110);
or U15810 (N_15810,N_15443,N_15460);
xnor U15811 (N_15811,N_15386,N_15261);
and U15812 (N_15812,N_15099,N_15327);
xnor U15813 (N_15813,N_15246,N_15302);
and U15814 (N_15814,N_15398,N_15301);
nor U15815 (N_15815,N_15429,N_15096);
and U15816 (N_15816,N_15072,N_15235);
nor U15817 (N_15817,N_15198,N_15328);
nand U15818 (N_15818,N_15341,N_15403);
nor U15819 (N_15819,N_15402,N_15080);
xnor U15820 (N_15820,N_15158,N_15273);
xnor U15821 (N_15821,N_15224,N_15396);
nand U15822 (N_15822,N_15128,N_15413);
nand U15823 (N_15823,N_15054,N_15273);
nor U15824 (N_15824,N_15372,N_15261);
and U15825 (N_15825,N_15080,N_15380);
xnor U15826 (N_15826,N_15012,N_15469);
nand U15827 (N_15827,N_15494,N_15298);
xnor U15828 (N_15828,N_15006,N_15389);
and U15829 (N_15829,N_15203,N_15493);
and U15830 (N_15830,N_15196,N_15293);
xor U15831 (N_15831,N_15268,N_15384);
or U15832 (N_15832,N_15084,N_15388);
xor U15833 (N_15833,N_15349,N_15299);
xor U15834 (N_15834,N_15302,N_15311);
xor U15835 (N_15835,N_15027,N_15117);
or U15836 (N_15836,N_15113,N_15009);
or U15837 (N_15837,N_15207,N_15097);
nand U15838 (N_15838,N_15093,N_15196);
xnor U15839 (N_15839,N_15289,N_15142);
and U15840 (N_15840,N_15131,N_15440);
and U15841 (N_15841,N_15358,N_15110);
nor U15842 (N_15842,N_15371,N_15441);
xor U15843 (N_15843,N_15195,N_15489);
nor U15844 (N_15844,N_15413,N_15142);
nor U15845 (N_15845,N_15321,N_15093);
and U15846 (N_15846,N_15381,N_15194);
and U15847 (N_15847,N_15259,N_15436);
nand U15848 (N_15848,N_15358,N_15323);
nor U15849 (N_15849,N_15260,N_15299);
and U15850 (N_15850,N_15391,N_15342);
nor U15851 (N_15851,N_15279,N_15248);
nor U15852 (N_15852,N_15028,N_15092);
nand U15853 (N_15853,N_15441,N_15033);
or U15854 (N_15854,N_15431,N_15370);
xnor U15855 (N_15855,N_15326,N_15426);
xnor U15856 (N_15856,N_15196,N_15363);
nand U15857 (N_15857,N_15336,N_15210);
nand U15858 (N_15858,N_15225,N_15319);
xor U15859 (N_15859,N_15032,N_15197);
nor U15860 (N_15860,N_15058,N_15433);
and U15861 (N_15861,N_15041,N_15087);
xor U15862 (N_15862,N_15277,N_15255);
nor U15863 (N_15863,N_15353,N_15019);
nor U15864 (N_15864,N_15369,N_15420);
nand U15865 (N_15865,N_15072,N_15026);
xnor U15866 (N_15866,N_15365,N_15097);
xnor U15867 (N_15867,N_15449,N_15265);
and U15868 (N_15868,N_15236,N_15200);
and U15869 (N_15869,N_15341,N_15446);
xnor U15870 (N_15870,N_15071,N_15003);
and U15871 (N_15871,N_15172,N_15229);
xnor U15872 (N_15872,N_15283,N_15041);
or U15873 (N_15873,N_15102,N_15419);
nand U15874 (N_15874,N_15192,N_15139);
xor U15875 (N_15875,N_15119,N_15495);
nand U15876 (N_15876,N_15288,N_15395);
nand U15877 (N_15877,N_15241,N_15211);
nor U15878 (N_15878,N_15116,N_15205);
or U15879 (N_15879,N_15055,N_15046);
nor U15880 (N_15880,N_15495,N_15157);
nor U15881 (N_15881,N_15346,N_15088);
or U15882 (N_15882,N_15070,N_15116);
nor U15883 (N_15883,N_15222,N_15004);
and U15884 (N_15884,N_15274,N_15223);
or U15885 (N_15885,N_15163,N_15391);
nand U15886 (N_15886,N_15149,N_15031);
or U15887 (N_15887,N_15262,N_15032);
and U15888 (N_15888,N_15165,N_15347);
nand U15889 (N_15889,N_15192,N_15477);
or U15890 (N_15890,N_15079,N_15154);
and U15891 (N_15891,N_15179,N_15186);
or U15892 (N_15892,N_15252,N_15333);
nand U15893 (N_15893,N_15339,N_15207);
xnor U15894 (N_15894,N_15144,N_15300);
nand U15895 (N_15895,N_15141,N_15375);
nand U15896 (N_15896,N_15066,N_15272);
nand U15897 (N_15897,N_15213,N_15165);
xor U15898 (N_15898,N_15449,N_15037);
nor U15899 (N_15899,N_15407,N_15467);
nor U15900 (N_15900,N_15205,N_15415);
or U15901 (N_15901,N_15124,N_15482);
nor U15902 (N_15902,N_15189,N_15313);
nor U15903 (N_15903,N_15180,N_15371);
and U15904 (N_15904,N_15061,N_15372);
nand U15905 (N_15905,N_15252,N_15476);
nand U15906 (N_15906,N_15113,N_15363);
xor U15907 (N_15907,N_15088,N_15187);
nand U15908 (N_15908,N_15488,N_15314);
nor U15909 (N_15909,N_15300,N_15274);
nand U15910 (N_15910,N_15399,N_15387);
and U15911 (N_15911,N_15324,N_15188);
nor U15912 (N_15912,N_15218,N_15487);
and U15913 (N_15913,N_15307,N_15241);
and U15914 (N_15914,N_15138,N_15168);
nor U15915 (N_15915,N_15331,N_15000);
xnor U15916 (N_15916,N_15193,N_15120);
or U15917 (N_15917,N_15363,N_15370);
or U15918 (N_15918,N_15082,N_15335);
or U15919 (N_15919,N_15337,N_15047);
nand U15920 (N_15920,N_15334,N_15060);
nor U15921 (N_15921,N_15455,N_15307);
and U15922 (N_15922,N_15464,N_15325);
xnor U15923 (N_15923,N_15097,N_15211);
nor U15924 (N_15924,N_15495,N_15444);
xnor U15925 (N_15925,N_15307,N_15070);
nand U15926 (N_15926,N_15186,N_15096);
nor U15927 (N_15927,N_15396,N_15435);
nand U15928 (N_15928,N_15326,N_15202);
nor U15929 (N_15929,N_15114,N_15338);
and U15930 (N_15930,N_15053,N_15284);
xnor U15931 (N_15931,N_15107,N_15496);
and U15932 (N_15932,N_15131,N_15492);
nand U15933 (N_15933,N_15185,N_15239);
nor U15934 (N_15934,N_15330,N_15206);
nor U15935 (N_15935,N_15401,N_15000);
and U15936 (N_15936,N_15373,N_15111);
nor U15937 (N_15937,N_15309,N_15268);
nand U15938 (N_15938,N_15205,N_15037);
nor U15939 (N_15939,N_15284,N_15223);
nand U15940 (N_15940,N_15095,N_15098);
nand U15941 (N_15941,N_15431,N_15122);
and U15942 (N_15942,N_15372,N_15386);
nor U15943 (N_15943,N_15079,N_15081);
xor U15944 (N_15944,N_15196,N_15477);
or U15945 (N_15945,N_15176,N_15234);
nor U15946 (N_15946,N_15055,N_15479);
and U15947 (N_15947,N_15479,N_15119);
and U15948 (N_15948,N_15115,N_15070);
nor U15949 (N_15949,N_15414,N_15007);
nor U15950 (N_15950,N_15331,N_15264);
xnor U15951 (N_15951,N_15429,N_15452);
nor U15952 (N_15952,N_15356,N_15120);
xnor U15953 (N_15953,N_15200,N_15145);
or U15954 (N_15954,N_15322,N_15280);
nand U15955 (N_15955,N_15306,N_15463);
nor U15956 (N_15956,N_15093,N_15490);
and U15957 (N_15957,N_15135,N_15025);
nand U15958 (N_15958,N_15411,N_15143);
xnor U15959 (N_15959,N_15456,N_15153);
nand U15960 (N_15960,N_15201,N_15447);
nand U15961 (N_15961,N_15427,N_15167);
and U15962 (N_15962,N_15362,N_15048);
or U15963 (N_15963,N_15178,N_15327);
and U15964 (N_15964,N_15377,N_15440);
xor U15965 (N_15965,N_15431,N_15295);
xor U15966 (N_15966,N_15482,N_15161);
nor U15967 (N_15967,N_15113,N_15455);
or U15968 (N_15968,N_15488,N_15352);
nand U15969 (N_15969,N_15317,N_15285);
nor U15970 (N_15970,N_15311,N_15281);
and U15971 (N_15971,N_15485,N_15089);
nor U15972 (N_15972,N_15291,N_15377);
or U15973 (N_15973,N_15022,N_15206);
xnor U15974 (N_15974,N_15314,N_15437);
nor U15975 (N_15975,N_15155,N_15009);
nor U15976 (N_15976,N_15121,N_15452);
nor U15977 (N_15977,N_15344,N_15400);
and U15978 (N_15978,N_15133,N_15031);
nand U15979 (N_15979,N_15173,N_15249);
and U15980 (N_15980,N_15286,N_15078);
or U15981 (N_15981,N_15046,N_15065);
and U15982 (N_15982,N_15464,N_15479);
or U15983 (N_15983,N_15472,N_15097);
xor U15984 (N_15984,N_15290,N_15404);
xnor U15985 (N_15985,N_15369,N_15464);
nand U15986 (N_15986,N_15012,N_15136);
nand U15987 (N_15987,N_15318,N_15090);
nor U15988 (N_15988,N_15353,N_15084);
nor U15989 (N_15989,N_15251,N_15167);
nor U15990 (N_15990,N_15190,N_15266);
or U15991 (N_15991,N_15480,N_15287);
nor U15992 (N_15992,N_15116,N_15245);
and U15993 (N_15993,N_15253,N_15109);
nor U15994 (N_15994,N_15334,N_15189);
nor U15995 (N_15995,N_15209,N_15293);
nand U15996 (N_15996,N_15478,N_15097);
nand U15997 (N_15997,N_15113,N_15377);
and U15998 (N_15998,N_15055,N_15209);
and U15999 (N_15999,N_15475,N_15008);
nand U16000 (N_16000,N_15862,N_15704);
xnor U16001 (N_16001,N_15760,N_15971);
nand U16002 (N_16002,N_15961,N_15608);
nand U16003 (N_16003,N_15908,N_15929);
nand U16004 (N_16004,N_15810,N_15831);
nor U16005 (N_16005,N_15906,N_15772);
nor U16006 (N_16006,N_15545,N_15999);
nand U16007 (N_16007,N_15617,N_15668);
nor U16008 (N_16008,N_15719,N_15991);
nor U16009 (N_16009,N_15875,N_15866);
xnor U16010 (N_16010,N_15652,N_15599);
xnor U16011 (N_16011,N_15918,N_15634);
nor U16012 (N_16012,N_15843,N_15542);
xor U16013 (N_16013,N_15680,N_15824);
or U16014 (N_16014,N_15664,N_15882);
and U16015 (N_16015,N_15763,N_15820);
and U16016 (N_16016,N_15586,N_15839);
xnor U16017 (N_16017,N_15658,N_15636);
and U16018 (N_16018,N_15770,N_15960);
and U16019 (N_16019,N_15932,N_15534);
or U16020 (N_16020,N_15877,N_15907);
nand U16021 (N_16021,N_15565,N_15830);
nor U16022 (N_16022,N_15854,N_15757);
xnor U16023 (N_16023,N_15879,N_15611);
or U16024 (N_16024,N_15792,N_15793);
or U16025 (N_16025,N_15712,N_15524);
nand U16026 (N_16026,N_15989,N_15963);
nor U16027 (N_16027,N_15616,N_15627);
and U16028 (N_16028,N_15531,N_15937);
nor U16029 (N_16029,N_15525,N_15596);
or U16030 (N_16030,N_15728,N_15613);
nand U16031 (N_16031,N_15628,N_15642);
nand U16032 (N_16032,N_15694,N_15501);
or U16033 (N_16033,N_15519,N_15859);
nand U16034 (N_16034,N_15836,N_15709);
or U16035 (N_16035,N_15602,N_15701);
and U16036 (N_16036,N_15548,N_15997);
or U16037 (N_16037,N_15902,N_15729);
nand U16038 (N_16038,N_15746,N_15603);
and U16039 (N_16039,N_15646,N_15780);
nand U16040 (N_16040,N_15752,N_15953);
or U16041 (N_16041,N_15607,N_15923);
and U16042 (N_16042,N_15696,N_15789);
or U16043 (N_16043,N_15678,N_15853);
or U16044 (N_16044,N_15576,N_15969);
or U16045 (N_16045,N_15684,N_15523);
or U16046 (N_16046,N_15822,N_15884);
or U16047 (N_16047,N_15503,N_15685);
or U16048 (N_16048,N_15919,N_15865);
xor U16049 (N_16049,N_15732,N_15869);
or U16050 (N_16050,N_15972,N_15952);
and U16051 (N_16051,N_15895,N_15549);
nor U16052 (N_16052,N_15625,N_15957);
or U16053 (N_16053,N_15977,N_15687);
xnor U16054 (N_16054,N_15659,N_15816);
nor U16055 (N_16055,N_15814,N_15842);
or U16056 (N_16056,N_15676,N_15898);
and U16057 (N_16057,N_15921,N_15914);
nand U16058 (N_16058,N_15809,N_15964);
xnor U16059 (N_16059,N_15554,N_15618);
and U16060 (N_16060,N_15691,N_15753);
nand U16061 (N_16061,N_15858,N_15569);
and U16062 (N_16062,N_15871,N_15594);
and U16063 (N_16063,N_15744,N_15716);
xnor U16064 (N_16064,N_15748,N_15689);
nor U16065 (N_16065,N_15801,N_15837);
nor U16066 (N_16066,N_15825,N_15998);
nand U16067 (N_16067,N_15551,N_15868);
or U16068 (N_16068,N_15773,N_15638);
and U16069 (N_16069,N_15890,N_15720);
nor U16070 (N_16070,N_15734,N_15872);
nor U16071 (N_16071,N_15873,N_15841);
nor U16072 (N_16072,N_15870,N_15894);
xnor U16073 (N_16073,N_15813,N_15582);
nand U16074 (N_16074,N_15624,N_15899);
xor U16075 (N_16075,N_15940,N_15537);
nor U16076 (N_16076,N_15555,N_15591);
or U16077 (N_16077,N_15677,N_15727);
or U16078 (N_16078,N_15718,N_15821);
and U16079 (N_16079,N_15572,N_15891);
nand U16080 (N_16080,N_15955,N_15665);
xor U16081 (N_16081,N_15754,N_15568);
nand U16082 (N_16082,N_15775,N_15897);
and U16083 (N_16083,N_15838,N_15946);
or U16084 (N_16084,N_15654,N_15769);
xor U16085 (N_16085,N_15896,N_15833);
nand U16086 (N_16086,N_15550,N_15776);
or U16087 (N_16087,N_15655,N_15571);
and U16088 (N_16088,N_15751,N_15553);
nand U16089 (N_16089,N_15818,N_15578);
nor U16090 (N_16090,N_15745,N_15847);
xnor U16091 (N_16091,N_15970,N_15788);
nor U16092 (N_16092,N_15812,N_15823);
nor U16093 (N_16093,N_15798,N_15924);
nor U16094 (N_16094,N_15768,N_15593);
nand U16095 (N_16095,N_15679,N_15826);
or U16096 (N_16096,N_15736,N_15543);
xnor U16097 (N_16097,N_15700,N_15533);
nor U16098 (N_16098,N_15583,N_15855);
or U16099 (N_16099,N_15589,N_15947);
xor U16100 (N_16100,N_15850,N_15620);
xnor U16101 (N_16101,N_15885,N_15633);
nand U16102 (N_16102,N_15771,N_15962);
and U16103 (N_16103,N_15874,N_15883);
xnor U16104 (N_16104,N_15673,N_15614);
nor U16105 (N_16105,N_15755,N_15632);
or U16106 (N_16106,N_15990,N_15721);
xor U16107 (N_16107,N_15939,N_15669);
xor U16108 (N_16108,N_15817,N_15804);
nor U16109 (N_16109,N_15764,N_15925);
xor U16110 (N_16110,N_15711,N_15693);
or U16111 (N_16111,N_15791,N_15705);
and U16112 (N_16112,N_15723,N_15795);
nand U16113 (N_16113,N_15520,N_15640);
and U16114 (N_16114,N_15735,N_15560);
or U16115 (N_16115,N_15846,N_15592);
xor U16116 (N_16116,N_15856,N_15819);
and U16117 (N_16117,N_15861,N_15522);
nand U16118 (N_16118,N_15767,N_15922);
nor U16119 (N_16119,N_15845,N_15670);
nor U16120 (N_16120,N_15504,N_15892);
nor U16121 (N_16121,N_15889,N_15913);
or U16122 (N_16122,N_15710,N_15660);
or U16123 (N_16123,N_15852,N_15546);
xor U16124 (N_16124,N_15849,N_15597);
nand U16125 (N_16125,N_15725,N_15781);
nor U16126 (N_16126,N_15917,N_15815);
nor U16127 (N_16127,N_15623,N_15629);
nand U16128 (N_16128,N_15888,N_15994);
and U16129 (N_16129,N_15948,N_15790);
nand U16130 (N_16130,N_15967,N_15564);
or U16131 (N_16131,N_15695,N_15581);
xor U16132 (N_16132,N_15675,N_15797);
nor U16133 (N_16133,N_15510,N_15527);
xnor U16134 (N_16134,N_15714,N_15517);
nor U16135 (N_16135,N_15979,N_15794);
nor U16136 (N_16136,N_15615,N_15552);
nand U16137 (N_16137,N_15762,N_15686);
nand U16138 (N_16138,N_15683,N_15784);
nand U16139 (N_16139,N_15577,N_15635);
or U16140 (N_16140,N_15749,N_15667);
nor U16141 (N_16141,N_15706,N_15600);
xnor U16142 (N_16142,N_15807,N_15742);
or U16143 (N_16143,N_15730,N_15834);
and U16144 (N_16144,N_15645,N_15938);
nand U16145 (N_16145,N_15766,N_15587);
and U16146 (N_16146,N_15876,N_15502);
and U16147 (N_16147,N_15713,N_15828);
or U16148 (N_16148,N_15765,N_15648);
nand U16149 (N_16149,N_15561,N_15911);
nor U16150 (N_16150,N_15738,N_15909);
nor U16151 (N_16151,N_15787,N_15905);
nor U16152 (N_16152,N_15521,N_15530);
nand U16153 (N_16153,N_15777,N_15500);
or U16154 (N_16154,N_15563,N_15604);
nor U16155 (N_16155,N_15848,N_15556);
xor U16156 (N_16156,N_15631,N_15987);
nand U16157 (N_16157,N_15860,N_15547);
and U16158 (N_16158,N_15539,N_15538);
or U16159 (N_16159,N_15980,N_15681);
and U16160 (N_16160,N_15944,N_15993);
nor U16161 (N_16161,N_15630,N_15590);
nor U16162 (N_16162,N_15863,N_15936);
or U16163 (N_16163,N_15601,N_15799);
nor U16164 (N_16164,N_15880,N_15942);
or U16165 (N_16165,N_15786,N_15573);
or U16166 (N_16166,N_15513,N_15647);
nand U16167 (N_16167,N_15536,N_15605);
nor U16168 (N_16168,N_15509,N_15579);
xnor U16169 (N_16169,N_15697,N_15674);
or U16170 (N_16170,N_15698,N_15912);
or U16171 (N_16171,N_15619,N_15878);
nor U16172 (N_16172,N_15835,N_15506);
or U16173 (N_16173,N_15759,N_15639);
xor U16174 (N_16174,N_15988,N_15945);
or U16175 (N_16175,N_15588,N_15900);
and U16176 (N_16176,N_15887,N_15951);
and U16177 (N_16177,N_15796,N_15805);
and U16178 (N_16178,N_15622,N_15950);
nand U16179 (N_16179,N_15644,N_15926);
nor U16180 (N_16180,N_15933,N_15982);
xnor U16181 (N_16181,N_15731,N_15692);
nand U16182 (N_16182,N_15558,N_15935);
and U16183 (N_16183,N_15934,N_15965);
and U16184 (N_16184,N_15996,N_15575);
xor U16185 (N_16185,N_15682,N_15507);
and U16186 (N_16186,N_15661,N_15761);
and U16187 (N_16187,N_15505,N_15584);
and U16188 (N_16188,N_15832,N_15840);
or U16189 (N_16189,N_15881,N_15612);
xnor U16190 (N_16190,N_15528,N_15785);
or U16191 (N_16191,N_15928,N_15574);
nand U16192 (N_16192,N_15904,N_15983);
nor U16193 (N_16193,N_15978,N_15708);
and U16194 (N_16194,N_15741,N_15740);
or U16195 (N_16195,N_15756,N_15956);
xnor U16196 (N_16196,N_15702,N_15526);
or U16197 (N_16197,N_15782,N_15920);
or U16198 (N_16198,N_15915,N_15653);
and U16199 (N_16199,N_15610,N_15974);
nor U16200 (N_16200,N_15535,N_15690);
xor U16201 (N_16201,N_15518,N_15540);
xor U16202 (N_16202,N_15717,N_15949);
or U16203 (N_16203,N_15808,N_15585);
nor U16204 (N_16204,N_15570,N_15910);
or U16205 (N_16205,N_15606,N_15774);
and U16206 (N_16206,N_15515,N_15943);
nand U16207 (N_16207,N_15778,N_15566);
nand U16208 (N_16208,N_15688,N_15511);
xor U16209 (N_16209,N_15722,N_15986);
nand U16210 (N_16210,N_15995,N_15626);
xor U16211 (N_16211,N_15637,N_15886);
or U16212 (N_16212,N_15671,N_15802);
or U16213 (N_16213,N_15739,N_15643);
nand U16214 (N_16214,N_15544,N_15609);
and U16215 (N_16215,N_15514,N_15743);
nor U16216 (N_16216,N_15985,N_15975);
xor U16217 (N_16217,N_15595,N_15901);
xor U16218 (N_16218,N_15529,N_15779);
nand U16219 (N_16219,N_15541,N_15783);
nor U16220 (N_16220,N_15973,N_15981);
and U16221 (N_16221,N_15703,N_15747);
xor U16222 (N_16222,N_15567,N_15984);
or U16223 (N_16223,N_15829,N_15666);
and U16224 (N_16224,N_15893,N_15656);
and U16225 (N_16225,N_15508,N_15532);
xor U16226 (N_16226,N_15737,N_15844);
xor U16227 (N_16227,N_15966,N_15724);
or U16228 (N_16228,N_15516,N_15959);
xor U16229 (N_16229,N_15707,N_15657);
nand U16230 (N_16230,N_15954,N_15851);
xnor U16231 (N_16231,N_15916,N_15976);
nor U16232 (N_16232,N_15857,N_15650);
xor U16233 (N_16233,N_15931,N_15699);
or U16234 (N_16234,N_15733,N_15559);
or U16235 (N_16235,N_15750,N_15715);
and U16236 (N_16236,N_15649,N_15811);
nor U16237 (N_16237,N_15927,N_15580);
nand U16238 (N_16238,N_15598,N_15672);
nand U16239 (N_16239,N_15562,N_15512);
xor U16240 (N_16240,N_15903,N_15641);
and U16241 (N_16241,N_15800,N_15557);
nor U16242 (N_16242,N_15651,N_15621);
and U16243 (N_16243,N_15941,N_15758);
xor U16244 (N_16244,N_15726,N_15992);
and U16245 (N_16245,N_15806,N_15958);
nor U16246 (N_16246,N_15864,N_15803);
and U16247 (N_16247,N_15968,N_15827);
nor U16248 (N_16248,N_15930,N_15663);
or U16249 (N_16249,N_15662,N_15867);
nand U16250 (N_16250,N_15980,N_15734);
xor U16251 (N_16251,N_15924,N_15609);
or U16252 (N_16252,N_15918,N_15830);
xor U16253 (N_16253,N_15972,N_15966);
and U16254 (N_16254,N_15892,N_15919);
nor U16255 (N_16255,N_15970,N_15822);
xnor U16256 (N_16256,N_15899,N_15862);
or U16257 (N_16257,N_15855,N_15924);
or U16258 (N_16258,N_15665,N_15996);
nand U16259 (N_16259,N_15978,N_15889);
and U16260 (N_16260,N_15877,N_15501);
and U16261 (N_16261,N_15587,N_15673);
nand U16262 (N_16262,N_15778,N_15915);
nor U16263 (N_16263,N_15765,N_15913);
nor U16264 (N_16264,N_15806,N_15851);
and U16265 (N_16265,N_15884,N_15924);
and U16266 (N_16266,N_15927,N_15547);
xnor U16267 (N_16267,N_15640,N_15554);
xor U16268 (N_16268,N_15972,N_15983);
nor U16269 (N_16269,N_15650,N_15646);
xnor U16270 (N_16270,N_15535,N_15937);
xnor U16271 (N_16271,N_15813,N_15745);
or U16272 (N_16272,N_15772,N_15524);
and U16273 (N_16273,N_15854,N_15733);
xnor U16274 (N_16274,N_15794,N_15739);
or U16275 (N_16275,N_15583,N_15531);
and U16276 (N_16276,N_15980,N_15744);
or U16277 (N_16277,N_15743,N_15798);
and U16278 (N_16278,N_15916,N_15512);
nor U16279 (N_16279,N_15595,N_15978);
nor U16280 (N_16280,N_15991,N_15557);
xor U16281 (N_16281,N_15505,N_15767);
or U16282 (N_16282,N_15569,N_15825);
nor U16283 (N_16283,N_15688,N_15535);
xnor U16284 (N_16284,N_15675,N_15602);
and U16285 (N_16285,N_15711,N_15953);
and U16286 (N_16286,N_15798,N_15943);
nand U16287 (N_16287,N_15901,N_15564);
and U16288 (N_16288,N_15945,N_15710);
nor U16289 (N_16289,N_15985,N_15628);
or U16290 (N_16290,N_15858,N_15592);
or U16291 (N_16291,N_15825,N_15925);
and U16292 (N_16292,N_15865,N_15632);
and U16293 (N_16293,N_15567,N_15991);
nand U16294 (N_16294,N_15756,N_15534);
and U16295 (N_16295,N_15862,N_15596);
nand U16296 (N_16296,N_15909,N_15747);
nor U16297 (N_16297,N_15945,N_15560);
or U16298 (N_16298,N_15817,N_15556);
nor U16299 (N_16299,N_15909,N_15625);
xor U16300 (N_16300,N_15857,N_15861);
xnor U16301 (N_16301,N_15668,N_15951);
and U16302 (N_16302,N_15841,N_15556);
xnor U16303 (N_16303,N_15666,N_15693);
xnor U16304 (N_16304,N_15507,N_15698);
nor U16305 (N_16305,N_15691,N_15660);
nand U16306 (N_16306,N_15835,N_15781);
xor U16307 (N_16307,N_15952,N_15888);
or U16308 (N_16308,N_15775,N_15627);
or U16309 (N_16309,N_15625,N_15986);
and U16310 (N_16310,N_15717,N_15640);
nor U16311 (N_16311,N_15777,N_15721);
xor U16312 (N_16312,N_15874,N_15971);
and U16313 (N_16313,N_15835,N_15981);
xor U16314 (N_16314,N_15870,N_15973);
or U16315 (N_16315,N_15895,N_15946);
nand U16316 (N_16316,N_15599,N_15879);
nand U16317 (N_16317,N_15768,N_15884);
nor U16318 (N_16318,N_15684,N_15965);
nand U16319 (N_16319,N_15719,N_15886);
nor U16320 (N_16320,N_15811,N_15837);
nor U16321 (N_16321,N_15578,N_15634);
xnor U16322 (N_16322,N_15634,N_15523);
nand U16323 (N_16323,N_15849,N_15755);
xor U16324 (N_16324,N_15637,N_15802);
and U16325 (N_16325,N_15723,N_15777);
or U16326 (N_16326,N_15925,N_15820);
or U16327 (N_16327,N_15942,N_15749);
xor U16328 (N_16328,N_15785,N_15614);
and U16329 (N_16329,N_15518,N_15888);
nor U16330 (N_16330,N_15607,N_15513);
or U16331 (N_16331,N_15746,N_15821);
nor U16332 (N_16332,N_15559,N_15720);
nor U16333 (N_16333,N_15713,N_15899);
or U16334 (N_16334,N_15554,N_15648);
or U16335 (N_16335,N_15771,N_15645);
and U16336 (N_16336,N_15922,N_15662);
and U16337 (N_16337,N_15901,N_15952);
and U16338 (N_16338,N_15642,N_15901);
or U16339 (N_16339,N_15670,N_15781);
xnor U16340 (N_16340,N_15794,N_15909);
nand U16341 (N_16341,N_15520,N_15864);
nor U16342 (N_16342,N_15861,N_15736);
nand U16343 (N_16343,N_15579,N_15893);
nor U16344 (N_16344,N_15811,N_15782);
nand U16345 (N_16345,N_15955,N_15587);
and U16346 (N_16346,N_15954,N_15831);
and U16347 (N_16347,N_15801,N_15666);
nor U16348 (N_16348,N_15575,N_15521);
nor U16349 (N_16349,N_15829,N_15705);
nand U16350 (N_16350,N_15652,N_15777);
or U16351 (N_16351,N_15864,N_15555);
nand U16352 (N_16352,N_15562,N_15567);
and U16353 (N_16353,N_15797,N_15584);
nand U16354 (N_16354,N_15859,N_15967);
nor U16355 (N_16355,N_15831,N_15981);
nor U16356 (N_16356,N_15694,N_15525);
nor U16357 (N_16357,N_15702,N_15761);
nor U16358 (N_16358,N_15985,N_15870);
or U16359 (N_16359,N_15641,N_15969);
nand U16360 (N_16360,N_15918,N_15502);
nand U16361 (N_16361,N_15965,N_15875);
nor U16362 (N_16362,N_15884,N_15896);
nand U16363 (N_16363,N_15574,N_15693);
xor U16364 (N_16364,N_15804,N_15725);
xnor U16365 (N_16365,N_15805,N_15685);
nand U16366 (N_16366,N_15588,N_15637);
or U16367 (N_16367,N_15730,N_15733);
nand U16368 (N_16368,N_15997,N_15809);
nor U16369 (N_16369,N_15597,N_15896);
and U16370 (N_16370,N_15742,N_15821);
nand U16371 (N_16371,N_15582,N_15945);
xor U16372 (N_16372,N_15807,N_15898);
xor U16373 (N_16373,N_15747,N_15527);
nand U16374 (N_16374,N_15896,N_15827);
or U16375 (N_16375,N_15563,N_15597);
nor U16376 (N_16376,N_15882,N_15666);
and U16377 (N_16377,N_15623,N_15898);
nor U16378 (N_16378,N_15855,N_15666);
and U16379 (N_16379,N_15734,N_15994);
xor U16380 (N_16380,N_15951,N_15730);
nand U16381 (N_16381,N_15913,N_15891);
xnor U16382 (N_16382,N_15561,N_15546);
xor U16383 (N_16383,N_15596,N_15626);
xnor U16384 (N_16384,N_15589,N_15615);
xor U16385 (N_16385,N_15693,N_15686);
nand U16386 (N_16386,N_15768,N_15674);
xor U16387 (N_16387,N_15555,N_15644);
and U16388 (N_16388,N_15846,N_15812);
xnor U16389 (N_16389,N_15876,N_15878);
xor U16390 (N_16390,N_15934,N_15673);
and U16391 (N_16391,N_15595,N_15946);
and U16392 (N_16392,N_15831,N_15568);
or U16393 (N_16393,N_15754,N_15550);
nand U16394 (N_16394,N_15684,N_15829);
nor U16395 (N_16395,N_15763,N_15561);
nor U16396 (N_16396,N_15511,N_15768);
nor U16397 (N_16397,N_15574,N_15877);
xor U16398 (N_16398,N_15596,N_15529);
nand U16399 (N_16399,N_15905,N_15844);
nand U16400 (N_16400,N_15645,N_15964);
nor U16401 (N_16401,N_15554,N_15582);
nand U16402 (N_16402,N_15773,N_15785);
nor U16403 (N_16403,N_15646,N_15661);
xor U16404 (N_16404,N_15631,N_15540);
xnor U16405 (N_16405,N_15708,N_15936);
and U16406 (N_16406,N_15646,N_15578);
xor U16407 (N_16407,N_15739,N_15761);
nand U16408 (N_16408,N_15702,N_15810);
and U16409 (N_16409,N_15576,N_15951);
and U16410 (N_16410,N_15525,N_15763);
and U16411 (N_16411,N_15598,N_15836);
nor U16412 (N_16412,N_15905,N_15828);
or U16413 (N_16413,N_15914,N_15952);
xor U16414 (N_16414,N_15581,N_15948);
nor U16415 (N_16415,N_15633,N_15916);
or U16416 (N_16416,N_15560,N_15814);
nor U16417 (N_16417,N_15769,N_15893);
xnor U16418 (N_16418,N_15616,N_15677);
and U16419 (N_16419,N_15875,N_15767);
or U16420 (N_16420,N_15522,N_15649);
nand U16421 (N_16421,N_15551,N_15959);
or U16422 (N_16422,N_15529,N_15917);
or U16423 (N_16423,N_15900,N_15736);
nand U16424 (N_16424,N_15822,N_15588);
nand U16425 (N_16425,N_15827,N_15788);
and U16426 (N_16426,N_15813,N_15837);
or U16427 (N_16427,N_15564,N_15809);
or U16428 (N_16428,N_15602,N_15952);
xor U16429 (N_16429,N_15679,N_15798);
or U16430 (N_16430,N_15895,N_15503);
nor U16431 (N_16431,N_15563,N_15608);
nand U16432 (N_16432,N_15721,N_15607);
or U16433 (N_16433,N_15590,N_15860);
or U16434 (N_16434,N_15950,N_15653);
nor U16435 (N_16435,N_15964,N_15935);
nor U16436 (N_16436,N_15963,N_15665);
or U16437 (N_16437,N_15705,N_15701);
and U16438 (N_16438,N_15760,N_15642);
or U16439 (N_16439,N_15961,N_15763);
nor U16440 (N_16440,N_15809,N_15548);
nor U16441 (N_16441,N_15780,N_15664);
or U16442 (N_16442,N_15558,N_15672);
nand U16443 (N_16443,N_15956,N_15561);
and U16444 (N_16444,N_15522,N_15920);
nor U16445 (N_16445,N_15779,N_15549);
or U16446 (N_16446,N_15573,N_15803);
and U16447 (N_16447,N_15810,N_15672);
nor U16448 (N_16448,N_15501,N_15720);
nand U16449 (N_16449,N_15700,N_15656);
and U16450 (N_16450,N_15579,N_15835);
nor U16451 (N_16451,N_15523,N_15841);
nand U16452 (N_16452,N_15811,N_15817);
and U16453 (N_16453,N_15558,N_15646);
xor U16454 (N_16454,N_15578,N_15964);
nor U16455 (N_16455,N_15611,N_15825);
nand U16456 (N_16456,N_15998,N_15936);
or U16457 (N_16457,N_15739,N_15903);
nand U16458 (N_16458,N_15580,N_15592);
xor U16459 (N_16459,N_15646,N_15996);
nor U16460 (N_16460,N_15704,N_15866);
xnor U16461 (N_16461,N_15597,N_15535);
or U16462 (N_16462,N_15910,N_15918);
and U16463 (N_16463,N_15710,N_15921);
nand U16464 (N_16464,N_15546,N_15930);
xor U16465 (N_16465,N_15959,N_15848);
nand U16466 (N_16466,N_15999,N_15965);
xor U16467 (N_16467,N_15893,N_15739);
xor U16468 (N_16468,N_15838,N_15600);
nor U16469 (N_16469,N_15886,N_15733);
and U16470 (N_16470,N_15810,N_15545);
nor U16471 (N_16471,N_15738,N_15544);
nor U16472 (N_16472,N_15731,N_15801);
and U16473 (N_16473,N_15773,N_15649);
nand U16474 (N_16474,N_15807,N_15945);
nand U16475 (N_16475,N_15907,N_15916);
nor U16476 (N_16476,N_15654,N_15741);
or U16477 (N_16477,N_15766,N_15916);
nand U16478 (N_16478,N_15939,N_15738);
and U16479 (N_16479,N_15645,N_15887);
nor U16480 (N_16480,N_15660,N_15555);
or U16481 (N_16481,N_15572,N_15929);
nand U16482 (N_16482,N_15506,N_15718);
nand U16483 (N_16483,N_15918,N_15692);
and U16484 (N_16484,N_15956,N_15892);
or U16485 (N_16485,N_15971,N_15841);
and U16486 (N_16486,N_15889,N_15518);
xnor U16487 (N_16487,N_15566,N_15971);
nand U16488 (N_16488,N_15508,N_15511);
nor U16489 (N_16489,N_15992,N_15978);
or U16490 (N_16490,N_15825,N_15526);
or U16491 (N_16491,N_15780,N_15728);
and U16492 (N_16492,N_15663,N_15755);
nand U16493 (N_16493,N_15612,N_15972);
and U16494 (N_16494,N_15792,N_15656);
nand U16495 (N_16495,N_15888,N_15853);
xor U16496 (N_16496,N_15639,N_15500);
xor U16497 (N_16497,N_15588,N_15539);
or U16498 (N_16498,N_15767,N_15965);
xnor U16499 (N_16499,N_15808,N_15541);
xnor U16500 (N_16500,N_16435,N_16058);
nand U16501 (N_16501,N_16031,N_16196);
and U16502 (N_16502,N_16133,N_16256);
and U16503 (N_16503,N_16291,N_16010);
xor U16504 (N_16504,N_16056,N_16459);
or U16505 (N_16505,N_16287,N_16330);
nand U16506 (N_16506,N_16345,N_16228);
nand U16507 (N_16507,N_16407,N_16036);
and U16508 (N_16508,N_16447,N_16308);
nor U16509 (N_16509,N_16357,N_16394);
nor U16510 (N_16510,N_16293,N_16311);
xor U16511 (N_16511,N_16427,N_16367);
nor U16512 (N_16512,N_16085,N_16245);
nand U16513 (N_16513,N_16443,N_16192);
nand U16514 (N_16514,N_16377,N_16009);
nand U16515 (N_16515,N_16301,N_16038);
and U16516 (N_16516,N_16296,N_16168);
or U16517 (N_16517,N_16231,N_16257);
nor U16518 (N_16518,N_16103,N_16346);
nand U16519 (N_16519,N_16139,N_16398);
nand U16520 (N_16520,N_16260,N_16277);
nor U16521 (N_16521,N_16000,N_16079);
and U16522 (N_16522,N_16267,N_16481);
nor U16523 (N_16523,N_16077,N_16131);
and U16524 (N_16524,N_16210,N_16057);
xnor U16525 (N_16525,N_16014,N_16097);
nand U16526 (N_16526,N_16033,N_16483);
or U16527 (N_16527,N_16471,N_16195);
nor U16528 (N_16528,N_16408,N_16326);
and U16529 (N_16529,N_16400,N_16446);
or U16530 (N_16530,N_16290,N_16107);
nand U16531 (N_16531,N_16083,N_16404);
nor U16532 (N_16532,N_16122,N_16166);
xnor U16533 (N_16533,N_16233,N_16414);
xnor U16534 (N_16534,N_16453,N_16302);
xnor U16535 (N_16535,N_16485,N_16282);
nor U16536 (N_16536,N_16149,N_16387);
and U16537 (N_16537,N_16395,N_16055);
nor U16538 (N_16538,N_16188,N_16121);
xnor U16539 (N_16539,N_16300,N_16240);
nor U16540 (N_16540,N_16418,N_16163);
xor U16541 (N_16541,N_16436,N_16136);
and U16542 (N_16542,N_16223,N_16349);
and U16543 (N_16543,N_16468,N_16070);
xor U16544 (N_16544,N_16189,N_16424);
xor U16545 (N_16545,N_16348,N_16109);
and U16546 (N_16546,N_16433,N_16324);
or U16547 (N_16547,N_16042,N_16399);
nor U16548 (N_16548,N_16239,N_16305);
nand U16549 (N_16549,N_16323,N_16132);
or U16550 (N_16550,N_16489,N_16297);
or U16551 (N_16551,N_16299,N_16177);
nor U16552 (N_16552,N_16384,N_16266);
nand U16553 (N_16553,N_16087,N_16072);
nor U16554 (N_16554,N_16007,N_16281);
nand U16555 (N_16555,N_16355,N_16120);
nor U16556 (N_16556,N_16371,N_16047);
or U16557 (N_16557,N_16295,N_16315);
or U16558 (N_16558,N_16250,N_16434);
and U16559 (N_16559,N_16337,N_16099);
and U16560 (N_16560,N_16202,N_16059);
nand U16561 (N_16561,N_16096,N_16265);
xor U16562 (N_16562,N_16352,N_16432);
nand U16563 (N_16563,N_16458,N_16279);
xnor U16564 (N_16564,N_16159,N_16187);
nand U16565 (N_16565,N_16126,N_16116);
xnor U16566 (N_16566,N_16452,N_16440);
or U16567 (N_16567,N_16431,N_16444);
nand U16568 (N_16568,N_16439,N_16309);
xor U16569 (N_16569,N_16235,N_16154);
nand U16570 (N_16570,N_16358,N_16181);
nor U16571 (N_16571,N_16455,N_16191);
xnor U16572 (N_16572,N_16006,N_16381);
nand U16573 (N_16573,N_16422,N_16197);
or U16574 (N_16574,N_16494,N_16227);
nor U16575 (N_16575,N_16340,N_16173);
nor U16576 (N_16576,N_16331,N_16319);
nor U16577 (N_16577,N_16135,N_16125);
and U16578 (N_16578,N_16252,N_16024);
nand U16579 (N_16579,N_16198,N_16270);
xor U16580 (N_16580,N_16288,N_16425);
or U16581 (N_16581,N_16220,N_16183);
nor U16582 (N_16582,N_16093,N_16338);
and U16583 (N_16583,N_16492,N_16380);
nor U16584 (N_16584,N_16030,N_16463);
nand U16585 (N_16585,N_16247,N_16128);
nand U16586 (N_16586,N_16449,N_16470);
xnor U16587 (N_16587,N_16495,N_16152);
xnor U16588 (N_16588,N_16115,N_16019);
or U16589 (N_16589,N_16334,N_16268);
xnor U16590 (N_16590,N_16382,N_16480);
or U16591 (N_16591,N_16075,N_16118);
nand U16592 (N_16592,N_16236,N_16062);
or U16593 (N_16593,N_16376,N_16406);
nor U16594 (N_16594,N_16137,N_16130);
xor U16595 (N_16595,N_16065,N_16264);
or U16596 (N_16596,N_16336,N_16158);
or U16597 (N_16597,N_16071,N_16332);
xnor U16598 (N_16598,N_16061,N_16221);
nor U16599 (N_16599,N_16386,N_16318);
xor U16600 (N_16600,N_16428,N_16273);
nor U16601 (N_16601,N_16230,N_16150);
nand U16602 (N_16602,N_16388,N_16496);
and U16603 (N_16603,N_16328,N_16066);
or U16604 (N_16604,N_16214,N_16285);
nand U16605 (N_16605,N_16207,N_16243);
or U16606 (N_16606,N_16094,N_16232);
nor U16607 (N_16607,N_16478,N_16110);
or U16608 (N_16608,N_16205,N_16088);
nor U16609 (N_16609,N_16016,N_16020);
and U16610 (N_16610,N_16383,N_16410);
or U16611 (N_16611,N_16484,N_16401);
or U16612 (N_16612,N_16144,N_16178);
or U16613 (N_16613,N_16204,N_16460);
xor U16614 (N_16614,N_16419,N_16089);
and U16615 (N_16615,N_16465,N_16375);
or U16616 (N_16616,N_16353,N_16325);
or U16617 (N_16617,N_16054,N_16498);
or U16618 (N_16618,N_16262,N_16373);
nand U16619 (N_16619,N_16403,N_16335);
or U16620 (N_16620,N_16015,N_16317);
nor U16621 (N_16621,N_16450,N_16027);
and U16622 (N_16622,N_16185,N_16316);
and U16623 (N_16623,N_16184,N_16350);
or U16624 (N_16624,N_16362,N_16186);
nor U16625 (N_16625,N_16343,N_16063);
xor U16626 (N_16626,N_16167,N_16175);
or U16627 (N_16627,N_16162,N_16224);
or U16628 (N_16628,N_16461,N_16155);
nor U16629 (N_16629,N_16312,N_16298);
nor U16630 (N_16630,N_16080,N_16246);
nand U16631 (N_16631,N_16102,N_16095);
or U16632 (N_16632,N_16438,N_16147);
nor U16633 (N_16633,N_16341,N_16164);
nand U16634 (N_16634,N_16364,N_16124);
xor U16635 (N_16635,N_16229,N_16105);
or U16636 (N_16636,N_16005,N_16251);
and U16637 (N_16637,N_16322,N_16078);
and U16638 (N_16638,N_16176,N_16397);
xor U16639 (N_16639,N_16476,N_16451);
nor U16640 (N_16640,N_16028,N_16157);
xor U16641 (N_16641,N_16004,N_16156);
or U16642 (N_16642,N_16025,N_16477);
and U16643 (N_16643,N_16112,N_16307);
and U16644 (N_16644,N_16361,N_16194);
nor U16645 (N_16645,N_16011,N_16248);
nand U16646 (N_16646,N_16034,N_16049);
or U16647 (N_16647,N_16420,N_16421);
nor U16648 (N_16648,N_16051,N_16263);
or U16649 (N_16649,N_16253,N_16486);
or U16650 (N_16650,N_16012,N_16368);
or U16651 (N_16651,N_16342,N_16379);
or U16652 (N_16652,N_16234,N_16190);
and U16653 (N_16653,N_16212,N_16129);
nand U16654 (N_16654,N_16101,N_16351);
or U16655 (N_16655,N_16359,N_16469);
or U16656 (N_16656,N_16487,N_16490);
nand U16657 (N_16657,N_16148,N_16151);
nor U16658 (N_16658,N_16050,N_16032);
or U16659 (N_16659,N_16292,N_16499);
and U16660 (N_16660,N_16117,N_16286);
nand U16661 (N_16661,N_16275,N_16416);
and U16662 (N_16662,N_16200,N_16064);
and U16663 (N_16663,N_16437,N_16213);
xnor U16664 (N_16664,N_16145,N_16203);
nand U16665 (N_16665,N_16442,N_16225);
and U16666 (N_16666,N_16199,N_16320);
nand U16667 (N_16667,N_16052,N_16321);
or U16668 (N_16668,N_16206,N_16249);
nand U16669 (N_16669,N_16073,N_16216);
or U16670 (N_16670,N_16276,N_16374);
xnor U16671 (N_16671,N_16053,N_16430);
nor U16672 (N_16672,N_16497,N_16026);
or U16673 (N_16673,N_16278,N_16160);
or U16674 (N_16674,N_16048,N_16037);
and U16675 (N_16675,N_16372,N_16411);
and U16676 (N_16676,N_16113,N_16493);
xor U16677 (N_16677,N_16356,N_16022);
nor U16678 (N_16678,N_16363,N_16413);
xor U16679 (N_16679,N_16365,N_16218);
nor U16680 (N_16680,N_16366,N_16043);
xnor U16681 (N_16681,N_16426,N_16114);
xor U16682 (N_16682,N_16165,N_16304);
and U16683 (N_16683,N_16313,N_16171);
nor U16684 (N_16684,N_16391,N_16226);
nand U16685 (N_16685,N_16172,N_16044);
nor U16686 (N_16686,N_16074,N_16069);
nor U16687 (N_16687,N_16211,N_16271);
and U16688 (N_16688,N_16182,N_16002);
xnor U16689 (N_16689,N_16385,N_16423);
and U16690 (N_16690,N_16378,N_16098);
nand U16691 (N_16691,N_16215,N_16310);
xor U16692 (N_16692,N_16369,N_16390);
xnor U16693 (N_16693,N_16018,N_16179);
nand U16694 (N_16694,N_16314,N_16039);
nand U16695 (N_16695,N_16108,N_16474);
and U16696 (N_16696,N_16219,N_16209);
and U16697 (N_16697,N_16429,N_16217);
nand U16698 (N_16698,N_16146,N_16142);
nand U16699 (N_16699,N_16344,N_16396);
or U16700 (N_16700,N_16269,N_16003);
nand U16701 (N_16701,N_16180,N_16169);
or U16702 (N_16702,N_16412,N_16140);
and U16703 (N_16703,N_16141,N_16457);
xnor U16704 (N_16704,N_16242,N_16347);
nor U16705 (N_16705,N_16491,N_16161);
or U16706 (N_16706,N_16360,N_16001);
and U16707 (N_16707,N_16405,N_16303);
xor U16708 (N_16708,N_16479,N_16090);
and U16709 (N_16709,N_16448,N_16409);
or U16710 (N_16710,N_16254,N_16272);
or U16711 (N_16711,N_16258,N_16104);
xnor U16712 (N_16712,N_16327,N_16100);
nand U16713 (N_16713,N_16111,N_16441);
xor U16714 (N_16714,N_16475,N_16106);
nor U16715 (N_16715,N_16127,N_16280);
and U16716 (N_16716,N_16086,N_16329);
and U16717 (N_16717,N_16084,N_16415);
nor U16718 (N_16718,N_16464,N_16029);
nand U16719 (N_16719,N_16306,N_16046);
nor U16720 (N_16720,N_16060,N_16138);
nor U16721 (N_16721,N_16040,N_16402);
xor U16722 (N_16722,N_16255,N_16222);
nor U16723 (N_16723,N_16170,N_16208);
xnor U16724 (N_16724,N_16174,N_16244);
nand U16725 (N_16725,N_16370,N_16092);
and U16726 (N_16726,N_16333,N_16091);
and U16727 (N_16727,N_16294,N_16045);
nand U16728 (N_16728,N_16274,N_16017);
or U16729 (N_16729,N_16119,N_16467);
xnor U16730 (N_16730,N_16023,N_16389);
and U16731 (N_16731,N_16082,N_16041);
and U16732 (N_16732,N_16201,N_16076);
xnor U16733 (N_16733,N_16067,N_16456);
nor U16734 (N_16734,N_16134,N_16289);
nand U16735 (N_16735,N_16081,N_16143);
xor U16736 (N_16736,N_16393,N_16153);
nor U16737 (N_16737,N_16454,N_16259);
and U16738 (N_16738,N_16482,N_16472);
nand U16739 (N_16739,N_16354,N_16473);
and U16740 (N_16740,N_16193,N_16488);
xor U16741 (N_16741,N_16013,N_16445);
xnor U16742 (N_16742,N_16417,N_16466);
nand U16743 (N_16743,N_16241,N_16008);
nand U16744 (N_16744,N_16392,N_16261);
nand U16745 (N_16745,N_16283,N_16284);
xnor U16746 (N_16746,N_16237,N_16035);
nand U16747 (N_16747,N_16068,N_16462);
and U16748 (N_16748,N_16021,N_16238);
and U16749 (N_16749,N_16339,N_16123);
nor U16750 (N_16750,N_16178,N_16302);
and U16751 (N_16751,N_16374,N_16015);
and U16752 (N_16752,N_16424,N_16007);
nor U16753 (N_16753,N_16310,N_16299);
nand U16754 (N_16754,N_16192,N_16240);
and U16755 (N_16755,N_16194,N_16446);
nor U16756 (N_16756,N_16253,N_16009);
nand U16757 (N_16757,N_16488,N_16078);
or U16758 (N_16758,N_16090,N_16324);
or U16759 (N_16759,N_16022,N_16299);
nor U16760 (N_16760,N_16350,N_16366);
nor U16761 (N_16761,N_16440,N_16226);
or U16762 (N_16762,N_16361,N_16183);
nand U16763 (N_16763,N_16410,N_16180);
nand U16764 (N_16764,N_16488,N_16173);
or U16765 (N_16765,N_16198,N_16264);
xor U16766 (N_16766,N_16448,N_16070);
xor U16767 (N_16767,N_16068,N_16398);
and U16768 (N_16768,N_16219,N_16325);
nand U16769 (N_16769,N_16060,N_16086);
and U16770 (N_16770,N_16230,N_16250);
nand U16771 (N_16771,N_16095,N_16044);
or U16772 (N_16772,N_16022,N_16305);
nand U16773 (N_16773,N_16419,N_16049);
nor U16774 (N_16774,N_16175,N_16116);
and U16775 (N_16775,N_16066,N_16275);
xor U16776 (N_16776,N_16397,N_16374);
or U16777 (N_16777,N_16346,N_16192);
nand U16778 (N_16778,N_16110,N_16178);
nand U16779 (N_16779,N_16353,N_16251);
xor U16780 (N_16780,N_16171,N_16356);
or U16781 (N_16781,N_16265,N_16487);
xnor U16782 (N_16782,N_16491,N_16226);
nor U16783 (N_16783,N_16455,N_16007);
xnor U16784 (N_16784,N_16108,N_16110);
or U16785 (N_16785,N_16351,N_16315);
nand U16786 (N_16786,N_16465,N_16332);
or U16787 (N_16787,N_16106,N_16003);
xor U16788 (N_16788,N_16281,N_16098);
nand U16789 (N_16789,N_16326,N_16323);
and U16790 (N_16790,N_16085,N_16479);
xor U16791 (N_16791,N_16032,N_16454);
xnor U16792 (N_16792,N_16302,N_16494);
and U16793 (N_16793,N_16116,N_16419);
nand U16794 (N_16794,N_16243,N_16291);
or U16795 (N_16795,N_16396,N_16102);
and U16796 (N_16796,N_16158,N_16345);
and U16797 (N_16797,N_16491,N_16308);
nor U16798 (N_16798,N_16423,N_16014);
nor U16799 (N_16799,N_16084,N_16225);
or U16800 (N_16800,N_16281,N_16476);
and U16801 (N_16801,N_16038,N_16066);
xnor U16802 (N_16802,N_16326,N_16279);
or U16803 (N_16803,N_16406,N_16415);
or U16804 (N_16804,N_16400,N_16355);
nor U16805 (N_16805,N_16490,N_16084);
or U16806 (N_16806,N_16016,N_16491);
and U16807 (N_16807,N_16279,N_16421);
xnor U16808 (N_16808,N_16303,N_16453);
or U16809 (N_16809,N_16256,N_16190);
or U16810 (N_16810,N_16360,N_16072);
xnor U16811 (N_16811,N_16286,N_16070);
or U16812 (N_16812,N_16484,N_16462);
nor U16813 (N_16813,N_16135,N_16284);
and U16814 (N_16814,N_16058,N_16328);
and U16815 (N_16815,N_16312,N_16410);
nor U16816 (N_16816,N_16098,N_16174);
nor U16817 (N_16817,N_16136,N_16122);
nand U16818 (N_16818,N_16299,N_16484);
and U16819 (N_16819,N_16283,N_16495);
or U16820 (N_16820,N_16416,N_16248);
nand U16821 (N_16821,N_16238,N_16485);
or U16822 (N_16822,N_16351,N_16155);
or U16823 (N_16823,N_16347,N_16435);
nand U16824 (N_16824,N_16011,N_16227);
nand U16825 (N_16825,N_16113,N_16158);
or U16826 (N_16826,N_16058,N_16463);
xnor U16827 (N_16827,N_16332,N_16211);
xor U16828 (N_16828,N_16030,N_16070);
nor U16829 (N_16829,N_16051,N_16281);
and U16830 (N_16830,N_16105,N_16382);
xnor U16831 (N_16831,N_16386,N_16232);
nand U16832 (N_16832,N_16188,N_16276);
and U16833 (N_16833,N_16219,N_16467);
or U16834 (N_16834,N_16436,N_16162);
or U16835 (N_16835,N_16331,N_16435);
xnor U16836 (N_16836,N_16462,N_16466);
and U16837 (N_16837,N_16471,N_16149);
and U16838 (N_16838,N_16296,N_16181);
and U16839 (N_16839,N_16364,N_16407);
and U16840 (N_16840,N_16155,N_16202);
nor U16841 (N_16841,N_16174,N_16309);
or U16842 (N_16842,N_16179,N_16178);
and U16843 (N_16843,N_16330,N_16437);
nand U16844 (N_16844,N_16344,N_16357);
nor U16845 (N_16845,N_16258,N_16384);
and U16846 (N_16846,N_16086,N_16446);
xnor U16847 (N_16847,N_16160,N_16041);
nand U16848 (N_16848,N_16250,N_16291);
or U16849 (N_16849,N_16408,N_16228);
xor U16850 (N_16850,N_16400,N_16208);
nand U16851 (N_16851,N_16082,N_16391);
and U16852 (N_16852,N_16462,N_16167);
xor U16853 (N_16853,N_16124,N_16344);
xor U16854 (N_16854,N_16375,N_16155);
nor U16855 (N_16855,N_16420,N_16106);
nor U16856 (N_16856,N_16451,N_16006);
xor U16857 (N_16857,N_16264,N_16484);
nand U16858 (N_16858,N_16271,N_16060);
xnor U16859 (N_16859,N_16094,N_16296);
and U16860 (N_16860,N_16136,N_16191);
and U16861 (N_16861,N_16322,N_16296);
and U16862 (N_16862,N_16485,N_16407);
or U16863 (N_16863,N_16388,N_16144);
nand U16864 (N_16864,N_16050,N_16484);
nor U16865 (N_16865,N_16486,N_16369);
or U16866 (N_16866,N_16184,N_16029);
nor U16867 (N_16867,N_16314,N_16255);
nor U16868 (N_16868,N_16042,N_16141);
nand U16869 (N_16869,N_16230,N_16478);
nand U16870 (N_16870,N_16061,N_16404);
xor U16871 (N_16871,N_16112,N_16471);
nand U16872 (N_16872,N_16420,N_16210);
nor U16873 (N_16873,N_16381,N_16343);
and U16874 (N_16874,N_16457,N_16195);
nand U16875 (N_16875,N_16070,N_16494);
nor U16876 (N_16876,N_16039,N_16372);
or U16877 (N_16877,N_16187,N_16456);
and U16878 (N_16878,N_16370,N_16043);
and U16879 (N_16879,N_16390,N_16349);
nand U16880 (N_16880,N_16467,N_16109);
nand U16881 (N_16881,N_16057,N_16223);
nor U16882 (N_16882,N_16063,N_16311);
and U16883 (N_16883,N_16114,N_16267);
nand U16884 (N_16884,N_16013,N_16498);
and U16885 (N_16885,N_16318,N_16246);
nand U16886 (N_16886,N_16061,N_16421);
nand U16887 (N_16887,N_16177,N_16196);
xnor U16888 (N_16888,N_16079,N_16465);
xor U16889 (N_16889,N_16188,N_16438);
and U16890 (N_16890,N_16076,N_16372);
nand U16891 (N_16891,N_16330,N_16363);
nor U16892 (N_16892,N_16326,N_16292);
nor U16893 (N_16893,N_16410,N_16389);
or U16894 (N_16894,N_16318,N_16489);
nor U16895 (N_16895,N_16166,N_16471);
and U16896 (N_16896,N_16201,N_16064);
nor U16897 (N_16897,N_16406,N_16353);
nand U16898 (N_16898,N_16188,N_16263);
nor U16899 (N_16899,N_16080,N_16041);
and U16900 (N_16900,N_16173,N_16288);
and U16901 (N_16901,N_16117,N_16247);
nor U16902 (N_16902,N_16247,N_16047);
or U16903 (N_16903,N_16218,N_16135);
or U16904 (N_16904,N_16217,N_16440);
or U16905 (N_16905,N_16480,N_16159);
or U16906 (N_16906,N_16357,N_16052);
and U16907 (N_16907,N_16443,N_16366);
xor U16908 (N_16908,N_16199,N_16469);
or U16909 (N_16909,N_16200,N_16234);
or U16910 (N_16910,N_16315,N_16402);
xnor U16911 (N_16911,N_16390,N_16393);
or U16912 (N_16912,N_16345,N_16150);
and U16913 (N_16913,N_16413,N_16343);
xor U16914 (N_16914,N_16128,N_16005);
xor U16915 (N_16915,N_16049,N_16228);
xor U16916 (N_16916,N_16422,N_16048);
nand U16917 (N_16917,N_16128,N_16475);
nor U16918 (N_16918,N_16332,N_16206);
nor U16919 (N_16919,N_16297,N_16322);
or U16920 (N_16920,N_16428,N_16464);
and U16921 (N_16921,N_16122,N_16180);
nand U16922 (N_16922,N_16132,N_16015);
xnor U16923 (N_16923,N_16160,N_16326);
and U16924 (N_16924,N_16154,N_16254);
xnor U16925 (N_16925,N_16479,N_16477);
xnor U16926 (N_16926,N_16154,N_16439);
or U16927 (N_16927,N_16042,N_16402);
or U16928 (N_16928,N_16233,N_16249);
nand U16929 (N_16929,N_16228,N_16384);
nor U16930 (N_16930,N_16386,N_16275);
nand U16931 (N_16931,N_16199,N_16007);
nor U16932 (N_16932,N_16332,N_16425);
or U16933 (N_16933,N_16296,N_16101);
nand U16934 (N_16934,N_16132,N_16354);
nand U16935 (N_16935,N_16130,N_16185);
xnor U16936 (N_16936,N_16218,N_16276);
nand U16937 (N_16937,N_16217,N_16015);
nand U16938 (N_16938,N_16154,N_16445);
and U16939 (N_16939,N_16491,N_16333);
nor U16940 (N_16940,N_16018,N_16173);
nand U16941 (N_16941,N_16342,N_16408);
nand U16942 (N_16942,N_16182,N_16462);
xor U16943 (N_16943,N_16105,N_16288);
and U16944 (N_16944,N_16085,N_16281);
xnor U16945 (N_16945,N_16134,N_16152);
nand U16946 (N_16946,N_16438,N_16279);
and U16947 (N_16947,N_16141,N_16472);
and U16948 (N_16948,N_16446,N_16376);
and U16949 (N_16949,N_16033,N_16408);
nor U16950 (N_16950,N_16437,N_16342);
nor U16951 (N_16951,N_16299,N_16172);
nor U16952 (N_16952,N_16062,N_16023);
xor U16953 (N_16953,N_16389,N_16057);
nand U16954 (N_16954,N_16255,N_16443);
and U16955 (N_16955,N_16074,N_16099);
nor U16956 (N_16956,N_16022,N_16066);
nor U16957 (N_16957,N_16477,N_16176);
and U16958 (N_16958,N_16286,N_16035);
nor U16959 (N_16959,N_16124,N_16231);
nor U16960 (N_16960,N_16340,N_16449);
or U16961 (N_16961,N_16147,N_16196);
or U16962 (N_16962,N_16474,N_16291);
and U16963 (N_16963,N_16452,N_16470);
nand U16964 (N_16964,N_16034,N_16111);
nor U16965 (N_16965,N_16130,N_16021);
nand U16966 (N_16966,N_16012,N_16393);
and U16967 (N_16967,N_16020,N_16204);
and U16968 (N_16968,N_16466,N_16335);
and U16969 (N_16969,N_16059,N_16413);
or U16970 (N_16970,N_16287,N_16314);
xor U16971 (N_16971,N_16455,N_16470);
nand U16972 (N_16972,N_16322,N_16032);
and U16973 (N_16973,N_16258,N_16058);
nand U16974 (N_16974,N_16237,N_16001);
and U16975 (N_16975,N_16120,N_16182);
and U16976 (N_16976,N_16033,N_16414);
or U16977 (N_16977,N_16347,N_16102);
and U16978 (N_16978,N_16014,N_16407);
nand U16979 (N_16979,N_16233,N_16404);
nand U16980 (N_16980,N_16466,N_16213);
xnor U16981 (N_16981,N_16396,N_16357);
nor U16982 (N_16982,N_16453,N_16345);
and U16983 (N_16983,N_16461,N_16490);
nand U16984 (N_16984,N_16071,N_16154);
xor U16985 (N_16985,N_16131,N_16177);
nor U16986 (N_16986,N_16391,N_16071);
nor U16987 (N_16987,N_16006,N_16496);
and U16988 (N_16988,N_16125,N_16275);
xor U16989 (N_16989,N_16169,N_16081);
and U16990 (N_16990,N_16358,N_16188);
or U16991 (N_16991,N_16163,N_16381);
or U16992 (N_16992,N_16194,N_16132);
or U16993 (N_16993,N_16493,N_16196);
and U16994 (N_16994,N_16146,N_16198);
or U16995 (N_16995,N_16076,N_16100);
or U16996 (N_16996,N_16148,N_16296);
and U16997 (N_16997,N_16217,N_16034);
nand U16998 (N_16998,N_16473,N_16313);
and U16999 (N_16999,N_16447,N_16325);
xnor U17000 (N_17000,N_16802,N_16768);
and U17001 (N_17001,N_16586,N_16597);
nand U17002 (N_17002,N_16773,N_16736);
xnor U17003 (N_17003,N_16934,N_16713);
and U17004 (N_17004,N_16737,N_16551);
or U17005 (N_17005,N_16609,N_16649);
xnor U17006 (N_17006,N_16905,N_16995);
nor U17007 (N_17007,N_16519,N_16552);
or U17008 (N_17008,N_16941,N_16815);
or U17009 (N_17009,N_16879,N_16801);
and U17010 (N_17010,N_16796,N_16919);
nand U17011 (N_17011,N_16527,N_16953);
xnor U17012 (N_17012,N_16897,N_16760);
or U17013 (N_17013,N_16863,N_16892);
xor U17014 (N_17014,N_16672,N_16780);
nand U17015 (N_17015,N_16891,N_16817);
and U17016 (N_17016,N_16833,N_16744);
or U17017 (N_17017,N_16762,N_16547);
nor U17018 (N_17018,N_16683,N_16793);
nor U17019 (N_17019,N_16738,N_16671);
and U17020 (N_17020,N_16991,N_16948);
nand U17021 (N_17021,N_16625,N_16741);
xor U17022 (N_17022,N_16579,N_16602);
nand U17023 (N_17023,N_16935,N_16984);
nor U17024 (N_17024,N_16732,N_16701);
nor U17025 (N_17025,N_16613,N_16510);
or U17026 (N_17026,N_16533,N_16917);
xor U17027 (N_17027,N_16924,N_16593);
nor U17028 (N_17028,N_16629,N_16858);
nand U17029 (N_17029,N_16662,N_16652);
xor U17030 (N_17030,N_16960,N_16557);
nand U17031 (N_17031,N_16926,N_16781);
and U17032 (N_17032,N_16733,N_16657);
nand U17033 (N_17033,N_16877,N_16665);
or U17034 (N_17034,N_16767,N_16631);
xor U17035 (N_17035,N_16871,N_16987);
nand U17036 (N_17036,N_16803,N_16911);
xnor U17037 (N_17037,N_16968,N_16835);
or U17038 (N_17038,N_16813,N_16699);
and U17039 (N_17039,N_16635,N_16689);
or U17040 (N_17040,N_16655,N_16661);
and U17041 (N_17041,N_16711,N_16918);
nand U17042 (N_17042,N_16676,N_16507);
nand U17043 (N_17043,N_16511,N_16537);
xnor U17044 (N_17044,N_16962,N_16814);
or U17045 (N_17045,N_16618,N_16639);
nand U17046 (N_17046,N_16806,N_16616);
and U17047 (N_17047,N_16585,N_16873);
and U17048 (N_17048,N_16816,N_16834);
nand U17049 (N_17049,N_16577,N_16660);
and U17050 (N_17050,N_16681,N_16598);
xnor U17051 (N_17051,N_16502,N_16986);
nand U17052 (N_17052,N_16809,N_16846);
xor U17053 (N_17053,N_16868,N_16853);
xnor U17054 (N_17054,N_16989,N_16811);
and U17055 (N_17055,N_16500,N_16983);
nor U17056 (N_17056,N_16979,N_16964);
xnor U17057 (N_17057,N_16644,N_16560);
nor U17058 (N_17058,N_16828,N_16578);
and U17059 (N_17059,N_16969,N_16772);
nand U17060 (N_17060,N_16821,N_16893);
and U17061 (N_17061,N_16620,N_16993);
nor U17062 (N_17062,N_16854,N_16686);
nor U17063 (N_17063,N_16734,N_16615);
and U17064 (N_17064,N_16883,N_16679);
nand U17065 (N_17065,N_16977,N_16610);
or U17066 (N_17066,N_16930,N_16538);
nor U17067 (N_17067,N_16932,N_16722);
nand U17068 (N_17068,N_16912,N_16745);
xnor U17069 (N_17069,N_16571,N_16687);
nand U17070 (N_17070,N_16723,N_16955);
xnor U17071 (N_17071,N_16970,N_16855);
xor U17072 (N_17072,N_16888,N_16943);
xnor U17073 (N_17073,N_16563,N_16994);
or U17074 (N_17074,N_16789,N_16503);
nor U17075 (N_17075,N_16797,N_16668);
xnor U17076 (N_17076,N_16886,N_16604);
xnor U17077 (N_17077,N_16637,N_16517);
and U17078 (N_17078,N_16561,N_16724);
or U17079 (N_17079,N_16965,N_16531);
and U17080 (N_17080,N_16600,N_16501);
nor U17081 (N_17081,N_16641,N_16626);
and U17082 (N_17082,N_16716,N_16592);
and U17083 (N_17083,N_16509,N_16752);
and U17084 (N_17084,N_16812,N_16518);
and U17085 (N_17085,N_16851,N_16574);
nand U17086 (N_17086,N_16727,N_16743);
or U17087 (N_17087,N_16808,N_16534);
xor U17088 (N_17088,N_16849,N_16513);
and U17089 (N_17089,N_16847,N_16971);
nor U17090 (N_17090,N_16838,N_16922);
xnor U17091 (N_17091,N_16712,N_16669);
and U17092 (N_17092,N_16785,N_16691);
nand U17093 (N_17093,N_16558,N_16862);
xnor U17094 (N_17094,N_16601,N_16908);
nand U17095 (N_17095,N_16820,N_16728);
nand U17096 (N_17096,N_16875,N_16735);
nand U17097 (N_17097,N_16647,N_16636);
xor U17098 (N_17098,N_16810,N_16582);
and U17099 (N_17099,N_16522,N_16946);
nor U17100 (N_17100,N_16895,N_16766);
or U17101 (N_17101,N_16524,N_16915);
or U17102 (N_17102,N_16795,N_16581);
and U17103 (N_17103,N_16865,N_16778);
nand U17104 (N_17104,N_16978,N_16562);
nor U17105 (N_17105,N_16696,N_16857);
and U17106 (N_17106,N_16758,N_16836);
xor U17107 (N_17107,N_16718,N_16539);
nand U17108 (N_17108,N_16944,N_16914);
nor U17109 (N_17109,N_16949,N_16685);
nor U17110 (N_17110,N_16695,N_16881);
nand U17111 (N_17111,N_16638,N_16623);
xnor U17112 (N_17112,N_16938,N_16933);
nand U17113 (N_17113,N_16512,N_16748);
nand U17114 (N_17114,N_16514,N_16937);
nand U17115 (N_17115,N_16872,N_16966);
nand U17116 (N_17116,N_16929,N_16876);
xor U17117 (N_17117,N_16988,N_16974);
xnor U17118 (N_17118,N_16945,N_16628);
nand U17119 (N_17119,N_16645,N_16697);
or U17120 (N_17120,N_16996,N_16887);
nand U17121 (N_17121,N_16859,N_16684);
or U17122 (N_17122,N_16516,N_16632);
xnor U17123 (N_17123,N_16902,N_16869);
and U17124 (N_17124,N_16554,N_16643);
or U17125 (N_17125,N_16931,N_16750);
or U17126 (N_17126,N_16666,N_16791);
nor U17127 (N_17127,N_16587,N_16575);
and U17128 (N_17128,N_16536,N_16916);
and U17129 (N_17129,N_16899,N_16800);
xor U17130 (N_17130,N_16614,N_16698);
xnor U17131 (N_17131,N_16640,N_16927);
and U17132 (N_17132,N_16505,N_16565);
nor U17133 (N_17133,N_16621,N_16588);
nor U17134 (N_17134,N_16589,N_16622);
nor U17135 (N_17135,N_16976,N_16923);
nor U17136 (N_17136,N_16526,N_16757);
nand U17137 (N_17137,N_16650,N_16546);
nor U17138 (N_17138,N_16981,N_16990);
xor U17139 (N_17139,N_16825,N_16627);
or U17140 (N_17140,N_16920,N_16909);
nor U17141 (N_17141,N_16824,N_16827);
and U17142 (N_17142,N_16951,N_16939);
and U17143 (N_17143,N_16559,N_16680);
nand U17144 (N_17144,N_16771,N_16947);
nand U17145 (N_17145,N_16594,N_16704);
nor U17146 (N_17146,N_16700,N_16548);
xor U17147 (N_17147,N_16599,N_16651);
nand U17148 (N_17148,N_16832,N_16694);
or U17149 (N_17149,N_16769,N_16659);
nor U17150 (N_17150,N_16894,N_16982);
and U17151 (N_17151,N_16831,N_16532);
xnor U17152 (N_17152,N_16870,N_16515);
or U17153 (N_17153,N_16787,N_16528);
and U17154 (N_17154,N_16707,N_16573);
nor U17155 (N_17155,N_16761,N_16880);
nand U17156 (N_17156,N_16749,N_16710);
nor U17157 (N_17157,N_16682,N_16544);
nand U17158 (N_17158,N_16692,N_16867);
and U17159 (N_17159,N_16726,N_16742);
xnor U17160 (N_17160,N_16717,N_16670);
xor U17161 (N_17161,N_16545,N_16731);
and U17162 (N_17162,N_16550,N_16913);
or U17163 (N_17163,N_16608,N_16942);
and U17164 (N_17164,N_16753,N_16568);
and U17165 (N_17165,N_16779,N_16763);
nand U17166 (N_17166,N_16782,N_16611);
nor U17167 (N_17167,N_16709,N_16861);
nor U17168 (N_17168,N_16940,N_16885);
nand U17169 (N_17169,N_16720,N_16841);
nand U17170 (N_17170,N_16997,N_16619);
or U17171 (N_17171,N_16607,N_16950);
or U17172 (N_17172,N_16958,N_16952);
nor U17173 (N_17173,N_16542,N_16756);
nand U17174 (N_17174,N_16878,N_16755);
nor U17175 (N_17175,N_16826,N_16882);
nand U17176 (N_17176,N_16606,N_16936);
xnor U17177 (N_17177,N_16856,N_16819);
nand U17178 (N_17178,N_16850,N_16673);
xor U17179 (N_17179,N_16729,N_16799);
and U17180 (N_17180,N_16928,N_16792);
xnor U17181 (N_17181,N_16693,N_16754);
nor U17182 (N_17182,N_16896,N_16900);
and U17183 (N_17183,N_16907,N_16543);
xor U17184 (N_17184,N_16654,N_16529);
and U17185 (N_17185,N_16830,N_16992);
and U17186 (N_17186,N_16617,N_16764);
xnor U17187 (N_17187,N_16590,N_16569);
or U17188 (N_17188,N_16975,N_16525);
nor U17189 (N_17189,N_16540,N_16798);
nor U17190 (N_17190,N_16583,N_16746);
nor U17191 (N_17191,N_16852,N_16642);
nor U17192 (N_17192,N_16624,N_16864);
nand U17193 (N_17193,N_16566,N_16903);
or U17194 (N_17194,N_16702,N_16706);
or U17195 (N_17195,N_16549,N_16818);
xor U17196 (N_17196,N_16521,N_16790);
or U17197 (N_17197,N_16751,N_16570);
and U17198 (N_17198,N_16985,N_16506);
nand U17199 (N_17199,N_16591,N_16972);
and U17200 (N_17200,N_16898,N_16690);
or U17201 (N_17201,N_16656,N_16630);
or U17202 (N_17202,N_16954,N_16580);
nand U17203 (N_17203,N_16794,N_16667);
xnor U17204 (N_17204,N_16634,N_16555);
nand U17205 (N_17205,N_16788,N_16805);
nand U17206 (N_17206,N_16703,N_16963);
nand U17207 (N_17207,N_16504,N_16664);
nor U17208 (N_17208,N_16823,N_16739);
or U17209 (N_17209,N_16860,N_16845);
nand U17210 (N_17210,N_16775,N_16715);
and U17211 (N_17211,N_16956,N_16961);
nand U17212 (N_17212,N_16646,N_16901);
and U17213 (N_17213,N_16523,N_16829);
or U17214 (N_17214,N_16804,N_16910);
and U17215 (N_17215,N_16714,N_16648);
nand U17216 (N_17216,N_16999,N_16957);
xnor U17217 (N_17217,N_16747,N_16677);
and U17218 (N_17218,N_16612,N_16674);
xnor U17219 (N_17219,N_16837,N_16844);
or U17220 (N_17220,N_16904,N_16719);
and U17221 (N_17221,N_16807,N_16603);
nor U17222 (N_17222,N_16973,N_16784);
nor U17223 (N_17223,N_16842,N_16508);
xor U17224 (N_17224,N_16998,N_16783);
xnor U17225 (N_17225,N_16866,N_16889);
and U17226 (N_17226,N_16584,N_16556);
nor U17227 (N_17227,N_16576,N_16925);
nand U17228 (N_17228,N_16564,N_16520);
xor U17229 (N_17229,N_16553,N_16633);
or U17230 (N_17230,N_16759,N_16740);
nor U17231 (N_17231,N_16721,N_16874);
xnor U17232 (N_17232,N_16595,N_16663);
and U17233 (N_17233,N_16678,N_16884);
nand U17234 (N_17234,N_16906,N_16921);
xnor U17235 (N_17235,N_16596,N_16530);
or U17236 (N_17236,N_16839,N_16840);
and U17237 (N_17237,N_16980,N_16843);
and U17238 (N_17238,N_16730,N_16653);
and U17239 (N_17239,N_16675,N_16959);
xor U17240 (N_17240,N_16848,N_16725);
and U17241 (N_17241,N_16822,N_16774);
xor U17242 (N_17242,N_16535,N_16658);
and U17243 (N_17243,N_16776,N_16786);
and U17244 (N_17244,N_16765,N_16572);
or U17245 (N_17245,N_16890,N_16708);
nor U17246 (N_17246,N_16605,N_16688);
xor U17247 (N_17247,N_16567,N_16770);
or U17248 (N_17248,N_16777,N_16705);
xor U17249 (N_17249,N_16967,N_16541);
or U17250 (N_17250,N_16676,N_16904);
and U17251 (N_17251,N_16876,N_16730);
or U17252 (N_17252,N_16569,N_16932);
nand U17253 (N_17253,N_16774,N_16686);
xor U17254 (N_17254,N_16988,N_16939);
nand U17255 (N_17255,N_16734,N_16966);
nor U17256 (N_17256,N_16843,N_16656);
xnor U17257 (N_17257,N_16993,N_16510);
xnor U17258 (N_17258,N_16978,N_16560);
xnor U17259 (N_17259,N_16856,N_16632);
nor U17260 (N_17260,N_16829,N_16870);
and U17261 (N_17261,N_16965,N_16676);
xnor U17262 (N_17262,N_16954,N_16675);
or U17263 (N_17263,N_16851,N_16557);
nand U17264 (N_17264,N_16627,N_16802);
xnor U17265 (N_17265,N_16653,N_16795);
xor U17266 (N_17266,N_16957,N_16880);
xnor U17267 (N_17267,N_16864,N_16523);
nor U17268 (N_17268,N_16751,N_16933);
and U17269 (N_17269,N_16557,N_16544);
nor U17270 (N_17270,N_16790,N_16635);
nand U17271 (N_17271,N_16741,N_16690);
xnor U17272 (N_17272,N_16651,N_16565);
xnor U17273 (N_17273,N_16728,N_16865);
nor U17274 (N_17274,N_16848,N_16880);
xor U17275 (N_17275,N_16761,N_16535);
and U17276 (N_17276,N_16837,N_16761);
or U17277 (N_17277,N_16943,N_16641);
or U17278 (N_17278,N_16764,N_16872);
and U17279 (N_17279,N_16918,N_16670);
and U17280 (N_17280,N_16662,N_16534);
xnor U17281 (N_17281,N_16813,N_16745);
xnor U17282 (N_17282,N_16803,N_16550);
xnor U17283 (N_17283,N_16733,N_16770);
nor U17284 (N_17284,N_16872,N_16679);
xnor U17285 (N_17285,N_16538,N_16573);
xnor U17286 (N_17286,N_16900,N_16512);
and U17287 (N_17287,N_16630,N_16831);
xnor U17288 (N_17288,N_16875,N_16739);
nor U17289 (N_17289,N_16500,N_16536);
xor U17290 (N_17290,N_16831,N_16793);
nor U17291 (N_17291,N_16910,N_16756);
nand U17292 (N_17292,N_16580,N_16808);
nor U17293 (N_17293,N_16529,N_16698);
or U17294 (N_17294,N_16885,N_16841);
nor U17295 (N_17295,N_16698,N_16890);
and U17296 (N_17296,N_16856,N_16837);
nor U17297 (N_17297,N_16780,N_16582);
nand U17298 (N_17298,N_16731,N_16702);
and U17299 (N_17299,N_16811,N_16925);
xor U17300 (N_17300,N_16933,N_16793);
xnor U17301 (N_17301,N_16974,N_16863);
xnor U17302 (N_17302,N_16601,N_16678);
xor U17303 (N_17303,N_16810,N_16925);
nand U17304 (N_17304,N_16814,N_16792);
and U17305 (N_17305,N_16722,N_16760);
xnor U17306 (N_17306,N_16699,N_16791);
and U17307 (N_17307,N_16981,N_16960);
xnor U17308 (N_17308,N_16587,N_16747);
or U17309 (N_17309,N_16920,N_16933);
or U17310 (N_17310,N_16632,N_16604);
xnor U17311 (N_17311,N_16879,N_16627);
or U17312 (N_17312,N_16619,N_16739);
nand U17313 (N_17313,N_16684,N_16764);
or U17314 (N_17314,N_16876,N_16850);
nor U17315 (N_17315,N_16626,N_16542);
and U17316 (N_17316,N_16740,N_16777);
or U17317 (N_17317,N_16701,N_16643);
or U17318 (N_17318,N_16575,N_16577);
and U17319 (N_17319,N_16959,N_16935);
nand U17320 (N_17320,N_16714,N_16561);
and U17321 (N_17321,N_16568,N_16761);
or U17322 (N_17322,N_16838,N_16647);
xnor U17323 (N_17323,N_16745,N_16519);
and U17324 (N_17324,N_16613,N_16553);
nor U17325 (N_17325,N_16891,N_16585);
nand U17326 (N_17326,N_16632,N_16504);
nand U17327 (N_17327,N_16571,N_16851);
or U17328 (N_17328,N_16916,N_16534);
or U17329 (N_17329,N_16965,N_16827);
xor U17330 (N_17330,N_16822,N_16731);
nand U17331 (N_17331,N_16576,N_16795);
or U17332 (N_17332,N_16910,N_16560);
nand U17333 (N_17333,N_16532,N_16800);
and U17334 (N_17334,N_16550,N_16956);
nand U17335 (N_17335,N_16787,N_16930);
nand U17336 (N_17336,N_16689,N_16855);
nor U17337 (N_17337,N_16734,N_16720);
or U17338 (N_17338,N_16790,N_16982);
xor U17339 (N_17339,N_16578,N_16661);
or U17340 (N_17340,N_16660,N_16981);
or U17341 (N_17341,N_16561,N_16730);
nand U17342 (N_17342,N_16601,N_16576);
or U17343 (N_17343,N_16628,N_16934);
and U17344 (N_17344,N_16636,N_16615);
xor U17345 (N_17345,N_16688,N_16570);
xnor U17346 (N_17346,N_16762,N_16619);
xnor U17347 (N_17347,N_16905,N_16847);
or U17348 (N_17348,N_16947,N_16845);
nor U17349 (N_17349,N_16714,N_16629);
nand U17350 (N_17350,N_16865,N_16784);
or U17351 (N_17351,N_16556,N_16726);
xnor U17352 (N_17352,N_16876,N_16670);
nand U17353 (N_17353,N_16679,N_16924);
nor U17354 (N_17354,N_16665,N_16660);
xor U17355 (N_17355,N_16572,N_16745);
nor U17356 (N_17356,N_16707,N_16861);
nor U17357 (N_17357,N_16864,N_16804);
nand U17358 (N_17358,N_16575,N_16777);
nand U17359 (N_17359,N_16970,N_16911);
nor U17360 (N_17360,N_16625,N_16575);
nor U17361 (N_17361,N_16931,N_16909);
nor U17362 (N_17362,N_16531,N_16814);
or U17363 (N_17363,N_16679,N_16631);
or U17364 (N_17364,N_16897,N_16767);
and U17365 (N_17365,N_16980,N_16626);
nor U17366 (N_17366,N_16871,N_16571);
nand U17367 (N_17367,N_16934,N_16590);
or U17368 (N_17368,N_16744,N_16989);
nand U17369 (N_17369,N_16885,N_16631);
xor U17370 (N_17370,N_16629,N_16667);
nor U17371 (N_17371,N_16898,N_16856);
nand U17372 (N_17372,N_16995,N_16533);
nand U17373 (N_17373,N_16621,N_16672);
and U17374 (N_17374,N_16559,N_16562);
nand U17375 (N_17375,N_16571,N_16631);
nand U17376 (N_17376,N_16648,N_16694);
xnor U17377 (N_17377,N_16572,N_16893);
nand U17378 (N_17378,N_16550,N_16652);
nor U17379 (N_17379,N_16676,N_16738);
or U17380 (N_17380,N_16673,N_16556);
xnor U17381 (N_17381,N_16794,N_16853);
xor U17382 (N_17382,N_16543,N_16547);
and U17383 (N_17383,N_16774,N_16942);
nand U17384 (N_17384,N_16742,N_16672);
nand U17385 (N_17385,N_16800,N_16552);
or U17386 (N_17386,N_16645,N_16734);
and U17387 (N_17387,N_16752,N_16614);
nor U17388 (N_17388,N_16613,N_16572);
and U17389 (N_17389,N_16648,N_16565);
xor U17390 (N_17390,N_16867,N_16587);
or U17391 (N_17391,N_16594,N_16829);
and U17392 (N_17392,N_16510,N_16911);
xor U17393 (N_17393,N_16925,N_16557);
nand U17394 (N_17394,N_16982,N_16933);
nand U17395 (N_17395,N_16680,N_16542);
or U17396 (N_17396,N_16711,N_16589);
xor U17397 (N_17397,N_16748,N_16915);
and U17398 (N_17398,N_16715,N_16855);
nor U17399 (N_17399,N_16791,N_16761);
nor U17400 (N_17400,N_16939,N_16662);
xor U17401 (N_17401,N_16959,N_16558);
xor U17402 (N_17402,N_16879,N_16687);
nor U17403 (N_17403,N_16762,N_16671);
xor U17404 (N_17404,N_16536,N_16929);
xor U17405 (N_17405,N_16681,N_16995);
or U17406 (N_17406,N_16595,N_16950);
nor U17407 (N_17407,N_16898,N_16557);
and U17408 (N_17408,N_16911,N_16989);
xor U17409 (N_17409,N_16672,N_16518);
and U17410 (N_17410,N_16576,N_16989);
nand U17411 (N_17411,N_16721,N_16990);
nor U17412 (N_17412,N_16944,N_16718);
nand U17413 (N_17413,N_16789,N_16971);
nor U17414 (N_17414,N_16690,N_16725);
nor U17415 (N_17415,N_16593,N_16657);
xnor U17416 (N_17416,N_16835,N_16654);
nand U17417 (N_17417,N_16782,N_16762);
nor U17418 (N_17418,N_16682,N_16624);
nand U17419 (N_17419,N_16612,N_16874);
nor U17420 (N_17420,N_16527,N_16571);
nand U17421 (N_17421,N_16918,N_16890);
nand U17422 (N_17422,N_16714,N_16545);
and U17423 (N_17423,N_16528,N_16505);
nand U17424 (N_17424,N_16555,N_16671);
nor U17425 (N_17425,N_16785,N_16708);
nor U17426 (N_17426,N_16650,N_16573);
or U17427 (N_17427,N_16683,N_16819);
xor U17428 (N_17428,N_16907,N_16565);
nor U17429 (N_17429,N_16509,N_16982);
xor U17430 (N_17430,N_16839,N_16605);
nor U17431 (N_17431,N_16630,N_16538);
nand U17432 (N_17432,N_16633,N_16754);
nor U17433 (N_17433,N_16848,N_16713);
nor U17434 (N_17434,N_16990,N_16773);
nor U17435 (N_17435,N_16630,N_16861);
nor U17436 (N_17436,N_16562,N_16556);
xor U17437 (N_17437,N_16746,N_16570);
nor U17438 (N_17438,N_16787,N_16786);
xnor U17439 (N_17439,N_16696,N_16792);
and U17440 (N_17440,N_16981,N_16932);
nand U17441 (N_17441,N_16575,N_16584);
or U17442 (N_17442,N_16533,N_16845);
nor U17443 (N_17443,N_16580,N_16961);
and U17444 (N_17444,N_16835,N_16581);
nand U17445 (N_17445,N_16652,N_16791);
xnor U17446 (N_17446,N_16514,N_16986);
xor U17447 (N_17447,N_16704,N_16709);
nor U17448 (N_17448,N_16851,N_16918);
nand U17449 (N_17449,N_16697,N_16768);
xnor U17450 (N_17450,N_16895,N_16959);
and U17451 (N_17451,N_16596,N_16552);
xnor U17452 (N_17452,N_16825,N_16559);
or U17453 (N_17453,N_16792,N_16760);
nor U17454 (N_17454,N_16552,N_16850);
and U17455 (N_17455,N_16845,N_16892);
xor U17456 (N_17456,N_16859,N_16581);
and U17457 (N_17457,N_16841,N_16599);
nand U17458 (N_17458,N_16795,N_16703);
and U17459 (N_17459,N_16706,N_16678);
nand U17460 (N_17460,N_16596,N_16913);
xor U17461 (N_17461,N_16918,N_16995);
nor U17462 (N_17462,N_16980,N_16999);
nand U17463 (N_17463,N_16643,N_16577);
or U17464 (N_17464,N_16929,N_16550);
or U17465 (N_17465,N_16647,N_16909);
or U17466 (N_17466,N_16686,N_16548);
and U17467 (N_17467,N_16969,N_16884);
nor U17468 (N_17468,N_16980,N_16719);
nor U17469 (N_17469,N_16742,N_16612);
nor U17470 (N_17470,N_16960,N_16545);
nor U17471 (N_17471,N_16901,N_16859);
xor U17472 (N_17472,N_16834,N_16799);
or U17473 (N_17473,N_16889,N_16576);
nor U17474 (N_17474,N_16728,N_16831);
and U17475 (N_17475,N_16975,N_16832);
nand U17476 (N_17476,N_16978,N_16651);
and U17477 (N_17477,N_16982,N_16577);
and U17478 (N_17478,N_16862,N_16591);
nor U17479 (N_17479,N_16989,N_16556);
nand U17480 (N_17480,N_16924,N_16755);
xnor U17481 (N_17481,N_16768,N_16824);
nor U17482 (N_17482,N_16928,N_16891);
nor U17483 (N_17483,N_16610,N_16640);
and U17484 (N_17484,N_16652,N_16685);
and U17485 (N_17485,N_16992,N_16942);
or U17486 (N_17486,N_16557,N_16834);
or U17487 (N_17487,N_16744,N_16731);
xnor U17488 (N_17488,N_16623,N_16579);
or U17489 (N_17489,N_16966,N_16976);
nand U17490 (N_17490,N_16665,N_16571);
or U17491 (N_17491,N_16675,N_16781);
nand U17492 (N_17492,N_16650,N_16695);
nor U17493 (N_17493,N_16617,N_16634);
and U17494 (N_17494,N_16977,N_16549);
nor U17495 (N_17495,N_16740,N_16933);
xor U17496 (N_17496,N_16880,N_16531);
and U17497 (N_17497,N_16584,N_16895);
nor U17498 (N_17498,N_16652,N_16932);
nand U17499 (N_17499,N_16913,N_16929);
or U17500 (N_17500,N_17291,N_17188);
xnor U17501 (N_17501,N_17235,N_17178);
xnor U17502 (N_17502,N_17071,N_17465);
or U17503 (N_17503,N_17162,N_17443);
xnor U17504 (N_17504,N_17313,N_17428);
xnor U17505 (N_17505,N_17077,N_17266);
nor U17506 (N_17506,N_17308,N_17249);
nand U17507 (N_17507,N_17305,N_17419);
nand U17508 (N_17508,N_17418,N_17052);
xor U17509 (N_17509,N_17415,N_17068);
nor U17510 (N_17510,N_17348,N_17247);
nor U17511 (N_17511,N_17282,N_17218);
nand U17512 (N_17512,N_17391,N_17490);
nor U17513 (N_17513,N_17021,N_17283);
nand U17514 (N_17514,N_17211,N_17070);
and U17515 (N_17515,N_17216,N_17194);
and U17516 (N_17516,N_17227,N_17464);
xor U17517 (N_17517,N_17397,N_17110);
or U17518 (N_17518,N_17297,N_17217);
nand U17519 (N_17519,N_17050,N_17384);
nor U17520 (N_17520,N_17011,N_17019);
and U17521 (N_17521,N_17163,N_17461);
and U17522 (N_17522,N_17060,N_17112);
nand U17523 (N_17523,N_17375,N_17251);
nor U17524 (N_17524,N_17481,N_17335);
nor U17525 (N_17525,N_17134,N_17451);
xor U17526 (N_17526,N_17399,N_17136);
or U17527 (N_17527,N_17425,N_17377);
nor U17528 (N_17528,N_17458,N_17173);
nand U17529 (N_17529,N_17454,N_17103);
nor U17530 (N_17530,N_17484,N_17259);
nand U17531 (N_17531,N_17347,N_17031);
nor U17532 (N_17532,N_17044,N_17219);
nor U17533 (N_17533,N_17439,N_17195);
xnor U17534 (N_17534,N_17098,N_17299);
nand U17535 (N_17535,N_17378,N_17099);
xor U17536 (N_17536,N_17013,N_17318);
and U17537 (N_17537,N_17404,N_17483);
nor U17538 (N_17538,N_17426,N_17226);
nor U17539 (N_17539,N_17317,N_17223);
nand U17540 (N_17540,N_17156,N_17165);
or U17541 (N_17541,N_17485,N_17158);
and U17542 (N_17542,N_17088,N_17414);
and U17543 (N_17543,N_17369,N_17301);
or U17544 (N_17544,N_17328,N_17101);
xnor U17545 (N_17545,N_17316,N_17017);
nand U17546 (N_17546,N_17444,N_17148);
or U17547 (N_17547,N_17180,N_17124);
xnor U17548 (N_17548,N_17323,N_17385);
and U17549 (N_17549,N_17286,N_17248);
nand U17550 (N_17550,N_17344,N_17135);
nand U17551 (N_17551,N_17491,N_17038);
or U17552 (N_17552,N_17466,N_17224);
or U17553 (N_17553,N_17062,N_17125);
xnor U17554 (N_17554,N_17142,N_17267);
or U17555 (N_17555,N_17287,N_17117);
and U17556 (N_17556,N_17141,N_17241);
and U17557 (N_17557,N_17460,N_17438);
xor U17558 (N_17558,N_17132,N_17175);
and U17559 (N_17559,N_17482,N_17288);
and U17560 (N_17560,N_17421,N_17154);
and U17561 (N_17561,N_17076,N_17370);
nor U17562 (N_17562,N_17215,N_17326);
nor U17563 (N_17563,N_17036,N_17091);
and U17564 (N_17564,N_17006,N_17392);
nor U17565 (N_17565,N_17368,N_17321);
nand U17566 (N_17566,N_17295,N_17113);
nor U17567 (N_17567,N_17222,N_17394);
nand U17568 (N_17568,N_17354,N_17236);
xnor U17569 (N_17569,N_17203,N_17284);
xor U17570 (N_17570,N_17055,N_17208);
and U17571 (N_17571,N_17420,N_17300);
and U17572 (N_17572,N_17280,N_17355);
xor U17573 (N_17573,N_17073,N_17167);
nand U17574 (N_17574,N_17272,N_17447);
nor U17575 (N_17575,N_17151,N_17127);
nand U17576 (N_17576,N_17493,N_17107);
or U17577 (N_17577,N_17057,N_17015);
xnor U17578 (N_17578,N_17005,N_17089);
xnor U17579 (N_17579,N_17410,N_17213);
nor U17580 (N_17580,N_17345,N_17176);
nand U17581 (N_17581,N_17403,N_17097);
or U17582 (N_17582,N_17309,N_17054);
nand U17583 (N_17583,N_17078,N_17435);
xnor U17584 (N_17584,N_17452,N_17225);
nand U17585 (N_17585,N_17168,N_17357);
xor U17586 (N_17586,N_17431,N_17085);
xnor U17587 (N_17587,N_17152,N_17450);
xor U17588 (N_17588,N_17095,N_17153);
nor U17589 (N_17589,N_17333,N_17413);
and U17590 (N_17590,N_17310,N_17043);
xor U17591 (N_17591,N_17379,N_17014);
and U17592 (N_17592,N_17207,N_17277);
or U17593 (N_17593,N_17059,N_17094);
nand U17594 (N_17594,N_17489,N_17026);
nand U17595 (N_17595,N_17325,N_17197);
nand U17596 (N_17596,N_17353,N_17022);
or U17597 (N_17597,N_17463,N_17367);
or U17598 (N_17598,N_17164,N_17398);
xnor U17599 (N_17599,N_17486,N_17030);
or U17600 (N_17600,N_17147,N_17276);
or U17601 (N_17601,N_17433,N_17246);
or U17602 (N_17602,N_17114,N_17408);
nand U17603 (N_17603,N_17193,N_17032);
and U17604 (N_17604,N_17007,N_17477);
nor U17605 (N_17605,N_17037,N_17093);
xor U17606 (N_17606,N_17170,N_17279);
and U17607 (N_17607,N_17473,N_17363);
and U17608 (N_17608,N_17358,N_17232);
and U17609 (N_17609,N_17100,N_17417);
and U17610 (N_17610,N_17494,N_17339);
nand U17611 (N_17611,N_17229,N_17183);
nor U17612 (N_17612,N_17067,N_17002);
and U17613 (N_17613,N_17075,N_17411);
nand U17614 (N_17614,N_17233,N_17122);
nor U17615 (N_17615,N_17471,N_17065);
or U17616 (N_17616,N_17159,N_17315);
nand U17617 (N_17617,N_17273,N_17496);
and U17618 (N_17618,N_17220,N_17427);
or U17619 (N_17619,N_17221,N_17035);
or U17620 (N_17620,N_17041,N_17437);
xnor U17621 (N_17621,N_17319,N_17462);
and U17622 (N_17622,N_17184,N_17109);
and U17623 (N_17623,N_17327,N_17240);
or U17624 (N_17624,N_17388,N_17406);
or U17625 (N_17625,N_17239,N_17245);
and U17626 (N_17626,N_17145,N_17008);
or U17627 (N_17627,N_17064,N_17047);
xor U17628 (N_17628,N_17372,N_17268);
nand U17629 (N_17629,N_17293,N_17105);
nor U17630 (N_17630,N_17474,N_17260);
xnor U17631 (N_17631,N_17289,N_17080);
nor U17632 (N_17632,N_17459,N_17129);
nand U17633 (N_17633,N_17262,N_17479);
nor U17634 (N_17634,N_17412,N_17387);
xnor U17635 (N_17635,N_17177,N_17296);
nor U17636 (N_17636,N_17340,N_17228);
and U17637 (N_17637,N_17243,N_17028);
and U17638 (N_17638,N_17209,N_17432);
nor U17639 (N_17639,N_17204,N_17079);
nand U17640 (N_17640,N_17373,N_17343);
nor U17641 (N_17641,N_17441,N_17254);
nor U17642 (N_17642,N_17468,N_17256);
and U17643 (N_17643,N_17445,N_17090);
and U17644 (N_17644,N_17402,N_17448);
nor U17645 (N_17645,N_17131,N_17237);
nor U17646 (N_17646,N_17478,N_17128);
or U17647 (N_17647,N_17390,N_17029);
nor U17648 (N_17648,N_17096,N_17341);
nand U17649 (N_17649,N_17169,N_17407);
nand U17650 (N_17650,N_17270,N_17409);
nor U17651 (N_17651,N_17265,N_17382);
nand U17652 (N_17652,N_17039,N_17389);
nor U17653 (N_17653,N_17386,N_17275);
nor U17654 (N_17654,N_17307,N_17115);
xor U17655 (N_17655,N_17274,N_17049);
or U17656 (N_17656,N_17250,N_17012);
nand U17657 (N_17657,N_17422,N_17130);
or U17658 (N_17658,N_17139,N_17189);
nor U17659 (N_17659,N_17269,N_17230);
nor U17660 (N_17660,N_17116,N_17051);
nor U17661 (N_17661,N_17499,N_17498);
or U17662 (N_17662,N_17359,N_17087);
or U17663 (N_17663,N_17242,N_17074);
nand U17664 (N_17664,N_17118,N_17469);
nor U17665 (N_17665,N_17104,N_17205);
or U17666 (N_17666,N_17192,N_17133);
and U17667 (N_17667,N_17362,N_17042);
or U17668 (N_17668,N_17395,N_17281);
and U17669 (N_17669,N_17033,N_17476);
or U17670 (N_17670,N_17449,N_17058);
nor U17671 (N_17671,N_17186,N_17004);
nand U17672 (N_17672,N_17330,N_17119);
nor U17673 (N_17673,N_17081,N_17253);
and U17674 (N_17674,N_17423,N_17048);
or U17675 (N_17675,N_17252,N_17185);
or U17676 (N_17676,N_17056,N_17111);
or U17677 (N_17677,N_17371,N_17082);
or U17678 (N_17678,N_17336,N_17108);
nand U17679 (N_17679,N_17155,N_17264);
or U17680 (N_17680,N_17027,N_17383);
nor U17681 (N_17681,N_17334,N_17430);
nor U17682 (N_17682,N_17434,N_17034);
nor U17683 (N_17683,N_17200,N_17102);
and U17684 (N_17684,N_17338,N_17332);
and U17685 (N_17685,N_17214,N_17010);
xor U17686 (N_17686,N_17003,N_17455);
nor U17687 (N_17687,N_17312,N_17198);
nor U17688 (N_17688,N_17053,N_17187);
and U17689 (N_17689,N_17424,N_17171);
or U17690 (N_17690,N_17381,N_17126);
nand U17691 (N_17691,N_17066,N_17244);
nand U17692 (N_17692,N_17196,N_17446);
xnor U17693 (N_17693,N_17456,N_17016);
nand U17694 (N_17694,N_17201,N_17364);
xnor U17695 (N_17695,N_17255,N_17120);
or U17696 (N_17696,N_17149,N_17457);
and U17697 (N_17697,N_17488,N_17429);
nand U17698 (N_17698,N_17238,N_17023);
nand U17699 (N_17699,N_17063,N_17292);
xor U17700 (N_17700,N_17306,N_17150);
nand U17701 (N_17701,N_17140,N_17181);
nand U17702 (N_17702,N_17401,N_17024);
xnor U17703 (N_17703,N_17314,N_17174);
and U17704 (N_17704,N_17000,N_17361);
nand U17705 (N_17705,N_17487,N_17137);
nor U17706 (N_17706,N_17322,N_17160);
or U17707 (N_17707,N_17298,N_17261);
and U17708 (N_17708,N_17380,N_17138);
nor U17709 (N_17709,N_17234,N_17349);
xnor U17710 (N_17710,N_17442,N_17199);
nand U17711 (N_17711,N_17086,N_17092);
nor U17712 (N_17712,N_17475,N_17020);
nor U17713 (N_17713,N_17144,N_17084);
and U17714 (N_17714,N_17146,N_17258);
and U17715 (N_17715,N_17356,N_17072);
nand U17716 (N_17716,N_17166,N_17182);
and U17717 (N_17717,N_17157,N_17342);
and U17718 (N_17718,N_17495,N_17470);
and U17719 (N_17719,N_17271,N_17278);
and U17720 (N_17720,N_17350,N_17352);
or U17721 (N_17721,N_17001,N_17061);
nand U17722 (N_17722,N_17294,N_17436);
nor U17723 (N_17723,N_17400,N_17083);
or U17724 (N_17724,N_17143,N_17202);
xnor U17725 (N_17725,N_17106,N_17467);
and U17726 (N_17726,N_17123,N_17472);
and U17727 (N_17727,N_17257,N_17416);
or U17728 (N_17728,N_17351,N_17302);
nor U17729 (N_17729,N_17337,N_17161);
xnor U17730 (N_17730,N_17210,N_17303);
and U17731 (N_17731,N_17320,N_17190);
nand U17732 (N_17732,N_17329,N_17346);
and U17733 (N_17733,N_17374,N_17331);
nor U17734 (N_17734,N_17285,N_17045);
xnor U17735 (N_17735,N_17121,N_17365);
or U17736 (N_17736,N_17405,N_17393);
xor U17737 (N_17737,N_17009,N_17018);
nor U17738 (N_17738,N_17480,N_17311);
xnor U17739 (N_17739,N_17440,N_17366);
or U17740 (N_17740,N_17191,N_17396);
nand U17741 (N_17741,N_17497,N_17263);
nor U17742 (N_17742,N_17040,N_17492);
nand U17743 (N_17743,N_17069,N_17172);
nand U17744 (N_17744,N_17179,N_17453);
nand U17745 (N_17745,N_17290,N_17376);
nand U17746 (N_17746,N_17304,N_17046);
xnor U17747 (N_17747,N_17360,N_17212);
xor U17748 (N_17748,N_17324,N_17025);
nand U17749 (N_17749,N_17231,N_17206);
nand U17750 (N_17750,N_17257,N_17057);
xnor U17751 (N_17751,N_17046,N_17371);
and U17752 (N_17752,N_17381,N_17260);
xnor U17753 (N_17753,N_17013,N_17114);
nor U17754 (N_17754,N_17329,N_17158);
or U17755 (N_17755,N_17228,N_17412);
nand U17756 (N_17756,N_17038,N_17343);
or U17757 (N_17757,N_17193,N_17147);
or U17758 (N_17758,N_17266,N_17188);
and U17759 (N_17759,N_17272,N_17343);
xor U17760 (N_17760,N_17179,N_17363);
or U17761 (N_17761,N_17464,N_17129);
nor U17762 (N_17762,N_17276,N_17355);
or U17763 (N_17763,N_17007,N_17114);
nor U17764 (N_17764,N_17446,N_17418);
and U17765 (N_17765,N_17057,N_17029);
nand U17766 (N_17766,N_17051,N_17232);
xor U17767 (N_17767,N_17491,N_17076);
and U17768 (N_17768,N_17388,N_17342);
and U17769 (N_17769,N_17276,N_17027);
xnor U17770 (N_17770,N_17202,N_17231);
xnor U17771 (N_17771,N_17080,N_17206);
xnor U17772 (N_17772,N_17484,N_17258);
nor U17773 (N_17773,N_17378,N_17072);
nand U17774 (N_17774,N_17174,N_17293);
nand U17775 (N_17775,N_17409,N_17072);
or U17776 (N_17776,N_17446,N_17168);
nor U17777 (N_17777,N_17203,N_17015);
nand U17778 (N_17778,N_17121,N_17458);
nor U17779 (N_17779,N_17458,N_17339);
nand U17780 (N_17780,N_17182,N_17089);
or U17781 (N_17781,N_17428,N_17193);
xnor U17782 (N_17782,N_17300,N_17140);
and U17783 (N_17783,N_17348,N_17456);
nor U17784 (N_17784,N_17009,N_17123);
or U17785 (N_17785,N_17328,N_17118);
or U17786 (N_17786,N_17478,N_17387);
and U17787 (N_17787,N_17393,N_17383);
and U17788 (N_17788,N_17092,N_17365);
or U17789 (N_17789,N_17320,N_17040);
nor U17790 (N_17790,N_17429,N_17443);
xnor U17791 (N_17791,N_17275,N_17136);
nand U17792 (N_17792,N_17150,N_17462);
nor U17793 (N_17793,N_17112,N_17282);
and U17794 (N_17794,N_17391,N_17075);
and U17795 (N_17795,N_17258,N_17404);
nand U17796 (N_17796,N_17453,N_17483);
xor U17797 (N_17797,N_17371,N_17018);
xor U17798 (N_17798,N_17385,N_17416);
xnor U17799 (N_17799,N_17450,N_17131);
nor U17800 (N_17800,N_17403,N_17054);
nor U17801 (N_17801,N_17177,N_17485);
or U17802 (N_17802,N_17360,N_17259);
or U17803 (N_17803,N_17030,N_17073);
xor U17804 (N_17804,N_17293,N_17457);
and U17805 (N_17805,N_17265,N_17158);
xor U17806 (N_17806,N_17306,N_17434);
nand U17807 (N_17807,N_17353,N_17031);
and U17808 (N_17808,N_17418,N_17322);
or U17809 (N_17809,N_17110,N_17452);
and U17810 (N_17810,N_17427,N_17232);
and U17811 (N_17811,N_17175,N_17496);
or U17812 (N_17812,N_17161,N_17292);
or U17813 (N_17813,N_17253,N_17219);
or U17814 (N_17814,N_17207,N_17143);
nor U17815 (N_17815,N_17466,N_17102);
nand U17816 (N_17816,N_17127,N_17482);
and U17817 (N_17817,N_17152,N_17182);
nor U17818 (N_17818,N_17475,N_17013);
nor U17819 (N_17819,N_17080,N_17153);
or U17820 (N_17820,N_17141,N_17162);
nor U17821 (N_17821,N_17321,N_17457);
or U17822 (N_17822,N_17097,N_17094);
nand U17823 (N_17823,N_17497,N_17162);
nor U17824 (N_17824,N_17443,N_17126);
and U17825 (N_17825,N_17495,N_17322);
and U17826 (N_17826,N_17382,N_17326);
xor U17827 (N_17827,N_17299,N_17309);
xnor U17828 (N_17828,N_17372,N_17326);
or U17829 (N_17829,N_17220,N_17009);
nand U17830 (N_17830,N_17380,N_17409);
nand U17831 (N_17831,N_17181,N_17184);
xnor U17832 (N_17832,N_17284,N_17355);
nand U17833 (N_17833,N_17467,N_17498);
nor U17834 (N_17834,N_17015,N_17241);
or U17835 (N_17835,N_17415,N_17435);
and U17836 (N_17836,N_17331,N_17198);
or U17837 (N_17837,N_17461,N_17296);
and U17838 (N_17838,N_17188,N_17381);
and U17839 (N_17839,N_17120,N_17139);
nand U17840 (N_17840,N_17091,N_17217);
nand U17841 (N_17841,N_17209,N_17180);
nand U17842 (N_17842,N_17155,N_17391);
xnor U17843 (N_17843,N_17103,N_17254);
nand U17844 (N_17844,N_17491,N_17253);
or U17845 (N_17845,N_17401,N_17349);
or U17846 (N_17846,N_17308,N_17296);
or U17847 (N_17847,N_17182,N_17083);
xnor U17848 (N_17848,N_17247,N_17335);
nor U17849 (N_17849,N_17328,N_17395);
nand U17850 (N_17850,N_17206,N_17115);
xnor U17851 (N_17851,N_17277,N_17253);
nand U17852 (N_17852,N_17446,N_17074);
nor U17853 (N_17853,N_17183,N_17196);
or U17854 (N_17854,N_17026,N_17313);
and U17855 (N_17855,N_17263,N_17350);
nor U17856 (N_17856,N_17478,N_17017);
nand U17857 (N_17857,N_17106,N_17223);
and U17858 (N_17858,N_17457,N_17151);
nand U17859 (N_17859,N_17272,N_17015);
nand U17860 (N_17860,N_17227,N_17144);
or U17861 (N_17861,N_17450,N_17195);
nor U17862 (N_17862,N_17170,N_17314);
nor U17863 (N_17863,N_17203,N_17312);
xnor U17864 (N_17864,N_17223,N_17049);
nand U17865 (N_17865,N_17236,N_17267);
nor U17866 (N_17866,N_17242,N_17225);
or U17867 (N_17867,N_17053,N_17232);
or U17868 (N_17868,N_17429,N_17355);
nor U17869 (N_17869,N_17040,N_17139);
xor U17870 (N_17870,N_17419,N_17354);
and U17871 (N_17871,N_17297,N_17171);
or U17872 (N_17872,N_17434,N_17218);
and U17873 (N_17873,N_17275,N_17264);
xnor U17874 (N_17874,N_17280,N_17200);
xor U17875 (N_17875,N_17385,N_17428);
nor U17876 (N_17876,N_17109,N_17495);
and U17877 (N_17877,N_17026,N_17244);
nand U17878 (N_17878,N_17274,N_17369);
nor U17879 (N_17879,N_17399,N_17296);
nand U17880 (N_17880,N_17175,N_17084);
nand U17881 (N_17881,N_17218,N_17407);
nand U17882 (N_17882,N_17129,N_17394);
or U17883 (N_17883,N_17424,N_17034);
nor U17884 (N_17884,N_17035,N_17036);
or U17885 (N_17885,N_17409,N_17395);
nand U17886 (N_17886,N_17449,N_17425);
or U17887 (N_17887,N_17194,N_17234);
and U17888 (N_17888,N_17062,N_17271);
nor U17889 (N_17889,N_17364,N_17475);
xnor U17890 (N_17890,N_17484,N_17263);
and U17891 (N_17891,N_17201,N_17193);
and U17892 (N_17892,N_17224,N_17262);
nor U17893 (N_17893,N_17148,N_17296);
nand U17894 (N_17894,N_17384,N_17304);
or U17895 (N_17895,N_17304,N_17192);
and U17896 (N_17896,N_17442,N_17004);
and U17897 (N_17897,N_17191,N_17291);
nand U17898 (N_17898,N_17174,N_17289);
xor U17899 (N_17899,N_17107,N_17289);
nor U17900 (N_17900,N_17284,N_17167);
or U17901 (N_17901,N_17420,N_17167);
nand U17902 (N_17902,N_17167,N_17102);
or U17903 (N_17903,N_17176,N_17026);
or U17904 (N_17904,N_17257,N_17139);
nand U17905 (N_17905,N_17111,N_17133);
nor U17906 (N_17906,N_17047,N_17085);
and U17907 (N_17907,N_17252,N_17021);
nand U17908 (N_17908,N_17455,N_17489);
nor U17909 (N_17909,N_17268,N_17109);
or U17910 (N_17910,N_17248,N_17428);
and U17911 (N_17911,N_17257,N_17455);
nor U17912 (N_17912,N_17487,N_17109);
nor U17913 (N_17913,N_17331,N_17094);
and U17914 (N_17914,N_17396,N_17455);
nand U17915 (N_17915,N_17395,N_17465);
nor U17916 (N_17916,N_17447,N_17264);
nor U17917 (N_17917,N_17388,N_17394);
or U17918 (N_17918,N_17214,N_17477);
nor U17919 (N_17919,N_17431,N_17081);
and U17920 (N_17920,N_17189,N_17462);
and U17921 (N_17921,N_17442,N_17383);
nand U17922 (N_17922,N_17334,N_17342);
nand U17923 (N_17923,N_17195,N_17428);
nor U17924 (N_17924,N_17367,N_17356);
and U17925 (N_17925,N_17415,N_17126);
nand U17926 (N_17926,N_17385,N_17171);
and U17927 (N_17927,N_17399,N_17366);
or U17928 (N_17928,N_17281,N_17102);
nor U17929 (N_17929,N_17479,N_17103);
and U17930 (N_17930,N_17467,N_17233);
xor U17931 (N_17931,N_17492,N_17056);
nor U17932 (N_17932,N_17453,N_17383);
nand U17933 (N_17933,N_17029,N_17111);
or U17934 (N_17934,N_17393,N_17476);
and U17935 (N_17935,N_17340,N_17023);
nor U17936 (N_17936,N_17413,N_17340);
and U17937 (N_17937,N_17002,N_17489);
and U17938 (N_17938,N_17328,N_17013);
or U17939 (N_17939,N_17371,N_17107);
or U17940 (N_17940,N_17298,N_17135);
and U17941 (N_17941,N_17038,N_17031);
xnor U17942 (N_17942,N_17013,N_17011);
and U17943 (N_17943,N_17157,N_17386);
and U17944 (N_17944,N_17394,N_17254);
nand U17945 (N_17945,N_17431,N_17435);
and U17946 (N_17946,N_17302,N_17159);
nor U17947 (N_17947,N_17491,N_17232);
or U17948 (N_17948,N_17326,N_17455);
or U17949 (N_17949,N_17045,N_17036);
and U17950 (N_17950,N_17181,N_17172);
and U17951 (N_17951,N_17417,N_17283);
nor U17952 (N_17952,N_17017,N_17195);
and U17953 (N_17953,N_17212,N_17308);
nor U17954 (N_17954,N_17338,N_17005);
xor U17955 (N_17955,N_17072,N_17475);
xor U17956 (N_17956,N_17192,N_17315);
or U17957 (N_17957,N_17489,N_17289);
nor U17958 (N_17958,N_17056,N_17317);
and U17959 (N_17959,N_17471,N_17206);
and U17960 (N_17960,N_17393,N_17170);
and U17961 (N_17961,N_17008,N_17044);
nand U17962 (N_17962,N_17436,N_17103);
xor U17963 (N_17963,N_17400,N_17316);
nand U17964 (N_17964,N_17276,N_17298);
and U17965 (N_17965,N_17303,N_17398);
and U17966 (N_17966,N_17467,N_17110);
nand U17967 (N_17967,N_17001,N_17051);
nand U17968 (N_17968,N_17225,N_17477);
or U17969 (N_17969,N_17142,N_17416);
or U17970 (N_17970,N_17023,N_17121);
or U17971 (N_17971,N_17415,N_17104);
xnor U17972 (N_17972,N_17426,N_17216);
and U17973 (N_17973,N_17074,N_17171);
nand U17974 (N_17974,N_17378,N_17429);
nor U17975 (N_17975,N_17482,N_17194);
nand U17976 (N_17976,N_17436,N_17357);
and U17977 (N_17977,N_17115,N_17378);
xor U17978 (N_17978,N_17076,N_17268);
and U17979 (N_17979,N_17245,N_17123);
nor U17980 (N_17980,N_17311,N_17108);
nand U17981 (N_17981,N_17342,N_17497);
nand U17982 (N_17982,N_17158,N_17422);
and U17983 (N_17983,N_17459,N_17266);
xnor U17984 (N_17984,N_17168,N_17360);
or U17985 (N_17985,N_17190,N_17464);
xor U17986 (N_17986,N_17421,N_17035);
or U17987 (N_17987,N_17109,N_17031);
or U17988 (N_17988,N_17434,N_17437);
xor U17989 (N_17989,N_17399,N_17287);
and U17990 (N_17990,N_17289,N_17095);
or U17991 (N_17991,N_17413,N_17149);
and U17992 (N_17992,N_17298,N_17034);
or U17993 (N_17993,N_17408,N_17279);
xor U17994 (N_17994,N_17275,N_17189);
and U17995 (N_17995,N_17238,N_17235);
nor U17996 (N_17996,N_17394,N_17244);
xnor U17997 (N_17997,N_17128,N_17240);
and U17998 (N_17998,N_17154,N_17007);
nor U17999 (N_17999,N_17163,N_17035);
and U18000 (N_18000,N_17772,N_17813);
nand U18001 (N_18001,N_17684,N_17636);
nand U18002 (N_18002,N_17640,N_17539);
nand U18003 (N_18003,N_17719,N_17723);
or U18004 (N_18004,N_17818,N_17965);
nor U18005 (N_18005,N_17710,N_17972);
nor U18006 (N_18006,N_17987,N_17588);
and U18007 (N_18007,N_17552,N_17509);
nor U18008 (N_18008,N_17675,N_17532);
or U18009 (N_18009,N_17561,N_17897);
nor U18010 (N_18010,N_17597,N_17716);
xor U18011 (N_18011,N_17760,N_17769);
xor U18012 (N_18012,N_17942,N_17519);
or U18013 (N_18013,N_17696,N_17872);
or U18014 (N_18014,N_17649,N_17614);
nor U18015 (N_18015,N_17590,N_17858);
nor U18016 (N_18016,N_17547,N_17889);
xor U18017 (N_18017,N_17944,N_17919);
nand U18018 (N_18018,N_17725,N_17850);
and U18019 (N_18019,N_17827,N_17974);
xor U18020 (N_18020,N_17817,N_17903);
or U18021 (N_18021,N_17578,N_17888);
xnor U18022 (N_18022,N_17984,N_17671);
xor U18023 (N_18023,N_17514,N_17855);
nor U18024 (N_18024,N_17607,N_17749);
nand U18025 (N_18025,N_17816,N_17791);
nor U18026 (N_18026,N_17873,N_17574);
nor U18027 (N_18027,N_17924,N_17704);
or U18028 (N_18028,N_17608,N_17633);
and U18029 (N_18029,N_17580,N_17811);
nand U18030 (N_18030,N_17925,N_17737);
or U18031 (N_18031,N_17799,N_17567);
nand U18032 (N_18032,N_17798,N_17999);
xnor U18033 (N_18033,N_17551,N_17908);
xnor U18034 (N_18034,N_17976,N_17709);
nand U18035 (N_18035,N_17927,N_17862);
nor U18036 (N_18036,N_17535,N_17893);
nand U18037 (N_18037,N_17836,N_17576);
nor U18038 (N_18038,N_17996,N_17500);
xor U18039 (N_18039,N_17910,N_17928);
or U18040 (N_18040,N_17786,N_17650);
xor U18041 (N_18041,N_17644,N_17613);
xnor U18042 (N_18042,N_17515,N_17602);
xnor U18043 (N_18043,N_17831,N_17544);
nor U18044 (N_18044,N_17657,N_17624);
and U18045 (N_18045,N_17529,N_17881);
nand U18046 (N_18046,N_17524,N_17978);
nor U18047 (N_18047,N_17992,N_17525);
nand U18048 (N_18048,N_17705,N_17842);
or U18049 (N_18049,N_17792,N_17592);
and U18050 (N_18050,N_17993,N_17587);
or U18051 (N_18051,N_17979,N_17689);
nand U18052 (N_18052,N_17936,N_17755);
or U18053 (N_18053,N_17700,N_17933);
and U18054 (N_18054,N_17963,N_17609);
nor U18055 (N_18055,N_17665,N_17546);
nand U18056 (N_18056,N_17534,N_17840);
and U18057 (N_18057,N_17711,N_17727);
nand U18058 (N_18058,N_17618,N_17807);
or U18059 (N_18059,N_17822,N_17651);
nor U18060 (N_18060,N_17680,N_17914);
or U18061 (N_18061,N_17594,N_17566);
and U18062 (N_18062,N_17983,N_17788);
or U18063 (N_18063,N_17681,N_17643);
xor U18064 (N_18064,N_17774,N_17756);
and U18065 (N_18065,N_17685,N_17593);
xnor U18066 (N_18066,N_17859,N_17692);
nor U18067 (N_18067,N_17701,N_17517);
nor U18068 (N_18068,N_17646,N_17948);
nor U18069 (N_18069,N_17967,N_17635);
or U18070 (N_18070,N_17875,N_17991);
and U18071 (N_18071,N_17629,N_17596);
nor U18072 (N_18072,N_17631,N_17707);
or U18073 (N_18073,N_17516,N_17664);
or U18074 (N_18074,N_17935,N_17776);
xor U18075 (N_18075,N_17502,N_17853);
or U18076 (N_18076,N_17528,N_17703);
and U18077 (N_18077,N_17956,N_17748);
or U18078 (N_18078,N_17896,N_17726);
and U18079 (N_18079,N_17601,N_17898);
nor U18080 (N_18080,N_17829,N_17950);
or U18081 (N_18081,N_17615,N_17848);
xor U18082 (N_18082,N_17878,N_17915);
or U18083 (N_18083,N_17804,N_17724);
and U18084 (N_18084,N_17513,N_17584);
nand U18085 (N_18085,N_17797,N_17966);
nor U18086 (N_18086,N_17874,N_17958);
and U18087 (N_18087,N_17672,N_17708);
nor U18088 (N_18088,N_17720,N_17523);
nand U18089 (N_18089,N_17834,N_17885);
and U18090 (N_18090,N_17638,N_17503);
and U18091 (N_18091,N_17789,N_17600);
xor U18092 (N_18092,N_17860,N_17639);
nor U18093 (N_18093,N_17536,N_17731);
nor U18094 (N_18094,N_17803,N_17621);
nand U18095 (N_18095,N_17746,N_17530);
nor U18096 (N_18096,N_17905,N_17663);
nor U18097 (N_18097,N_17877,N_17954);
xor U18098 (N_18098,N_17728,N_17501);
xnor U18099 (N_18099,N_17538,N_17922);
or U18100 (N_18100,N_17911,N_17619);
and U18101 (N_18101,N_17995,N_17603);
or U18102 (N_18102,N_17931,N_17863);
xnor U18103 (N_18103,N_17790,N_17985);
xor U18104 (N_18104,N_17895,N_17989);
xnor U18105 (N_18105,N_17913,N_17870);
nand U18106 (N_18106,N_17674,N_17645);
nand U18107 (N_18107,N_17962,N_17718);
nor U18108 (N_18108,N_17879,N_17548);
nor U18109 (N_18109,N_17808,N_17990);
xnor U18110 (N_18110,N_17821,N_17861);
nor U18111 (N_18111,N_17982,N_17697);
and U18112 (N_18112,N_17997,N_17845);
and U18113 (N_18113,N_17557,N_17955);
or U18114 (N_18114,N_17653,N_17570);
xnor U18115 (N_18115,N_17864,N_17655);
or U18116 (N_18116,N_17951,N_17775);
nor U18117 (N_18117,N_17814,N_17785);
and U18118 (N_18118,N_17658,N_17626);
or U18119 (N_18119,N_17761,N_17959);
or U18120 (N_18120,N_17986,N_17980);
xor U18121 (N_18121,N_17768,N_17975);
or U18122 (N_18122,N_17691,N_17752);
and U18123 (N_18123,N_17952,N_17662);
nand U18124 (N_18124,N_17867,N_17506);
nand U18125 (N_18125,N_17637,N_17510);
xnor U18126 (N_18126,N_17642,N_17838);
nand U18127 (N_18127,N_17964,N_17577);
nor U18128 (N_18128,N_17932,N_17605);
nor U18129 (N_18129,N_17627,N_17949);
nand U18130 (N_18130,N_17902,N_17533);
xnor U18131 (N_18131,N_17656,N_17698);
nand U18132 (N_18132,N_17632,N_17504);
or U18133 (N_18133,N_17679,N_17564);
xnor U18134 (N_18134,N_17521,N_17736);
nand U18135 (N_18135,N_17743,N_17682);
or U18136 (N_18136,N_17880,N_17540);
or U18137 (N_18137,N_17738,N_17851);
and U18138 (N_18138,N_17695,N_17690);
nand U18139 (N_18139,N_17599,N_17634);
xnor U18140 (N_18140,N_17505,N_17545);
nor U18141 (N_18141,N_17666,N_17777);
xor U18142 (N_18142,N_17941,N_17563);
and U18143 (N_18143,N_17543,N_17939);
and U18144 (N_18144,N_17825,N_17699);
nand U18145 (N_18145,N_17654,N_17556);
nand U18146 (N_18146,N_17953,N_17869);
xor U18147 (N_18147,N_17843,N_17583);
nand U18148 (N_18148,N_17542,N_17960);
xor U18149 (N_18149,N_17733,N_17886);
nor U18150 (N_18150,N_17766,N_17926);
xor U18151 (N_18151,N_17806,N_17961);
xnor U18152 (N_18152,N_17751,N_17883);
and U18153 (N_18153,N_17907,N_17735);
xor U18154 (N_18154,N_17899,N_17706);
or U18155 (N_18155,N_17809,N_17668);
nand U18156 (N_18156,N_17591,N_17630);
xor U18157 (N_18157,N_17713,N_17764);
nor U18158 (N_18158,N_17661,N_17930);
nor U18159 (N_18159,N_17659,N_17890);
and U18160 (N_18160,N_17652,N_17616);
nor U18161 (N_18161,N_17667,N_17508);
or U18162 (N_18162,N_17957,N_17796);
nor U18163 (N_18163,N_17669,N_17841);
and U18164 (N_18164,N_17744,N_17891);
and U18165 (N_18165,N_17921,N_17969);
xor U18166 (N_18166,N_17839,N_17904);
or U18167 (N_18167,N_17541,N_17917);
or U18168 (N_18168,N_17740,N_17887);
nor U18169 (N_18169,N_17520,N_17712);
and U18170 (N_18170,N_17894,N_17522);
nand U18171 (N_18171,N_17779,N_17968);
nor U18172 (N_18172,N_17604,N_17832);
nor U18173 (N_18173,N_17598,N_17846);
nand U18174 (N_18174,N_17625,N_17800);
nor U18175 (N_18175,N_17729,N_17526);
and U18176 (N_18176,N_17623,N_17824);
or U18177 (N_18177,N_17611,N_17909);
nor U18178 (N_18178,N_17783,N_17571);
or U18179 (N_18179,N_17871,N_17586);
or U18180 (N_18180,N_17550,N_17901);
or U18181 (N_18181,N_17741,N_17730);
or U18182 (N_18182,N_17765,N_17866);
xnor U18183 (N_18183,N_17812,N_17763);
and U18184 (N_18184,N_17820,N_17773);
xor U18185 (N_18185,N_17687,N_17676);
nand U18186 (N_18186,N_17802,N_17660);
nor U18187 (N_18187,N_17884,N_17946);
and U18188 (N_18188,N_17531,N_17753);
xnor U18189 (N_18189,N_17518,N_17854);
or U18190 (N_18190,N_17945,N_17787);
nor U18191 (N_18191,N_17606,N_17826);
xnor U18192 (N_18192,N_17579,N_17929);
nor U18193 (N_18193,N_17673,N_17833);
or U18194 (N_18194,N_17549,N_17981);
nor U18195 (N_18195,N_17757,N_17569);
and U18196 (N_18196,N_17694,N_17648);
or U18197 (N_18197,N_17555,N_17937);
nand U18198 (N_18198,N_17849,N_17617);
nand U18199 (N_18199,N_17781,N_17670);
nor U18200 (N_18200,N_17947,N_17784);
nand U18201 (N_18201,N_17585,N_17573);
and U18202 (N_18202,N_17582,N_17553);
or U18203 (N_18203,N_17830,N_17868);
or U18204 (N_18204,N_17865,N_17844);
and U18205 (N_18205,N_17977,N_17537);
or U18206 (N_18206,N_17810,N_17900);
or U18207 (N_18207,N_17562,N_17923);
xnor U18208 (N_18208,N_17793,N_17620);
nor U18209 (N_18209,N_17837,N_17794);
nand U18210 (N_18210,N_17823,N_17767);
or U18211 (N_18211,N_17938,N_17916);
and U18212 (N_18212,N_17759,N_17778);
or U18213 (N_18213,N_17507,N_17847);
and U18214 (N_18214,N_17702,N_17819);
or U18215 (N_18215,N_17686,N_17714);
nand U18216 (N_18216,N_17988,N_17565);
xor U18217 (N_18217,N_17994,N_17581);
or U18218 (N_18218,N_17750,N_17717);
nand U18219 (N_18219,N_17912,N_17747);
xnor U18220 (N_18220,N_17693,N_17512);
nand U18221 (N_18221,N_17721,N_17876);
nor U18222 (N_18222,N_17882,N_17677);
nand U18223 (N_18223,N_17575,N_17568);
xnor U18224 (N_18224,N_17795,N_17828);
xnor U18225 (N_18225,N_17732,N_17641);
xnor U18226 (N_18226,N_17754,N_17595);
nand U18227 (N_18227,N_17805,N_17801);
nand U18228 (N_18228,N_17688,N_17815);
or U18229 (N_18229,N_17970,N_17856);
nor U18230 (N_18230,N_17683,N_17722);
and U18231 (N_18231,N_17742,N_17572);
nand U18232 (N_18232,N_17612,N_17857);
or U18233 (N_18233,N_17558,N_17762);
nor U18234 (N_18234,N_17647,N_17560);
nor U18235 (N_18235,N_17998,N_17734);
or U18236 (N_18236,N_17906,N_17770);
nor U18237 (N_18237,N_17511,N_17835);
or U18238 (N_18238,N_17918,N_17758);
nand U18239 (N_18239,N_17715,N_17920);
and U18240 (N_18240,N_17852,N_17973);
xnor U18241 (N_18241,N_17892,N_17589);
or U18242 (N_18242,N_17771,N_17527);
nor U18243 (N_18243,N_17782,N_17610);
and U18244 (N_18244,N_17628,N_17943);
or U18245 (N_18245,N_17739,N_17780);
nor U18246 (N_18246,N_17971,N_17554);
xnor U18247 (N_18247,N_17940,N_17622);
and U18248 (N_18248,N_17559,N_17934);
and U18249 (N_18249,N_17678,N_17745);
xnor U18250 (N_18250,N_17534,N_17513);
nor U18251 (N_18251,N_17786,N_17617);
xor U18252 (N_18252,N_17821,N_17779);
nand U18253 (N_18253,N_17671,N_17741);
and U18254 (N_18254,N_17654,N_17926);
and U18255 (N_18255,N_17723,N_17672);
or U18256 (N_18256,N_17595,N_17839);
nand U18257 (N_18257,N_17746,N_17889);
and U18258 (N_18258,N_17880,N_17854);
and U18259 (N_18259,N_17612,N_17775);
and U18260 (N_18260,N_17759,N_17890);
xnor U18261 (N_18261,N_17807,N_17792);
xor U18262 (N_18262,N_17842,N_17530);
xnor U18263 (N_18263,N_17505,N_17702);
xor U18264 (N_18264,N_17578,N_17740);
xnor U18265 (N_18265,N_17774,N_17933);
xor U18266 (N_18266,N_17547,N_17852);
nand U18267 (N_18267,N_17871,N_17875);
and U18268 (N_18268,N_17888,N_17625);
xor U18269 (N_18269,N_17697,N_17979);
xnor U18270 (N_18270,N_17609,N_17702);
nand U18271 (N_18271,N_17504,N_17680);
and U18272 (N_18272,N_17778,N_17943);
nor U18273 (N_18273,N_17943,N_17702);
xnor U18274 (N_18274,N_17789,N_17708);
xnor U18275 (N_18275,N_17693,N_17528);
and U18276 (N_18276,N_17914,N_17954);
and U18277 (N_18277,N_17724,N_17979);
nand U18278 (N_18278,N_17782,N_17586);
nor U18279 (N_18279,N_17820,N_17513);
xnor U18280 (N_18280,N_17802,N_17750);
and U18281 (N_18281,N_17862,N_17859);
nand U18282 (N_18282,N_17845,N_17930);
nor U18283 (N_18283,N_17853,N_17963);
and U18284 (N_18284,N_17642,N_17679);
xnor U18285 (N_18285,N_17981,N_17847);
or U18286 (N_18286,N_17683,N_17608);
nor U18287 (N_18287,N_17821,N_17938);
nand U18288 (N_18288,N_17812,N_17621);
or U18289 (N_18289,N_17982,N_17640);
or U18290 (N_18290,N_17952,N_17532);
nand U18291 (N_18291,N_17755,N_17821);
and U18292 (N_18292,N_17831,N_17906);
xnor U18293 (N_18293,N_17528,N_17913);
nor U18294 (N_18294,N_17798,N_17716);
nand U18295 (N_18295,N_17544,N_17536);
xnor U18296 (N_18296,N_17773,N_17860);
xor U18297 (N_18297,N_17882,N_17594);
and U18298 (N_18298,N_17634,N_17594);
or U18299 (N_18299,N_17634,N_17877);
and U18300 (N_18300,N_17624,N_17836);
nand U18301 (N_18301,N_17905,N_17936);
or U18302 (N_18302,N_17554,N_17676);
or U18303 (N_18303,N_17863,N_17576);
nand U18304 (N_18304,N_17791,N_17649);
xnor U18305 (N_18305,N_17703,N_17689);
nand U18306 (N_18306,N_17922,N_17883);
and U18307 (N_18307,N_17894,N_17768);
nor U18308 (N_18308,N_17735,N_17896);
xor U18309 (N_18309,N_17643,N_17601);
nand U18310 (N_18310,N_17865,N_17640);
nand U18311 (N_18311,N_17739,N_17825);
xnor U18312 (N_18312,N_17758,N_17644);
xor U18313 (N_18313,N_17620,N_17796);
or U18314 (N_18314,N_17781,N_17535);
or U18315 (N_18315,N_17694,N_17900);
or U18316 (N_18316,N_17793,N_17940);
xor U18317 (N_18317,N_17944,N_17543);
nor U18318 (N_18318,N_17909,N_17793);
nor U18319 (N_18319,N_17559,N_17702);
nor U18320 (N_18320,N_17970,N_17865);
nand U18321 (N_18321,N_17566,N_17829);
or U18322 (N_18322,N_17959,N_17998);
nand U18323 (N_18323,N_17569,N_17970);
xor U18324 (N_18324,N_17749,N_17560);
and U18325 (N_18325,N_17873,N_17526);
and U18326 (N_18326,N_17645,N_17962);
nor U18327 (N_18327,N_17633,N_17622);
xnor U18328 (N_18328,N_17824,N_17989);
and U18329 (N_18329,N_17958,N_17810);
nand U18330 (N_18330,N_17692,N_17916);
nand U18331 (N_18331,N_17916,N_17817);
or U18332 (N_18332,N_17558,N_17604);
nand U18333 (N_18333,N_17999,N_17591);
and U18334 (N_18334,N_17897,N_17765);
nand U18335 (N_18335,N_17548,N_17882);
nand U18336 (N_18336,N_17512,N_17740);
nor U18337 (N_18337,N_17987,N_17772);
xor U18338 (N_18338,N_17880,N_17957);
and U18339 (N_18339,N_17519,N_17802);
nor U18340 (N_18340,N_17731,N_17696);
nand U18341 (N_18341,N_17603,N_17764);
nand U18342 (N_18342,N_17579,N_17933);
and U18343 (N_18343,N_17552,N_17807);
and U18344 (N_18344,N_17897,N_17862);
nor U18345 (N_18345,N_17966,N_17653);
and U18346 (N_18346,N_17612,N_17708);
or U18347 (N_18347,N_17903,N_17692);
nand U18348 (N_18348,N_17997,N_17965);
xnor U18349 (N_18349,N_17654,N_17797);
or U18350 (N_18350,N_17571,N_17927);
nand U18351 (N_18351,N_17806,N_17740);
or U18352 (N_18352,N_17598,N_17531);
nor U18353 (N_18353,N_17632,N_17514);
and U18354 (N_18354,N_17837,N_17922);
or U18355 (N_18355,N_17877,N_17729);
or U18356 (N_18356,N_17722,N_17568);
nand U18357 (N_18357,N_17731,N_17676);
and U18358 (N_18358,N_17550,N_17736);
nand U18359 (N_18359,N_17763,N_17732);
and U18360 (N_18360,N_17833,N_17520);
nand U18361 (N_18361,N_17738,N_17737);
nand U18362 (N_18362,N_17683,N_17674);
or U18363 (N_18363,N_17897,N_17610);
xnor U18364 (N_18364,N_17955,N_17977);
xnor U18365 (N_18365,N_17615,N_17759);
and U18366 (N_18366,N_17609,N_17635);
or U18367 (N_18367,N_17506,N_17831);
and U18368 (N_18368,N_17912,N_17718);
or U18369 (N_18369,N_17676,N_17615);
xnor U18370 (N_18370,N_17642,N_17639);
and U18371 (N_18371,N_17988,N_17884);
xnor U18372 (N_18372,N_17814,N_17644);
nor U18373 (N_18373,N_17510,N_17533);
or U18374 (N_18374,N_17934,N_17902);
nor U18375 (N_18375,N_17573,N_17525);
xor U18376 (N_18376,N_17675,N_17814);
nor U18377 (N_18377,N_17556,N_17865);
xnor U18378 (N_18378,N_17661,N_17784);
xor U18379 (N_18379,N_17687,N_17955);
nor U18380 (N_18380,N_17611,N_17557);
or U18381 (N_18381,N_17867,N_17704);
xnor U18382 (N_18382,N_17940,N_17701);
xor U18383 (N_18383,N_17907,N_17881);
or U18384 (N_18384,N_17994,N_17618);
and U18385 (N_18385,N_17690,N_17615);
or U18386 (N_18386,N_17555,N_17547);
and U18387 (N_18387,N_17782,N_17990);
nand U18388 (N_18388,N_17637,N_17680);
nand U18389 (N_18389,N_17744,N_17655);
or U18390 (N_18390,N_17801,N_17954);
nand U18391 (N_18391,N_17835,N_17713);
nand U18392 (N_18392,N_17537,N_17669);
xor U18393 (N_18393,N_17580,N_17561);
nand U18394 (N_18394,N_17925,N_17745);
and U18395 (N_18395,N_17977,N_17604);
nand U18396 (N_18396,N_17618,N_17770);
and U18397 (N_18397,N_17667,N_17950);
nor U18398 (N_18398,N_17715,N_17526);
and U18399 (N_18399,N_17693,N_17580);
nor U18400 (N_18400,N_17691,N_17605);
nor U18401 (N_18401,N_17626,N_17856);
xor U18402 (N_18402,N_17847,N_17777);
nor U18403 (N_18403,N_17755,N_17999);
nand U18404 (N_18404,N_17910,N_17754);
and U18405 (N_18405,N_17695,N_17564);
or U18406 (N_18406,N_17768,N_17898);
nand U18407 (N_18407,N_17770,N_17594);
xor U18408 (N_18408,N_17838,N_17786);
and U18409 (N_18409,N_17557,N_17944);
and U18410 (N_18410,N_17908,N_17833);
nand U18411 (N_18411,N_17691,N_17979);
nand U18412 (N_18412,N_17712,N_17859);
xor U18413 (N_18413,N_17648,N_17936);
or U18414 (N_18414,N_17781,N_17734);
xor U18415 (N_18415,N_17964,N_17533);
nand U18416 (N_18416,N_17838,N_17548);
nand U18417 (N_18417,N_17515,N_17970);
or U18418 (N_18418,N_17748,N_17734);
or U18419 (N_18419,N_17562,N_17634);
and U18420 (N_18420,N_17936,N_17857);
xnor U18421 (N_18421,N_17679,N_17901);
xor U18422 (N_18422,N_17610,N_17972);
or U18423 (N_18423,N_17723,N_17580);
and U18424 (N_18424,N_17809,N_17825);
or U18425 (N_18425,N_17611,N_17857);
nor U18426 (N_18426,N_17873,N_17555);
or U18427 (N_18427,N_17861,N_17519);
nand U18428 (N_18428,N_17834,N_17757);
nand U18429 (N_18429,N_17581,N_17660);
and U18430 (N_18430,N_17827,N_17951);
nor U18431 (N_18431,N_17588,N_17720);
xor U18432 (N_18432,N_17812,N_17912);
or U18433 (N_18433,N_17923,N_17552);
nand U18434 (N_18434,N_17787,N_17831);
xor U18435 (N_18435,N_17804,N_17814);
nor U18436 (N_18436,N_17652,N_17704);
or U18437 (N_18437,N_17757,N_17809);
or U18438 (N_18438,N_17693,N_17769);
nand U18439 (N_18439,N_17647,N_17759);
or U18440 (N_18440,N_17842,N_17719);
and U18441 (N_18441,N_17551,N_17682);
nand U18442 (N_18442,N_17505,N_17651);
xor U18443 (N_18443,N_17686,N_17632);
or U18444 (N_18444,N_17860,N_17652);
and U18445 (N_18445,N_17644,N_17743);
nand U18446 (N_18446,N_17862,N_17637);
or U18447 (N_18447,N_17520,N_17515);
or U18448 (N_18448,N_17685,N_17573);
nor U18449 (N_18449,N_17614,N_17759);
nand U18450 (N_18450,N_17813,N_17778);
and U18451 (N_18451,N_17545,N_17756);
nand U18452 (N_18452,N_17860,N_17512);
or U18453 (N_18453,N_17690,N_17700);
xnor U18454 (N_18454,N_17601,N_17682);
nor U18455 (N_18455,N_17769,N_17935);
nand U18456 (N_18456,N_17631,N_17914);
nor U18457 (N_18457,N_17697,N_17589);
nand U18458 (N_18458,N_17563,N_17674);
xor U18459 (N_18459,N_17866,N_17916);
nand U18460 (N_18460,N_17880,N_17583);
xor U18461 (N_18461,N_17795,N_17815);
and U18462 (N_18462,N_17938,N_17507);
or U18463 (N_18463,N_17779,N_17544);
or U18464 (N_18464,N_17659,N_17999);
xnor U18465 (N_18465,N_17549,N_17907);
and U18466 (N_18466,N_17714,N_17734);
xnor U18467 (N_18467,N_17523,N_17921);
and U18468 (N_18468,N_17593,N_17505);
nand U18469 (N_18469,N_17502,N_17609);
and U18470 (N_18470,N_17705,N_17936);
and U18471 (N_18471,N_17638,N_17684);
nor U18472 (N_18472,N_17611,N_17658);
xnor U18473 (N_18473,N_17968,N_17830);
nor U18474 (N_18474,N_17733,N_17556);
and U18475 (N_18475,N_17973,N_17798);
nand U18476 (N_18476,N_17873,N_17742);
or U18477 (N_18477,N_17878,N_17614);
and U18478 (N_18478,N_17775,N_17862);
xnor U18479 (N_18479,N_17884,N_17501);
or U18480 (N_18480,N_17709,N_17739);
nor U18481 (N_18481,N_17658,N_17970);
xnor U18482 (N_18482,N_17996,N_17622);
xnor U18483 (N_18483,N_17997,N_17975);
xnor U18484 (N_18484,N_17986,N_17864);
nor U18485 (N_18485,N_17569,N_17706);
xnor U18486 (N_18486,N_17917,N_17514);
xor U18487 (N_18487,N_17847,N_17735);
xor U18488 (N_18488,N_17726,N_17622);
and U18489 (N_18489,N_17566,N_17628);
nor U18490 (N_18490,N_17516,N_17712);
or U18491 (N_18491,N_17541,N_17858);
nor U18492 (N_18492,N_17580,N_17852);
and U18493 (N_18493,N_17634,N_17611);
and U18494 (N_18494,N_17641,N_17808);
nand U18495 (N_18495,N_17547,N_17864);
and U18496 (N_18496,N_17537,N_17946);
or U18497 (N_18497,N_17742,N_17961);
nor U18498 (N_18498,N_17770,N_17713);
nor U18499 (N_18499,N_17528,N_17601);
nor U18500 (N_18500,N_18361,N_18410);
or U18501 (N_18501,N_18433,N_18370);
and U18502 (N_18502,N_18440,N_18258);
or U18503 (N_18503,N_18356,N_18055);
xnor U18504 (N_18504,N_18204,N_18305);
nor U18505 (N_18505,N_18363,N_18067);
or U18506 (N_18506,N_18398,N_18143);
and U18507 (N_18507,N_18111,N_18409);
nand U18508 (N_18508,N_18183,N_18148);
and U18509 (N_18509,N_18252,N_18051);
nand U18510 (N_18510,N_18322,N_18181);
nor U18511 (N_18511,N_18100,N_18401);
and U18512 (N_18512,N_18493,N_18019);
nand U18513 (N_18513,N_18281,N_18288);
nand U18514 (N_18514,N_18229,N_18109);
nand U18515 (N_18515,N_18166,N_18053);
or U18516 (N_18516,N_18466,N_18395);
nor U18517 (N_18517,N_18479,N_18415);
nand U18518 (N_18518,N_18221,N_18414);
nand U18519 (N_18519,N_18133,N_18357);
nand U18520 (N_18520,N_18056,N_18187);
or U18521 (N_18521,N_18323,N_18169);
xnor U18522 (N_18522,N_18317,N_18303);
and U18523 (N_18523,N_18245,N_18113);
or U18524 (N_18524,N_18249,N_18329);
xnor U18525 (N_18525,N_18330,N_18309);
and U18526 (N_18526,N_18435,N_18304);
or U18527 (N_18527,N_18441,N_18134);
nor U18528 (N_18528,N_18485,N_18428);
nor U18529 (N_18529,N_18394,N_18349);
nand U18530 (N_18530,N_18348,N_18200);
or U18531 (N_18531,N_18327,N_18460);
nand U18532 (N_18532,N_18312,N_18465);
nand U18533 (N_18533,N_18332,N_18117);
or U18534 (N_18534,N_18475,N_18246);
nor U18535 (N_18535,N_18197,N_18144);
and U18536 (N_18536,N_18066,N_18346);
nor U18537 (N_18537,N_18145,N_18037);
nor U18538 (N_18538,N_18264,N_18343);
nor U18539 (N_18539,N_18175,N_18426);
nand U18540 (N_18540,N_18017,N_18400);
nand U18541 (N_18541,N_18020,N_18368);
and U18542 (N_18542,N_18146,N_18225);
nor U18543 (N_18543,N_18129,N_18034);
xor U18544 (N_18544,N_18456,N_18052);
nand U18545 (N_18545,N_18238,N_18006);
nand U18546 (N_18546,N_18021,N_18198);
nor U18547 (N_18547,N_18339,N_18495);
and U18548 (N_18548,N_18326,N_18098);
or U18549 (N_18549,N_18116,N_18282);
nand U18550 (N_18550,N_18230,N_18096);
or U18551 (N_18551,N_18344,N_18074);
nand U18552 (N_18552,N_18242,N_18172);
or U18553 (N_18553,N_18408,N_18499);
xnor U18554 (N_18554,N_18075,N_18489);
and U18555 (N_18555,N_18022,N_18331);
and U18556 (N_18556,N_18217,N_18110);
and U18557 (N_18557,N_18285,N_18399);
nand U18558 (N_18558,N_18259,N_18419);
xnor U18559 (N_18559,N_18418,N_18201);
nor U18560 (N_18560,N_18027,N_18023);
or U18561 (N_18561,N_18379,N_18089);
nor U18562 (N_18562,N_18417,N_18091);
xor U18563 (N_18563,N_18284,N_18255);
nor U18564 (N_18564,N_18454,N_18464);
and U18565 (N_18565,N_18068,N_18458);
xnor U18566 (N_18566,N_18371,N_18218);
nand U18567 (N_18567,N_18035,N_18293);
and U18568 (N_18568,N_18373,N_18459);
xor U18569 (N_18569,N_18468,N_18234);
xnor U18570 (N_18570,N_18267,N_18412);
or U18571 (N_18571,N_18321,N_18397);
and U18572 (N_18572,N_18380,N_18286);
nor U18573 (N_18573,N_18083,N_18290);
or U18574 (N_18574,N_18029,N_18248);
nor U18575 (N_18575,N_18140,N_18112);
or U18576 (N_18576,N_18353,N_18277);
nor U18577 (N_18577,N_18043,N_18271);
nand U18578 (N_18578,N_18061,N_18093);
xnor U18579 (N_18579,N_18260,N_18173);
nor U18580 (N_18580,N_18351,N_18488);
or U18581 (N_18581,N_18478,N_18388);
or U18582 (N_18582,N_18168,N_18461);
or U18583 (N_18583,N_18208,N_18250);
or U18584 (N_18584,N_18064,N_18270);
xor U18585 (N_18585,N_18039,N_18220);
xnor U18586 (N_18586,N_18231,N_18206);
and U18587 (N_18587,N_18185,N_18387);
nor U18588 (N_18588,N_18085,N_18265);
or U18589 (N_18589,N_18384,N_18236);
or U18590 (N_18590,N_18097,N_18115);
xor U18591 (N_18591,N_18307,N_18196);
nor U18592 (N_18592,N_18268,N_18429);
nand U18593 (N_18593,N_18421,N_18184);
nand U18594 (N_18594,N_18299,N_18287);
xor U18595 (N_18595,N_18060,N_18416);
or U18596 (N_18596,N_18158,N_18030);
or U18597 (N_18597,N_18124,N_18448);
or U18598 (N_18598,N_18063,N_18391);
xnor U18599 (N_18599,N_18015,N_18192);
nand U18600 (N_18600,N_18136,N_18130);
or U18601 (N_18601,N_18223,N_18228);
and U18602 (N_18602,N_18182,N_18033);
and U18603 (N_18603,N_18247,N_18402);
nor U18604 (N_18604,N_18011,N_18310);
and U18605 (N_18605,N_18237,N_18072);
or U18606 (N_18606,N_18390,N_18233);
or U18607 (N_18607,N_18362,N_18407);
xor U18608 (N_18608,N_18154,N_18057);
xnor U18609 (N_18609,N_18449,N_18122);
or U18610 (N_18610,N_18123,N_18420);
or U18611 (N_18611,N_18202,N_18383);
nand U18612 (N_18612,N_18498,N_18194);
nor U18613 (N_18613,N_18308,N_18472);
nor U18614 (N_18614,N_18040,N_18207);
and U18615 (N_18615,N_18215,N_18147);
and U18616 (N_18616,N_18241,N_18012);
nand U18617 (N_18617,N_18014,N_18107);
nor U18618 (N_18618,N_18275,N_18048);
nand U18619 (N_18619,N_18090,N_18176);
nand U18620 (N_18620,N_18151,N_18278);
nor U18621 (N_18621,N_18203,N_18396);
nand U18622 (N_18622,N_18024,N_18199);
nor U18623 (N_18623,N_18337,N_18177);
nand U18624 (N_18624,N_18046,N_18452);
xnor U18625 (N_18625,N_18491,N_18497);
nor U18626 (N_18626,N_18354,N_18073);
and U18627 (N_18627,N_18009,N_18042);
nand U18628 (N_18628,N_18381,N_18222);
nand U18629 (N_18629,N_18347,N_18018);
and U18630 (N_18630,N_18077,N_18125);
nor U18631 (N_18631,N_18119,N_18050);
nor U18632 (N_18632,N_18439,N_18150);
and U18633 (N_18633,N_18082,N_18432);
and U18634 (N_18634,N_18101,N_18316);
or U18635 (N_18635,N_18405,N_18374);
and U18636 (N_18636,N_18224,N_18069);
nor U18637 (N_18637,N_18137,N_18131);
xnor U18638 (N_18638,N_18164,N_18477);
or U18639 (N_18639,N_18126,N_18302);
xor U18640 (N_18640,N_18049,N_18434);
and U18641 (N_18641,N_18128,N_18291);
xnor U18642 (N_18642,N_18360,N_18062);
or U18643 (N_18643,N_18045,N_18080);
or U18644 (N_18644,N_18179,N_18191);
xor U18645 (N_18645,N_18445,N_18438);
xnor U18646 (N_18646,N_18104,N_18422);
and U18647 (N_18647,N_18482,N_18295);
or U18648 (N_18648,N_18094,N_18254);
xor U18649 (N_18649,N_18494,N_18292);
and U18650 (N_18650,N_18319,N_18139);
and U18651 (N_18651,N_18423,N_18372);
nor U18652 (N_18652,N_18274,N_18078);
and U18653 (N_18653,N_18002,N_18451);
or U18654 (N_18654,N_18219,N_18135);
nand U18655 (N_18655,N_18016,N_18364);
or U18656 (N_18656,N_18365,N_18038);
nor U18657 (N_18657,N_18359,N_18257);
or U18658 (N_18658,N_18340,N_18335);
nor U18659 (N_18659,N_18272,N_18296);
and U18660 (N_18660,N_18232,N_18193);
and U18661 (N_18661,N_18160,N_18403);
nor U18662 (N_18662,N_18141,N_18484);
xor U18663 (N_18663,N_18178,N_18496);
or U18664 (N_18664,N_18032,N_18079);
or U18665 (N_18665,N_18092,N_18081);
nand U18666 (N_18666,N_18411,N_18457);
or U18667 (N_18667,N_18437,N_18188);
nand U18668 (N_18668,N_18358,N_18386);
nand U18669 (N_18669,N_18476,N_18306);
or U18670 (N_18670,N_18297,N_18253);
nand U18671 (N_18671,N_18120,N_18328);
or U18672 (N_18672,N_18350,N_18474);
or U18673 (N_18673,N_18086,N_18480);
nor U18674 (N_18674,N_18318,N_18031);
nand U18675 (N_18675,N_18070,N_18170);
nand U18676 (N_18676,N_18008,N_18443);
or U18677 (N_18677,N_18369,N_18171);
xor U18678 (N_18678,N_18167,N_18161);
or U18679 (N_18679,N_18156,N_18262);
nor U18680 (N_18680,N_18084,N_18453);
and U18681 (N_18681,N_18481,N_18470);
or U18682 (N_18682,N_18393,N_18367);
nor U18683 (N_18683,N_18149,N_18324);
nor U18684 (N_18684,N_18342,N_18054);
and U18685 (N_18685,N_18382,N_18446);
xnor U18686 (N_18686,N_18355,N_18243);
nor U18687 (N_18687,N_18256,N_18462);
and U18688 (N_18688,N_18471,N_18280);
and U18689 (N_18689,N_18121,N_18235);
nand U18690 (N_18690,N_18162,N_18044);
nand U18691 (N_18691,N_18026,N_18138);
nand U18692 (N_18692,N_18376,N_18186);
nor U18693 (N_18693,N_18025,N_18430);
and U18694 (N_18694,N_18227,N_18283);
and U18695 (N_18695,N_18320,N_18406);
or U18696 (N_18696,N_18102,N_18276);
nand U18697 (N_18697,N_18240,N_18311);
or U18698 (N_18698,N_18004,N_18298);
nand U18699 (N_18699,N_18279,N_18028);
nand U18700 (N_18700,N_18076,N_18180);
or U18701 (N_18701,N_18157,N_18103);
xnor U18702 (N_18702,N_18490,N_18333);
xnor U18703 (N_18703,N_18263,N_18105);
nand U18704 (N_18704,N_18071,N_18338);
xnor U18705 (N_18705,N_18239,N_18226);
nand U18706 (N_18706,N_18189,N_18013);
or U18707 (N_18707,N_18289,N_18155);
nand U18708 (N_18708,N_18244,N_18377);
or U18709 (N_18709,N_18294,N_18261);
xnor U18710 (N_18710,N_18214,N_18152);
or U18711 (N_18711,N_18467,N_18487);
xnor U18712 (N_18712,N_18132,N_18392);
nor U18713 (N_18713,N_18007,N_18486);
or U18714 (N_18714,N_18450,N_18425);
xor U18715 (N_18715,N_18216,N_18003);
nand U18716 (N_18716,N_18127,N_18047);
xnor U18717 (N_18717,N_18345,N_18036);
xor U18718 (N_18718,N_18389,N_18174);
and U18719 (N_18719,N_18251,N_18142);
xor U18720 (N_18720,N_18114,N_18315);
nand U18721 (N_18721,N_18404,N_18483);
and U18722 (N_18722,N_18473,N_18001);
nor U18723 (N_18723,N_18336,N_18041);
nor U18724 (N_18724,N_18153,N_18444);
nor U18725 (N_18725,N_18301,N_18058);
and U18726 (N_18726,N_18266,N_18385);
or U18727 (N_18727,N_18269,N_18436);
or U18728 (N_18728,N_18108,N_18325);
or U18729 (N_18729,N_18212,N_18341);
xor U18730 (N_18730,N_18463,N_18059);
nor U18731 (N_18731,N_18099,N_18210);
nand U18732 (N_18732,N_18088,N_18334);
or U18733 (N_18733,N_18195,N_18314);
or U18734 (N_18734,N_18442,N_18163);
and U18735 (N_18735,N_18447,N_18492);
nor U18736 (N_18736,N_18366,N_18313);
nor U18737 (N_18737,N_18190,N_18209);
nand U18738 (N_18738,N_18087,N_18273);
and U18739 (N_18739,N_18431,N_18065);
and U18740 (N_18740,N_18469,N_18378);
and U18741 (N_18741,N_18424,N_18211);
nor U18742 (N_18742,N_18095,N_18010);
and U18743 (N_18743,N_18000,N_18213);
and U18744 (N_18744,N_18413,N_18427);
nor U18745 (N_18745,N_18352,N_18118);
and U18746 (N_18746,N_18455,N_18106);
and U18747 (N_18747,N_18159,N_18300);
and U18748 (N_18748,N_18165,N_18375);
nand U18749 (N_18749,N_18205,N_18005);
nor U18750 (N_18750,N_18410,N_18040);
or U18751 (N_18751,N_18455,N_18264);
xnor U18752 (N_18752,N_18051,N_18340);
or U18753 (N_18753,N_18294,N_18242);
nor U18754 (N_18754,N_18326,N_18284);
and U18755 (N_18755,N_18082,N_18154);
xor U18756 (N_18756,N_18338,N_18406);
or U18757 (N_18757,N_18000,N_18476);
and U18758 (N_18758,N_18430,N_18106);
xnor U18759 (N_18759,N_18181,N_18023);
or U18760 (N_18760,N_18418,N_18162);
xnor U18761 (N_18761,N_18088,N_18288);
xor U18762 (N_18762,N_18090,N_18403);
xnor U18763 (N_18763,N_18457,N_18203);
xor U18764 (N_18764,N_18000,N_18438);
or U18765 (N_18765,N_18206,N_18417);
nor U18766 (N_18766,N_18130,N_18014);
nor U18767 (N_18767,N_18019,N_18480);
or U18768 (N_18768,N_18088,N_18068);
and U18769 (N_18769,N_18034,N_18455);
or U18770 (N_18770,N_18357,N_18039);
and U18771 (N_18771,N_18125,N_18476);
xnor U18772 (N_18772,N_18138,N_18496);
nor U18773 (N_18773,N_18199,N_18156);
nand U18774 (N_18774,N_18202,N_18107);
xor U18775 (N_18775,N_18279,N_18090);
and U18776 (N_18776,N_18379,N_18055);
or U18777 (N_18777,N_18019,N_18332);
or U18778 (N_18778,N_18207,N_18122);
nand U18779 (N_18779,N_18311,N_18368);
nor U18780 (N_18780,N_18325,N_18037);
xor U18781 (N_18781,N_18093,N_18156);
and U18782 (N_18782,N_18447,N_18412);
and U18783 (N_18783,N_18021,N_18068);
xor U18784 (N_18784,N_18158,N_18093);
xor U18785 (N_18785,N_18141,N_18187);
xnor U18786 (N_18786,N_18373,N_18106);
xor U18787 (N_18787,N_18024,N_18371);
xnor U18788 (N_18788,N_18248,N_18176);
nand U18789 (N_18789,N_18005,N_18226);
nand U18790 (N_18790,N_18057,N_18386);
nand U18791 (N_18791,N_18249,N_18211);
nor U18792 (N_18792,N_18416,N_18192);
or U18793 (N_18793,N_18107,N_18018);
nand U18794 (N_18794,N_18280,N_18351);
nor U18795 (N_18795,N_18414,N_18256);
or U18796 (N_18796,N_18192,N_18351);
nand U18797 (N_18797,N_18052,N_18192);
xnor U18798 (N_18798,N_18135,N_18362);
nand U18799 (N_18799,N_18149,N_18178);
nand U18800 (N_18800,N_18413,N_18412);
xor U18801 (N_18801,N_18327,N_18194);
xor U18802 (N_18802,N_18210,N_18381);
xnor U18803 (N_18803,N_18267,N_18284);
and U18804 (N_18804,N_18237,N_18202);
xor U18805 (N_18805,N_18318,N_18235);
or U18806 (N_18806,N_18423,N_18153);
or U18807 (N_18807,N_18263,N_18001);
xnor U18808 (N_18808,N_18001,N_18305);
or U18809 (N_18809,N_18148,N_18354);
xor U18810 (N_18810,N_18396,N_18094);
and U18811 (N_18811,N_18460,N_18426);
xnor U18812 (N_18812,N_18347,N_18407);
nor U18813 (N_18813,N_18212,N_18492);
xnor U18814 (N_18814,N_18025,N_18127);
nand U18815 (N_18815,N_18448,N_18299);
or U18816 (N_18816,N_18463,N_18083);
nand U18817 (N_18817,N_18499,N_18411);
or U18818 (N_18818,N_18284,N_18116);
xor U18819 (N_18819,N_18218,N_18459);
nor U18820 (N_18820,N_18024,N_18294);
xor U18821 (N_18821,N_18117,N_18455);
xor U18822 (N_18822,N_18485,N_18360);
or U18823 (N_18823,N_18400,N_18462);
xor U18824 (N_18824,N_18352,N_18159);
or U18825 (N_18825,N_18343,N_18137);
and U18826 (N_18826,N_18042,N_18022);
xor U18827 (N_18827,N_18465,N_18244);
nand U18828 (N_18828,N_18187,N_18091);
or U18829 (N_18829,N_18306,N_18191);
and U18830 (N_18830,N_18430,N_18123);
nand U18831 (N_18831,N_18043,N_18077);
nor U18832 (N_18832,N_18127,N_18251);
or U18833 (N_18833,N_18286,N_18231);
xnor U18834 (N_18834,N_18403,N_18153);
nand U18835 (N_18835,N_18444,N_18468);
and U18836 (N_18836,N_18190,N_18403);
or U18837 (N_18837,N_18363,N_18236);
nor U18838 (N_18838,N_18206,N_18341);
nand U18839 (N_18839,N_18273,N_18239);
and U18840 (N_18840,N_18412,N_18045);
nand U18841 (N_18841,N_18192,N_18168);
or U18842 (N_18842,N_18419,N_18136);
or U18843 (N_18843,N_18390,N_18042);
or U18844 (N_18844,N_18259,N_18125);
nor U18845 (N_18845,N_18457,N_18432);
nand U18846 (N_18846,N_18364,N_18351);
xor U18847 (N_18847,N_18496,N_18314);
nor U18848 (N_18848,N_18105,N_18165);
and U18849 (N_18849,N_18342,N_18068);
or U18850 (N_18850,N_18430,N_18251);
or U18851 (N_18851,N_18055,N_18368);
nand U18852 (N_18852,N_18235,N_18022);
xnor U18853 (N_18853,N_18391,N_18305);
nor U18854 (N_18854,N_18251,N_18064);
nand U18855 (N_18855,N_18176,N_18027);
and U18856 (N_18856,N_18124,N_18371);
and U18857 (N_18857,N_18028,N_18403);
xor U18858 (N_18858,N_18493,N_18298);
xnor U18859 (N_18859,N_18486,N_18121);
xor U18860 (N_18860,N_18045,N_18332);
nor U18861 (N_18861,N_18290,N_18178);
or U18862 (N_18862,N_18052,N_18278);
xor U18863 (N_18863,N_18237,N_18060);
and U18864 (N_18864,N_18103,N_18094);
nor U18865 (N_18865,N_18090,N_18198);
nand U18866 (N_18866,N_18024,N_18462);
and U18867 (N_18867,N_18281,N_18034);
nor U18868 (N_18868,N_18073,N_18370);
nor U18869 (N_18869,N_18126,N_18495);
nor U18870 (N_18870,N_18068,N_18178);
nand U18871 (N_18871,N_18153,N_18359);
nor U18872 (N_18872,N_18081,N_18231);
and U18873 (N_18873,N_18087,N_18412);
xnor U18874 (N_18874,N_18365,N_18258);
and U18875 (N_18875,N_18383,N_18063);
or U18876 (N_18876,N_18233,N_18131);
xnor U18877 (N_18877,N_18313,N_18188);
nand U18878 (N_18878,N_18313,N_18147);
xnor U18879 (N_18879,N_18066,N_18212);
xor U18880 (N_18880,N_18420,N_18037);
and U18881 (N_18881,N_18302,N_18011);
nand U18882 (N_18882,N_18030,N_18096);
nor U18883 (N_18883,N_18400,N_18170);
nand U18884 (N_18884,N_18117,N_18237);
or U18885 (N_18885,N_18218,N_18034);
xnor U18886 (N_18886,N_18133,N_18321);
and U18887 (N_18887,N_18224,N_18072);
xor U18888 (N_18888,N_18077,N_18215);
and U18889 (N_18889,N_18447,N_18276);
and U18890 (N_18890,N_18162,N_18433);
and U18891 (N_18891,N_18016,N_18040);
or U18892 (N_18892,N_18168,N_18496);
nand U18893 (N_18893,N_18044,N_18055);
or U18894 (N_18894,N_18027,N_18175);
nand U18895 (N_18895,N_18100,N_18275);
nor U18896 (N_18896,N_18489,N_18448);
and U18897 (N_18897,N_18257,N_18052);
xnor U18898 (N_18898,N_18204,N_18015);
and U18899 (N_18899,N_18274,N_18105);
nand U18900 (N_18900,N_18218,N_18373);
and U18901 (N_18901,N_18417,N_18066);
nor U18902 (N_18902,N_18096,N_18016);
xor U18903 (N_18903,N_18077,N_18089);
xnor U18904 (N_18904,N_18387,N_18164);
and U18905 (N_18905,N_18260,N_18121);
nor U18906 (N_18906,N_18193,N_18083);
or U18907 (N_18907,N_18007,N_18452);
and U18908 (N_18908,N_18138,N_18215);
or U18909 (N_18909,N_18423,N_18481);
or U18910 (N_18910,N_18369,N_18248);
nor U18911 (N_18911,N_18159,N_18161);
and U18912 (N_18912,N_18018,N_18210);
nor U18913 (N_18913,N_18345,N_18363);
nand U18914 (N_18914,N_18453,N_18118);
and U18915 (N_18915,N_18007,N_18433);
nor U18916 (N_18916,N_18067,N_18298);
nand U18917 (N_18917,N_18339,N_18096);
nor U18918 (N_18918,N_18336,N_18146);
or U18919 (N_18919,N_18251,N_18327);
xnor U18920 (N_18920,N_18437,N_18006);
nor U18921 (N_18921,N_18443,N_18438);
nand U18922 (N_18922,N_18408,N_18117);
nor U18923 (N_18923,N_18157,N_18387);
or U18924 (N_18924,N_18384,N_18209);
xor U18925 (N_18925,N_18291,N_18175);
or U18926 (N_18926,N_18321,N_18494);
nor U18927 (N_18927,N_18001,N_18108);
or U18928 (N_18928,N_18160,N_18431);
and U18929 (N_18929,N_18410,N_18359);
or U18930 (N_18930,N_18300,N_18330);
or U18931 (N_18931,N_18075,N_18198);
and U18932 (N_18932,N_18448,N_18084);
nor U18933 (N_18933,N_18330,N_18364);
xor U18934 (N_18934,N_18055,N_18244);
xnor U18935 (N_18935,N_18246,N_18347);
and U18936 (N_18936,N_18008,N_18201);
nor U18937 (N_18937,N_18031,N_18480);
or U18938 (N_18938,N_18019,N_18280);
and U18939 (N_18939,N_18257,N_18209);
or U18940 (N_18940,N_18089,N_18432);
nand U18941 (N_18941,N_18467,N_18155);
nor U18942 (N_18942,N_18039,N_18112);
nand U18943 (N_18943,N_18362,N_18265);
nand U18944 (N_18944,N_18351,N_18161);
nor U18945 (N_18945,N_18140,N_18336);
and U18946 (N_18946,N_18450,N_18307);
nor U18947 (N_18947,N_18144,N_18097);
and U18948 (N_18948,N_18063,N_18309);
and U18949 (N_18949,N_18322,N_18260);
nor U18950 (N_18950,N_18084,N_18151);
or U18951 (N_18951,N_18336,N_18165);
nand U18952 (N_18952,N_18126,N_18371);
nor U18953 (N_18953,N_18312,N_18200);
nand U18954 (N_18954,N_18042,N_18182);
nand U18955 (N_18955,N_18215,N_18165);
nand U18956 (N_18956,N_18111,N_18005);
xor U18957 (N_18957,N_18166,N_18238);
and U18958 (N_18958,N_18159,N_18170);
nand U18959 (N_18959,N_18295,N_18137);
nand U18960 (N_18960,N_18462,N_18305);
xnor U18961 (N_18961,N_18462,N_18041);
nand U18962 (N_18962,N_18403,N_18436);
nand U18963 (N_18963,N_18233,N_18331);
and U18964 (N_18964,N_18152,N_18200);
xor U18965 (N_18965,N_18237,N_18386);
nand U18966 (N_18966,N_18492,N_18089);
and U18967 (N_18967,N_18049,N_18377);
nand U18968 (N_18968,N_18248,N_18322);
xnor U18969 (N_18969,N_18034,N_18124);
nor U18970 (N_18970,N_18114,N_18139);
or U18971 (N_18971,N_18344,N_18050);
or U18972 (N_18972,N_18485,N_18338);
xor U18973 (N_18973,N_18162,N_18310);
nand U18974 (N_18974,N_18181,N_18054);
xor U18975 (N_18975,N_18499,N_18468);
nor U18976 (N_18976,N_18122,N_18089);
nand U18977 (N_18977,N_18330,N_18048);
nor U18978 (N_18978,N_18112,N_18180);
or U18979 (N_18979,N_18391,N_18384);
nor U18980 (N_18980,N_18028,N_18081);
nor U18981 (N_18981,N_18197,N_18162);
xor U18982 (N_18982,N_18425,N_18333);
xnor U18983 (N_18983,N_18168,N_18076);
nor U18984 (N_18984,N_18237,N_18246);
nand U18985 (N_18985,N_18203,N_18271);
xnor U18986 (N_18986,N_18352,N_18024);
nor U18987 (N_18987,N_18015,N_18102);
nor U18988 (N_18988,N_18273,N_18125);
nor U18989 (N_18989,N_18083,N_18496);
and U18990 (N_18990,N_18088,N_18080);
nor U18991 (N_18991,N_18393,N_18263);
and U18992 (N_18992,N_18367,N_18039);
or U18993 (N_18993,N_18070,N_18204);
and U18994 (N_18994,N_18168,N_18199);
and U18995 (N_18995,N_18138,N_18301);
xnor U18996 (N_18996,N_18103,N_18091);
xnor U18997 (N_18997,N_18332,N_18277);
and U18998 (N_18998,N_18416,N_18142);
and U18999 (N_18999,N_18454,N_18408);
xor U19000 (N_19000,N_18935,N_18625);
or U19001 (N_19001,N_18794,N_18995);
nand U19002 (N_19002,N_18706,N_18890);
and U19003 (N_19003,N_18659,N_18901);
nand U19004 (N_19004,N_18926,N_18673);
nand U19005 (N_19005,N_18723,N_18754);
or U19006 (N_19006,N_18806,N_18899);
or U19007 (N_19007,N_18676,N_18656);
and U19008 (N_19008,N_18830,N_18955);
or U19009 (N_19009,N_18593,N_18562);
xnor U19010 (N_19010,N_18699,N_18517);
or U19011 (N_19011,N_18936,N_18829);
xnor U19012 (N_19012,N_18916,N_18712);
nor U19013 (N_19013,N_18972,N_18558);
nor U19014 (N_19014,N_18951,N_18559);
nor U19015 (N_19015,N_18502,N_18866);
xor U19016 (N_19016,N_18848,N_18822);
or U19017 (N_19017,N_18708,N_18937);
nand U19018 (N_19018,N_18949,N_18819);
and U19019 (N_19019,N_18931,N_18568);
nand U19020 (N_19020,N_18629,N_18545);
nand U19021 (N_19021,N_18898,N_18869);
xor U19022 (N_19022,N_18883,N_18617);
nor U19023 (N_19023,N_18698,N_18628);
nor U19024 (N_19024,N_18770,N_18504);
nand U19025 (N_19025,N_18792,N_18594);
xor U19026 (N_19026,N_18624,N_18555);
nand U19027 (N_19027,N_18726,N_18897);
and U19028 (N_19028,N_18560,N_18549);
nand U19029 (N_19029,N_18824,N_18700);
or U19030 (N_19030,N_18732,N_18881);
xor U19031 (N_19031,N_18574,N_18648);
xnor U19032 (N_19032,N_18512,N_18727);
nand U19033 (N_19033,N_18679,N_18613);
xnor U19034 (N_19034,N_18839,N_18932);
or U19035 (N_19035,N_18515,N_18831);
and U19036 (N_19036,N_18983,N_18526);
and U19037 (N_19037,N_18683,N_18705);
nor U19038 (N_19038,N_18996,N_18618);
or U19039 (N_19039,N_18967,N_18713);
nand U19040 (N_19040,N_18752,N_18561);
and U19041 (N_19041,N_18587,N_18685);
xor U19042 (N_19042,N_18525,N_18510);
nand U19043 (N_19043,N_18777,N_18841);
and U19044 (N_19044,N_18544,N_18785);
nor U19045 (N_19045,N_18578,N_18507);
or U19046 (N_19046,N_18772,N_18760);
nand U19047 (N_19047,N_18579,N_18582);
and U19048 (N_19048,N_18636,N_18532);
and U19049 (N_19049,N_18882,N_18756);
nor U19050 (N_19050,N_18720,N_18704);
nor U19051 (N_19051,N_18791,N_18552);
nor U19052 (N_19052,N_18500,N_18827);
xor U19053 (N_19053,N_18680,N_18787);
xnor U19054 (N_19054,N_18971,N_18516);
or U19055 (N_19055,N_18590,N_18646);
or U19056 (N_19056,N_18803,N_18854);
or U19057 (N_19057,N_18766,N_18759);
and U19058 (N_19058,N_18661,N_18911);
and U19059 (N_19059,N_18860,N_18797);
xor U19060 (N_19060,N_18779,N_18811);
nand U19061 (N_19061,N_18880,N_18874);
or U19062 (N_19062,N_18736,N_18551);
nor U19063 (N_19063,N_18832,N_18891);
and U19064 (N_19064,N_18722,N_18608);
nand U19065 (N_19065,N_18952,N_18564);
xnor U19066 (N_19066,N_18998,N_18573);
nand U19067 (N_19067,N_18684,N_18592);
or U19068 (N_19068,N_18817,N_18533);
and U19069 (N_19069,N_18924,N_18858);
nand U19070 (N_19070,N_18630,N_18609);
nand U19071 (N_19071,N_18658,N_18614);
and U19072 (N_19072,N_18553,N_18762);
and U19073 (N_19073,N_18912,N_18687);
nand U19074 (N_19074,N_18838,N_18847);
and U19075 (N_19075,N_18994,N_18538);
nand U19076 (N_19076,N_18585,N_18671);
and U19077 (N_19077,N_18729,N_18653);
or U19078 (N_19078,N_18634,N_18719);
nor U19079 (N_19079,N_18511,N_18984);
nand U19080 (N_19080,N_18980,N_18767);
nand U19081 (N_19081,N_18902,N_18690);
and U19082 (N_19082,N_18733,N_18796);
and U19083 (N_19083,N_18715,N_18765);
or U19084 (N_19084,N_18607,N_18521);
or U19085 (N_19085,N_18668,N_18606);
or U19086 (N_19086,N_18850,N_18725);
or U19087 (N_19087,N_18793,N_18818);
nor U19088 (N_19088,N_18600,N_18744);
nand U19089 (N_19089,N_18966,N_18844);
or U19090 (N_19090,N_18523,N_18695);
xor U19091 (N_19091,N_18776,N_18737);
or U19092 (N_19092,N_18717,N_18851);
nor U19093 (N_19093,N_18825,N_18710);
or U19094 (N_19094,N_18637,N_18993);
nor U19095 (N_19095,N_18989,N_18954);
and U19096 (N_19096,N_18863,N_18666);
xnor U19097 (N_19097,N_18519,N_18927);
and U19098 (N_19098,N_18997,N_18864);
nand U19099 (N_19099,N_18821,N_18669);
and U19100 (N_19100,N_18755,N_18815);
and U19101 (N_19101,N_18859,N_18893);
xnor U19102 (N_19102,N_18780,N_18612);
nor U19103 (N_19103,N_18900,N_18694);
xor U19104 (N_19104,N_18651,N_18702);
xor U19105 (N_19105,N_18978,N_18915);
xnor U19106 (N_19106,N_18956,N_18627);
xor U19107 (N_19107,N_18716,N_18662);
or U19108 (N_19108,N_18742,N_18670);
and U19109 (N_19109,N_18639,N_18961);
and U19110 (N_19110,N_18960,N_18657);
and U19111 (N_19111,N_18745,N_18513);
nand U19112 (N_19112,N_18878,N_18746);
xor U19113 (N_19113,N_18773,N_18524);
nand U19114 (N_19114,N_18784,N_18798);
or U19115 (N_19115,N_18789,N_18686);
and U19116 (N_19116,N_18988,N_18535);
xnor U19117 (N_19117,N_18758,N_18743);
xnor U19118 (N_19118,N_18906,N_18539);
nand U19119 (N_19119,N_18718,N_18801);
nand U19120 (N_19120,N_18570,N_18734);
xor U19121 (N_19121,N_18580,N_18596);
or U19122 (N_19122,N_18509,N_18833);
nand U19123 (N_19123,N_18884,N_18853);
nand U19124 (N_19124,N_18977,N_18922);
and U19125 (N_19125,N_18693,N_18649);
nor U19126 (N_19126,N_18944,N_18602);
and U19127 (N_19127,N_18923,N_18976);
or U19128 (N_19128,N_18595,N_18805);
and U19129 (N_19129,N_18885,N_18692);
or U19130 (N_19130,N_18855,N_18589);
and U19131 (N_19131,N_18871,N_18810);
nand U19132 (N_19132,N_18753,N_18808);
xor U19133 (N_19133,N_18632,N_18599);
nor U19134 (N_19134,N_18527,N_18550);
and U19135 (N_19135,N_18938,N_18642);
and U19136 (N_19136,N_18862,N_18540);
and U19137 (N_19137,N_18894,N_18514);
nand U19138 (N_19138,N_18774,N_18873);
and U19139 (N_19139,N_18925,N_18889);
or U19140 (N_19140,N_18775,N_18541);
and U19141 (N_19141,N_18895,N_18849);
xor U19142 (N_19142,N_18645,N_18908);
xor U19143 (N_19143,N_18748,N_18888);
nand U19144 (N_19144,N_18800,N_18728);
and U19145 (N_19145,N_18957,N_18750);
and U19146 (N_19146,N_18751,N_18667);
and U19147 (N_19147,N_18799,N_18530);
and U19148 (N_19148,N_18741,N_18528);
and U19149 (N_19149,N_18577,N_18531);
nor U19150 (N_19150,N_18586,N_18962);
and U19151 (N_19151,N_18857,N_18946);
and U19152 (N_19152,N_18826,N_18563);
nand U19153 (N_19153,N_18677,N_18761);
nor U19154 (N_19154,N_18622,N_18747);
nand U19155 (N_19155,N_18782,N_18868);
nand U19156 (N_19156,N_18730,N_18537);
or U19157 (N_19157,N_18711,N_18681);
or U19158 (N_19158,N_18663,N_18764);
and U19159 (N_19159,N_18616,N_18768);
nand U19160 (N_19160,N_18929,N_18975);
and U19161 (N_19161,N_18876,N_18992);
xnor U19162 (N_19162,N_18974,N_18964);
or U19163 (N_19163,N_18940,N_18979);
or U19164 (N_19164,N_18757,N_18739);
xnor U19165 (N_19165,N_18626,N_18565);
nand U19166 (N_19166,N_18566,N_18675);
xor U19167 (N_19167,N_18837,N_18620);
nor U19168 (N_19168,N_18875,N_18691);
nor U19169 (N_19169,N_18583,N_18548);
and U19170 (N_19170,N_18968,N_18852);
xnor U19171 (N_19171,N_18917,N_18856);
xor U19172 (N_19172,N_18763,N_18571);
xnor U19173 (N_19173,N_18603,N_18921);
xnor U19174 (N_19174,N_18543,N_18892);
nor U19175 (N_19175,N_18913,N_18598);
nand U19176 (N_19176,N_18534,N_18999);
nor U19177 (N_19177,N_18556,N_18738);
or U19178 (N_19178,N_18947,N_18572);
xor U19179 (N_19179,N_18814,N_18865);
xnor U19180 (N_19180,N_18790,N_18861);
and U19181 (N_19181,N_18807,N_18591);
xor U19182 (N_19182,N_18621,N_18703);
nand U19183 (N_19183,N_18945,N_18778);
and U19184 (N_19184,N_18641,N_18948);
nand U19185 (N_19185,N_18554,N_18879);
and U19186 (N_19186,N_18633,N_18678);
xor U19187 (N_19187,N_18689,N_18816);
nand U19188 (N_19188,N_18836,N_18547);
xor U19189 (N_19189,N_18597,N_18652);
and U19190 (N_19190,N_18877,N_18735);
and U19191 (N_19191,N_18781,N_18820);
xnor U19192 (N_19192,N_18887,N_18843);
nand U19193 (N_19193,N_18963,N_18542);
xnor U19194 (N_19194,N_18520,N_18605);
nor U19195 (N_19195,N_18982,N_18501);
and U19196 (N_19196,N_18688,N_18672);
nand U19197 (N_19197,N_18985,N_18828);
nor U19198 (N_19198,N_18909,N_18958);
and U19199 (N_19199,N_18953,N_18904);
nand U19200 (N_19200,N_18508,N_18886);
nand U19201 (N_19201,N_18804,N_18584);
or U19202 (N_19202,N_18823,N_18990);
nand U19203 (N_19203,N_18987,N_18802);
xor U19204 (N_19204,N_18918,N_18867);
nand U19205 (N_19205,N_18788,N_18522);
nand U19206 (N_19206,N_18576,N_18575);
nor U19207 (N_19207,N_18569,N_18943);
nor U19208 (N_19208,N_18934,N_18601);
xor U19209 (N_19209,N_18795,N_18655);
and U19210 (N_19210,N_18643,N_18834);
nand U19211 (N_19211,N_18872,N_18812);
nor U19212 (N_19212,N_18682,N_18503);
or U19213 (N_19213,N_18870,N_18939);
nand U19214 (N_19214,N_18644,N_18840);
nor U19215 (N_19215,N_18986,N_18950);
nand U19216 (N_19216,N_18933,N_18707);
or U19217 (N_19217,N_18506,N_18635);
and U19218 (N_19218,N_18709,N_18674);
nor U19219 (N_19219,N_18959,N_18981);
and U19220 (N_19220,N_18623,N_18665);
and U19221 (N_19221,N_18941,N_18905);
xor U19222 (N_19222,N_18965,N_18610);
xor U19223 (N_19223,N_18647,N_18697);
and U19224 (N_19224,N_18611,N_18724);
and U19225 (N_19225,N_18567,N_18638);
and U19226 (N_19226,N_18581,N_18546);
and U19227 (N_19227,N_18664,N_18910);
xor U19228 (N_19228,N_18604,N_18518);
or U19229 (N_19229,N_18615,N_18701);
xnor U19230 (N_19230,N_18650,N_18973);
and U19231 (N_19231,N_18557,N_18845);
or U19232 (N_19232,N_18930,N_18536);
nand U19233 (N_19233,N_18896,N_18588);
and U19234 (N_19234,N_18942,N_18505);
and U19235 (N_19235,N_18991,N_18970);
nand U19236 (N_19236,N_18928,N_18631);
and U19237 (N_19237,N_18919,N_18809);
xnor U19238 (N_19238,N_18769,N_18846);
or U19239 (N_19239,N_18740,N_18721);
and U19240 (N_19240,N_18920,N_18731);
and U19241 (N_19241,N_18640,N_18619);
xor U19242 (N_19242,N_18654,N_18813);
xor U19243 (N_19243,N_18660,N_18749);
and U19244 (N_19244,N_18907,N_18529);
and U19245 (N_19245,N_18914,N_18696);
and U19246 (N_19246,N_18969,N_18903);
and U19247 (N_19247,N_18786,N_18714);
nand U19248 (N_19248,N_18783,N_18842);
and U19249 (N_19249,N_18835,N_18771);
xnor U19250 (N_19250,N_18554,N_18585);
nor U19251 (N_19251,N_18854,N_18518);
or U19252 (N_19252,N_18945,N_18811);
nand U19253 (N_19253,N_18795,N_18692);
nand U19254 (N_19254,N_18744,N_18882);
and U19255 (N_19255,N_18988,N_18690);
or U19256 (N_19256,N_18632,N_18930);
nor U19257 (N_19257,N_18653,N_18619);
nand U19258 (N_19258,N_18993,N_18810);
xor U19259 (N_19259,N_18955,N_18506);
nand U19260 (N_19260,N_18686,N_18572);
xor U19261 (N_19261,N_18820,N_18949);
and U19262 (N_19262,N_18689,N_18671);
and U19263 (N_19263,N_18654,N_18851);
nand U19264 (N_19264,N_18632,N_18543);
or U19265 (N_19265,N_18688,N_18705);
xor U19266 (N_19266,N_18546,N_18630);
nor U19267 (N_19267,N_18748,N_18728);
or U19268 (N_19268,N_18955,N_18954);
or U19269 (N_19269,N_18555,N_18793);
nand U19270 (N_19270,N_18512,N_18608);
nand U19271 (N_19271,N_18690,N_18711);
nand U19272 (N_19272,N_18523,N_18970);
and U19273 (N_19273,N_18679,N_18718);
nand U19274 (N_19274,N_18565,N_18599);
and U19275 (N_19275,N_18996,N_18973);
and U19276 (N_19276,N_18954,N_18613);
or U19277 (N_19277,N_18617,N_18958);
or U19278 (N_19278,N_18619,N_18870);
nand U19279 (N_19279,N_18754,N_18627);
nand U19280 (N_19280,N_18592,N_18631);
or U19281 (N_19281,N_18888,N_18686);
or U19282 (N_19282,N_18645,N_18546);
xnor U19283 (N_19283,N_18845,N_18948);
nand U19284 (N_19284,N_18574,N_18674);
nor U19285 (N_19285,N_18941,N_18903);
xor U19286 (N_19286,N_18898,N_18657);
nand U19287 (N_19287,N_18967,N_18640);
nor U19288 (N_19288,N_18667,N_18561);
xnor U19289 (N_19289,N_18958,N_18605);
and U19290 (N_19290,N_18582,N_18776);
nor U19291 (N_19291,N_18656,N_18876);
nand U19292 (N_19292,N_18824,N_18565);
nand U19293 (N_19293,N_18677,N_18798);
nor U19294 (N_19294,N_18980,N_18719);
xor U19295 (N_19295,N_18693,N_18958);
nor U19296 (N_19296,N_18596,N_18871);
xor U19297 (N_19297,N_18850,N_18835);
or U19298 (N_19298,N_18678,N_18844);
nand U19299 (N_19299,N_18990,N_18677);
and U19300 (N_19300,N_18724,N_18650);
nand U19301 (N_19301,N_18911,N_18683);
nand U19302 (N_19302,N_18860,N_18727);
nand U19303 (N_19303,N_18811,N_18744);
and U19304 (N_19304,N_18968,N_18956);
xor U19305 (N_19305,N_18596,N_18725);
xnor U19306 (N_19306,N_18705,N_18891);
xor U19307 (N_19307,N_18646,N_18618);
xor U19308 (N_19308,N_18641,N_18741);
xnor U19309 (N_19309,N_18991,N_18914);
and U19310 (N_19310,N_18581,N_18744);
or U19311 (N_19311,N_18965,N_18678);
or U19312 (N_19312,N_18696,N_18786);
xor U19313 (N_19313,N_18780,N_18534);
nand U19314 (N_19314,N_18813,N_18993);
xor U19315 (N_19315,N_18511,N_18761);
xor U19316 (N_19316,N_18875,N_18839);
nor U19317 (N_19317,N_18986,N_18866);
or U19318 (N_19318,N_18743,N_18510);
or U19319 (N_19319,N_18515,N_18747);
nand U19320 (N_19320,N_18627,N_18614);
or U19321 (N_19321,N_18552,N_18794);
xor U19322 (N_19322,N_18760,N_18792);
and U19323 (N_19323,N_18881,N_18590);
nand U19324 (N_19324,N_18540,N_18781);
nor U19325 (N_19325,N_18958,N_18724);
nor U19326 (N_19326,N_18744,N_18617);
and U19327 (N_19327,N_18975,N_18774);
nand U19328 (N_19328,N_18548,N_18816);
and U19329 (N_19329,N_18890,N_18643);
xor U19330 (N_19330,N_18807,N_18924);
xor U19331 (N_19331,N_18710,N_18598);
nor U19332 (N_19332,N_18886,N_18717);
xnor U19333 (N_19333,N_18529,N_18879);
nand U19334 (N_19334,N_18852,N_18800);
nand U19335 (N_19335,N_18852,N_18669);
or U19336 (N_19336,N_18804,N_18695);
xnor U19337 (N_19337,N_18555,N_18866);
or U19338 (N_19338,N_18513,N_18690);
and U19339 (N_19339,N_18923,N_18940);
nor U19340 (N_19340,N_18999,N_18820);
or U19341 (N_19341,N_18755,N_18663);
xnor U19342 (N_19342,N_18660,N_18706);
nand U19343 (N_19343,N_18603,N_18778);
xor U19344 (N_19344,N_18632,N_18980);
nor U19345 (N_19345,N_18650,N_18940);
or U19346 (N_19346,N_18741,N_18867);
nand U19347 (N_19347,N_18661,N_18503);
or U19348 (N_19348,N_18536,N_18701);
xnor U19349 (N_19349,N_18512,N_18780);
nand U19350 (N_19350,N_18885,N_18502);
or U19351 (N_19351,N_18569,N_18701);
nor U19352 (N_19352,N_18846,N_18501);
xnor U19353 (N_19353,N_18601,N_18839);
or U19354 (N_19354,N_18727,N_18814);
nand U19355 (N_19355,N_18651,N_18970);
and U19356 (N_19356,N_18503,N_18612);
nand U19357 (N_19357,N_18826,N_18534);
nor U19358 (N_19358,N_18700,N_18733);
xnor U19359 (N_19359,N_18837,N_18746);
or U19360 (N_19360,N_18910,N_18854);
or U19361 (N_19361,N_18962,N_18652);
nor U19362 (N_19362,N_18630,N_18981);
xnor U19363 (N_19363,N_18952,N_18808);
xor U19364 (N_19364,N_18654,N_18959);
nand U19365 (N_19365,N_18946,N_18967);
xnor U19366 (N_19366,N_18546,N_18789);
xnor U19367 (N_19367,N_18639,N_18780);
nor U19368 (N_19368,N_18597,N_18894);
nand U19369 (N_19369,N_18867,N_18510);
nor U19370 (N_19370,N_18894,N_18906);
nor U19371 (N_19371,N_18971,N_18614);
xor U19372 (N_19372,N_18881,N_18561);
xor U19373 (N_19373,N_18969,N_18997);
and U19374 (N_19374,N_18999,N_18573);
and U19375 (N_19375,N_18646,N_18601);
and U19376 (N_19376,N_18596,N_18616);
xor U19377 (N_19377,N_18679,N_18658);
nand U19378 (N_19378,N_18659,N_18862);
nor U19379 (N_19379,N_18818,N_18733);
nand U19380 (N_19380,N_18943,N_18793);
or U19381 (N_19381,N_18523,N_18900);
xor U19382 (N_19382,N_18953,N_18800);
xnor U19383 (N_19383,N_18989,N_18605);
nand U19384 (N_19384,N_18580,N_18645);
xor U19385 (N_19385,N_18923,N_18844);
xnor U19386 (N_19386,N_18947,N_18716);
nor U19387 (N_19387,N_18526,N_18688);
or U19388 (N_19388,N_18889,N_18669);
nor U19389 (N_19389,N_18788,N_18653);
nand U19390 (N_19390,N_18554,N_18679);
or U19391 (N_19391,N_18613,N_18937);
nand U19392 (N_19392,N_18779,N_18795);
or U19393 (N_19393,N_18966,N_18665);
xor U19394 (N_19394,N_18693,N_18857);
or U19395 (N_19395,N_18754,N_18875);
or U19396 (N_19396,N_18570,N_18739);
nor U19397 (N_19397,N_18671,N_18595);
nand U19398 (N_19398,N_18599,N_18834);
and U19399 (N_19399,N_18731,N_18648);
xnor U19400 (N_19400,N_18784,N_18708);
xnor U19401 (N_19401,N_18532,N_18736);
and U19402 (N_19402,N_18850,N_18971);
nor U19403 (N_19403,N_18649,N_18779);
xnor U19404 (N_19404,N_18866,N_18826);
xnor U19405 (N_19405,N_18714,N_18925);
and U19406 (N_19406,N_18732,N_18646);
nor U19407 (N_19407,N_18745,N_18719);
nor U19408 (N_19408,N_18554,N_18670);
xnor U19409 (N_19409,N_18704,N_18596);
and U19410 (N_19410,N_18531,N_18878);
and U19411 (N_19411,N_18876,N_18914);
or U19412 (N_19412,N_18590,N_18665);
or U19413 (N_19413,N_18900,N_18783);
nor U19414 (N_19414,N_18737,N_18616);
nor U19415 (N_19415,N_18954,N_18980);
or U19416 (N_19416,N_18769,N_18939);
nand U19417 (N_19417,N_18947,N_18983);
xnor U19418 (N_19418,N_18971,N_18598);
or U19419 (N_19419,N_18734,N_18579);
xnor U19420 (N_19420,N_18992,N_18868);
xor U19421 (N_19421,N_18997,N_18803);
nor U19422 (N_19422,N_18579,N_18687);
or U19423 (N_19423,N_18778,N_18994);
nand U19424 (N_19424,N_18639,N_18606);
nand U19425 (N_19425,N_18801,N_18767);
or U19426 (N_19426,N_18827,N_18514);
nand U19427 (N_19427,N_18619,N_18710);
nand U19428 (N_19428,N_18712,N_18682);
xnor U19429 (N_19429,N_18912,N_18756);
nand U19430 (N_19430,N_18911,N_18749);
or U19431 (N_19431,N_18599,N_18601);
and U19432 (N_19432,N_18794,N_18836);
xnor U19433 (N_19433,N_18564,N_18925);
xnor U19434 (N_19434,N_18770,N_18637);
and U19435 (N_19435,N_18827,N_18993);
xnor U19436 (N_19436,N_18717,N_18545);
nor U19437 (N_19437,N_18846,N_18545);
xor U19438 (N_19438,N_18823,N_18754);
nor U19439 (N_19439,N_18828,N_18892);
or U19440 (N_19440,N_18552,N_18742);
and U19441 (N_19441,N_18880,N_18578);
and U19442 (N_19442,N_18685,N_18701);
nand U19443 (N_19443,N_18563,N_18777);
xor U19444 (N_19444,N_18821,N_18503);
nand U19445 (N_19445,N_18926,N_18717);
nor U19446 (N_19446,N_18578,N_18576);
and U19447 (N_19447,N_18796,N_18710);
and U19448 (N_19448,N_18754,N_18554);
and U19449 (N_19449,N_18507,N_18965);
xor U19450 (N_19450,N_18502,N_18994);
nor U19451 (N_19451,N_18516,N_18928);
or U19452 (N_19452,N_18602,N_18631);
xor U19453 (N_19453,N_18534,N_18719);
xnor U19454 (N_19454,N_18817,N_18531);
and U19455 (N_19455,N_18869,N_18516);
xnor U19456 (N_19456,N_18546,N_18634);
xor U19457 (N_19457,N_18972,N_18621);
nor U19458 (N_19458,N_18994,N_18763);
nor U19459 (N_19459,N_18811,N_18813);
nand U19460 (N_19460,N_18570,N_18562);
nand U19461 (N_19461,N_18947,N_18636);
xnor U19462 (N_19462,N_18687,N_18500);
or U19463 (N_19463,N_18682,N_18561);
nor U19464 (N_19464,N_18918,N_18742);
nor U19465 (N_19465,N_18534,N_18813);
or U19466 (N_19466,N_18688,N_18676);
or U19467 (N_19467,N_18508,N_18648);
xor U19468 (N_19468,N_18630,N_18834);
xor U19469 (N_19469,N_18654,N_18590);
nand U19470 (N_19470,N_18633,N_18838);
xnor U19471 (N_19471,N_18500,N_18931);
nor U19472 (N_19472,N_18699,N_18545);
xor U19473 (N_19473,N_18779,N_18532);
or U19474 (N_19474,N_18929,N_18966);
xor U19475 (N_19475,N_18848,N_18992);
xor U19476 (N_19476,N_18542,N_18927);
nand U19477 (N_19477,N_18993,N_18513);
or U19478 (N_19478,N_18932,N_18583);
xnor U19479 (N_19479,N_18711,N_18579);
xnor U19480 (N_19480,N_18509,N_18737);
nand U19481 (N_19481,N_18630,N_18536);
xnor U19482 (N_19482,N_18914,N_18724);
and U19483 (N_19483,N_18942,N_18668);
nor U19484 (N_19484,N_18780,N_18835);
or U19485 (N_19485,N_18651,N_18893);
and U19486 (N_19486,N_18926,N_18509);
nor U19487 (N_19487,N_18809,N_18665);
nand U19488 (N_19488,N_18762,N_18670);
and U19489 (N_19489,N_18637,N_18788);
nand U19490 (N_19490,N_18880,N_18634);
and U19491 (N_19491,N_18803,N_18873);
xor U19492 (N_19492,N_18630,N_18991);
xor U19493 (N_19493,N_18641,N_18866);
nand U19494 (N_19494,N_18749,N_18872);
and U19495 (N_19495,N_18822,N_18869);
and U19496 (N_19496,N_18710,N_18827);
nor U19497 (N_19497,N_18951,N_18577);
and U19498 (N_19498,N_18696,N_18769);
or U19499 (N_19499,N_18929,N_18796);
nor U19500 (N_19500,N_19263,N_19027);
nor U19501 (N_19501,N_19240,N_19399);
xnor U19502 (N_19502,N_19129,N_19260);
or U19503 (N_19503,N_19214,N_19119);
or U19504 (N_19504,N_19287,N_19018);
and U19505 (N_19505,N_19438,N_19433);
xor U19506 (N_19506,N_19203,N_19123);
and U19507 (N_19507,N_19396,N_19460);
nand U19508 (N_19508,N_19454,N_19485);
nor U19509 (N_19509,N_19209,N_19207);
nor U19510 (N_19510,N_19335,N_19418);
nand U19511 (N_19511,N_19405,N_19345);
xor U19512 (N_19512,N_19417,N_19033);
xnor U19513 (N_19513,N_19217,N_19420);
or U19514 (N_19514,N_19053,N_19140);
or U19515 (N_19515,N_19308,N_19486);
and U19516 (N_19516,N_19480,N_19302);
or U19517 (N_19517,N_19491,N_19012);
nor U19518 (N_19518,N_19303,N_19450);
xnor U19519 (N_19519,N_19011,N_19488);
and U19520 (N_19520,N_19430,N_19205);
xnor U19521 (N_19521,N_19296,N_19178);
xor U19522 (N_19522,N_19333,N_19259);
xor U19523 (N_19523,N_19111,N_19481);
and U19524 (N_19524,N_19092,N_19061);
nor U19525 (N_19525,N_19023,N_19139);
nand U19526 (N_19526,N_19134,N_19466);
and U19527 (N_19527,N_19472,N_19327);
nand U19528 (N_19528,N_19367,N_19187);
and U19529 (N_19529,N_19400,N_19414);
nor U19530 (N_19530,N_19162,N_19191);
nand U19531 (N_19531,N_19198,N_19342);
and U19532 (N_19532,N_19106,N_19483);
xor U19533 (N_19533,N_19247,N_19250);
nor U19534 (N_19534,N_19320,N_19306);
nor U19535 (N_19535,N_19297,N_19397);
xnor U19536 (N_19536,N_19494,N_19238);
and U19537 (N_19537,N_19182,N_19300);
nand U19538 (N_19538,N_19341,N_19143);
and U19539 (N_19539,N_19257,N_19120);
and U19540 (N_19540,N_19432,N_19457);
nor U19541 (N_19541,N_19468,N_19368);
nor U19542 (N_19542,N_19299,N_19069);
and U19543 (N_19543,N_19019,N_19274);
or U19544 (N_19544,N_19422,N_19099);
and U19545 (N_19545,N_19394,N_19065);
nand U19546 (N_19546,N_19177,N_19313);
or U19547 (N_19547,N_19455,N_19412);
or U19548 (N_19548,N_19153,N_19361);
or U19549 (N_19549,N_19116,N_19073);
nand U19550 (N_19550,N_19163,N_19040);
nor U19551 (N_19551,N_19358,N_19426);
or U19552 (N_19552,N_19445,N_19141);
and U19553 (N_19553,N_19072,N_19464);
xnor U19554 (N_19554,N_19431,N_19379);
or U19555 (N_19555,N_19050,N_19314);
and U19556 (N_19556,N_19088,N_19102);
nor U19557 (N_19557,N_19015,N_19301);
nand U19558 (N_19558,N_19444,N_19046);
nor U19559 (N_19559,N_19070,N_19309);
nor U19560 (N_19560,N_19463,N_19210);
nor U19561 (N_19561,N_19315,N_19227);
or U19562 (N_19562,N_19490,N_19125);
and U19563 (N_19563,N_19117,N_19068);
or U19564 (N_19564,N_19272,N_19062);
and U19565 (N_19565,N_19336,N_19453);
nor U19566 (N_19566,N_19470,N_19326);
or U19567 (N_19567,N_19028,N_19035);
nor U19568 (N_19568,N_19077,N_19363);
or U19569 (N_19569,N_19482,N_19475);
and U19570 (N_19570,N_19183,N_19293);
or U19571 (N_19571,N_19271,N_19378);
or U19572 (N_19572,N_19041,N_19280);
xor U19573 (N_19573,N_19221,N_19126);
xnor U19574 (N_19574,N_19108,N_19498);
or U19575 (N_19575,N_19132,N_19168);
and U19576 (N_19576,N_19038,N_19044);
xor U19577 (N_19577,N_19144,N_19366);
xnor U19578 (N_19578,N_19478,N_19093);
and U19579 (N_19579,N_19419,N_19042);
or U19580 (N_19580,N_19157,N_19246);
or U19581 (N_19581,N_19305,N_19310);
or U19582 (N_19582,N_19404,N_19265);
xor U19583 (N_19583,N_19356,N_19376);
xnor U19584 (N_19584,N_19415,N_19323);
and U19585 (N_19585,N_19359,N_19014);
and U19586 (N_19586,N_19135,N_19186);
or U19587 (N_19587,N_19322,N_19152);
nor U19588 (N_19588,N_19115,N_19109);
or U19589 (N_19589,N_19442,N_19121);
or U19590 (N_19590,N_19059,N_19031);
and U19591 (N_19591,N_19022,N_19000);
and U19592 (N_19592,N_19085,N_19286);
nand U19593 (N_19593,N_19087,N_19131);
nor U19594 (N_19594,N_19461,N_19383);
nand U19595 (N_19595,N_19262,N_19202);
and U19596 (N_19596,N_19146,N_19372);
nand U19597 (N_19597,N_19278,N_19055);
and U19598 (N_19598,N_19057,N_19136);
nor U19599 (N_19599,N_19094,N_19199);
and U19600 (N_19600,N_19413,N_19312);
xnor U19601 (N_19601,N_19304,N_19288);
and U19602 (N_19602,N_19337,N_19197);
and U19603 (N_19603,N_19452,N_19316);
nor U19604 (N_19604,N_19066,N_19446);
xor U19605 (N_19605,N_19078,N_19492);
and U19606 (N_19606,N_19175,N_19155);
nor U19607 (N_19607,N_19034,N_19266);
nor U19608 (N_19608,N_19231,N_19456);
xor U19609 (N_19609,N_19007,N_19317);
nand U19610 (N_19610,N_19357,N_19017);
or U19611 (N_19611,N_19392,N_19244);
and U19612 (N_19612,N_19101,N_19098);
xnor U19613 (N_19613,N_19024,N_19346);
and U19614 (N_19614,N_19324,N_19104);
and U19615 (N_19615,N_19295,N_19159);
nand U19616 (N_19616,N_19393,N_19484);
nand U19617 (N_19617,N_19332,N_19100);
and U19618 (N_19618,N_19499,N_19124);
nand U19619 (N_19619,N_19473,N_19084);
nor U19620 (N_19620,N_19190,N_19355);
and U19621 (N_19621,N_19167,N_19200);
and U19622 (N_19622,N_19234,N_19381);
xor U19623 (N_19623,N_19292,N_19459);
and U19624 (N_19624,N_19462,N_19060);
xor U19625 (N_19625,N_19429,N_19439);
nor U19626 (N_19626,N_19003,N_19273);
and U19627 (N_19627,N_19147,N_19074);
and U19628 (N_19628,N_19403,N_19290);
or U19629 (N_19629,N_19387,N_19275);
xor U19630 (N_19630,N_19171,N_19281);
and U19631 (N_19631,N_19476,N_19174);
and U19632 (N_19632,N_19408,N_19172);
nor U19633 (N_19633,N_19370,N_19064);
and U19634 (N_19634,N_19496,N_19477);
nand U19635 (N_19635,N_19267,N_19213);
and U19636 (N_19636,N_19090,N_19165);
or U19637 (N_19637,N_19170,N_19364);
nand U19638 (N_19638,N_19201,N_19375);
nor U19639 (N_19639,N_19307,N_19402);
nand U19640 (N_19640,N_19192,N_19122);
nor U19641 (N_19641,N_19369,N_19344);
nand U19642 (N_19642,N_19043,N_19401);
nor U19643 (N_19643,N_19130,N_19242);
nor U19644 (N_19644,N_19254,N_19321);
and U19645 (N_19645,N_19371,N_19052);
nor U19646 (N_19646,N_19193,N_19021);
and U19647 (N_19647,N_19268,N_19009);
nand U19648 (N_19648,N_19164,N_19425);
nand U19649 (N_19649,N_19283,N_19264);
xnor U19650 (N_19650,N_19339,N_19091);
xnor U19651 (N_19651,N_19349,N_19330);
and U19652 (N_19652,N_19020,N_19360);
and U19653 (N_19653,N_19113,N_19056);
nand U19654 (N_19654,N_19239,N_19252);
nand U19655 (N_19655,N_19215,N_19421);
nor U19656 (N_19656,N_19142,N_19185);
nor U19657 (N_19657,N_19105,N_19351);
or U19658 (N_19658,N_19071,N_19443);
nor U19659 (N_19659,N_19008,N_19235);
and U19660 (N_19660,N_19365,N_19289);
xnor U19661 (N_19661,N_19347,N_19237);
nor U19662 (N_19662,N_19277,N_19045);
or U19663 (N_19663,N_19410,N_19243);
and U19664 (N_19664,N_19225,N_19435);
and U19665 (N_19665,N_19352,N_19270);
nand U19666 (N_19666,N_19127,N_19229);
nor U19667 (N_19667,N_19424,N_19382);
and U19668 (N_19668,N_19437,N_19228);
nand U19669 (N_19669,N_19013,N_19169);
or U19670 (N_19670,N_19005,N_19158);
or U19671 (N_19671,N_19386,N_19016);
or U19672 (N_19672,N_19373,N_19075);
nor U19673 (N_19673,N_19469,N_19039);
xor U19674 (N_19674,N_19082,N_19407);
or U19675 (N_19675,N_19318,N_19493);
xnor U19676 (N_19676,N_19331,N_19047);
and U19677 (N_19677,N_19001,N_19282);
nand U19678 (N_19678,N_19248,N_19095);
nand U19679 (N_19679,N_19233,N_19416);
xor U19680 (N_19680,N_19118,N_19133);
xor U19681 (N_19681,N_19110,N_19002);
nand U19682 (N_19682,N_19440,N_19058);
and U19683 (N_19683,N_19223,N_19096);
and U19684 (N_19684,N_19030,N_19334);
xnor U19685 (N_19685,N_19436,N_19226);
xnor U19686 (N_19686,N_19465,N_19049);
and U19687 (N_19687,N_19026,N_19241);
or U19688 (N_19688,N_19189,N_19184);
or U19689 (N_19689,N_19195,N_19089);
or U19690 (N_19690,N_19103,N_19329);
or U19691 (N_19691,N_19353,N_19249);
nand U19692 (N_19692,N_19441,N_19427);
or U19693 (N_19693,N_19285,N_19145);
or U19694 (N_19694,N_19173,N_19385);
xnor U19695 (N_19695,N_19208,N_19284);
nand U19696 (N_19696,N_19220,N_19294);
nor U19697 (N_19697,N_19390,N_19256);
nand U19698 (N_19698,N_19048,N_19398);
xor U19699 (N_19699,N_19154,N_19389);
nand U19700 (N_19700,N_19374,N_19114);
xor U19701 (N_19701,N_19449,N_19251);
nand U19702 (N_19702,N_19380,N_19311);
nand U19703 (N_19703,N_19279,N_19325);
nor U19704 (N_19704,N_19362,N_19343);
nand U19705 (N_19705,N_19086,N_19388);
or U19706 (N_19706,N_19276,N_19076);
and U19707 (N_19707,N_19479,N_19204);
nor U19708 (N_19708,N_19206,N_19338);
and U19709 (N_19709,N_19236,N_19148);
xor U19710 (N_19710,N_19032,N_19212);
or U19711 (N_19711,N_19406,N_19149);
nand U19712 (N_19712,N_19224,N_19261);
or U19713 (N_19713,N_19188,N_19253);
nor U19714 (N_19714,N_19151,N_19150);
nor U19715 (N_19715,N_19471,N_19218);
and U19716 (N_19716,N_19451,N_19211);
or U19717 (N_19717,N_19010,N_19161);
and U19718 (N_19718,N_19298,N_19409);
xor U19719 (N_19719,N_19128,N_19447);
nor U19720 (N_19720,N_19029,N_19348);
xor U19721 (N_19721,N_19328,N_19181);
and U19722 (N_19722,N_19051,N_19230);
xor U19723 (N_19723,N_19081,N_19222);
xnor U19724 (N_19724,N_19216,N_19340);
nand U19725 (N_19725,N_19395,N_19025);
xnor U19726 (N_19726,N_19080,N_19156);
nor U19727 (N_19727,N_19107,N_19160);
or U19728 (N_19728,N_19434,N_19423);
nand U19729 (N_19729,N_19350,N_19219);
nand U19730 (N_19730,N_19487,N_19319);
or U19731 (N_19731,N_19377,N_19079);
nand U19732 (N_19732,N_19269,N_19138);
and U19733 (N_19733,N_19037,N_19054);
nand U19734 (N_19734,N_19006,N_19194);
or U19735 (N_19735,N_19196,N_19428);
and U19736 (N_19736,N_19258,N_19384);
xnor U19737 (N_19737,N_19291,N_19474);
and U19738 (N_19738,N_19255,N_19391);
xnor U19739 (N_19739,N_19448,N_19176);
nor U19740 (N_19740,N_19467,N_19489);
nor U19741 (N_19741,N_19067,N_19411);
or U19742 (N_19742,N_19004,N_19245);
or U19743 (N_19743,N_19112,N_19137);
xor U19744 (N_19744,N_19497,N_19097);
xor U19745 (N_19745,N_19083,N_19180);
xnor U19746 (N_19746,N_19495,N_19063);
xnor U19747 (N_19747,N_19458,N_19354);
nand U19748 (N_19748,N_19232,N_19166);
nor U19749 (N_19749,N_19036,N_19179);
xnor U19750 (N_19750,N_19493,N_19006);
xnor U19751 (N_19751,N_19003,N_19385);
or U19752 (N_19752,N_19342,N_19266);
or U19753 (N_19753,N_19343,N_19467);
nor U19754 (N_19754,N_19199,N_19411);
or U19755 (N_19755,N_19416,N_19344);
xor U19756 (N_19756,N_19190,N_19014);
xnor U19757 (N_19757,N_19060,N_19030);
xnor U19758 (N_19758,N_19338,N_19427);
nand U19759 (N_19759,N_19421,N_19352);
nor U19760 (N_19760,N_19403,N_19032);
nor U19761 (N_19761,N_19188,N_19477);
or U19762 (N_19762,N_19013,N_19116);
xnor U19763 (N_19763,N_19432,N_19395);
nor U19764 (N_19764,N_19422,N_19335);
nand U19765 (N_19765,N_19037,N_19060);
and U19766 (N_19766,N_19279,N_19400);
nand U19767 (N_19767,N_19027,N_19191);
nand U19768 (N_19768,N_19180,N_19061);
nand U19769 (N_19769,N_19409,N_19423);
and U19770 (N_19770,N_19122,N_19372);
xnor U19771 (N_19771,N_19178,N_19139);
and U19772 (N_19772,N_19487,N_19351);
and U19773 (N_19773,N_19232,N_19230);
nor U19774 (N_19774,N_19202,N_19354);
xnor U19775 (N_19775,N_19030,N_19245);
nand U19776 (N_19776,N_19498,N_19340);
nand U19777 (N_19777,N_19194,N_19200);
and U19778 (N_19778,N_19006,N_19009);
nand U19779 (N_19779,N_19204,N_19354);
nand U19780 (N_19780,N_19111,N_19410);
nor U19781 (N_19781,N_19091,N_19329);
nor U19782 (N_19782,N_19136,N_19126);
or U19783 (N_19783,N_19424,N_19047);
xnor U19784 (N_19784,N_19264,N_19463);
nor U19785 (N_19785,N_19130,N_19284);
and U19786 (N_19786,N_19117,N_19013);
xnor U19787 (N_19787,N_19472,N_19457);
or U19788 (N_19788,N_19197,N_19258);
nand U19789 (N_19789,N_19343,N_19295);
nor U19790 (N_19790,N_19051,N_19346);
and U19791 (N_19791,N_19245,N_19329);
or U19792 (N_19792,N_19078,N_19183);
or U19793 (N_19793,N_19466,N_19399);
nand U19794 (N_19794,N_19143,N_19270);
and U19795 (N_19795,N_19209,N_19462);
nand U19796 (N_19796,N_19004,N_19438);
xor U19797 (N_19797,N_19132,N_19209);
xor U19798 (N_19798,N_19205,N_19283);
xor U19799 (N_19799,N_19409,N_19156);
and U19800 (N_19800,N_19207,N_19130);
or U19801 (N_19801,N_19318,N_19481);
and U19802 (N_19802,N_19495,N_19376);
xnor U19803 (N_19803,N_19332,N_19236);
and U19804 (N_19804,N_19363,N_19424);
nor U19805 (N_19805,N_19340,N_19177);
and U19806 (N_19806,N_19398,N_19244);
xnor U19807 (N_19807,N_19435,N_19001);
nor U19808 (N_19808,N_19270,N_19489);
nand U19809 (N_19809,N_19130,N_19076);
xnor U19810 (N_19810,N_19392,N_19406);
nand U19811 (N_19811,N_19429,N_19361);
nand U19812 (N_19812,N_19013,N_19407);
nand U19813 (N_19813,N_19132,N_19017);
nor U19814 (N_19814,N_19088,N_19358);
and U19815 (N_19815,N_19499,N_19279);
nand U19816 (N_19816,N_19337,N_19452);
and U19817 (N_19817,N_19195,N_19339);
or U19818 (N_19818,N_19276,N_19188);
or U19819 (N_19819,N_19258,N_19347);
xor U19820 (N_19820,N_19274,N_19182);
or U19821 (N_19821,N_19445,N_19178);
nand U19822 (N_19822,N_19097,N_19465);
nand U19823 (N_19823,N_19100,N_19349);
nor U19824 (N_19824,N_19014,N_19128);
nor U19825 (N_19825,N_19013,N_19071);
xnor U19826 (N_19826,N_19320,N_19287);
xnor U19827 (N_19827,N_19322,N_19188);
or U19828 (N_19828,N_19314,N_19110);
xor U19829 (N_19829,N_19331,N_19166);
and U19830 (N_19830,N_19341,N_19343);
nand U19831 (N_19831,N_19402,N_19442);
xor U19832 (N_19832,N_19224,N_19375);
nor U19833 (N_19833,N_19234,N_19314);
or U19834 (N_19834,N_19234,N_19200);
and U19835 (N_19835,N_19188,N_19492);
nor U19836 (N_19836,N_19410,N_19095);
nor U19837 (N_19837,N_19161,N_19173);
nand U19838 (N_19838,N_19449,N_19428);
nand U19839 (N_19839,N_19037,N_19091);
and U19840 (N_19840,N_19261,N_19169);
xor U19841 (N_19841,N_19450,N_19143);
or U19842 (N_19842,N_19117,N_19280);
and U19843 (N_19843,N_19276,N_19118);
nand U19844 (N_19844,N_19244,N_19097);
nor U19845 (N_19845,N_19440,N_19110);
and U19846 (N_19846,N_19169,N_19342);
nand U19847 (N_19847,N_19225,N_19325);
xor U19848 (N_19848,N_19126,N_19148);
xor U19849 (N_19849,N_19249,N_19216);
nand U19850 (N_19850,N_19202,N_19249);
and U19851 (N_19851,N_19439,N_19492);
nand U19852 (N_19852,N_19309,N_19123);
and U19853 (N_19853,N_19190,N_19224);
nand U19854 (N_19854,N_19130,N_19092);
and U19855 (N_19855,N_19149,N_19073);
xnor U19856 (N_19856,N_19079,N_19014);
xor U19857 (N_19857,N_19393,N_19071);
xnor U19858 (N_19858,N_19121,N_19167);
and U19859 (N_19859,N_19387,N_19413);
xnor U19860 (N_19860,N_19205,N_19471);
or U19861 (N_19861,N_19281,N_19208);
nand U19862 (N_19862,N_19240,N_19396);
nand U19863 (N_19863,N_19323,N_19244);
xnor U19864 (N_19864,N_19494,N_19354);
or U19865 (N_19865,N_19128,N_19053);
or U19866 (N_19866,N_19476,N_19306);
and U19867 (N_19867,N_19322,N_19345);
and U19868 (N_19868,N_19152,N_19014);
nor U19869 (N_19869,N_19464,N_19358);
nor U19870 (N_19870,N_19393,N_19133);
nand U19871 (N_19871,N_19429,N_19049);
nor U19872 (N_19872,N_19241,N_19161);
or U19873 (N_19873,N_19322,N_19165);
nor U19874 (N_19874,N_19098,N_19048);
and U19875 (N_19875,N_19031,N_19000);
nor U19876 (N_19876,N_19387,N_19283);
nor U19877 (N_19877,N_19490,N_19135);
or U19878 (N_19878,N_19057,N_19344);
nor U19879 (N_19879,N_19113,N_19317);
nand U19880 (N_19880,N_19402,N_19453);
nand U19881 (N_19881,N_19174,N_19044);
and U19882 (N_19882,N_19297,N_19360);
and U19883 (N_19883,N_19392,N_19479);
or U19884 (N_19884,N_19301,N_19041);
and U19885 (N_19885,N_19147,N_19261);
xnor U19886 (N_19886,N_19276,N_19146);
nor U19887 (N_19887,N_19320,N_19227);
or U19888 (N_19888,N_19354,N_19356);
or U19889 (N_19889,N_19475,N_19108);
xor U19890 (N_19890,N_19494,N_19345);
nor U19891 (N_19891,N_19470,N_19431);
and U19892 (N_19892,N_19388,N_19273);
or U19893 (N_19893,N_19375,N_19037);
or U19894 (N_19894,N_19191,N_19111);
xnor U19895 (N_19895,N_19196,N_19271);
and U19896 (N_19896,N_19383,N_19470);
xnor U19897 (N_19897,N_19400,N_19116);
xor U19898 (N_19898,N_19285,N_19470);
nor U19899 (N_19899,N_19067,N_19480);
and U19900 (N_19900,N_19020,N_19246);
nand U19901 (N_19901,N_19480,N_19466);
nand U19902 (N_19902,N_19479,N_19186);
nand U19903 (N_19903,N_19131,N_19096);
nor U19904 (N_19904,N_19463,N_19496);
nor U19905 (N_19905,N_19344,N_19361);
or U19906 (N_19906,N_19474,N_19085);
nand U19907 (N_19907,N_19059,N_19010);
nor U19908 (N_19908,N_19248,N_19328);
xor U19909 (N_19909,N_19122,N_19280);
and U19910 (N_19910,N_19253,N_19160);
or U19911 (N_19911,N_19258,N_19312);
xor U19912 (N_19912,N_19402,N_19139);
nand U19913 (N_19913,N_19232,N_19047);
xnor U19914 (N_19914,N_19406,N_19360);
and U19915 (N_19915,N_19226,N_19353);
or U19916 (N_19916,N_19198,N_19197);
and U19917 (N_19917,N_19182,N_19483);
and U19918 (N_19918,N_19407,N_19400);
nor U19919 (N_19919,N_19410,N_19440);
or U19920 (N_19920,N_19021,N_19115);
or U19921 (N_19921,N_19089,N_19344);
nor U19922 (N_19922,N_19454,N_19046);
nor U19923 (N_19923,N_19428,N_19330);
xor U19924 (N_19924,N_19031,N_19116);
and U19925 (N_19925,N_19083,N_19039);
or U19926 (N_19926,N_19169,N_19135);
and U19927 (N_19927,N_19053,N_19496);
and U19928 (N_19928,N_19222,N_19402);
and U19929 (N_19929,N_19062,N_19085);
and U19930 (N_19930,N_19268,N_19330);
xor U19931 (N_19931,N_19476,N_19197);
or U19932 (N_19932,N_19021,N_19078);
nand U19933 (N_19933,N_19441,N_19175);
nor U19934 (N_19934,N_19448,N_19211);
and U19935 (N_19935,N_19061,N_19449);
nor U19936 (N_19936,N_19130,N_19426);
nor U19937 (N_19937,N_19344,N_19373);
nand U19938 (N_19938,N_19474,N_19068);
or U19939 (N_19939,N_19241,N_19081);
and U19940 (N_19940,N_19232,N_19060);
nor U19941 (N_19941,N_19271,N_19434);
xnor U19942 (N_19942,N_19119,N_19000);
nor U19943 (N_19943,N_19018,N_19222);
nand U19944 (N_19944,N_19239,N_19194);
nand U19945 (N_19945,N_19109,N_19401);
xor U19946 (N_19946,N_19042,N_19190);
or U19947 (N_19947,N_19123,N_19375);
nand U19948 (N_19948,N_19201,N_19141);
nand U19949 (N_19949,N_19458,N_19469);
xnor U19950 (N_19950,N_19098,N_19045);
nand U19951 (N_19951,N_19156,N_19002);
nand U19952 (N_19952,N_19489,N_19420);
nand U19953 (N_19953,N_19209,N_19115);
xnor U19954 (N_19954,N_19360,N_19023);
xnor U19955 (N_19955,N_19132,N_19035);
or U19956 (N_19956,N_19461,N_19230);
nor U19957 (N_19957,N_19485,N_19481);
nand U19958 (N_19958,N_19418,N_19278);
nand U19959 (N_19959,N_19062,N_19353);
xor U19960 (N_19960,N_19371,N_19280);
nand U19961 (N_19961,N_19427,N_19214);
and U19962 (N_19962,N_19169,N_19003);
and U19963 (N_19963,N_19243,N_19399);
nor U19964 (N_19964,N_19454,N_19474);
and U19965 (N_19965,N_19358,N_19055);
nand U19966 (N_19966,N_19202,N_19415);
or U19967 (N_19967,N_19283,N_19474);
nand U19968 (N_19968,N_19274,N_19327);
and U19969 (N_19969,N_19428,N_19154);
or U19970 (N_19970,N_19225,N_19141);
xnor U19971 (N_19971,N_19494,N_19179);
nand U19972 (N_19972,N_19231,N_19006);
or U19973 (N_19973,N_19465,N_19214);
nor U19974 (N_19974,N_19032,N_19271);
xor U19975 (N_19975,N_19095,N_19380);
and U19976 (N_19976,N_19208,N_19115);
and U19977 (N_19977,N_19415,N_19055);
or U19978 (N_19978,N_19446,N_19401);
and U19979 (N_19979,N_19170,N_19428);
xor U19980 (N_19980,N_19248,N_19393);
and U19981 (N_19981,N_19414,N_19252);
nand U19982 (N_19982,N_19167,N_19395);
nand U19983 (N_19983,N_19040,N_19007);
and U19984 (N_19984,N_19484,N_19276);
nor U19985 (N_19985,N_19029,N_19096);
nor U19986 (N_19986,N_19180,N_19106);
nor U19987 (N_19987,N_19273,N_19349);
and U19988 (N_19988,N_19102,N_19421);
xor U19989 (N_19989,N_19365,N_19069);
nand U19990 (N_19990,N_19005,N_19177);
or U19991 (N_19991,N_19065,N_19461);
and U19992 (N_19992,N_19030,N_19100);
xnor U19993 (N_19993,N_19252,N_19167);
nand U19994 (N_19994,N_19162,N_19195);
and U19995 (N_19995,N_19433,N_19208);
nand U19996 (N_19996,N_19493,N_19168);
nor U19997 (N_19997,N_19389,N_19252);
xnor U19998 (N_19998,N_19387,N_19224);
or U19999 (N_19999,N_19199,N_19075);
and UO_0 (O_0,N_19702,N_19801);
xor UO_1 (O_1,N_19617,N_19689);
or UO_2 (O_2,N_19934,N_19872);
and UO_3 (O_3,N_19746,N_19862);
nor UO_4 (O_4,N_19873,N_19697);
and UO_5 (O_5,N_19879,N_19928);
and UO_6 (O_6,N_19667,N_19940);
nor UO_7 (O_7,N_19803,N_19683);
and UO_8 (O_8,N_19882,N_19728);
nor UO_9 (O_9,N_19500,N_19608);
or UO_10 (O_10,N_19751,N_19810);
or UO_11 (O_11,N_19591,N_19826);
nand UO_12 (O_12,N_19626,N_19755);
or UO_13 (O_13,N_19527,N_19551);
nand UO_14 (O_14,N_19630,N_19641);
xor UO_15 (O_15,N_19696,N_19650);
nand UO_16 (O_16,N_19831,N_19548);
nor UO_17 (O_17,N_19596,N_19605);
nand UO_18 (O_18,N_19804,N_19656);
nand UO_19 (O_19,N_19578,N_19681);
xor UO_20 (O_20,N_19682,N_19999);
and UO_21 (O_21,N_19526,N_19558);
or UO_22 (O_22,N_19542,N_19592);
and UO_23 (O_23,N_19902,N_19890);
or UO_24 (O_24,N_19530,N_19645);
xnor UO_25 (O_25,N_19658,N_19983);
and UO_26 (O_26,N_19567,N_19936);
or UO_27 (O_27,N_19508,N_19564);
or UO_28 (O_28,N_19986,N_19788);
nand UO_29 (O_29,N_19834,N_19783);
nand UO_30 (O_30,N_19708,N_19501);
nor UO_31 (O_31,N_19997,N_19993);
or UO_32 (O_32,N_19620,N_19917);
xnor UO_33 (O_33,N_19741,N_19833);
nor UO_34 (O_34,N_19857,N_19970);
or UO_35 (O_35,N_19758,N_19868);
xor UO_36 (O_36,N_19623,N_19759);
xor UO_37 (O_37,N_19737,N_19557);
and UO_38 (O_38,N_19972,N_19732);
xor UO_39 (O_39,N_19524,N_19780);
nand UO_40 (O_40,N_19733,N_19984);
nor UO_41 (O_41,N_19808,N_19739);
or UO_42 (O_42,N_19786,N_19622);
or UO_43 (O_43,N_19865,N_19633);
xor UO_44 (O_44,N_19646,N_19600);
and UO_45 (O_45,N_19721,N_19980);
nor UO_46 (O_46,N_19824,N_19680);
nor UO_47 (O_47,N_19653,N_19504);
nand UO_48 (O_48,N_19580,N_19976);
or UO_49 (O_49,N_19760,N_19821);
nor UO_50 (O_50,N_19669,N_19877);
xor UO_51 (O_51,N_19919,N_19540);
or UO_52 (O_52,N_19965,N_19503);
nor UO_53 (O_53,N_19543,N_19654);
xnor UO_54 (O_54,N_19866,N_19714);
xor UO_55 (O_55,N_19718,N_19762);
and UO_56 (O_56,N_19546,N_19581);
nand UO_57 (O_57,N_19687,N_19560);
and UO_58 (O_58,N_19561,N_19756);
or UO_59 (O_59,N_19719,N_19609);
or UO_60 (O_60,N_19966,N_19793);
xor UO_61 (O_61,N_19789,N_19675);
nor UO_62 (O_62,N_19555,N_19914);
xnor UO_63 (O_63,N_19659,N_19853);
xnor UO_64 (O_64,N_19878,N_19674);
nand UO_65 (O_65,N_19782,N_19898);
or UO_66 (O_66,N_19943,N_19693);
nand UO_67 (O_67,N_19601,N_19948);
xor UO_68 (O_68,N_19937,N_19846);
nand UO_69 (O_69,N_19973,N_19598);
and UO_70 (O_70,N_19664,N_19707);
and UO_71 (O_71,N_19894,N_19790);
nand UO_72 (O_72,N_19992,N_19875);
nor UO_73 (O_73,N_19812,N_19842);
nor UO_74 (O_74,N_19807,N_19671);
nor UO_75 (O_75,N_19761,N_19549);
nor UO_76 (O_76,N_19507,N_19797);
or UO_77 (O_77,N_19825,N_19946);
nand UO_78 (O_78,N_19676,N_19638);
nor UO_79 (O_79,N_19534,N_19796);
nor UO_80 (O_80,N_19896,N_19847);
nand UO_81 (O_81,N_19864,N_19811);
and UO_82 (O_82,N_19515,N_19985);
nor UO_83 (O_83,N_19536,N_19805);
xor UO_84 (O_84,N_19647,N_19722);
nor UO_85 (O_85,N_19691,N_19749);
nand UO_86 (O_86,N_19962,N_19899);
xor UO_87 (O_87,N_19539,N_19860);
nor UO_88 (O_88,N_19684,N_19705);
xnor UO_89 (O_89,N_19514,N_19552);
and UO_90 (O_90,N_19566,N_19660);
nand UO_91 (O_91,N_19665,N_19517);
or UO_92 (O_92,N_19951,N_19883);
and UO_93 (O_93,N_19744,N_19612);
xor UO_94 (O_94,N_19969,N_19963);
xor UO_95 (O_95,N_19513,N_19640);
or UO_96 (O_96,N_19672,N_19520);
xor UO_97 (O_97,N_19794,N_19925);
nand UO_98 (O_98,N_19938,N_19795);
and UO_99 (O_99,N_19677,N_19624);
nand UO_100 (O_100,N_19798,N_19785);
or UO_101 (O_101,N_19979,N_19929);
or UO_102 (O_102,N_19909,N_19799);
nor UO_103 (O_103,N_19932,N_19611);
nand UO_104 (O_104,N_19800,N_19767);
nand UO_105 (O_105,N_19629,N_19613);
or UO_106 (O_106,N_19974,N_19852);
nand UO_107 (O_107,N_19886,N_19918);
and UO_108 (O_108,N_19631,N_19518);
nor UO_109 (O_109,N_19636,N_19690);
nand UO_110 (O_110,N_19784,N_19774);
or UO_111 (O_111,N_19961,N_19933);
nand UO_112 (O_112,N_19582,N_19519);
and UO_113 (O_113,N_19634,N_19643);
nand UO_114 (O_114,N_19856,N_19547);
or UO_115 (O_115,N_19982,N_19945);
or UO_116 (O_116,N_19935,N_19829);
and UO_117 (O_117,N_19678,N_19532);
nand UO_118 (O_118,N_19571,N_19538);
nor UO_119 (O_119,N_19977,N_19625);
nand UO_120 (O_120,N_19791,N_19991);
nand UO_121 (O_121,N_19509,N_19729);
and UO_122 (O_122,N_19603,N_19569);
nand UO_123 (O_123,N_19688,N_19610);
or UO_124 (O_124,N_19848,N_19743);
nand UO_125 (O_125,N_19648,N_19736);
and UO_126 (O_126,N_19816,N_19698);
or UO_127 (O_127,N_19731,N_19738);
xnor UO_128 (O_128,N_19644,N_19818);
or UO_129 (O_129,N_19924,N_19740);
and UO_130 (O_130,N_19770,N_19900);
nor UO_131 (O_131,N_19942,N_19837);
nand UO_132 (O_132,N_19576,N_19577);
and UO_133 (O_133,N_19944,N_19891);
nand UO_134 (O_134,N_19850,N_19832);
and UO_135 (O_135,N_19709,N_19892);
nor UO_136 (O_136,N_19628,N_19779);
nor UO_137 (O_137,N_19615,N_19716);
nand UO_138 (O_138,N_19787,N_19817);
and UO_139 (O_139,N_19655,N_19606);
nand UO_140 (O_140,N_19927,N_19544);
and UO_141 (O_141,N_19637,N_19968);
or UO_142 (O_142,N_19754,N_19588);
nor UO_143 (O_143,N_19642,N_19957);
xnor UO_144 (O_144,N_19627,N_19712);
or UO_145 (O_145,N_19960,N_19911);
nand UO_146 (O_146,N_19747,N_19828);
or UO_147 (O_147,N_19954,N_19996);
nor UO_148 (O_148,N_19981,N_19988);
or UO_149 (O_149,N_19735,N_19750);
nor UO_150 (O_150,N_19823,N_19521);
nand UO_151 (O_151,N_19859,N_19913);
nand UO_152 (O_152,N_19772,N_19745);
nand UO_153 (O_153,N_19904,N_19710);
or UO_154 (O_154,N_19512,N_19584);
and UO_155 (O_155,N_19769,N_19621);
nor UO_156 (O_156,N_19533,N_19727);
or UO_157 (O_157,N_19777,N_19773);
or UO_158 (O_158,N_19563,N_19679);
nand UO_159 (O_159,N_19916,N_19956);
nor UO_160 (O_160,N_19673,N_19836);
xnor UO_161 (O_161,N_19931,N_19553);
nand UO_162 (O_162,N_19947,N_19704);
xnor UO_163 (O_163,N_19887,N_19851);
nor UO_164 (O_164,N_19863,N_19867);
or UO_165 (O_165,N_19595,N_19967);
xor UO_166 (O_166,N_19742,N_19895);
or UO_167 (O_167,N_19830,N_19923);
nor UO_168 (O_168,N_19941,N_19858);
and UO_169 (O_169,N_19870,N_19775);
nor UO_170 (O_170,N_19910,N_19994);
nor UO_171 (O_171,N_19670,N_19550);
or UO_172 (O_172,N_19599,N_19713);
nand UO_173 (O_173,N_19989,N_19706);
nor UO_174 (O_174,N_19881,N_19570);
xor UO_175 (O_175,N_19901,N_19562);
nor UO_176 (O_176,N_19725,N_19871);
nor UO_177 (O_177,N_19978,N_19995);
nand UO_178 (O_178,N_19531,N_19661);
and UO_179 (O_179,N_19699,N_19586);
nand UO_180 (O_180,N_19903,N_19845);
xor UO_181 (O_181,N_19921,N_19639);
or UO_182 (O_182,N_19651,N_19556);
xor UO_183 (O_183,N_19594,N_19619);
nand UO_184 (O_184,N_19694,N_19559);
nor UO_185 (O_185,N_19700,N_19579);
nand UO_186 (O_186,N_19666,N_19815);
or UO_187 (O_187,N_19939,N_19545);
xor UO_188 (O_188,N_19930,N_19876);
nand UO_189 (O_189,N_19583,N_19955);
or UO_190 (O_190,N_19516,N_19975);
xnor UO_191 (O_191,N_19802,N_19987);
nand UO_192 (O_192,N_19915,N_19502);
nor UO_193 (O_193,N_19964,N_19575);
nand UO_194 (O_194,N_19888,N_19568);
or UO_195 (O_195,N_19781,N_19734);
xor UO_196 (O_196,N_19726,N_19505);
nor UO_197 (O_197,N_19602,N_19776);
nor UO_198 (O_198,N_19572,N_19953);
and UO_199 (O_199,N_19908,N_19748);
or UO_200 (O_200,N_19528,N_19841);
nand UO_201 (O_201,N_19529,N_19885);
and UO_202 (O_202,N_19510,N_19554);
nor UO_203 (O_203,N_19587,N_19950);
or UO_204 (O_204,N_19537,N_19616);
and UO_205 (O_205,N_19685,N_19843);
xor UO_206 (O_206,N_19912,N_19695);
nand UO_207 (O_207,N_19854,N_19668);
and UO_208 (O_208,N_19792,N_19778);
nor UO_209 (O_209,N_19839,N_19663);
nor UO_210 (O_210,N_19765,N_19607);
xnor UO_211 (O_211,N_19590,N_19764);
and UO_212 (O_212,N_19724,N_19565);
xor UO_213 (O_213,N_19771,N_19893);
or UO_214 (O_214,N_19753,N_19880);
xnor UO_215 (O_215,N_19813,N_19819);
nand UO_216 (O_216,N_19525,N_19589);
or UO_217 (O_217,N_19597,N_19766);
nor UO_218 (O_218,N_19827,N_19998);
xnor UO_219 (O_219,N_19952,N_19506);
xor UO_220 (O_220,N_19897,N_19715);
nand UO_221 (O_221,N_19861,N_19686);
and UO_222 (O_222,N_19822,N_19585);
and UO_223 (O_223,N_19593,N_19523);
nand UO_224 (O_224,N_19717,N_19949);
and UO_225 (O_225,N_19535,N_19752);
xnor UO_226 (O_226,N_19768,N_19662);
xor UO_227 (O_227,N_19926,N_19869);
xnor UO_228 (O_228,N_19763,N_19840);
nand UO_229 (O_229,N_19838,N_19905);
nand UO_230 (O_230,N_19632,N_19959);
nor UO_231 (O_231,N_19844,N_19958);
nor UO_232 (O_232,N_19806,N_19884);
xnor UO_233 (O_233,N_19820,N_19723);
or UO_234 (O_234,N_19906,N_19990);
nand UO_235 (O_235,N_19855,N_19920);
or UO_236 (O_236,N_19573,N_19835);
xnor UO_237 (O_237,N_19614,N_19720);
nor UO_238 (O_238,N_19874,N_19511);
nand UO_239 (O_239,N_19889,N_19757);
nand UO_240 (O_240,N_19649,N_19907);
and UO_241 (O_241,N_19730,N_19809);
xor UO_242 (O_242,N_19703,N_19701);
and UO_243 (O_243,N_19574,N_19692);
nand UO_244 (O_244,N_19604,N_19635);
nand UO_245 (O_245,N_19522,N_19618);
nor UO_246 (O_246,N_19849,N_19541);
nand UO_247 (O_247,N_19657,N_19922);
nor UO_248 (O_248,N_19971,N_19814);
and UO_249 (O_249,N_19652,N_19711);
or UO_250 (O_250,N_19928,N_19598);
or UO_251 (O_251,N_19631,N_19629);
nand UO_252 (O_252,N_19729,N_19546);
and UO_253 (O_253,N_19904,N_19758);
and UO_254 (O_254,N_19698,N_19900);
xor UO_255 (O_255,N_19687,N_19569);
nand UO_256 (O_256,N_19953,N_19792);
or UO_257 (O_257,N_19570,N_19818);
or UO_258 (O_258,N_19619,N_19628);
nor UO_259 (O_259,N_19708,N_19874);
nor UO_260 (O_260,N_19723,N_19831);
and UO_261 (O_261,N_19956,N_19814);
xnor UO_262 (O_262,N_19629,N_19846);
xor UO_263 (O_263,N_19840,N_19543);
xnor UO_264 (O_264,N_19831,N_19799);
and UO_265 (O_265,N_19529,N_19610);
xnor UO_266 (O_266,N_19919,N_19743);
nor UO_267 (O_267,N_19984,N_19972);
nor UO_268 (O_268,N_19634,N_19859);
or UO_269 (O_269,N_19621,N_19682);
and UO_270 (O_270,N_19938,N_19617);
xnor UO_271 (O_271,N_19851,N_19867);
and UO_272 (O_272,N_19717,N_19534);
or UO_273 (O_273,N_19629,N_19601);
nor UO_274 (O_274,N_19572,N_19853);
nand UO_275 (O_275,N_19766,N_19829);
or UO_276 (O_276,N_19815,N_19898);
and UO_277 (O_277,N_19923,N_19722);
and UO_278 (O_278,N_19894,N_19639);
and UO_279 (O_279,N_19993,N_19543);
nor UO_280 (O_280,N_19775,N_19724);
xnor UO_281 (O_281,N_19905,N_19973);
or UO_282 (O_282,N_19900,N_19651);
nor UO_283 (O_283,N_19649,N_19698);
xor UO_284 (O_284,N_19866,N_19509);
nand UO_285 (O_285,N_19884,N_19551);
nor UO_286 (O_286,N_19962,N_19618);
nand UO_287 (O_287,N_19680,N_19988);
xnor UO_288 (O_288,N_19544,N_19872);
nor UO_289 (O_289,N_19683,N_19875);
and UO_290 (O_290,N_19635,N_19529);
nand UO_291 (O_291,N_19539,N_19635);
and UO_292 (O_292,N_19874,N_19640);
xnor UO_293 (O_293,N_19585,N_19917);
nand UO_294 (O_294,N_19781,N_19887);
nand UO_295 (O_295,N_19765,N_19670);
or UO_296 (O_296,N_19752,N_19914);
xor UO_297 (O_297,N_19647,N_19745);
nand UO_298 (O_298,N_19648,N_19636);
or UO_299 (O_299,N_19895,N_19856);
or UO_300 (O_300,N_19976,N_19547);
nand UO_301 (O_301,N_19516,N_19525);
nor UO_302 (O_302,N_19501,N_19612);
nor UO_303 (O_303,N_19694,N_19659);
nor UO_304 (O_304,N_19954,N_19669);
xnor UO_305 (O_305,N_19565,N_19907);
nand UO_306 (O_306,N_19584,N_19974);
nor UO_307 (O_307,N_19979,N_19695);
and UO_308 (O_308,N_19614,N_19599);
or UO_309 (O_309,N_19837,N_19610);
nand UO_310 (O_310,N_19670,N_19517);
nand UO_311 (O_311,N_19922,N_19585);
and UO_312 (O_312,N_19594,N_19687);
and UO_313 (O_313,N_19527,N_19949);
xnor UO_314 (O_314,N_19834,N_19500);
nand UO_315 (O_315,N_19630,N_19612);
nand UO_316 (O_316,N_19550,N_19714);
xnor UO_317 (O_317,N_19708,N_19505);
xor UO_318 (O_318,N_19907,N_19940);
xor UO_319 (O_319,N_19546,N_19521);
nand UO_320 (O_320,N_19894,N_19571);
or UO_321 (O_321,N_19838,N_19794);
xor UO_322 (O_322,N_19526,N_19784);
xor UO_323 (O_323,N_19685,N_19741);
nor UO_324 (O_324,N_19893,N_19619);
nor UO_325 (O_325,N_19921,N_19579);
nor UO_326 (O_326,N_19854,N_19644);
nand UO_327 (O_327,N_19737,N_19933);
or UO_328 (O_328,N_19799,N_19688);
nand UO_329 (O_329,N_19630,N_19652);
and UO_330 (O_330,N_19993,N_19887);
or UO_331 (O_331,N_19730,N_19900);
or UO_332 (O_332,N_19779,N_19857);
xnor UO_333 (O_333,N_19658,N_19777);
nand UO_334 (O_334,N_19781,N_19812);
or UO_335 (O_335,N_19651,N_19686);
nor UO_336 (O_336,N_19873,N_19921);
and UO_337 (O_337,N_19503,N_19851);
or UO_338 (O_338,N_19752,N_19683);
and UO_339 (O_339,N_19640,N_19614);
nor UO_340 (O_340,N_19851,N_19918);
and UO_341 (O_341,N_19558,N_19998);
nor UO_342 (O_342,N_19627,N_19799);
nand UO_343 (O_343,N_19717,N_19702);
or UO_344 (O_344,N_19946,N_19922);
nor UO_345 (O_345,N_19568,N_19795);
xnor UO_346 (O_346,N_19541,N_19955);
and UO_347 (O_347,N_19804,N_19654);
nor UO_348 (O_348,N_19689,N_19961);
nor UO_349 (O_349,N_19559,N_19710);
nand UO_350 (O_350,N_19514,N_19760);
or UO_351 (O_351,N_19608,N_19782);
nor UO_352 (O_352,N_19530,N_19599);
and UO_353 (O_353,N_19689,N_19590);
or UO_354 (O_354,N_19559,N_19832);
or UO_355 (O_355,N_19975,N_19572);
nor UO_356 (O_356,N_19745,N_19901);
nor UO_357 (O_357,N_19851,N_19552);
and UO_358 (O_358,N_19934,N_19593);
and UO_359 (O_359,N_19695,N_19933);
xor UO_360 (O_360,N_19596,N_19976);
xnor UO_361 (O_361,N_19962,N_19946);
xnor UO_362 (O_362,N_19537,N_19699);
xor UO_363 (O_363,N_19802,N_19791);
or UO_364 (O_364,N_19964,N_19891);
or UO_365 (O_365,N_19836,N_19945);
nor UO_366 (O_366,N_19930,N_19897);
nor UO_367 (O_367,N_19985,N_19902);
xnor UO_368 (O_368,N_19761,N_19720);
nand UO_369 (O_369,N_19952,N_19646);
nand UO_370 (O_370,N_19883,N_19956);
and UO_371 (O_371,N_19803,N_19767);
xnor UO_372 (O_372,N_19719,N_19845);
nor UO_373 (O_373,N_19944,N_19875);
xor UO_374 (O_374,N_19580,N_19501);
nand UO_375 (O_375,N_19740,N_19963);
xnor UO_376 (O_376,N_19907,N_19601);
and UO_377 (O_377,N_19620,N_19705);
xor UO_378 (O_378,N_19656,N_19841);
or UO_379 (O_379,N_19657,N_19578);
or UO_380 (O_380,N_19621,N_19993);
nor UO_381 (O_381,N_19882,N_19960);
or UO_382 (O_382,N_19671,N_19539);
nand UO_383 (O_383,N_19809,N_19925);
xor UO_384 (O_384,N_19797,N_19876);
and UO_385 (O_385,N_19783,N_19627);
or UO_386 (O_386,N_19888,N_19932);
or UO_387 (O_387,N_19916,N_19669);
nor UO_388 (O_388,N_19739,N_19604);
nand UO_389 (O_389,N_19934,N_19996);
or UO_390 (O_390,N_19883,N_19763);
xor UO_391 (O_391,N_19977,N_19896);
xnor UO_392 (O_392,N_19964,N_19940);
xnor UO_393 (O_393,N_19777,N_19858);
nor UO_394 (O_394,N_19606,N_19522);
and UO_395 (O_395,N_19914,N_19610);
nand UO_396 (O_396,N_19770,N_19720);
nand UO_397 (O_397,N_19778,N_19714);
or UO_398 (O_398,N_19948,N_19808);
xor UO_399 (O_399,N_19960,N_19537);
nand UO_400 (O_400,N_19781,N_19565);
and UO_401 (O_401,N_19868,N_19904);
nand UO_402 (O_402,N_19753,N_19536);
or UO_403 (O_403,N_19664,N_19865);
xnor UO_404 (O_404,N_19928,N_19889);
or UO_405 (O_405,N_19796,N_19840);
or UO_406 (O_406,N_19603,N_19894);
xnor UO_407 (O_407,N_19680,N_19766);
xnor UO_408 (O_408,N_19737,N_19886);
or UO_409 (O_409,N_19711,N_19552);
and UO_410 (O_410,N_19897,N_19596);
nor UO_411 (O_411,N_19511,N_19818);
xor UO_412 (O_412,N_19795,N_19543);
nor UO_413 (O_413,N_19805,N_19931);
nor UO_414 (O_414,N_19560,N_19559);
xor UO_415 (O_415,N_19770,N_19527);
xor UO_416 (O_416,N_19511,N_19681);
and UO_417 (O_417,N_19582,N_19982);
and UO_418 (O_418,N_19970,N_19939);
or UO_419 (O_419,N_19605,N_19600);
xnor UO_420 (O_420,N_19644,N_19535);
and UO_421 (O_421,N_19751,N_19649);
or UO_422 (O_422,N_19500,N_19606);
or UO_423 (O_423,N_19587,N_19597);
and UO_424 (O_424,N_19830,N_19863);
xnor UO_425 (O_425,N_19639,N_19707);
and UO_426 (O_426,N_19777,N_19632);
nor UO_427 (O_427,N_19643,N_19629);
and UO_428 (O_428,N_19595,N_19886);
xnor UO_429 (O_429,N_19929,N_19523);
xnor UO_430 (O_430,N_19766,N_19927);
nand UO_431 (O_431,N_19966,N_19716);
nand UO_432 (O_432,N_19934,N_19680);
nand UO_433 (O_433,N_19630,N_19526);
nor UO_434 (O_434,N_19842,N_19568);
nor UO_435 (O_435,N_19935,N_19930);
xor UO_436 (O_436,N_19666,N_19682);
or UO_437 (O_437,N_19955,N_19907);
xnor UO_438 (O_438,N_19953,N_19820);
xnor UO_439 (O_439,N_19962,N_19621);
or UO_440 (O_440,N_19538,N_19879);
nand UO_441 (O_441,N_19630,N_19521);
xnor UO_442 (O_442,N_19824,N_19991);
or UO_443 (O_443,N_19873,N_19661);
xnor UO_444 (O_444,N_19635,N_19739);
and UO_445 (O_445,N_19761,N_19569);
xnor UO_446 (O_446,N_19594,N_19519);
nand UO_447 (O_447,N_19540,N_19653);
and UO_448 (O_448,N_19724,N_19979);
xnor UO_449 (O_449,N_19840,N_19679);
xnor UO_450 (O_450,N_19743,N_19999);
nand UO_451 (O_451,N_19770,N_19890);
xnor UO_452 (O_452,N_19599,N_19603);
or UO_453 (O_453,N_19505,N_19503);
or UO_454 (O_454,N_19801,N_19761);
or UO_455 (O_455,N_19616,N_19626);
or UO_456 (O_456,N_19830,N_19507);
nand UO_457 (O_457,N_19860,N_19766);
xor UO_458 (O_458,N_19863,N_19622);
nand UO_459 (O_459,N_19565,N_19562);
xor UO_460 (O_460,N_19510,N_19529);
xor UO_461 (O_461,N_19769,N_19608);
xor UO_462 (O_462,N_19728,N_19501);
nand UO_463 (O_463,N_19752,N_19892);
or UO_464 (O_464,N_19566,N_19833);
and UO_465 (O_465,N_19771,N_19909);
and UO_466 (O_466,N_19869,N_19606);
nand UO_467 (O_467,N_19950,N_19653);
and UO_468 (O_468,N_19635,N_19979);
nor UO_469 (O_469,N_19913,N_19980);
and UO_470 (O_470,N_19870,N_19882);
and UO_471 (O_471,N_19689,N_19621);
xnor UO_472 (O_472,N_19844,N_19777);
and UO_473 (O_473,N_19800,N_19717);
or UO_474 (O_474,N_19535,N_19552);
and UO_475 (O_475,N_19573,N_19960);
xor UO_476 (O_476,N_19943,N_19851);
or UO_477 (O_477,N_19548,N_19979);
and UO_478 (O_478,N_19527,N_19855);
and UO_479 (O_479,N_19790,N_19548);
or UO_480 (O_480,N_19674,N_19755);
or UO_481 (O_481,N_19534,N_19711);
nand UO_482 (O_482,N_19585,N_19823);
nor UO_483 (O_483,N_19524,N_19963);
xor UO_484 (O_484,N_19841,N_19650);
xnor UO_485 (O_485,N_19643,N_19874);
or UO_486 (O_486,N_19888,N_19837);
nor UO_487 (O_487,N_19523,N_19957);
nand UO_488 (O_488,N_19792,N_19969);
nand UO_489 (O_489,N_19990,N_19959);
nand UO_490 (O_490,N_19930,N_19917);
nand UO_491 (O_491,N_19607,N_19557);
or UO_492 (O_492,N_19760,N_19956);
xnor UO_493 (O_493,N_19651,N_19949);
nand UO_494 (O_494,N_19743,N_19651);
xor UO_495 (O_495,N_19850,N_19931);
or UO_496 (O_496,N_19554,N_19514);
nand UO_497 (O_497,N_19995,N_19793);
or UO_498 (O_498,N_19584,N_19852);
xnor UO_499 (O_499,N_19549,N_19779);
nor UO_500 (O_500,N_19680,N_19687);
nor UO_501 (O_501,N_19800,N_19855);
and UO_502 (O_502,N_19519,N_19577);
xnor UO_503 (O_503,N_19917,N_19937);
nor UO_504 (O_504,N_19629,N_19801);
nand UO_505 (O_505,N_19786,N_19866);
nand UO_506 (O_506,N_19978,N_19852);
and UO_507 (O_507,N_19862,N_19946);
or UO_508 (O_508,N_19759,N_19987);
xor UO_509 (O_509,N_19764,N_19513);
xor UO_510 (O_510,N_19502,N_19763);
and UO_511 (O_511,N_19540,N_19575);
or UO_512 (O_512,N_19704,N_19624);
xnor UO_513 (O_513,N_19757,N_19600);
nand UO_514 (O_514,N_19548,N_19969);
nand UO_515 (O_515,N_19726,N_19749);
and UO_516 (O_516,N_19997,N_19798);
xor UO_517 (O_517,N_19900,N_19857);
nand UO_518 (O_518,N_19836,N_19695);
nor UO_519 (O_519,N_19897,N_19581);
nand UO_520 (O_520,N_19856,N_19985);
xnor UO_521 (O_521,N_19641,N_19551);
nand UO_522 (O_522,N_19968,N_19959);
or UO_523 (O_523,N_19573,N_19726);
xor UO_524 (O_524,N_19578,N_19859);
nor UO_525 (O_525,N_19720,N_19782);
and UO_526 (O_526,N_19680,N_19679);
xnor UO_527 (O_527,N_19552,N_19822);
or UO_528 (O_528,N_19623,N_19674);
nor UO_529 (O_529,N_19821,N_19542);
or UO_530 (O_530,N_19818,N_19604);
and UO_531 (O_531,N_19521,N_19561);
xor UO_532 (O_532,N_19669,N_19721);
nor UO_533 (O_533,N_19586,N_19925);
xnor UO_534 (O_534,N_19523,N_19948);
or UO_535 (O_535,N_19676,N_19672);
xnor UO_536 (O_536,N_19804,N_19990);
nand UO_537 (O_537,N_19964,N_19905);
nand UO_538 (O_538,N_19835,N_19720);
nor UO_539 (O_539,N_19694,N_19817);
and UO_540 (O_540,N_19705,N_19667);
xnor UO_541 (O_541,N_19873,N_19885);
or UO_542 (O_542,N_19983,N_19731);
nand UO_543 (O_543,N_19798,N_19612);
nor UO_544 (O_544,N_19833,N_19726);
xnor UO_545 (O_545,N_19691,N_19592);
or UO_546 (O_546,N_19922,N_19790);
xor UO_547 (O_547,N_19678,N_19595);
and UO_548 (O_548,N_19778,N_19632);
xnor UO_549 (O_549,N_19961,N_19789);
xor UO_550 (O_550,N_19805,N_19901);
or UO_551 (O_551,N_19602,N_19889);
nand UO_552 (O_552,N_19675,N_19828);
or UO_553 (O_553,N_19531,N_19757);
and UO_554 (O_554,N_19638,N_19691);
nor UO_555 (O_555,N_19785,N_19996);
nand UO_556 (O_556,N_19568,N_19510);
or UO_557 (O_557,N_19650,N_19878);
xnor UO_558 (O_558,N_19736,N_19546);
nor UO_559 (O_559,N_19687,N_19954);
and UO_560 (O_560,N_19856,N_19646);
nor UO_561 (O_561,N_19810,N_19584);
nand UO_562 (O_562,N_19961,N_19920);
nand UO_563 (O_563,N_19859,N_19515);
nand UO_564 (O_564,N_19556,N_19924);
nand UO_565 (O_565,N_19730,N_19532);
nor UO_566 (O_566,N_19511,N_19899);
or UO_567 (O_567,N_19512,N_19612);
or UO_568 (O_568,N_19864,N_19701);
and UO_569 (O_569,N_19571,N_19521);
and UO_570 (O_570,N_19651,N_19588);
nand UO_571 (O_571,N_19729,N_19995);
or UO_572 (O_572,N_19510,N_19546);
nor UO_573 (O_573,N_19813,N_19834);
nor UO_574 (O_574,N_19604,N_19675);
nand UO_575 (O_575,N_19772,N_19524);
nand UO_576 (O_576,N_19820,N_19893);
or UO_577 (O_577,N_19781,N_19558);
xnor UO_578 (O_578,N_19895,N_19947);
and UO_579 (O_579,N_19562,N_19585);
and UO_580 (O_580,N_19559,N_19665);
and UO_581 (O_581,N_19570,N_19583);
and UO_582 (O_582,N_19500,N_19716);
or UO_583 (O_583,N_19708,N_19585);
nand UO_584 (O_584,N_19631,N_19707);
and UO_585 (O_585,N_19885,N_19759);
nand UO_586 (O_586,N_19663,N_19830);
nor UO_587 (O_587,N_19602,N_19728);
or UO_588 (O_588,N_19536,N_19942);
and UO_589 (O_589,N_19535,N_19961);
xor UO_590 (O_590,N_19765,N_19929);
nor UO_591 (O_591,N_19996,N_19824);
nand UO_592 (O_592,N_19923,N_19856);
nand UO_593 (O_593,N_19664,N_19567);
or UO_594 (O_594,N_19789,N_19699);
xnor UO_595 (O_595,N_19549,N_19694);
nor UO_596 (O_596,N_19575,N_19946);
nor UO_597 (O_597,N_19875,N_19730);
xnor UO_598 (O_598,N_19566,N_19584);
xnor UO_599 (O_599,N_19903,N_19966);
and UO_600 (O_600,N_19674,N_19865);
nor UO_601 (O_601,N_19827,N_19563);
or UO_602 (O_602,N_19760,N_19604);
or UO_603 (O_603,N_19947,N_19740);
nand UO_604 (O_604,N_19883,N_19851);
or UO_605 (O_605,N_19902,N_19825);
nand UO_606 (O_606,N_19910,N_19546);
xor UO_607 (O_607,N_19687,N_19608);
xnor UO_608 (O_608,N_19912,N_19502);
nor UO_609 (O_609,N_19523,N_19915);
or UO_610 (O_610,N_19513,N_19692);
or UO_611 (O_611,N_19904,N_19703);
xnor UO_612 (O_612,N_19553,N_19932);
and UO_613 (O_613,N_19771,N_19868);
and UO_614 (O_614,N_19534,N_19680);
nand UO_615 (O_615,N_19669,N_19554);
and UO_616 (O_616,N_19753,N_19500);
nor UO_617 (O_617,N_19719,N_19962);
nor UO_618 (O_618,N_19966,N_19827);
and UO_619 (O_619,N_19879,N_19746);
nand UO_620 (O_620,N_19726,N_19834);
nand UO_621 (O_621,N_19572,N_19538);
nor UO_622 (O_622,N_19909,N_19544);
xnor UO_623 (O_623,N_19697,N_19925);
nor UO_624 (O_624,N_19878,N_19761);
nand UO_625 (O_625,N_19614,N_19813);
nor UO_626 (O_626,N_19782,N_19838);
xnor UO_627 (O_627,N_19683,N_19691);
nor UO_628 (O_628,N_19974,N_19860);
nand UO_629 (O_629,N_19753,N_19905);
or UO_630 (O_630,N_19856,N_19568);
xor UO_631 (O_631,N_19934,N_19542);
or UO_632 (O_632,N_19951,N_19913);
and UO_633 (O_633,N_19523,N_19933);
nand UO_634 (O_634,N_19678,N_19567);
or UO_635 (O_635,N_19819,N_19784);
and UO_636 (O_636,N_19564,N_19595);
nand UO_637 (O_637,N_19596,N_19786);
or UO_638 (O_638,N_19714,N_19711);
nor UO_639 (O_639,N_19783,N_19970);
nand UO_640 (O_640,N_19659,N_19523);
xor UO_641 (O_641,N_19650,N_19772);
nand UO_642 (O_642,N_19712,N_19634);
and UO_643 (O_643,N_19767,N_19839);
or UO_644 (O_644,N_19733,N_19957);
nor UO_645 (O_645,N_19858,N_19808);
and UO_646 (O_646,N_19914,N_19834);
and UO_647 (O_647,N_19907,N_19791);
and UO_648 (O_648,N_19880,N_19689);
or UO_649 (O_649,N_19585,N_19858);
nand UO_650 (O_650,N_19909,N_19542);
xnor UO_651 (O_651,N_19603,N_19537);
nand UO_652 (O_652,N_19775,N_19940);
nor UO_653 (O_653,N_19667,N_19859);
and UO_654 (O_654,N_19648,N_19626);
xor UO_655 (O_655,N_19899,N_19742);
or UO_656 (O_656,N_19997,N_19703);
nor UO_657 (O_657,N_19891,N_19952);
nand UO_658 (O_658,N_19585,N_19819);
nor UO_659 (O_659,N_19690,N_19872);
nor UO_660 (O_660,N_19735,N_19654);
xnor UO_661 (O_661,N_19799,N_19716);
nor UO_662 (O_662,N_19554,N_19731);
nand UO_663 (O_663,N_19695,N_19892);
nor UO_664 (O_664,N_19995,N_19750);
nand UO_665 (O_665,N_19972,N_19813);
nor UO_666 (O_666,N_19867,N_19720);
xnor UO_667 (O_667,N_19946,N_19733);
nand UO_668 (O_668,N_19570,N_19510);
nor UO_669 (O_669,N_19638,N_19855);
nor UO_670 (O_670,N_19512,N_19930);
xnor UO_671 (O_671,N_19576,N_19956);
nand UO_672 (O_672,N_19874,N_19552);
or UO_673 (O_673,N_19504,N_19865);
nor UO_674 (O_674,N_19514,N_19800);
nand UO_675 (O_675,N_19683,N_19556);
or UO_676 (O_676,N_19948,N_19859);
or UO_677 (O_677,N_19532,N_19921);
or UO_678 (O_678,N_19714,N_19638);
and UO_679 (O_679,N_19743,N_19952);
nand UO_680 (O_680,N_19622,N_19744);
xnor UO_681 (O_681,N_19972,N_19956);
nor UO_682 (O_682,N_19509,N_19734);
or UO_683 (O_683,N_19936,N_19959);
xnor UO_684 (O_684,N_19600,N_19545);
and UO_685 (O_685,N_19941,N_19979);
and UO_686 (O_686,N_19700,N_19959);
nand UO_687 (O_687,N_19896,N_19996);
xor UO_688 (O_688,N_19798,N_19835);
xnor UO_689 (O_689,N_19748,N_19608);
and UO_690 (O_690,N_19846,N_19762);
nor UO_691 (O_691,N_19649,N_19686);
nor UO_692 (O_692,N_19933,N_19570);
nor UO_693 (O_693,N_19509,N_19673);
xnor UO_694 (O_694,N_19880,N_19929);
nor UO_695 (O_695,N_19535,N_19651);
xor UO_696 (O_696,N_19633,N_19771);
and UO_697 (O_697,N_19720,N_19563);
and UO_698 (O_698,N_19537,N_19503);
and UO_699 (O_699,N_19739,N_19999);
and UO_700 (O_700,N_19620,N_19791);
nand UO_701 (O_701,N_19550,N_19655);
and UO_702 (O_702,N_19570,N_19663);
nand UO_703 (O_703,N_19968,N_19522);
nand UO_704 (O_704,N_19870,N_19891);
nor UO_705 (O_705,N_19841,N_19598);
or UO_706 (O_706,N_19580,N_19943);
nand UO_707 (O_707,N_19609,N_19880);
and UO_708 (O_708,N_19943,N_19608);
nand UO_709 (O_709,N_19836,N_19782);
nor UO_710 (O_710,N_19629,N_19818);
xnor UO_711 (O_711,N_19761,N_19512);
or UO_712 (O_712,N_19529,N_19777);
nor UO_713 (O_713,N_19912,N_19590);
and UO_714 (O_714,N_19873,N_19817);
and UO_715 (O_715,N_19591,N_19620);
and UO_716 (O_716,N_19933,N_19917);
xnor UO_717 (O_717,N_19752,N_19515);
or UO_718 (O_718,N_19581,N_19849);
or UO_719 (O_719,N_19657,N_19557);
nor UO_720 (O_720,N_19518,N_19663);
and UO_721 (O_721,N_19966,N_19942);
nand UO_722 (O_722,N_19955,N_19789);
nor UO_723 (O_723,N_19905,N_19749);
xnor UO_724 (O_724,N_19719,N_19620);
nor UO_725 (O_725,N_19998,N_19668);
or UO_726 (O_726,N_19505,N_19713);
xnor UO_727 (O_727,N_19951,N_19755);
nor UO_728 (O_728,N_19944,N_19791);
xnor UO_729 (O_729,N_19818,N_19936);
and UO_730 (O_730,N_19640,N_19601);
nor UO_731 (O_731,N_19842,N_19612);
and UO_732 (O_732,N_19935,N_19552);
nand UO_733 (O_733,N_19911,N_19850);
xnor UO_734 (O_734,N_19657,N_19610);
or UO_735 (O_735,N_19824,N_19692);
and UO_736 (O_736,N_19638,N_19674);
and UO_737 (O_737,N_19742,N_19678);
nand UO_738 (O_738,N_19506,N_19755);
nand UO_739 (O_739,N_19617,N_19566);
and UO_740 (O_740,N_19764,N_19876);
and UO_741 (O_741,N_19961,N_19638);
and UO_742 (O_742,N_19759,N_19896);
nor UO_743 (O_743,N_19816,N_19997);
or UO_744 (O_744,N_19718,N_19839);
nand UO_745 (O_745,N_19961,N_19938);
or UO_746 (O_746,N_19990,N_19728);
xnor UO_747 (O_747,N_19878,N_19563);
nor UO_748 (O_748,N_19731,N_19684);
nand UO_749 (O_749,N_19590,N_19532);
and UO_750 (O_750,N_19765,N_19630);
nor UO_751 (O_751,N_19843,N_19557);
or UO_752 (O_752,N_19703,N_19568);
nand UO_753 (O_753,N_19724,N_19628);
xnor UO_754 (O_754,N_19754,N_19810);
or UO_755 (O_755,N_19739,N_19850);
nor UO_756 (O_756,N_19690,N_19739);
and UO_757 (O_757,N_19910,N_19936);
nor UO_758 (O_758,N_19805,N_19528);
and UO_759 (O_759,N_19565,N_19922);
and UO_760 (O_760,N_19981,N_19767);
and UO_761 (O_761,N_19565,N_19710);
xnor UO_762 (O_762,N_19992,N_19701);
nand UO_763 (O_763,N_19687,N_19590);
nor UO_764 (O_764,N_19760,N_19607);
and UO_765 (O_765,N_19903,N_19996);
and UO_766 (O_766,N_19721,N_19501);
nand UO_767 (O_767,N_19691,N_19601);
or UO_768 (O_768,N_19731,N_19560);
or UO_769 (O_769,N_19993,N_19756);
nor UO_770 (O_770,N_19674,N_19517);
xnor UO_771 (O_771,N_19620,N_19828);
nand UO_772 (O_772,N_19622,N_19860);
xor UO_773 (O_773,N_19759,N_19570);
nor UO_774 (O_774,N_19551,N_19804);
nand UO_775 (O_775,N_19507,N_19969);
and UO_776 (O_776,N_19557,N_19598);
nand UO_777 (O_777,N_19839,N_19745);
or UO_778 (O_778,N_19971,N_19567);
and UO_779 (O_779,N_19610,N_19732);
nor UO_780 (O_780,N_19759,N_19847);
xor UO_781 (O_781,N_19756,N_19666);
or UO_782 (O_782,N_19824,N_19594);
or UO_783 (O_783,N_19624,N_19943);
nand UO_784 (O_784,N_19710,N_19946);
nor UO_785 (O_785,N_19587,N_19833);
or UO_786 (O_786,N_19862,N_19517);
nor UO_787 (O_787,N_19602,N_19578);
or UO_788 (O_788,N_19915,N_19683);
nand UO_789 (O_789,N_19614,N_19629);
and UO_790 (O_790,N_19946,N_19753);
nor UO_791 (O_791,N_19902,N_19864);
xor UO_792 (O_792,N_19907,N_19885);
or UO_793 (O_793,N_19756,N_19514);
xnor UO_794 (O_794,N_19988,N_19796);
and UO_795 (O_795,N_19563,N_19800);
or UO_796 (O_796,N_19968,N_19759);
nor UO_797 (O_797,N_19541,N_19889);
or UO_798 (O_798,N_19982,N_19552);
nor UO_799 (O_799,N_19638,N_19963);
xnor UO_800 (O_800,N_19637,N_19806);
nor UO_801 (O_801,N_19512,N_19688);
and UO_802 (O_802,N_19952,N_19615);
or UO_803 (O_803,N_19663,N_19511);
or UO_804 (O_804,N_19924,N_19842);
and UO_805 (O_805,N_19545,N_19974);
and UO_806 (O_806,N_19669,N_19798);
nand UO_807 (O_807,N_19926,N_19501);
xor UO_808 (O_808,N_19922,N_19827);
nand UO_809 (O_809,N_19527,N_19580);
or UO_810 (O_810,N_19580,N_19599);
and UO_811 (O_811,N_19508,N_19957);
xor UO_812 (O_812,N_19956,N_19911);
and UO_813 (O_813,N_19722,N_19621);
and UO_814 (O_814,N_19635,N_19922);
and UO_815 (O_815,N_19571,N_19819);
or UO_816 (O_816,N_19672,N_19545);
and UO_817 (O_817,N_19721,N_19732);
nand UO_818 (O_818,N_19707,N_19671);
and UO_819 (O_819,N_19795,N_19709);
xnor UO_820 (O_820,N_19689,N_19915);
or UO_821 (O_821,N_19838,N_19816);
or UO_822 (O_822,N_19997,N_19846);
nand UO_823 (O_823,N_19802,N_19690);
nor UO_824 (O_824,N_19968,N_19829);
nand UO_825 (O_825,N_19500,N_19614);
or UO_826 (O_826,N_19577,N_19982);
nand UO_827 (O_827,N_19534,N_19787);
or UO_828 (O_828,N_19830,N_19724);
and UO_829 (O_829,N_19990,N_19701);
and UO_830 (O_830,N_19583,N_19778);
xnor UO_831 (O_831,N_19555,N_19619);
xnor UO_832 (O_832,N_19529,N_19854);
xnor UO_833 (O_833,N_19720,N_19671);
and UO_834 (O_834,N_19919,N_19761);
nand UO_835 (O_835,N_19761,N_19518);
xor UO_836 (O_836,N_19999,N_19584);
nor UO_837 (O_837,N_19888,N_19694);
nor UO_838 (O_838,N_19726,N_19597);
xnor UO_839 (O_839,N_19634,N_19869);
xor UO_840 (O_840,N_19990,N_19932);
nor UO_841 (O_841,N_19547,N_19632);
and UO_842 (O_842,N_19732,N_19826);
xnor UO_843 (O_843,N_19953,N_19565);
or UO_844 (O_844,N_19636,N_19903);
or UO_845 (O_845,N_19830,N_19520);
nand UO_846 (O_846,N_19599,N_19541);
and UO_847 (O_847,N_19699,N_19947);
xor UO_848 (O_848,N_19714,N_19518);
nand UO_849 (O_849,N_19808,N_19941);
nand UO_850 (O_850,N_19913,N_19648);
nor UO_851 (O_851,N_19926,N_19796);
and UO_852 (O_852,N_19672,N_19881);
xnor UO_853 (O_853,N_19514,N_19683);
or UO_854 (O_854,N_19743,N_19796);
nor UO_855 (O_855,N_19577,N_19663);
or UO_856 (O_856,N_19556,N_19846);
or UO_857 (O_857,N_19885,N_19923);
nand UO_858 (O_858,N_19754,N_19764);
nand UO_859 (O_859,N_19835,N_19993);
nor UO_860 (O_860,N_19691,N_19730);
or UO_861 (O_861,N_19904,N_19577);
nor UO_862 (O_862,N_19916,N_19920);
or UO_863 (O_863,N_19993,N_19708);
xor UO_864 (O_864,N_19848,N_19679);
nor UO_865 (O_865,N_19933,N_19688);
or UO_866 (O_866,N_19756,N_19827);
or UO_867 (O_867,N_19890,N_19819);
xor UO_868 (O_868,N_19770,N_19935);
nor UO_869 (O_869,N_19777,N_19930);
and UO_870 (O_870,N_19507,N_19940);
nor UO_871 (O_871,N_19683,N_19560);
xnor UO_872 (O_872,N_19750,N_19554);
and UO_873 (O_873,N_19600,N_19822);
xnor UO_874 (O_874,N_19697,N_19560);
nor UO_875 (O_875,N_19597,N_19684);
xnor UO_876 (O_876,N_19720,N_19860);
xnor UO_877 (O_877,N_19634,N_19912);
nand UO_878 (O_878,N_19645,N_19864);
nor UO_879 (O_879,N_19707,N_19730);
nand UO_880 (O_880,N_19853,N_19566);
and UO_881 (O_881,N_19823,N_19559);
or UO_882 (O_882,N_19828,N_19954);
or UO_883 (O_883,N_19613,N_19988);
or UO_884 (O_884,N_19726,N_19502);
or UO_885 (O_885,N_19881,N_19532);
nor UO_886 (O_886,N_19946,N_19882);
or UO_887 (O_887,N_19584,N_19642);
nand UO_888 (O_888,N_19695,N_19535);
nand UO_889 (O_889,N_19552,N_19958);
nand UO_890 (O_890,N_19861,N_19959);
xnor UO_891 (O_891,N_19503,N_19572);
and UO_892 (O_892,N_19959,N_19839);
nand UO_893 (O_893,N_19854,N_19620);
and UO_894 (O_894,N_19689,N_19813);
nor UO_895 (O_895,N_19525,N_19608);
nand UO_896 (O_896,N_19901,N_19997);
nand UO_897 (O_897,N_19748,N_19875);
or UO_898 (O_898,N_19727,N_19607);
xor UO_899 (O_899,N_19518,N_19810);
or UO_900 (O_900,N_19566,N_19777);
xnor UO_901 (O_901,N_19978,N_19879);
nor UO_902 (O_902,N_19794,N_19929);
nand UO_903 (O_903,N_19916,N_19821);
nor UO_904 (O_904,N_19830,N_19973);
nor UO_905 (O_905,N_19798,N_19972);
nor UO_906 (O_906,N_19548,N_19782);
or UO_907 (O_907,N_19700,N_19522);
nor UO_908 (O_908,N_19835,N_19816);
or UO_909 (O_909,N_19526,N_19512);
and UO_910 (O_910,N_19718,N_19672);
nand UO_911 (O_911,N_19969,N_19562);
nand UO_912 (O_912,N_19877,N_19913);
and UO_913 (O_913,N_19676,N_19512);
or UO_914 (O_914,N_19806,N_19743);
and UO_915 (O_915,N_19903,N_19847);
nor UO_916 (O_916,N_19577,N_19831);
xor UO_917 (O_917,N_19649,N_19986);
and UO_918 (O_918,N_19513,N_19660);
and UO_919 (O_919,N_19749,N_19953);
xor UO_920 (O_920,N_19915,N_19831);
nand UO_921 (O_921,N_19543,N_19905);
nand UO_922 (O_922,N_19852,N_19742);
nor UO_923 (O_923,N_19721,N_19690);
xor UO_924 (O_924,N_19600,N_19862);
xor UO_925 (O_925,N_19862,N_19646);
xor UO_926 (O_926,N_19621,N_19616);
xor UO_927 (O_927,N_19736,N_19607);
nor UO_928 (O_928,N_19873,N_19865);
xnor UO_929 (O_929,N_19848,N_19988);
xnor UO_930 (O_930,N_19923,N_19709);
nor UO_931 (O_931,N_19790,N_19736);
nand UO_932 (O_932,N_19858,N_19723);
nor UO_933 (O_933,N_19624,N_19979);
nand UO_934 (O_934,N_19884,N_19763);
nor UO_935 (O_935,N_19765,N_19987);
or UO_936 (O_936,N_19556,N_19900);
and UO_937 (O_937,N_19677,N_19920);
nand UO_938 (O_938,N_19584,N_19623);
nand UO_939 (O_939,N_19528,N_19924);
nor UO_940 (O_940,N_19536,N_19711);
and UO_941 (O_941,N_19938,N_19676);
nand UO_942 (O_942,N_19855,N_19909);
xnor UO_943 (O_943,N_19502,N_19643);
or UO_944 (O_944,N_19733,N_19830);
or UO_945 (O_945,N_19530,N_19667);
nand UO_946 (O_946,N_19897,N_19739);
or UO_947 (O_947,N_19544,N_19780);
nand UO_948 (O_948,N_19794,N_19581);
or UO_949 (O_949,N_19633,N_19590);
nand UO_950 (O_950,N_19532,N_19763);
nor UO_951 (O_951,N_19537,N_19978);
or UO_952 (O_952,N_19558,N_19614);
nand UO_953 (O_953,N_19556,N_19734);
nand UO_954 (O_954,N_19967,N_19719);
xor UO_955 (O_955,N_19568,N_19851);
nor UO_956 (O_956,N_19942,N_19748);
nand UO_957 (O_957,N_19523,N_19560);
nor UO_958 (O_958,N_19911,N_19932);
nand UO_959 (O_959,N_19600,N_19764);
nor UO_960 (O_960,N_19728,N_19918);
xnor UO_961 (O_961,N_19674,N_19696);
xor UO_962 (O_962,N_19746,N_19564);
or UO_963 (O_963,N_19504,N_19864);
and UO_964 (O_964,N_19843,N_19509);
xnor UO_965 (O_965,N_19536,N_19928);
xnor UO_966 (O_966,N_19925,N_19647);
nand UO_967 (O_967,N_19745,N_19992);
nor UO_968 (O_968,N_19932,N_19542);
or UO_969 (O_969,N_19560,N_19682);
or UO_970 (O_970,N_19967,N_19928);
xor UO_971 (O_971,N_19857,N_19712);
and UO_972 (O_972,N_19842,N_19547);
and UO_973 (O_973,N_19536,N_19692);
and UO_974 (O_974,N_19992,N_19865);
nand UO_975 (O_975,N_19560,N_19908);
or UO_976 (O_976,N_19783,N_19911);
or UO_977 (O_977,N_19575,N_19751);
nand UO_978 (O_978,N_19696,N_19752);
nor UO_979 (O_979,N_19920,N_19768);
or UO_980 (O_980,N_19893,N_19874);
xor UO_981 (O_981,N_19526,N_19886);
or UO_982 (O_982,N_19710,N_19966);
or UO_983 (O_983,N_19917,N_19656);
nor UO_984 (O_984,N_19527,N_19975);
nor UO_985 (O_985,N_19995,N_19541);
nand UO_986 (O_986,N_19908,N_19989);
or UO_987 (O_987,N_19513,N_19512);
xnor UO_988 (O_988,N_19688,N_19697);
or UO_989 (O_989,N_19602,N_19510);
or UO_990 (O_990,N_19781,N_19849);
nor UO_991 (O_991,N_19537,N_19963);
or UO_992 (O_992,N_19881,N_19595);
and UO_993 (O_993,N_19556,N_19971);
and UO_994 (O_994,N_19567,N_19690);
and UO_995 (O_995,N_19706,N_19534);
nor UO_996 (O_996,N_19818,N_19552);
or UO_997 (O_997,N_19529,N_19919);
or UO_998 (O_998,N_19858,N_19971);
and UO_999 (O_999,N_19593,N_19807);
nor UO_1000 (O_1000,N_19598,N_19845);
nand UO_1001 (O_1001,N_19815,N_19600);
nand UO_1002 (O_1002,N_19955,N_19950);
nand UO_1003 (O_1003,N_19823,N_19962);
nand UO_1004 (O_1004,N_19710,N_19979);
nand UO_1005 (O_1005,N_19976,N_19797);
nand UO_1006 (O_1006,N_19735,N_19539);
nand UO_1007 (O_1007,N_19685,N_19777);
xnor UO_1008 (O_1008,N_19927,N_19930);
and UO_1009 (O_1009,N_19914,N_19783);
nand UO_1010 (O_1010,N_19885,N_19855);
and UO_1011 (O_1011,N_19709,N_19627);
nand UO_1012 (O_1012,N_19550,N_19605);
xnor UO_1013 (O_1013,N_19616,N_19995);
xor UO_1014 (O_1014,N_19612,N_19906);
xnor UO_1015 (O_1015,N_19584,N_19593);
nand UO_1016 (O_1016,N_19934,N_19521);
xnor UO_1017 (O_1017,N_19594,N_19908);
and UO_1018 (O_1018,N_19878,N_19631);
nand UO_1019 (O_1019,N_19985,N_19923);
or UO_1020 (O_1020,N_19631,N_19935);
and UO_1021 (O_1021,N_19639,N_19718);
nor UO_1022 (O_1022,N_19731,N_19675);
nand UO_1023 (O_1023,N_19511,N_19746);
nor UO_1024 (O_1024,N_19778,N_19902);
nor UO_1025 (O_1025,N_19741,N_19708);
nand UO_1026 (O_1026,N_19866,N_19822);
xor UO_1027 (O_1027,N_19794,N_19748);
or UO_1028 (O_1028,N_19586,N_19556);
nand UO_1029 (O_1029,N_19527,N_19719);
nor UO_1030 (O_1030,N_19630,N_19911);
xor UO_1031 (O_1031,N_19645,N_19752);
nor UO_1032 (O_1032,N_19688,N_19962);
or UO_1033 (O_1033,N_19692,N_19831);
xor UO_1034 (O_1034,N_19947,N_19846);
and UO_1035 (O_1035,N_19664,N_19702);
nand UO_1036 (O_1036,N_19921,N_19512);
nor UO_1037 (O_1037,N_19597,N_19895);
or UO_1038 (O_1038,N_19631,N_19578);
xnor UO_1039 (O_1039,N_19827,N_19849);
and UO_1040 (O_1040,N_19742,N_19921);
nand UO_1041 (O_1041,N_19588,N_19973);
and UO_1042 (O_1042,N_19567,N_19638);
nand UO_1043 (O_1043,N_19943,N_19647);
nand UO_1044 (O_1044,N_19810,N_19965);
or UO_1045 (O_1045,N_19777,N_19812);
or UO_1046 (O_1046,N_19628,N_19911);
nor UO_1047 (O_1047,N_19930,N_19805);
nor UO_1048 (O_1048,N_19777,N_19785);
and UO_1049 (O_1049,N_19784,N_19776);
or UO_1050 (O_1050,N_19617,N_19730);
nor UO_1051 (O_1051,N_19735,N_19540);
nand UO_1052 (O_1052,N_19844,N_19873);
and UO_1053 (O_1053,N_19631,N_19924);
and UO_1054 (O_1054,N_19544,N_19795);
xor UO_1055 (O_1055,N_19964,N_19816);
nor UO_1056 (O_1056,N_19939,N_19929);
nand UO_1057 (O_1057,N_19874,N_19544);
and UO_1058 (O_1058,N_19821,N_19797);
nand UO_1059 (O_1059,N_19811,N_19630);
nor UO_1060 (O_1060,N_19682,N_19544);
and UO_1061 (O_1061,N_19539,N_19650);
xor UO_1062 (O_1062,N_19501,N_19506);
nand UO_1063 (O_1063,N_19643,N_19829);
nand UO_1064 (O_1064,N_19825,N_19792);
or UO_1065 (O_1065,N_19877,N_19738);
nand UO_1066 (O_1066,N_19857,N_19697);
nand UO_1067 (O_1067,N_19740,N_19574);
xor UO_1068 (O_1068,N_19577,N_19935);
and UO_1069 (O_1069,N_19625,N_19958);
and UO_1070 (O_1070,N_19512,N_19780);
nand UO_1071 (O_1071,N_19612,N_19776);
or UO_1072 (O_1072,N_19910,N_19911);
xnor UO_1073 (O_1073,N_19768,N_19652);
and UO_1074 (O_1074,N_19691,N_19826);
nor UO_1075 (O_1075,N_19580,N_19747);
nand UO_1076 (O_1076,N_19816,N_19706);
and UO_1077 (O_1077,N_19533,N_19657);
and UO_1078 (O_1078,N_19668,N_19612);
nor UO_1079 (O_1079,N_19905,N_19979);
or UO_1080 (O_1080,N_19697,N_19728);
nor UO_1081 (O_1081,N_19571,N_19760);
and UO_1082 (O_1082,N_19559,N_19952);
nor UO_1083 (O_1083,N_19524,N_19757);
and UO_1084 (O_1084,N_19911,N_19858);
or UO_1085 (O_1085,N_19906,N_19773);
and UO_1086 (O_1086,N_19645,N_19868);
xor UO_1087 (O_1087,N_19552,N_19751);
xnor UO_1088 (O_1088,N_19768,N_19909);
xor UO_1089 (O_1089,N_19851,N_19891);
and UO_1090 (O_1090,N_19826,N_19739);
nor UO_1091 (O_1091,N_19542,N_19957);
or UO_1092 (O_1092,N_19729,N_19507);
or UO_1093 (O_1093,N_19520,N_19595);
or UO_1094 (O_1094,N_19897,N_19722);
or UO_1095 (O_1095,N_19562,N_19672);
and UO_1096 (O_1096,N_19735,N_19552);
or UO_1097 (O_1097,N_19951,N_19622);
nand UO_1098 (O_1098,N_19845,N_19607);
nand UO_1099 (O_1099,N_19771,N_19842);
xor UO_1100 (O_1100,N_19837,N_19773);
nor UO_1101 (O_1101,N_19938,N_19848);
nand UO_1102 (O_1102,N_19710,N_19638);
nand UO_1103 (O_1103,N_19546,N_19927);
xnor UO_1104 (O_1104,N_19597,N_19851);
and UO_1105 (O_1105,N_19556,N_19566);
xor UO_1106 (O_1106,N_19668,N_19997);
or UO_1107 (O_1107,N_19987,N_19508);
or UO_1108 (O_1108,N_19875,N_19935);
nor UO_1109 (O_1109,N_19683,N_19748);
or UO_1110 (O_1110,N_19808,N_19771);
nor UO_1111 (O_1111,N_19667,N_19549);
or UO_1112 (O_1112,N_19823,N_19898);
nor UO_1113 (O_1113,N_19857,N_19968);
nand UO_1114 (O_1114,N_19704,N_19617);
and UO_1115 (O_1115,N_19799,N_19708);
or UO_1116 (O_1116,N_19759,N_19696);
or UO_1117 (O_1117,N_19949,N_19857);
xor UO_1118 (O_1118,N_19939,N_19913);
xor UO_1119 (O_1119,N_19525,N_19866);
nor UO_1120 (O_1120,N_19570,N_19687);
xor UO_1121 (O_1121,N_19811,N_19761);
and UO_1122 (O_1122,N_19956,N_19876);
xor UO_1123 (O_1123,N_19605,N_19976);
nand UO_1124 (O_1124,N_19526,N_19680);
or UO_1125 (O_1125,N_19611,N_19825);
nand UO_1126 (O_1126,N_19689,N_19766);
and UO_1127 (O_1127,N_19865,N_19877);
nor UO_1128 (O_1128,N_19689,N_19692);
or UO_1129 (O_1129,N_19954,N_19594);
nor UO_1130 (O_1130,N_19577,N_19955);
nor UO_1131 (O_1131,N_19734,N_19849);
nand UO_1132 (O_1132,N_19803,N_19520);
xnor UO_1133 (O_1133,N_19890,N_19822);
nor UO_1134 (O_1134,N_19503,N_19663);
xnor UO_1135 (O_1135,N_19538,N_19806);
nand UO_1136 (O_1136,N_19731,N_19587);
nor UO_1137 (O_1137,N_19846,N_19897);
or UO_1138 (O_1138,N_19928,N_19761);
and UO_1139 (O_1139,N_19748,N_19539);
nor UO_1140 (O_1140,N_19881,N_19892);
nand UO_1141 (O_1141,N_19867,N_19519);
nor UO_1142 (O_1142,N_19938,N_19981);
nor UO_1143 (O_1143,N_19983,N_19584);
xor UO_1144 (O_1144,N_19697,N_19804);
nand UO_1145 (O_1145,N_19985,N_19623);
nor UO_1146 (O_1146,N_19969,N_19502);
xnor UO_1147 (O_1147,N_19613,N_19953);
and UO_1148 (O_1148,N_19889,N_19733);
xor UO_1149 (O_1149,N_19606,N_19592);
nor UO_1150 (O_1150,N_19581,N_19782);
xnor UO_1151 (O_1151,N_19907,N_19943);
nor UO_1152 (O_1152,N_19890,N_19505);
nor UO_1153 (O_1153,N_19925,N_19839);
nand UO_1154 (O_1154,N_19968,N_19989);
or UO_1155 (O_1155,N_19573,N_19838);
nand UO_1156 (O_1156,N_19554,N_19930);
or UO_1157 (O_1157,N_19720,N_19604);
xor UO_1158 (O_1158,N_19871,N_19772);
xnor UO_1159 (O_1159,N_19861,N_19864);
nand UO_1160 (O_1160,N_19953,N_19935);
or UO_1161 (O_1161,N_19931,N_19623);
nor UO_1162 (O_1162,N_19697,N_19853);
xnor UO_1163 (O_1163,N_19901,N_19684);
and UO_1164 (O_1164,N_19964,N_19740);
nand UO_1165 (O_1165,N_19804,N_19545);
xor UO_1166 (O_1166,N_19905,N_19710);
nor UO_1167 (O_1167,N_19843,N_19684);
nor UO_1168 (O_1168,N_19922,N_19760);
xnor UO_1169 (O_1169,N_19914,N_19564);
and UO_1170 (O_1170,N_19640,N_19672);
or UO_1171 (O_1171,N_19876,N_19847);
or UO_1172 (O_1172,N_19830,N_19654);
or UO_1173 (O_1173,N_19984,N_19539);
nor UO_1174 (O_1174,N_19679,N_19831);
xor UO_1175 (O_1175,N_19866,N_19621);
nand UO_1176 (O_1176,N_19533,N_19532);
nand UO_1177 (O_1177,N_19635,N_19934);
nor UO_1178 (O_1178,N_19554,N_19722);
nand UO_1179 (O_1179,N_19551,N_19659);
nand UO_1180 (O_1180,N_19886,N_19702);
and UO_1181 (O_1181,N_19573,N_19690);
nand UO_1182 (O_1182,N_19757,N_19672);
nand UO_1183 (O_1183,N_19774,N_19628);
and UO_1184 (O_1184,N_19602,N_19687);
or UO_1185 (O_1185,N_19821,N_19773);
nor UO_1186 (O_1186,N_19621,N_19840);
nand UO_1187 (O_1187,N_19587,N_19606);
and UO_1188 (O_1188,N_19653,N_19695);
and UO_1189 (O_1189,N_19832,N_19574);
nor UO_1190 (O_1190,N_19824,N_19919);
nor UO_1191 (O_1191,N_19660,N_19743);
nand UO_1192 (O_1192,N_19694,N_19907);
nand UO_1193 (O_1193,N_19565,N_19725);
or UO_1194 (O_1194,N_19581,N_19609);
and UO_1195 (O_1195,N_19811,N_19837);
and UO_1196 (O_1196,N_19802,N_19676);
nand UO_1197 (O_1197,N_19901,N_19669);
xnor UO_1198 (O_1198,N_19668,N_19669);
or UO_1199 (O_1199,N_19770,N_19913);
and UO_1200 (O_1200,N_19966,N_19521);
xnor UO_1201 (O_1201,N_19503,N_19998);
nor UO_1202 (O_1202,N_19707,N_19821);
nor UO_1203 (O_1203,N_19566,N_19581);
or UO_1204 (O_1204,N_19851,N_19758);
nor UO_1205 (O_1205,N_19918,N_19938);
xnor UO_1206 (O_1206,N_19823,N_19685);
and UO_1207 (O_1207,N_19841,N_19961);
and UO_1208 (O_1208,N_19787,N_19799);
and UO_1209 (O_1209,N_19912,N_19837);
xor UO_1210 (O_1210,N_19500,N_19855);
and UO_1211 (O_1211,N_19512,N_19658);
nor UO_1212 (O_1212,N_19768,N_19541);
or UO_1213 (O_1213,N_19595,N_19941);
nand UO_1214 (O_1214,N_19905,N_19640);
xor UO_1215 (O_1215,N_19951,N_19782);
nor UO_1216 (O_1216,N_19942,N_19568);
nand UO_1217 (O_1217,N_19805,N_19945);
and UO_1218 (O_1218,N_19543,N_19996);
and UO_1219 (O_1219,N_19513,N_19525);
or UO_1220 (O_1220,N_19686,N_19970);
nand UO_1221 (O_1221,N_19796,N_19927);
nand UO_1222 (O_1222,N_19875,N_19769);
nand UO_1223 (O_1223,N_19925,N_19774);
xnor UO_1224 (O_1224,N_19522,N_19782);
nor UO_1225 (O_1225,N_19973,N_19855);
nor UO_1226 (O_1226,N_19896,N_19981);
nand UO_1227 (O_1227,N_19777,N_19788);
xnor UO_1228 (O_1228,N_19981,N_19696);
nand UO_1229 (O_1229,N_19982,N_19644);
xor UO_1230 (O_1230,N_19710,N_19508);
and UO_1231 (O_1231,N_19560,N_19765);
and UO_1232 (O_1232,N_19844,N_19883);
or UO_1233 (O_1233,N_19997,N_19833);
and UO_1234 (O_1234,N_19951,N_19843);
nor UO_1235 (O_1235,N_19765,N_19552);
or UO_1236 (O_1236,N_19540,N_19672);
nand UO_1237 (O_1237,N_19985,N_19953);
and UO_1238 (O_1238,N_19757,N_19526);
xor UO_1239 (O_1239,N_19839,N_19923);
or UO_1240 (O_1240,N_19657,N_19691);
and UO_1241 (O_1241,N_19902,N_19536);
or UO_1242 (O_1242,N_19682,N_19813);
nor UO_1243 (O_1243,N_19817,N_19540);
and UO_1244 (O_1244,N_19952,N_19808);
xor UO_1245 (O_1245,N_19529,N_19721);
nand UO_1246 (O_1246,N_19800,N_19694);
or UO_1247 (O_1247,N_19804,N_19983);
nand UO_1248 (O_1248,N_19504,N_19725);
nand UO_1249 (O_1249,N_19736,N_19965);
and UO_1250 (O_1250,N_19883,N_19724);
xnor UO_1251 (O_1251,N_19851,N_19995);
or UO_1252 (O_1252,N_19999,N_19706);
or UO_1253 (O_1253,N_19728,N_19541);
nor UO_1254 (O_1254,N_19928,N_19692);
or UO_1255 (O_1255,N_19736,N_19933);
nor UO_1256 (O_1256,N_19718,N_19887);
and UO_1257 (O_1257,N_19949,N_19930);
nand UO_1258 (O_1258,N_19981,N_19721);
and UO_1259 (O_1259,N_19902,N_19799);
or UO_1260 (O_1260,N_19722,N_19978);
nor UO_1261 (O_1261,N_19755,N_19757);
nor UO_1262 (O_1262,N_19826,N_19853);
or UO_1263 (O_1263,N_19578,N_19886);
and UO_1264 (O_1264,N_19609,N_19741);
and UO_1265 (O_1265,N_19517,N_19563);
nor UO_1266 (O_1266,N_19521,N_19884);
or UO_1267 (O_1267,N_19822,N_19640);
and UO_1268 (O_1268,N_19544,N_19960);
or UO_1269 (O_1269,N_19776,N_19638);
xor UO_1270 (O_1270,N_19564,N_19849);
or UO_1271 (O_1271,N_19870,N_19763);
and UO_1272 (O_1272,N_19571,N_19680);
nor UO_1273 (O_1273,N_19741,N_19813);
nand UO_1274 (O_1274,N_19971,N_19914);
nor UO_1275 (O_1275,N_19659,N_19531);
nand UO_1276 (O_1276,N_19741,N_19907);
xor UO_1277 (O_1277,N_19514,N_19953);
nand UO_1278 (O_1278,N_19646,N_19685);
nor UO_1279 (O_1279,N_19986,N_19619);
or UO_1280 (O_1280,N_19626,N_19960);
xnor UO_1281 (O_1281,N_19845,N_19923);
and UO_1282 (O_1282,N_19604,N_19690);
and UO_1283 (O_1283,N_19518,N_19509);
nor UO_1284 (O_1284,N_19767,N_19544);
and UO_1285 (O_1285,N_19607,N_19969);
nand UO_1286 (O_1286,N_19519,N_19555);
nor UO_1287 (O_1287,N_19908,N_19618);
and UO_1288 (O_1288,N_19641,N_19590);
nor UO_1289 (O_1289,N_19919,N_19789);
or UO_1290 (O_1290,N_19978,N_19563);
and UO_1291 (O_1291,N_19566,N_19914);
or UO_1292 (O_1292,N_19737,N_19802);
xnor UO_1293 (O_1293,N_19685,N_19787);
nor UO_1294 (O_1294,N_19651,N_19893);
and UO_1295 (O_1295,N_19657,N_19906);
nand UO_1296 (O_1296,N_19646,N_19742);
or UO_1297 (O_1297,N_19796,N_19873);
xor UO_1298 (O_1298,N_19643,N_19685);
nor UO_1299 (O_1299,N_19912,N_19793);
nand UO_1300 (O_1300,N_19532,N_19802);
xnor UO_1301 (O_1301,N_19820,N_19904);
nor UO_1302 (O_1302,N_19677,N_19864);
nor UO_1303 (O_1303,N_19674,N_19698);
nor UO_1304 (O_1304,N_19566,N_19531);
or UO_1305 (O_1305,N_19732,N_19915);
or UO_1306 (O_1306,N_19575,N_19694);
or UO_1307 (O_1307,N_19757,N_19607);
nand UO_1308 (O_1308,N_19843,N_19910);
nand UO_1309 (O_1309,N_19692,N_19515);
xnor UO_1310 (O_1310,N_19673,N_19580);
nor UO_1311 (O_1311,N_19610,N_19626);
and UO_1312 (O_1312,N_19896,N_19667);
and UO_1313 (O_1313,N_19806,N_19656);
or UO_1314 (O_1314,N_19770,N_19782);
nor UO_1315 (O_1315,N_19510,N_19521);
xor UO_1316 (O_1316,N_19973,N_19937);
xor UO_1317 (O_1317,N_19507,N_19709);
or UO_1318 (O_1318,N_19920,N_19579);
and UO_1319 (O_1319,N_19523,N_19623);
nand UO_1320 (O_1320,N_19968,N_19696);
and UO_1321 (O_1321,N_19571,N_19672);
and UO_1322 (O_1322,N_19732,N_19568);
xor UO_1323 (O_1323,N_19644,N_19737);
nor UO_1324 (O_1324,N_19626,N_19644);
xor UO_1325 (O_1325,N_19741,N_19842);
or UO_1326 (O_1326,N_19805,N_19565);
nor UO_1327 (O_1327,N_19673,N_19869);
or UO_1328 (O_1328,N_19893,N_19886);
or UO_1329 (O_1329,N_19678,N_19584);
nor UO_1330 (O_1330,N_19661,N_19953);
and UO_1331 (O_1331,N_19742,N_19508);
nor UO_1332 (O_1332,N_19839,N_19881);
and UO_1333 (O_1333,N_19903,N_19907);
nand UO_1334 (O_1334,N_19650,N_19939);
or UO_1335 (O_1335,N_19644,N_19617);
and UO_1336 (O_1336,N_19717,N_19659);
or UO_1337 (O_1337,N_19800,N_19688);
nand UO_1338 (O_1338,N_19930,N_19605);
or UO_1339 (O_1339,N_19634,N_19509);
and UO_1340 (O_1340,N_19650,N_19810);
and UO_1341 (O_1341,N_19606,N_19535);
xnor UO_1342 (O_1342,N_19987,N_19655);
or UO_1343 (O_1343,N_19760,N_19707);
and UO_1344 (O_1344,N_19852,N_19634);
nand UO_1345 (O_1345,N_19756,N_19975);
nor UO_1346 (O_1346,N_19946,N_19852);
xnor UO_1347 (O_1347,N_19803,N_19707);
or UO_1348 (O_1348,N_19936,N_19797);
nand UO_1349 (O_1349,N_19899,N_19568);
and UO_1350 (O_1350,N_19544,N_19718);
or UO_1351 (O_1351,N_19792,N_19701);
or UO_1352 (O_1352,N_19585,N_19594);
xnor UO_1353 (O_1353,N_19627,N_19562);
nand UO_1354 (O_1354,N_19803,N_19941);
or UO_1355 (O_1355,N_19691,N_19576);
nand UO_1356 (O_1356,N_19679,N_19642);
and UO_1357 (O_1357,N_19511,N_19648);
nor UO_1358 (O_1358,N_19726,N_19584);
or UO_1359 (O_1359,N_19645,N_19888);
nor UO_1360 (O_1360,N_19528,N_19979);
nor UO_1361 (O_1361,N_19560,N_19997);
or UO_1362 (O_1362,N_19587,N_19978);
and UO_1363 (O_1363,N_19863,N_19935);
nor UO_1364 (O_1364,N_19648,N_19823);
xnor UO_1365 (O_1365,N_19944,N_19857);
and UO_1366 (O_1366,N_19877,N_19717);
xnor UO_1367 (O_1367,N_19953,N_19880);
or UO_1368 (O_1368,N_19759,N_19575);
or UO_1369 (O_1369,N_19753,N_19534);
and UO_1370 (O_1370,N_19790,N_19803);
nor UO_1371 (O_1371,N_19773,N_19592);
nand UO_1372 (O_1372,N_19686,N_19900);
xor UO_1373 (O_1373,N_19794,N_19866);
xor UO_1374 (O_1374,N_19766,N_19710);
or UO_1375 (O_1375,N_19928,N_19674);
xnor UO_1376 (O_1376,N_19528,N_19648);
xnor UO_1377 (O_1377,N_19665,N_19534);
xor UO_1378 (O_1378,N_19914,N_19536);
nand UO_1379 (O_1379,N_19823,N_19566);
or UO_1380 (O_1380,N_19891,N_19666);
and UO_1381 (O_1381,N_19622,N_19789);
nor UO_1382 (O_1382,N_19980,N_19625);
xor UO_1383 (O_1383,N_19727,N_19803);
and UO_1384 (O_1384,N_19834,N_19581);
and UO_1385 (O_1385,N_19678,N_19889);
and UO_1386 (O_1386,N_19854,N_19655);
nand UO_1387 (O_1387,N_19903,N_19895);
and UO_1388 (O_1388,N_19775,N_19856);
or UO_1389 (O_1389,N_19684,N_19569);
and UO_1390 (O_1390,N_19898,N_19884);
or UO_1391 (O_1391,N_19610,N_19831);
and UO_1392 (O_1392,N_19854,N_19833);
or UO_1393 (O_1393,N_19542,N_19602);
and UO_1394 (O_1394,N_19815,N_19568);
or UO_1395 (O_1395,N_19819,N_19824);
and UO_1396 (O_1396,N_19817,N_19536);
nand UO_1397 (O_1397,N_19615,N_19954);
or UO_1398 (O_1398,N_19928,N_19734);
and UO_1399 (O_1399,N_19515,N_19666);
nor UO_1400 (O_1400,N_19641,N_19897);
xnor UO_1401 (O_1401,N_19708,N_19989);
or UO_1402 (O_1402,N_19591,N_19666);
or UO_1403 (O_1403,N_19748,N_19743);
xor UO_1404 (O_1404,N_19802,N_19675);
and UO_1405 (O_1405,N_19604,N_19701);
and UO_1406 (O_1406,N_19980,N_19730);
xor UO_1407 (O_1407,N_19909,N_19653);
xor UO_1408 (O_1408,N_19667,N_19658);
and UO_1409 (O_1409,N_19896,N_19552);
and UO_1410 (O_1410,N_19616,N_19743);
and UO_1411 (O_1411,N_19914,N_19563);
nand UO_1412 (O_1412,N_19528,N_19501);
nor UO_1413 (O_1413,N_19601,N_19567);
and UO_1414 (O_1414,N_19715,N_19986);
and UO_1415 (O_1415,N_19524,N_19693);
and UO_1416 (O_1416,N_19760,N_19591);
and UO_1417 (O_1417,N_19818,N_19605);
and UO_1418 (O_1418,N_19789,N_19794);
xor UO_1419 (O_1419,N_19960,N_19995);
nor UO_1420 (O_1420,N_19561,N_19625);
nand UO_1421 (O_1421,N_19853,N_19762);
nand UO_1422 (O_1422,N_19762,N_19955);
nand UO_1423 (O_1423,N_19503,N_19995);
and UO_1424 (O_1424,N_19983,N_19994);
and UO_1425 (O_1425,N_19791,N_19603);
nor UO_1426 (O_1426,N_19793,N_19979);
and UO_1427 (O_1427,N_19965,N_19637);
and UO_1428 (O_1428,N_19641,N_19668);
and UO_1429 (O_1429,N_19921,N_19842);
or UO_1430 (O_1430,N_19628,N_19958);
nor UO_1431 (O_1431,N_19615,N_19781);
nand UO_1432 (O_1432,N_19934,N_19733);
nand UO_1433 (O_1433,N_19644,N_19599);
nand UO_1434 (O_1434,N_19961,N_19991);
xnor UO_1435 (O_1435,N_19807,N_19936);
nor UO_1436 (O_1436,N_19799,N_19897);
nand UO_1437 (O_1437,N_19572,N_19779);
and UO_1438 (O_1438,N_19895,N_19704);
nand UO_1439 (O_1439,N_19698,N_19742);
or UO_1440 (O_1440,N_19955,N_19898);
or UO_1441 (O_1441,N_19715,N_19866);
nand UO_1442 (O_1442,N_19817,N_19875);
or UO_1443 (O_1443,N_19979,N_19560);
or UO_1444 (O_1444,N_19576,N_19898);
xor UO_1445 (O_1445,N_19598,N_19693);
xor UO_1446 (O_1446,N_19799,N_19757);
nor UO_1447 (O_1447,N_19965,N_19771);
and UO_1448 (O_1448,N_19900,N_19501);
xnor UO_1449 (O_1449,N_19576,N_19801);
and UO_1450 (O_1450,N_19815,N_19546);
and UO_1451 (O_1451,N_19859,N_19558);
nand UO_1452 (O_1452,N_19547,N_19875);
nand UO_1453 (O_1453,N_19961,N_19573);
nand UO_1454 (O_1454,N_19853,N_19526);
xnor UO_1455 (O_1455,N_19700,N_19960);
nand UO_1456 (O_1456,N_19650,N_19672);
and UO_1457 (O_1457,N_19851,N_19920);
nor UO_1458 (O_1458,N_19596,N_19849);
nor UO_1459 (O_1459,N_19831,N_19852);
nor UO_1460 (O_1460,N_19716,N_19705);
and UO_1461 (O_1461,N_19809,N_19779);
and UO_1462 (O_1462,N_19830,N_19993);
nand UO_1463 (O_1463,N_19566,N_19671);
xor UO_1464 (O_1464,N_19914,N_19647);
or UO_1465 (O_1465,N_19579,N_19719);
and UO_1466 (O_1466,N_19635,N_19908);
or UO_1467 (O_1467,N_19862,N_19537);
or UO_1468 (O_1468,N_19695,N_19905);
or UO_1469 (O_1469,N_19814,N_19921);
nor UO_1470 (O_1470,N_19509,N_19610);
or UO_1471 (O_1471,N_19704,N_19625);
nor UO_1472 (O_1472,N_19596,N_19932);
nor UO_1473 (O_1473,N_19699,N_19713);
and UO_1474 (O_1474,N_19971,N_19662);
nor UO_1475 (O_1475,N_19545,N_19857);
nand UO_1476 (O_1476,N_19548,N_19812);
or UO_1477 (O_1477,N_19620,N_19821);
xnor UO_1478 (O_1478,N_19525,N_19801);
xor UO_1479 (O_1479,N_19776,N_19910);
nor UO_1480 (O_1480,N_19745,N_19728);
xor UO_1481 (O_1481,N_19587,N_19672);
or UO_1482 (O_1482,N_19755,N_19855);
nor UO_1483 (O_1483,N_19721,N_19781);
and UO_1484 (O_1484,N_19812,N_19507);
and UO_1485 (O_1485,N_19522,N_19807);
xor UO_1486 (O_1486,N_19803,N_19792);
xnor UO_1487 (O_1487,N_19944,N_19584);
xnor UO_1488 (O_1488,N_19688,N_19809);
xor UO_1489 (O_1489,N_19800,N_19579);
nand UO_1490 (O_1490,N_19775,N_19830);
or UO_1491 (O_1491,N_19948,N_19854);
or UO_1492 (O_1492,N_19972,N_19657);
or UO_1493 (O_1493,N_19696,N_19519);
nor UO_1494 (O_1494,N_19932,N_19641);
or UO_1495 (O_1495,N_19771,N_19811);
nand UO_1496 (O_1496,N_19783,N_19531);
nand UO_1497 (O_1497,N_19545,N_19874);
xnor UO_1498 (O_1498,N_19758,N_19503);
and UO_1499 (O_1499,N_19511,N_19586);
or UO_1500 (O_1500,N_19831,N_19559);
and UO_1501 (O_1501,N_19848,N_19837);
or UO_1502 (O_1502,N_19614,N_19505);
nand UO_1503 (O_1503,N_19821,N_19782);
xnor UO_1504 (O_1504,N_19530,N_19604);
xor UO_1505 (O_1505,N_19966,N_19837);
nor UO_1506 (O_1506,N_19657,N_19666);
nand UO_1507 (O_1507,N_19593,N_19524);
xnor UO_1508 (O_1508,N_19711,N_19633);
and UO_1509 (O_1509,N_19721,N_19830);
xor UO_1510 (O_1510,N_19536,N_19693);
nor UO_1511 (O_1511,N_19503,N_19939);
nand UO_1512 (O_1512,N_19651,N_19562);
nor UO_1513 (O_1513,N_19812,N_19899);
xor UO_1514 (O_1514,N_19757,N_19956);
nor UO_1515 (O_1515,N_19768,N_19962);
nor UO_1516 (O_1516,N_19703,N_19734);
and UO_1517 (O_1517,N_19726,N_19570);
or UO_1518 (O_1518,N_19856,N_19805);
and UO_1519 (O_1519,N_19579,N_19519);
xor UO_1520 (O_1520,N_19531,N_19723);
nor UO_1521 (O_1521,N_19828,N_19934);
or UO_1522 (O_1522,N_19518,N_19569);
nor UO_1523 (O_1523,N_19777,N_19652);
or UO_1524 (O_1524,N_19950,N_19542);
xnor UO_1525 (O_1525,N_19975,N_19751);
or UO_1526 (O_1526,N_19513,N_19979);
nand UO_1527 (O_1527,N_19708,N_19587);
or UO_1528 (O_1528,N_19644,N_19867);
or UO_1529 (O_1529,N_19882,N_19970);
or UO_1530 (O_1530,N_19540,N_19539);
nand UO_1531 (O_1531,N_19783,N_19655);
xnor UO_1532 (O_1532,N_19517,N_19570);
nor UO_1533 (O_1533,N_19978,N_19969);
and UO_1534 (O_1534,N_19935,N_19820);
xnor UO_1535 (O_1535,N_19584,N_19723);
xnor UO_1536 (O_1536,N_19772,N_19886);
or UO_1537 (O_1537,N_19678,N_19712);
or UO_1538 (O_1538,N_19670,N_19937);
nand UO_1539 (O_1539,N_19685,N_19805);
nor UO_1540 (O_1540,N_19509,N_19748);
nand UO_1541 (O_1541,N_19708,N_19664);
and UO_1542 (O_1542,N_19934,N_19971);
nand UO_1543 (O_1543,N_19910,N_19658);
xnor UO_1544 (O_1544,N_19818,N_19710);
xnor UO_1545 (O_1545,N_19585,N_19898);
xor UO_1546 (O_1546,N_19683,N_19962);
and UO_1547 (O_1547,N_19747,N_19668);
and UO_1548 (O_1548,N_19740,N_19851);
nand UO_1549 (O_1549,N_19700,N_19610);
and UO_1550 (O_1550,N_19584,N_19956);
and UO_1551 (O_1551,N_19731,N_19780);
and UO_1552 (O_1552,N_19705,N_19803);
xnor UO_1553 (O_1553,N_19629,N_19805);
nor UO_1554 (O_1554,N_19659,N_19976);
nand UO_1555 (O_1555,N_19724,N_19722);
nand UO_1556 (O_1556,N_19589,N_19674);
and UO_1557 (O_1557,N_19905,N_19522);
nor UO_1558 (O_1558,N_19873,N_19576);
or UO_1559 (O_1559,N_19551,N_19997);
nand UO_1560 (O_1560,N_19586,N_19562);
nor UO_1561 (O_1561,N_19879,N_19843);
xnor UO_1562 (O_1562,N_19573,N_19616);
and UO_1563 (O_1563,N_19830,N_19536);
nor UO_1564 (O_1564,N_19872,N_19823);
and UO_1565 (O_1565,N_19748,N_19730);
or UO_1566 (O_1566,N_19574,N_19789);
or UO_1567 (O_1567,N_19943,N_19996);
nor UO_1568 (O_1568,N_19840,N_19587);
or UO_1569 (O_1569,N_19548,N_19985);
nand UO_1570 (O_1570,N_19537,N_19948);
and UO_1571 (O_1571,N_19883,N_19645);
or UO_1572 (O_1572,N_19711,N_19612);
nor UO_1573 (O_1573,N_19700,N_19557);
xnor UO_1574 (O_1574,N_19735,N_19946);
and UO_1575 (O_1575,N_19924,N_19663);
nor UO_1576 (O_1576,N_19622,N_19855);
nor UO_1577 (O_1577,N_19545,N_19530);
and UO_1578 (O_1578,N_19716,N_19948);
and UO_1579 (O_1579,N_19750,N_19721);
and UO_1580 (O_1580,N_19620,N_19888);
xor UO_1581 (O_1581,N_19880,N_19632);
xnor UO_1582 (O_1582,N_19637,N_19682);
nand UO_1583 (O_1583,N_19887,N_19511);
and UO_1584 (O_1584,N_19608,N_19645);
nor UO_1585 (O_1585,N_19813,N_19958);
xor UO_1586 (O_1586,N_19641,N_19657);
or UO_1587 (O_1587,N_19560,N_19616);
nor UO_1588 (O_1588,N_19503,N_19929);
xnor UO_1589 (O_1589,N_19709,N_19700);
nand UO_1590 (O_1590,N_19942,N_19863);
or UO_1591 (O_1591,N_19618,N_19509);
nand UO_1592 (O_1592,N_19539,N_19681);
nand UO_1593 (O_1593,N_19951,N_19915);
and UO_1594 (O_1594,N_19989,N_19615);
nand UO_1595 (O_1595,N_19680,N_19813);
nand UO_1596 (O_1596,N_19909,N_19659);
xnor UO_1597 (O_1597,N_19942,N_19542);
nor UO_1598 (O_1598,N_19578,N_19747);
nand UO_1599 (O_1599,N_19735,N_19587);
nand UO_1600 (O_1600,N_19710,N_19856);
and UO_1601 (O_1601,N_19655,N_19858);
or UO_1602 (O_1602,N_19749,N_19528);
nand UO_1603 (O_1603,N_19832,N_19953);
nor UO_1604 (O_1604,N_19897,N_19861);
nor UO_1605 (O_1605,N_19727,N_19891);
nand UO_1606 (O_1606,N_19881,N_19894);
nand UO_1607 (O_1607,N_19597,N_19599);
nand UO_1608 (O_1608,N_19985,N_19616);
or UO_1609 (O_1609,N_19868,N_19628);
or UO_1610 (O_1610,N_19516,N_19865);
xnor UO_1611 (O_1611,N_19839,N_19812);
nor UO_1612 (O_1612,N_19535,N_19600);
nor UO_1613 (O_1613,N_19913,N_19509);
nor UO_1614 (O_1614,N_19521,N_19917);
nand UO_1615 (O_1615,N_19520,N_19680);
xnor UO_1616 (O_1616,N_19973,N_19685);
nand UO_1617 (O_1617,N_19960,N_19982);
or UO_1618 (O_1618,N_19813,N_19592);
xor UO_1619 (O_1619,N_19801,N_19620);
and UO_1620 (O_1620,N_19504,N_19702);
nand UO_1621 (O_1621,N_19524,N_19750);
nor UO_1622 (O_1622,N_19738,N_19860);
nand UO_1623 (O_1623,N_19950,N_19806);
and UO_1624 (O_1624,N_19634,N_19560);
nor UO_1625 (O_1625,N_19945,N_19968);
nor UO_1626 (O_1626,N_19562,N_19581);
and UO_1627 (O_1627,N_19881,N_19784);
xnor UO_1628 (O_1628,N_19675,N_19609);
or UO_1629 (O_1629,N_19721,N_19704);
and UO_1630 (O_1630,N_19845,N_19566);
and UO_1631 (O_1631,N_19935,N_19605);
xnor UO_1632 (O_1632,N_19636,N_19502);
nand UO_1633 (O_1633,N_19933,N_19613);
and UO_1634 (O_1634,N_19542,N_19769);
xnor UO_1635 (O_1635,N_19975,N_19973);
nand UO_1636 (O_1636,N_19652,N_19564);
nand UO_1637 (O_1637,N_19734,N_19979);
nand UO_1638 (O_1638,N_19716,N_19665);
xor UO_1639 (O_1639,N_19589,N_19555);
nand UO_1640 (O_1640,N_19945,N_19893);
and UO_1641 (O_1641,N_19608,N_19722);
nor UO_1642 (O_1642,N_19852,N_19869);
and UO_1643 (O_1643,N_19962,N_19801);
and UO_1644 (O_1644,N_19588,N_19959);
and UO_1645 (O_1645,N_19598,N_19523);
and UO_1646 (O_1646,N_19896,N_19936);
or UO_1647 (O_1647,N_19866,N_19780);
xor UO_1648 (O_1648,N_19779,N_19960);
nand UO_1649 (O_1649,N_19946,N_19785);
nor UO_1650 (O_1650,N_19692,N_19545);
nand UO_1651 (O_1651,N_19530,N_19825);
and UO_1652 (O_1652,N_19976,N_19882);
or UO_1653 (O_1653,N_19943,N_19578);
nand UO_1654 (O_1654,N_19889,N_19952);
nand UO_1655 (O_1655,N_19773,N_19840);
nor UO_1656 (O_1656,N_19581,N_19573);
nor UO_1657 (O_1657,N_19824,N_19908);
nand UO_1658 (O_1658,N_19674,N_19566);
nor UO_1659 (O_1659,N_19565,N_19757);
nand UO_1660 (O_1660,N_19799,N_19919);
nand UO_1661 (O_1661,N_19619,N_19812);
nor UO_1662 (O_1662,N_19637,N_19652);
nand UO_1663 (O_1663,N_19668,N_19815);
xnor UO_1664 (O_1664,N_19796,N_19799);
nor UO_1665 (O_1665,N_19661,N_19764);
or UO_1666 (O_1666,N_19852,N_19784);
or UO_1667 (O_1667,N_19723,N_19805);
and UO_1668 (O_1668,N_19566,N_19702);
nand UO_1669 (O_1669,N_19641,N_19771);
and UO_1670 (O_1670,N_19550,N_19676);
nor UO_1671 (O_1671,N_19867,N_19998);
xnor UO_1672 (O_1672,N_19674,N_19663);
or UO_1673 (O_1673,N_19784,N_19536);
nor UO_1674 (O_1674,N_19552,N_19932);
nor UO_1675 (O_1675,N_19880,N_19571);
xor UO_1676 (O_1676,N_19817,N_19929);
or UO_1677 (O_1677,N_19983,N_19730);
xor UO_1678 (O_1678,N_19793,N_19843);
and UO_1679 (O_1679,N_19607,N_19876);
or UO_1680 (O_1680,N_19793,N_19888);
nor UO_1681 (O_1681,N_19814,N_19596);
and UO_1682 (O_1682,N_19627,N_19523);
and UO_1683 (O_1683,N_19514,N_19950);
and UO_1684 (O_1684,N_19653,N_19672);
and UO_1685 (O_1685,N_19877,N_19722);
or UO_1686 (O_1686,N_19751,N_19950);
nand UO_1687 (O_1687,N_19586,N_19527);
nand UO_1688 (O_1688,N_19747,N_19705);
nor UO_1689 (O_1689,N_19747,N_19704);
xnor UO_1690 (O_1690,N_19573,N_19504);
nand UO_1691 (O_1691,N_19552,N_19856);
or UO_1692 (O_1692,N_19994,N_19512);
or UO_1693 (O_1693,N_19925,N_19954);
nand UO_1694 (O_1694,N_19953,N_19538);
and UO_1695 (O_1695,N_19744,N_19841);
nand UO_1696 (O_1696,N_19855,N_19958);
nor UO_1697 (O_1697,N_19570,N_19676);
or UO_1698 (O_1698,N_19686,N_19935);
nor UO_1699 (O_1699,N_19547,N_19507);
and UO_1700 (O_1700,N_19961,N_19875);
or UO_1701 (O_1701,N_19831,N_19729);
xor UO_1702 (O_1702,N_19568,N_19526);
and UO_1703 (O_1703,N_19832,N_19909);
xor UO_1704 (O_1704,N_19743,N_19977);
or UO_1705 (O_1705,N_19609,N_19560);
xor UO_1706 (O_1706,N_19705,N_19810);
or UO_1707 (O_1707,N_19728,N_19855);
or UO_1708 (O_1708,N_19690,N_19523);
and UO_1709 (O_1709,N_19908,N_19615);
nor UO_1710 (O_1710,N_19850,N_19685);
or UO_1711 (O_1711,N_19721,N_19755);
nor UO_1712 (O_1712,N_19525,N_19822);
and UO_1713 (O_1713,N_19799,N_19650);
and UO_1714 (O_1714,N_19844,N_19604);
nand UO_1715 (O_1715,N_19665,N_19874);
and UO_1716 (O_1716,N_19850,N_19610);
or UO_1717 (O_1717,N_19604,N_19810);
and UO_1718 (O_1718,N_19948,N_19812);
or UO_1719 (O_1719,N_19638,N_19560);
or UO_1720 (O_1720,N_19886,N_19705);
xnor UO_1721 (O_1721,N_19557,N_19804);
nor UO_1722 (O_1722,N_19724,N_19810);
nand UO_1723 (O_1723,N_19788,N_19933);
nor UO_1724 (O_1724,N_19530,N_19565);
nand UO_1725 (O_1725,N_19883,N_19743);
and UO_1726 (O_1726,N_19810,N_19528);
nand UO_1727 (O_1727,N_19677,N_19588);
nand UO_1728 (O_1728,N_19507,N_19848);
or UO_1729 (O_1729,N_19660,N_19687);
nor UO_1730 (O_1730,N_19932,N_19808);
and UO_1731 (O_1731,N_19564,N_19585);
nor UO_1732 (O_1732,N_19574,N_19533);
or UO_1733 (O_1733,N_19651,N_19664);
or UO_1734 (O_1734,N_19834,N_19819);
nand UO_1735 (O_1735,N_19790,N_19514);
and UO_1736 (O_1736,N_19501,N_19810);
or UO_1737 (O_1737,N_19510,N_19605);
nand UO_1738 (O_1738,N_19510,N_19722);
or UO_1739 (O_1739,N_19505,N_19569);
nand UO_1740 (O_1740,N_19686,N_19752);
and UO_1741 (O_1741,N_19693,N_19682);
and UO_1742 (O_1742,N_19512,N_19888);
nand UO_1743 (O_1743,N_19736,N_19559);
and UO_1744 (O_1744,N_19615,N_19951);
nor UO_1745 (O_1745,N_19828,N_19551);
nand UO_1746 (O_1746,N_19924,N_19898);
nand UO_1747 (O_1747,N_19722,N_19596);
or UO_1748 (O_1748,N_19793,N_19820);
and UO_1749 (O_1749,N_19842,N_19644);
and UO_1750 (O_1750,N_19682,N_19690);
and UO_1751 (O_1751,N_19769,N_19704);
nor UO_1752 (O_1752,N_19797,N_19578);
xnor UO_1753 (O_1753,N_19896,N_19638);
or UO_1754 (O_1754,N_19707,N_19564);
xnor UO_1755 (O_1755,N_19967,N_19849);
or UO_1756 (O_1756,N_19820,N_19859);
nand UO_1757 (O_1757,N_19945,N_19737);
nor UO_1758 (O_1758,N_19657,N_19808);
nand UO_1759 (O_1759,N_19911,N_19844);
or UO_1760 (O_1760,N_19794,N_19719);
nand UO_1761 (O_1761,N_19789,N_19781);
nand UO_1762 (O_1762,N_19764,N_19546);
nand UO_1763 (O_1763,N_19872,N_19827);
and UO_1764 (O_1764,N_19857,N_19531);
and UO_1765 (O_1765,N_19701,N_19568);
nor UO_1766 (O_1766,N_19784,N_19755);
xor UO_1767 (O_1767,N_19763,N_19534);
nand UO_1768 (O_1768,N_19509,N_19976);
xnor UO_1769 (O_1769,N_19850,N_19898);
or UO_1770 (O_1770,N_19941,N_19565);
and UO_1771 (O_1771,N_19674,N_19905);
or UO_1772 (O_1772,N_19638,N_19967);
nand UO_1773 (O_1773,N_19566,N_19540);
nand UO_1774 (O_1774,N_19807,N_19552);
and UO_1775 (O_1775,N_19773,N_19580);
xnor UO_1776 (O_1776,N_19684,N_19603);
or UO_1777 (O_1777,N_19815,N_19608);
nand UO_1778 (O_1778,N_19604,N_19984);
nand UO_1779 (O_1779,N_19971,N_19744);
xor UO_1780 (O_1780,N_19895,N_19759);
nand UO_1781 (O_1781,N_19897,N_19977);
and UO_1782 (O_1782,N_19965,N_19589);
or UO_1783 (O_1783,N_19725,N_19551);
xnor UO_1784 (O_1784,N_19585,N_19601);
or UO_1785 (O_1785,N_19817,N_19756);
or UO_1786 (O_1786,N_19888,N_19545);
or UO_1787 (O_1787,N_19647,N_19894);
or UO_1788 (O_1788,N_19580,N_19972);
nand UO_1789 (O_1789,N_19984,N_19563);
nand UO_1790 (O_1790,N_19857,N_19514);
nor UO_1791 (O_1791,N_19715,N_19814);
xnor UO_1792 (O_1792,N_19605,N_19822);
nor UO_1793 (O_1793,N_19530,N_19917);
or UO_1794 (O_1794,N_19929,N_19960);
and UO_1795 (O_1795,N_19925,N_19557);
nor UO_1796 (O_1796,N_19970,N_19536);
nor UO_1797 (O_1797,N_19888,N_19569);
or UO_1798 (O_1798,N_19655,N_19937);
nor UO_1799 (O_1799,N_19987,N_19719);
nand UO_1800 (O_1800,N_19605,N_19720);
or UO_1801 (O_1801,N_19723,N_19961);
nand UO_1802 (O_1802,N_19528,N_19626);
nand UO_1803 (O_1803,N_19865,N_19547);
xnor UO_1804 (O_1804,N_19628,N_19893);
nand UO_1805 (O_1805,N_19804,N_19619);
and UO_1806 (O_1806,N_19718,N_19912);
or UO_1807 (O_1807,N_19544,N_19646);
and UO_1808 (O_1808,N_19564,N_19609);
nor UO_1809 (O_1809,N_19906,N_19764);
nor UO_1810 (O_1810,N_19847,N_19922);
or UO_1811 (O_1811,N_19714,N_19922);
or UO_1812 (O_1812,N_19587,N_19878);
and UO_1813 (O_1813,N_19905,N_19854);
nand UO_1814 (O_1814,N_19702,N_19570);
nor UO_1815 (O_1815,N_19663,N_19603);
nor UO_1816 (O_1816,N_19821,N_19507);
nand UO_1817 (O_1817,N_19723,N_19859);
or UO_1818 (O_1818,N_19599,N_19764);
and UO_1819 (O_1819,N_19690,N_19532);
or UO_1820 (O_1820,N_19560,N_19529);
xnor UO_1821 (O_1821,N_19811,N_19655);
nand UO_1822 (O_1822,N_19730,N_19616);
nand UO_1823 (O_1823,N_19811,N_19858);
nor UO_1824 (O_1824,N_19904,N_19934);
and UO_1825 (O_1825,N_19648,N_19762);
or UO_1826 (O_1826,N_19848,N_19877);
xor UO_1827 (O_1827,N_19991,N_19891);
nand UO_1828 (O_1828,N_19503,N_19836);
xor UO_1829 (O_1829,N_19531,N_19620);
or UO_1830 (O_1830,N_19956,N_19955);
nand UO_1831 (O_1831,N_19599,N_19994);
nand UO_1832 (O_1832,N_19840,N_19857);
and UO_1833 (O_1833,N_19564,N_19938);
nand UO_1834 (O_1834,N_19885,N_19525);
xnor UO_1835 (O_1835,N_19517,N_19791);
or UO_1836 (O_1836,N_19535,N_19938);
and UO_1837 (O_1837,N_19609,N_19974);
nor UO_1838 (O_1838,N_19861,N_19856);
or UO_1839 (O_1839,N_19700,N_19651);
and UO_1840 (O_1840,N_19546,N_19977);
nor UO_1841 (O_1841,N_19851,N_19542);
and UO_1842 (O_1842,N_19730,N_19544);
or UO_1843 (O_1843,N_19900,N_19690);
nand UO_1844 (O_1844,N_19558,N_19729);
nand UO_1845 (O_1845,N_19644,N_19900);
or UO_1846 (O_1846,N_19824,N_19504);
and UO_1847 (O_1847,N_19736,N_19640);
nand UO_1848 (O_1848,N_19723,N_19606);
nor UO_1849 (O_1849,N_19740,N_19772);
and UO_1850 (O_1850,N_19775,N_19596);
nor UO_1851 (O_1851,N_19501,N_19986);
xor UO_1852 (O_1852,N_19732,N_19695);
or UO_1853 (O_1853,N_19673,N_19607);
and UO_1854 (O_1854,N_19697,N_19738);
nand UO_1855 (O_1855,N_19512,N_19998);
nand UO_1856 (O_1856,N_19658,N_19729);
nor UO_1857 (O_1857,N_19572,N_19504);
and UO_1858 (O_1858,N_19958,N_19513);
nand UO_1859 (O_1859,N_19870,N_19818);
nand UO_1860 (O_1860,N_19596,N_19586);
or UO_1861 (O_1861,N_19859,N_19569);
nand UO_1862 (O_1862,N_19994,N_19724);
and UO_1863 (O_1863,N_19547,N_19678);
and UO_1864 (O_1864,N_19501,N_19774);
xnor UO_1865 (O_1865,N_19907,N_19962);
xor UO_1866 (O_1866,N_19678,N_19558);
and UO_1867 (O_1867,N_19934,N_19719);
xor UO_1868 (O_1868,N_19745,N_19986);
or UO_1869 (O_1869,N_19724,N_19595);
nor UO_1870 (O_1870,N_19806,N_19506);
nand UO_1871 (O_1871,N_19709,N_19819);
xor UO_1872 (O_1872,N_19853,N_19685);
nand UO_1873 (O_1873,N_19750,N_19704);
nand UO_1874 (O_1874,N_19559,N_19852);
or UO_1875 (O_1875,N_19548,N_19774);
nor UO_1876 (O_1876,N_19729,N_19764);
nand UO_1877 (O_1877,N_19941,N_19761);
or UO_1878 (O_1878,N_19923,N_19991);
nor UO_1879 (O_1879,N_19777,N_19691);
xor UO_1880 (O_1880,N_19817,N_19932);
nor UO_1881 (O_1881,N_19620,N_19606);
and UO_1882 (O_1882,N_19795,N_19729);
nand UO_1883 (O_1883,N_19717,N_19854);
or UO_1884 (O_1884,N_19562,N_19759);
nand UO_1885 (O_1885,N_19969,N_19691);
xor UO_1886 (O_1886,N_19564,N_19973);
nor UO_1887 (O_1887,N_19875,N_19507);
xnor UO_1888 (O_1888,N_19923,N_19593);
nand UO_1889 (O_1889,N_19753,N_19734);
and UO_1890 (O_1890,N_19961,N_19762);
and UO_1891 (O_1891,N_19728,N_19666);
nor UO_1892 (O_1892,N_19527,N_19844);
nand UO_1893 (O_1893,N_19800,N_19621);
and UO_1894 (O_1894,N_19515,N_19639);
or UO_1895 (O_1895,N_19709,N_19510);
nand UO_1896 (O_1896,N_19879,N_19639);
nor UO_1897 (O_1897,N_19873,N_19714);
and UO_1898 (O_1898,N_19540,N_19565);
nand UO_1899 (O_1899,N_19584,N_19815);
and UO_1900 (O_1900,N_19905,N_19578);
and UO_1901 (O_1901,N_19794,N_19676);
nand UO_1902 (O_1902,N_19512,N_19942);
nand UO_1903 (O_1903,N_19645,N_19535);
nand UO_1904 (O_1904,N_19568,N_19833);
or UO_1905 (O_1905,N_19710,N_19562);
xnor UO_1906 (O_1906,N_19993,N_19913);
or UO_1907 (O_1907,N_19663,N_19864);
xnor UO_1908 (O_1908,N_19633,N_19738);
and UO_1909 (O_1909,N_19912,N_19647);
nor UO_1910 (O_1910,N_19711,N_19922);
and UO_1911 (O_1911,N_19747,N_19506);
nand UO_1912 (O_1912,N_19855,N_19876);
and UO_1913 (O_1913,N_19566,N_19535);
nand UO_1914 (O_1914,N_19523,N_19785);
and UO_1915 (O_1915,N_19658,N_19952);
nand UO_1916 (O_1916,N_19773,N_19596);
or UO_1917 (O_1917,N_19536,N_19803);
and UO_1918 (O_1918,N_19856,N_19624);
nand UO_1919 (O_1919,N_19764,N_19678);
nor UO_1920 (O_1920,N_19843,N_19909);
nor UO_1921 (O_1921,N_19889,N_19968);
and UO_1922 (O_1922,N_19809,N_19655);
or UO_1923 (O_1923,N_19936,N_19969);
xor UO_1924 (O_1924,N_19878,N_19744);
nor UO_1925 (O_1925,N_19626,N_19929);
nand UO_1926 (O_1926,N_19792,N_19795);
nand UO_1927 (O_1927,N_19841,N_19743);
and UO_1928 (O_1928,N_19666,N_19762);
and UO_1929 (O_1929,N_19573,N_19925);
xnor UO_1930 (O_1930,N_19525,N_19717);
and UO_1931 (O_1931,N_19518,N_19528);
xor UO_1932 (O_1932,N_19695,N_19941);
xnor UO_1933 (O_1933,N_19940,N_19859);
nor UO_1934 (O_1934,N_19907,N_19630);
and UO_1935 (O_1935,N_19698,N_19660);
xor UO_1936 (O_1936,N_19664,N_19715);
or UO_1937 (O_1937,N_19686,N_19685);
or UO_1938 (O_1938,N_19970,N_19501);
nand UO_1939 (O_1939,N_19640,N_19713);
xor UO_1940 (O_1940,N_19751,N_19764);
nor UO_1941 (O_1941,N_19617,N_19649);
nor UO_1942 (O_1942,N_19816,N_19736);
nor UO_1943 (O_1943,N_19562,N_19923);
and UO_1944 (O_1944,N_19822,N_19796);
nor UO_1945 (O_1945,N_19942,N_19829);
and UO_1946 (O_1946,N_19590,N_19983);
nand UO_1947 (O_1947,N_19969,N_19829);
xor UO_1948 (O_1948,N_19860,N_19773);
xnor UO_1949 (O_1949,N_19701,N_19654);
or UO_1950 (O_1950,N_19691,N_19718);
xnor UO_1951 (O_1951,N_19788,N_19871);
or UO_1952 (O_1952,N_19606,N_19671);
and UO_1953 (O_1953,N_19661,N_19605);
xnor UO_1954 (O_1954,N_19616,N_19607);
xnor UO_1955 (O_1955,N_19900,N_19667);
xnor UO_1956 (O_1956,N_19668,N_19506);
or UO_1957 (O_1957,N_19577,N_19750);
xnor UO_1958 (O_1958,N_19958,N_19827);
or UO_1959 (O_1959,N_19939,N_19781);
or UO_1960 (O_1960,N_19746,N_19779);
nor UO_1961 (O_1961,N_19815,N_19629);
and UO_1962 (O_1962,N_19605,N_19852);
or UO_1963 (O_1963,N_19644,N_19549);
nand UO_1964 (O_1964,N_19587,N_19911);
nand UO_1965 (O_1965,N_19522,N_19718);
nand UO_1966 (O_1966,N_19591,N_19845);
or UO_1967 (O_1967,N_19860,N_19627);
xnor UO_1968 (O_1968,N_19573,N_19582);
and UO_1969 (O_1969,N_19787,N_19829);
nor UO_1970 (O_1970,N_19863,N_19780);
and UO_1971 (O_1971,N_19965,N_19849);
xnor UO_1972 (O_1972,N_19753,N_19554);
and UO_1973 (O_1973,N_19999,N_19627);
xor UO_1974 (O_1974,N_19686,N_19850);
nand UO_1975 (O_1975,N_19839,N_19832);
nor UO_1976 (O_1976,N_19561,N_19558);
nand UO_1977 (O_1977,N_19942,N_19778);
or UO_1978 (O_1978,N_19921,N_19902);
nor UO_1979 (O_1979,N_19911,N_19761);
nor UO_1980 (O_1980,N_19871,N_19977);
or UO_1981 (O_1981,N_19638,N_19642);
and UO_1982 (O_1982,N_19791,N_19634);
xor UO_1983 (O_1983,N_19509,N_19849);
xnor UO_1984 (O_1984,N_19889,N_19789);
or UO_1985 (O_1985,N_19643,N_19522);
and UO_1986 (O_1986,N_19945,N_19695);
and UO_1987 (O_1987,N_19785,N_19872);
xor UO_1988 (O_1988,N_19694,N_19998);
and UO_1989 (O_1989,N_19890,N_19801);
nand UO_1990 (O_1990,N_19755,N_19580);
nand UO_1991 (O_1991,N_19680,N_19607);
and UO_1992 (O_1992,N_19870,N_19752);
and UO_1993 (O_1993,N_19834,N_19713);
nor UO_1994 (O_1994,N_19976,N_19960);
nand UO_1995 (O_1995,N_19648,N_19994);
or UO_1996 (O_1996,N_19862,N_19618);
xor UO_1997 (O_1997,N_19914,N_19630);
nand UO_1998 (O_1998,N_19543,N_19559);
nor UO_1999 (O_1999,N_19725,N_19695);
xor UO_2000 (O_2000,N_19789,N_19953);
and UO_2001 (O_2001,N_19889,N_19835);
nor UO_2002 (O_2002,N_19639,N_19730);
and UO_2003 (O_2003,N_19793,N_19634);
nor UO_2004 (O_2004,N_19754,N_19935);
nor UO_2005 (O_2005,N_19731,N_19645);
xnor UO_2006 (O_2006,N_19579,N_19663);
or UO_2007 (O_2007,N_19812,N_19660);
and UO_2008 (O_2008,N_19837,N_19776);
and UO_2009 (O_2009,N_19757,N_19699);
xor UO_2010 (O_2010,N_19694,N_19990);
nand UO_2011 (O_2011,N_19556,N_19505);
nor UO_2012 (O_2012,N_19674,N_19787);
xnor UO_2013 (O_2013,N_19983,N_19688);
or UO_2014 (O_2014,N_19997,N_19582);
and UO_2015 (O_2015,N_19701,N_19625);
nand UO_2016 (O_2016,N_19701,N_19655);
nor UO_2017 (O_2017,N_19641,N_19848);
nand UO_2018 (O_2018,N_19917,N_19883);
and UO_2019 (O_2019,N_19731,N_19609);
nor UO_2020 (O_2020,N_19916,N_19672);
nand UO_2021 (O_2021,N_19568,N_19925);
or UO_2022 (O_2022,N_19778,N_19830);
nand UO_2023 (O_2023,N_19870,N_19859);
and UO_2024 (O_2024,N_19870,N_19824);
nor UO_2025 (O_2025,N_19945,N_19728);
or UO_2026 (O_2026,N_19869,N_19941);
nor UO_2027 (O_2027,N_19844,N_19587);
nand UO_2028 (O_2028,N_19939,N_19849);
or UO_2029 (O_2029,N_19988,N_19615);
nand UO_2030 (O_2030,N_19971,N_19999);
nor UO_2031 (O_2031,N_19645,N_19955);
or UO_2032 (O_2032,N_19747,N_19744);
and UO_2033 (O_2033,N_19683,N_19579);
and UO_2034 (O_2034,N_19664,N_19543);
or UO_2035 (O_2035,N_19768,N_19824);
or UO_2036 (O_2036,N_19687,N_19838);
and UO_2037 (O_2037,N_19603,N_19929);
or UO_2038 (O_2038,N_19980,N_19752);
nor UO_2039 (O_2039,N_19860,N_19985);
xor UO_2040 (O_2040,N_19728,N_19723);
or UO_2041 (O_2041,N_19631,N_19581);
and UO_2042 (O_2042,N_19725,N_19624);
and UO_2043 (O_2043,N_19917,N_19934);
xor UO_2044 (O_2044,N_19853,N_19854);
or UO_2045 (O_2045,N_19590,N_19681);
nor UO_2046 (O_2046,N_19750,N_19507);
and UO_2047 (O_2047,N_19729,N_19576);
and UO_2048 (O_2048,N_19912,N_19642);
and UO_2049 (O_2049,N_19633,N_19866);
and UO_2050 (O_2050,N_19632,N_19668);
or UO_2051 (O_2051,N_19675,N_19968);
nand UO_2052 (O_2052,N_19503,N_19974);
and UO_2053 (O_2053,N_19625,N_19996);
and UO_2054 (O_2054,N_19582,N_19987);
and UO_2055 (O_2055,N_19796,N_19504);
nor UO_2056 (O_2056,N_19737,N_19505);
nand UO_2057 (O_2057,N_19598,N_19588);
xnor UO_2058 (O_2058,N_19560,N_19768);
or UO_2059 (O_2059,N_19634,N_19672);
nand UO_2060 (O_2060,N_19608,N_19724);
nand UO_2061 (O_2061,N_19589,N_19759);
nor UO_2062 (O_2062,N_19548,N_19788);
and UO_2063 (O_2063,N_19802,N_19799);
and UO_2064 (O_2064,N_19965,N_19679);
or UO_2065 (O_2065,N_19690,N_19855);
and UO_2066 (O_2066,N_19881,N_19957);
or UO_2067 (O_2067,N_19509,N_19659);
nor UO_2068 (O_2068,N_19553,N_19915);
nand UO_2069 (O_2069,N_19833,N_19604);
and UO_2070 (O_2070,N_19996,N_19639);
nor UO_2071 (O_2071,N_19563,N_19564);
and UO_2072 (O_2072,N_19550,N_19886);
nand UO_2073 (O_2073,N_19673,N_19544);
xnor UO_2074 (O_2074,N_19598,N_19621);
xor UO_2075 (O_2075,N_19514,N_19518);
or UO_2076 (O_2076,N_19562,N_19955);
or UO_2077 (O_2077,N_19790,N_19814);
and UO_2078 (O_2078,N_19898,N_19985);
nor UO_2079 (O_2079,N_19524,N_19554);
nand UO_2080 (O_2080,N_19953,N_19688);
or UO_2081 (O_2081,N_19601,N_19755);
and UO_2082 (O_2082,N_19962,N_19739);
nor UO_2083 (O_2083,N_19642,N_19983);
nand UO_2084 (O_2084,N_19596,N_19944);
nor UO_2085 (O_2085,N_19681,N_19504);
and UO_2086 (O_2086,N_19980,N_19911);
or UO_2087 (O_2087,N_19649,N_19723);
nand UO_2088 (O_2088,N_19843,N_19678);
or UO_2089 (O_2089,N_19756,N_19657);
and UO_2090 (O_2090,N_19590,N_19520);
nand UO_2091 (O_2091,N_19729,N_19982);
and UO_2092 (O_2092,N_19528,N_19687);
nand UO_2093 (O_2093,N_19761,N_19790);
xnor UO_2094 (O_2094,N_19529,N_19780);
nand UO_2095 (O_2095,N_19705,N_19744);
and UO_2096 (O_2096,N_19933,N_19513);
nand UO_2097 (O_2097,N_19501,N_19517);
or UO_2098 (O_2098,N_19635,N_19634);
and UO_2099 (O_2099,N_19648,N_19664);
xor UO_2100 (O_2100,N_19857,N_19847);
nand UO_2101 (O_2101,N_19787,N_19736);
nand UO_2102 (O_2102,N_19987,N_19587);
and UO_2103 (O_2103,N_19919,N_19874);
nand UO_2104 (O_2104,N_19791,N_19781);
nor UO_2105 (O_2105,N_19654,N_19616);
xnor UO_2106 (O_2106,N_19855,N_19666);
xor UO_2107 (O_2107,N_19612,N_19554);
nor UO_2108 (O_2108,N_19590,N_19964);
or UO_2109 (O_2109,N_19694,N_19765);
nand UO_2110 (O_2110,N_19648,N_19867);
nor UO_2111 (O_2111,N_19548,N_19614);
xor UO_2112 (O_2112,N_19536,N_19990);
nand UO_2113 (O_2113,N_19582,N_19623);
xor UO_2114 (O_2114,N_19676,N_19637);
or UO_2115 (O_2115,N_19754,N_19584);
nand UO_2116 (O_2116,N_19746,N_19985);
nor UO_2117 (O_2117,N_19863,N_19963);
nand UO_2118 (O_2118,N_19825,N_19829);
and UO_2119 (O_2119,N_19549,N_19678);
nor UO_2120 (O_2120,N_19827,N_19974);
xor UO_2121 (O_2121,N_19654,N_19594);
or UO_2122 (O_2122,N_19647,N_19519);
nand UO_2123 (O_2123,N_19815,N_19604);
nand UO_2124 (O_2124,N_19840,N_19975);
or UO_2125 (O_2125,N_19666,N_19928);
nand UO_2126 (O_2126,N_19673,N_19502);
and UO_2127 (O_2127,N_19549,N_19905);
xnor UO_2128 (O_2128,N_19685,N_19635);
nor UO_2129 (O_2129,N_19884,N_19552);
nor UO_2130 (O_2130,N_19548,N_19847);
and UO_2131 (O_2131,N_19720,N_19544);
nor UO_2132 (O_2132,N_19504,N_19675);
nand UO_2133 (O_2133,N_19948,N_19611);
nand UO_2134 (O_2134,N_19667,N_19694);
and UO_2135 (O_2135,N_19543,N_19815);
or UO_2136 (O_2136,N_19696,N_19897);
xor UO_2137 (O_2137,N_19908,N_19777);
or UO_2138 (O_2138,N_19640,N_19563);
nor UO_2139 (O_2139,N_19937,N_19955);
nand UO_2140 (O_2140,N_19926,N_19740);
xor UO_2141 (O_2141,N_19740,N_19692);
or UO_2142 (O_2142,N_19888,N_19915);
nand UO_2143 (O_2143,N_19526,N_19987);
and UO_2144 (O_2144,N_19615,N_19608);
xor UO_2145 (O_2145,N_19823,N_19983);
xnor UO_2146 (O_2146,N_19654,N_19771);
nor UO_2147 (O_2147,N_19646,N_19950);
nor UO_2148 (O_2148,N_19827,N_19812);
nand UO_2149 (O_2149,N_19930,N_19630);
and UO_2150 (O_2150,N_19715,N_19590);
nand UO_2151 (O_2151,N_19850,N_19588);
xor UO_2152 (O_2152,N_19522,N_19571);
xnor UO_2153 (O_2153,N_19751,N_19859);
xor UO_2154 (O_2154,N_19829,N_19780);
and UO_2155 (O_2155,N_19949,N_19556);
nor UO_2156 (O_2156,N_19916,N_19732);
xnor UO_2157 (O_2157,N_19786,N_19973);
and UO_2158 (O_2158,N_19610,N_19972);
nand UO_2159 (O_2159,N_19867,N_19892);
xor UO_2160 (O_2160,N_19923,N_19915);
and UO_2161 (O_2161,N_19936,N_19722);
xor UO_2162 (O_2162,N_19848,N_19919);
xnor UO_2163 (O_2163,N_19895,N_19617);
and UO_2164 (O_2164,N_19524,N_19691);
xor UO_2165 (O_2165,N_19597,N_19871);
and UO_2166 (O_2166,N_19868,N_19789);
nor UO_2167 (O_2167,N_19963,N_19767);
and UO_2168 (O_2168,N_19527,N_19952);
and UO_2169 (O_2169,N_19741,N_19534);
or UO_2170 (O_2170,N_19699,N_19726);
or UO_2171 (O_2171,N_19627,N_19532);
nor UO_2172 (O_2172,N_19546,N_19543);
or UO_2173 (O_2173,N_19981,N_19814);
nor UO_2174 (O_2174,N_19631,N_19648);
and UO_2175 (O_2175,N_19569,N_19951);
and UO_2176 (O_2176,N_19544,N_19515);
and UO_2177 (O_2177,N_19920,N_19913);
nand UO_2178 (O_2178,N_19924,N_19755);
nand UO_2179 (O_2179,N_19635,N_19546);
and UO_2180 (O_2180,N_19572,N_19937);
or UO_2181 (O_2181,N_19678,N_19617);
xnor UO_2182 (O_2182,N_19698,N_19890);
nor UO_2183 (O_2183,N_19950,N_19791);
xor UO_2184 (O_2184,N_19586,N_19661);
or UO_2185 (O_2185,N_19607,N_19718);
and UO_2186 (O_2186,N_19922,N_19848);
xor UO_2187 (O_2187,N_19940,N_19647);
and UO_2188 (O_2188,N_19724,N_19742);
xnor UO_2189 (O_2189,N_19746,N_19542);
nand UO_2190 (O_2190,N_19571,N_19832);
or UO_2191 (O_2191,N_19976,N_19732);
nor UO_2192 (O_2192,N_19528,N_19963);
xor UO_2193 (O_2193,N_19828,N_19762);
and UO_2194 (O_2194,N_19930,N_19622);
or UO_2195 (O_2195,N_19543,N_19808);
and UO_2196 (O_2196,N_19798,N_19696);
nor UO_2197 (O_2197,N_19755,N_19878);
and UO_2198 (O_2198,N_19630,N_19651);
or UO_2199 (O_2199,N_19630,N_19572);
xnor UO_2200 (O_2200,N_19834,N_19563);
xnor UO_2201 (O_2201,N_19981,N_19789);
or UO_2202 (O_2202,N_19718,N_19565);
and UO_2203 (O_2203,N_19919,N_19527);
or UO_2204 (O_2204,N_19592,N_19723);
and UO_2205 (O_2205,N_19705,N_19507);
and UO_2206 (O_2206,N_19771,N_19845);
or UO_2207 (O_2207,N_19766,N_19793);
nor UO_2208 (O_2208,N_19647,N_19924);
nor UO_2209 (O_2209,N_19911,N_19823);
nor UO_2210 (O_2210,N_19577,N_19801);
or UO_2211 (O_2211,N_19718,N_19984);
xnor UO_2212 (O_2212,N_19946,N_19896);
nand UO_2213 (O_2213,N_19858,N_19801);
and UO_2214 (O_2214,N_19959,N_19979);
xor UO_2215 (O_2215,N_19950,N_19616);
nor UO_2216 (O_2216,N_19954,N_19604);
nor UO_2217 (O_2217,N_19691,N_19612);
nor UO_2218 (O_2218,N_19550,N_19987);
or UO_2219 (O_2219,N_19691,N_19676);
and UO_2220 (O_2220,N_19917,N_19788);
nor UO_2221 (O_2221,N_19686,N_19586);
and UO_2222 (O_2222,N_19817,N_19557);
nor UO_2223 (O_2223,N_19648,N_19953);
nor UO_2224 (O_2224,N_19879,N_19778);
and UO_2225 (O_2225,N_19760,N_19670);
nand UO_2226 (O_2226,N_19890,N_19592);
nand UO_2227 (O_2227,N_19569,N_19572);
and UO_2228 (O_2228,N_19796,N_19608);
or UO_2229 (O_2229,N_19743,N_19588);
and UO_2230 (O_2230,N_19947,N_19976);
xnor UO_2231 (O_2231,N_19869,N_19661);
nor UO_2232 (O_2232,N_19959,N_19549);
or UO_2233 (O_2233,N_19787,N_19649);
and UO_2234 (O_2234,N_19960,N_19780);
nor UO_2235 (O_2235,N_19901,N_19853);
nand UO_2236 (O_2236,N_19860,N_19858);
nor UO_2237 (O_2237,N_19968,N_19714);
xor UO_2238 (O_2238,N_19515,N_19686);
nor UO_2239 (O_2239,N_19687,N_19941);
nand UO_2240 (O_2240,N_19752,N_19621);
nand UO_2241 (O_2241,N_19832,N_19854);
nand UO_2242 (O_2242,N_19773,N_19839);
or UO_2243 (O_2243,N_19578,N_19658);
nand UO_2244 (O_2244,N_19663,N_19760);
xor UO_2245 (O_2245,N_19739,N_19732);
nor UO_2246 (O_2246,N_19664,N_19983);
nand UO_2247 (O_2247,N_19520,N_19979);
xnor UO_2248 (O_2248,N_19596,N_19804);
xor UO_2249 (O_2249,N_19707,N_19982);
nor UO_2250 (O_2250,N_19918,N_19680);
and UO_2251 (O_2251,N_19614,N_19526);
xnor UO_2252 (O_2252,N_19929,N_19910);
or UO_2253 (O_2253,N_19868,N_19806);
nand UO_2254 (O_2254,N_19856,N_19850);
xnor UO_2255 (O_2255,N_19972,N_19586);
and UO_2256 (O_2256,N_19832,N_19884);
nor UO_2257 (O_2257,N_19669,N_19888);
nor UO_2258 (O_2258,N_19693,N_19783);
xor UO_2259 (O_2259,N_19798,N_19941);
xnor UO_2260 (O_2260,N_19676,N_19714);
and UO_2261 (O_2261,N_19658,N_19727);
nor UO_2262 (O_2262,N_19899,N_19959);
or UO_2263 (O_2263,N_19996,N_19603);
and UO_2264 (O_2264,N_19649,N_19928);
and UO_2265 (O_2265,N_19629,N_19607);
nand UO_2266 (O_2266,N_19809,N_19927);
xor UO_2267 (O_2267,N_19700,N_19742);
and UO_2268 (O_2268,N_19888,N_19930);
nand UO_2269 (O_2269,N_19519,N_19733);
xnor UO_2270 (O_2270,N_19794,N_19637);
nand UO_2271 (O_2271,N_19645,N_19648);
nor UO_2272 (O_2272,N_19985,N_19832);
and UO_2273 (O_2273,N_19690,N_19649);
and UO_2274 (O_2274,N_19982,N_19943);
xor UO_2275 (O_2275,N_19839,N_19880);
xor UO_2276 (O_2276,N_19507,N_19918);
xnor UO_2277 (O_2277,N_19737,N_19862);
nand UO_2278 (O_2278,N_19721,N_19886);
xnor UO_2279 (O_2279,N_19566,N_19893);
xor UO_2280 (O_2280,N_19766,N_19505);
or UO_2281 (O_2281,N_19592,N_19608);
and UO_2282 (O_2282,N_19680,N_19799);
xor UO_2283 (O_2283,N_19973,N_19771);
or UO_2284 (O_2284,N_19756,N_19654);
nor UO_2285 (O_2285,N_19509,N_19607);
xnor UO_2286 (O_2286,N_19525,N_19668);
xor UO_2287 (O_2287,N_19597,N_19737);
nand UO_2288 (O_2288,N_19504,N_19860);
or UO_2289 (O_2289,N_19851,N_19924);
or UO_2290 (O_2290,N_19870,N_19943);
nor UO_2291 (O_2291,N_19570,N_19701);
nor UO_2292 (O_2292,N_19987,N_19712);
and UO_2293 (O_2293,N_19640,N_19801);
xnor UO_2294 (O_2294,N_19552,N_19622);
and UO_2295 (O_2295,N_19680,N_19561);
or UO_2296 (O_2296,N_19529,N_19893);
and UO_2297 (O_2297,N_19774,N_19619);
nor UO_2298 (O_2298,N_19533,N_19915);
and UO_2299 (O_2299,N_19866,N_19642);
and UO_2300 (O_2300,N_19533,N_19505);
nand UO_2301 (O_2301,N_19747,N_19712);
or UO_2302 (O_2302,N_19678,N_19582);
or UO_2303 (O_2303,N_19642,N_19993);
and UO_2304 (O_2304,N_19912,N_19890);
or UO_2305 (O_2305,N_19572,N_19995);
and UO_2306 (O_2306,N_19838,N_19662);
or UO_2307 (O_2307,N_19536,N_19519);
nand UO_2308 (O_2308,N_19986,N_19520);
or UO_2309 (O_2309,N_19579,N_19795);
and UO_2310 (O_2310,N_19951,N_19967);
nor UO_2311 (O_2311,N_19989,N_19701);
and UO_2312 (O_2312,N_19667,N_19708);
nand UO_2313 (O_2313,N_19690,N_19752);
nand UO_2314 (O_2314,N_19563,N_19886);
xnor UO_2315 (O_2315,N_19751,N_19836);
or UO_2316 (O_2316,N_19598,N_19831);
or UO_2317 (O_2317,N_19744,N_19918);
nand UO_2318 (O_2318,N_19660,N_19877);
and UO_2319 (O_2319,N_19573,N_19934);
and UO_2320 (O_2320,N_19636,N_19884);
and UO_2321 (O_2321,N_19744,N_19616);
xor UO_2322 (O_2322,N_19561,N_19518);
nor UO_2323 (O_2323,N_19748,N_19669);
nand UO_2324 (O_2324,N_19578,N_19902);
and UO_2325 (O_2325,N_19831,N_19829);
nand UO_2326 (O_2326,N_19708,N_19919);
nand UO_2327 (O_2327,N_19541,N_19918);
nor UO_2328 (O_2328,N_19742,N_19534);
or UO_2329 (O_2329,N_19681,N_19568);
and UO_2330 (O_2330,N_19767,N_19752);
nand UO_2331 (O_2331,N_19611,N_19694);
and UO_2332 (O_2332,N_19504,N_19661);
nor UO_2333 (O_2333,N_19889,N_19864);
nor UO_2334 (O_2334,N_19754,N_19988);
or UO_2335 (O_2335,N_19938,N_19738);
nand UO_2336 (O_2336,N_19527,N_19926);
nor UO_2337 (O_2337,N_19643,N_19702);
or UO_2338 (O_2338,N_19787,N_19511);
or UO_2339 (O_2339,N_19691,N_19757);
xnor UO_2340 (O_2340,N_19582,N_19925);
nor UO_2341 (O_2341,N_19552,N_19644);
nand UO_2342 (O_2342,N_19829,N_19775);
and UO_2343 (O_2343,N_19717,N_19683);
and UO_2344 (O_2344,N_19697,N_19616);
nor UO_2345 (O_2345,N_19856,N_19922);
nor UO_2346 (O_2346,N_19580,N_19739);
and UO_2347 (O_2347,N_19529,N_19888);
or UO_2348 (O_2348,N_19800,N_19928);
nor UO_2349 (O_2349,N_19936,N_19739);
and UO_2350 (O_2350,N_19557,N_19551);
xnor UO_2351 (O_2351,N_19870,N_19764);
xor UO_2352 (O_2352,N_19908,N_19658);
and UO_2353 (O_2353,N_19611,N_19882);
and UO_2354 (O_2354,N_19738,N_19850);
xnor UO_2355 (O_2355,N_19999,N_19789);
and UO_2356 (O_2356,N_19503,N_19845);
xnor UO_2357 (O_2357,N_19769,N_19855);
or UO_2358 (O_2358,N_19970,N_19841);
and UO_2359 (O_2359,N_19507,N_19825);
nand UO_2360 (O_2360,N_19629,N_19842);
nand UO_2361 (O_2361,N_19766,N_19937);
nor UO_2362 (O_2362,N_19643,N_19881);
and UO_2363 (O_2363,N_19826,N_19792);
or UO_2364 (O_2364,N_19855,N_19837);
nand UO_2365 (O_2365,N_19523,N_19840);
or UO_2366 (O_2366,N_19826,N_19911);
and UO_2367 (O_2367,N_19719,N_19858);
or UO_2368 (O_2368,N_19576,N_19914);
nand UO_2369 (O_2369,N_19705,N_19890);
nor UO_2370 (O_2370,N_19838,N_19918);
or UO_2371 (O_2371,N_19936,N_19983);
nand UO_2372 (O_2372,N_19712,N_19819);
nand UO_2373 (O_2373,N_19588,N_19911);
xor UO_2374 (O_2374,N_19837,N_19964);
xor UO_2375 (O_2375,N_19856,N_19909);
nand UO_2376 (O_2376,N_19724,N_19859);
nor UO_2377 (O_2377,N_19682,N_19762);
and UO_2378 (O_2378,N_19917,N_19990);
xnor UO_2379 (O_2379,N_19530,N_19501);
or UO_2380 (O_2380,N_19787,N_19550);
nand UO_2381 (O_2381,N_19870,N_19557);
and UO_2382 (O_2382,N_19651,N_19770);
and UO_2383 (O_2383,N_19578,N_19875);
nand UO_2384 (O_2384,N_19615,N_19515);
nor UO_2385 (O_2385,N_19530,N_19988);
nor UO_2386 (O_2386,N_19593,N_19905);
or UO_2387 (O_2387,N_19816,N_19594);
nand UO_2388 (O_2388,N_19782,N_19606);
nand UO_2389 (O_2389,N_19725,N_19939);
nor UO_2390 (O_2390,N_19970,N_19511);
or UO_2391 (O_2391,N_19995,N_19893);
nor UO_2392 (O_2392,N_19831,N_19943);
or UO_2393 (O_2393,N_19571,N_19656);
nand UO_2394 (O_2394,N_19915,N_19560);
xnor UO_2395 (O_2395,N_19986,N_19673);
nor UO_2396 (O_2396,N_19504,N_19592);
nor UO_2397 (O_2397,N_19765,N_19656);
and UO_2398 (O_2398,N_19679,N_19784);
xor UO_2399 (O_2399,N_19915,N_19536);
nor UO_2400 (O_2400,N_19671,N_19509);
nand UO_2401 (O_2401,N_19900,N_19719);
or UO_2402 (O_2402,N_19703,N_19618);
or UO_2403 (O_2403,N_19970,N_19971);
nor UO_2404 (O_2404,N_19828,N_19673);
or UO_2405 (O_2405,N_19662,N_19617);
nor UO_2406 (O_2406,N_19762,N_19746);
nor UO_2407 (O_2407,N_19932,N_19754);
nand UO_2408 (O_2408,N_19910,N_19722);
and UO_2409 (O_2409,N_19860,N_19975);
nor UO_2410 (O_2410,N_19679,N_19816);
and UO_2411 (O_2411,N_19803,N_19681);
or UO_2412 (O_2412,N_19643,N_19964);
nand UO_2413 (O_2413,N_19787,N_19850);
and UO_2414 (O_2414,N_19906,N_19770);
nor UO_2415 (O_2415,N_19653,N_19885);
xnor UO_2416 (O_2416,N_19622,N_19645);
and UO_2417 (O_2417,N_19865,N_19896);
nor UO_2418 (O_2418,N_19754,N_19683);
xor UO_2419 (O_2419,N_19753,N_19775);
or UO_2420 (O_2420,N_19774,N_19560);
xnor UO_2421 (O_2421,N_19704,N_19521);
nand UO_2422 (O_2422,N_19807,N_19919);
or UO_2423 (O_2423,N_19642,N_19734);
or UO_2424 (O_2424,N_19690,N_19906);
nor UO_2425 (O_2425,N_19530,N_19856);
nand UO_2426 (O_2426,N_19642,N_19896);
nor UO_2427 (O_2427,N_19538,N_19562);
xor UO_2428 (O_2428,N_19715,N_19571);
xor UO_2429 (O_2429,N_19870,N_19756);
xor UO_2430 (O_2430,N_19618,N_19593);
and UO_2431 (O_2431,N_19700,N_19597);
and UO_2432 (O_2432,N_19942,N_19744);
nand UO_2433 (O_2433,N_19549,N_19822);
and UO_2434 (O_2434,N_19857,N_19580);
nand UO_2435 (O_2435,N_19896,N_19815);
xor UO_2436 (O_2436,N_19766,N_19992);
nand UO_2437 (O_2437,N_19530,N_19566);
xnor UO_2438 (O_2438,N_19655,N_19871);
or UO_2439 (O_2439,N_19705,N_19864);
nand UO_2440 (O_2440,N_19630,N_19655);
or UO_2441 (O_2441,N_19987,N_19552);
or UO_2442 (O_2442,N_19795,N_19886);
nor UO_2443 (O_2443,N_19545,N_19615);
and UO_2444 (O_2444,N_19706,N_19733);
nand UO_2445 (O_2445,N_19503,N_19818);
and UO_2446 (O_2446,N_19716,N_19765);
xor UO_2447 (O_2447,N_19626,N_19771);
and UO_2448 (O_2448,N_19912,N_19735);
and UO_2449 (O_2449,N_19708,N_19972);
nand UO_2450 (O_2450,N_19743,N_19640);
xor UO_2451 (O_2451,N_19994,N_19777);
and UO_2452 (O_2452,N_19756,N_19878);
or UO_2453 (O_2453,N_19892,N_19876);
nand UO_2454 (O_2454,N_19960,N_19922);
or UO_2455 (O_2455,N_19865,N_19563);
or UO_2456 (O_2456,N_19876,N_19860);
xnor UO_2457 (O_2457,N_19974,N_19786);
and UO_2458 (O_2458,N_19542,N_19812);
and UO_2459 (O_2459,N_19832,N_19702);
xor UO_2460 (O_2460,N_19738,N_19728);
nor UO_2461 (O_2461,N_19874,N_19653);
xor UO_2462 (O_2462,N_19726,N_19665);
and UO_2463 (O_2463,N_19996,N_19885);
nand UO_2464 (O_2464,N_19617,N_19741);
xor UO_2465 (O_2465,N_19550,N_19932);
nor UO_2466 (O_2466,N_19970,N_19530);
nor UO_2467 (O_2467,N_19687,N_19955);
xor UO_2468 (O_2468,N_19692,N_19867);
nor UO_2469 (O_2469,N_19663,N_19931);
nand UO_2470 (O_2470,N_19991,N_19838);
nand UO_2471 (O_2471,N_19838,N_19655);
nand UO_2472 (O_2472,N_19699,N_19571);
or UO_2473 (O_2473,N_19813,N_19722);
xnor UO_2474 (O_2474,N_19543,N_19899);
or UO_2475 (O_2475,N_19738,N_19531);
nand UO_2476 (O_2476,N_19839,N_19596);
xnor UO_2477 (O_2477,N_19882,N_19595);
xnor UO_2478 (O_2478,N_19561,N_19513);
xnor UO_2479 (O_2479,N_19901,N_19592);
and UO_2480 (O_2480,N_19747,N_19765);
and UO_2481 (O_2481,N_19677,N_19702);
nor UO_2482 (O_2482,N_19941,N_19632);
or UO_2483 (O_2483,N_19592,N_19719);
xor UO_2484 (O_2484,N_19564,N_19812);
nand UO_2485 (O_2485,N_19524,N_19851);
nor UO_2486 (O_2486,N_19748,N_19910);
nor UO_2487 (O_2487,N_19598,N_19786);
and UO_2488 (O_2488,N_19881,N_19503);
xnor UO_2489 (O_2489,N_19918,N_19879);
nor UO_2490 (O_2490,N_19586,N_19659);
nor UO_2491 (O_2491,N_19633,N_19723);
xnor UO_2492 (O_2492,N_19711,N_19817);
or UO_2493 (O_2493,N_19784,N_19653);
or UO_2494 (O_2494,N_19640,N_19587);
nor UO_2495 (O_2495,N_19572,N_19838);
nand UO_2496 (O_2496,N_19659,N_19742);
nand UO_2497 (O_2497,N_19527,N_19939);
nand UO_2498 (O_2498,N_19597,N_19893);
nor UO_2499 (O_2499,N_19807,N_19806);
endmodule