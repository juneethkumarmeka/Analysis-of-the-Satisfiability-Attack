module basic_500_3000_500_5_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_23,In_60);
and U1 (N_1,In_3,In_340);
and U2 (N_2,In_469,In_35);
xor U3 (N_3,In_363,In_359);
xnor U4 (N_4,In_374,In_16);
nand U5 (N_5,In_241,In_314);
nor U6 (N_6,In_437,In_422);
nand U7 (N_7,In_85,In_4);
and U8 (N_8,In_13,In_455);
xor U9 (N_9,In_235,In_337);
xor U10 (N_10,In_398,In_321);
nor U11 (N_11,In_343,In_308);
nand U12 (N_12,In_388,In_458);
nor U13 (N_13,In_21,In_475);
and U14 (N_14,In_147,In_58);
xor U15 (N_15,In_394,In_356);
and U16 (N_16,In_223,In_200);
or U17 (N_17,In_297,In_492);
nand U18 (N_18,In_282,In_432);
xor U19 (N_19,In_357,In_375);
or U20 (N_20,In_38,In_79);
nand U21 (N_21,In_157,In_392);
nor U22 (N_22,In_336,In_345);
or U23 (N_23,In_73,In_350);
and U24 (N_24,In_248,In_286);
nand U25 (N_25,In_454,In_252);
and U26 (N_26,In_414,In_180);
and U27 (N_27,In_50,In_203);
nand U28 (N_28,In_197,In_333);
nor U29 (N_29,In_277,In_22);
xnor U30 (N_30,In_349,In_331);
and U31 (N_31,In_423,In_54);
or U32 (N_32,In_80,In_284);
and U33 (N_33,In_471,In_249);
xor U34 (N_34,In_225,In_191);
nand U35 (N_35,In_227,In_199);
xor U36 (N_36,In_364,In_419);
and U37 (N_37,In_353,In_450);
nor U38 (N_38,In_294,In_233);
and U39 (N_39,In_135,In_186);
xnor U40 (N_40,In_125,In_228);
or U41 (N_41,In_189,In_445);
xnor U42 (N_42,In_303,In_202);
xnor U43 (N_43,In_290,In_372);
or U44 (N_44,In_209,In_32);
nor U45 (N_45,In_236,In_92);
xor U46 (N_46,In_103,In_190);
xnor U47 (N_47,In_102,In_401);
nand U48 (N_48,In_255,In_481);
or U49 (N_49,In_212,In_399);
nor U50 (N_50,In_110,In_421);
and U51 (N_51,In_172,In_114);
nor U52 (N_52,In_55,In_376);
nand U53 (N_53,In_335,In_355);
nand U54 (N_54,In_330,In_63);
xor U55 (N_55,In_247,In_380);
xor U56 (N_56,In_149,In_497);
nor U57 (N_57,In_251,In_459);
nor U58 (N_58,In_90,In_354);
nand U59 (N_59,In_105,In_24);
nor U60 (N_60,In_461,In_295);
and U61 (N_61,In_265,In_438);
and U62 (N_62,In_358,In_31);
nand U63 (N_63,In_278,In_153);
or U64 (N_64,In_62,In_28);
nand U65 (N_65,In_178,In_325);
or U66 (N_66,In_317,In_442);
nor U67 (N_67,In_309,In_133);
nand U68 (N_68,In_8,In_86);
and U69 (N_69,In_107,In_371);
or U70 (N_70,In_74,In_47);
nor U71 (N_71,In_143,In_491);
nor U72 (N_72,In_395,In_166);
or U73 (N_73,In_272,In_379);
and U74 (N_74,In_45,In_118);
xor U75 (N_75,In_342,In_188);
nand U76 (N_76,In_232,In_257);
or U77 (N_77,In_390,In_430);
or U78 (N_78,In_222,In_307);
xor U79 (N_79,In_57,In_254);
and U80 (N_80,In_37,In_383);
and U81 (N_81,In_221,In_75);
xnor U82 (N_82,In_56,In_361);
and U83 (N_83,In_77,In_476);
nor U84 (N_84,In_96,In_88);
or U85 (N_85,In_283,In_44);
xnor U86 (N_86,In_391,In_453);
xor U87 (N_87,In_404,In_240);
nand U88 (N_88,In_245,In_39);
nand U89 (N_89,In_29,In_1);
nand U90 (N_90,In_387,In_137);
or U91 (N_91,In_216,In_368);
and U92 (N_92,In_348,In_490);
and U93 (N_93,In_229,In_250);
nand U94 (N_94,In_136,In_301);
nor U95 (N_95,In_402,In_464);
nor U96 (N_96,In_17,In_433);
nor U97 (N_97,In_279,In_385);
nor U98 (N_98,In_470,In_124);
and U99 (N_99,In_167,In_319);
nor U100 (N_100,In_264,In_488);
or U101 (N_101,In_129,In_381);
and U102 (N_102,In_489,In_367);
or U103 (N_103,In_195,In_138);
nor U104 (N_104,In_498,In_253);
or U105 (N_105,In_20,In_177);
and U106 (N_106,In_462,In_302);
nand U107 (N_107,In_465,In_448);
or U108 (N_108,In_121,In_169);
or U109 (N_109,In_292,In_425);
nand U110 (N_110,In_173,In_76);
or U111 (N_111,In_436,In_41);
nand U112 (N_112,In_256,In_494);
or U113 (N_113,In_420,In_408);
nand U114 (N_114,In_226,In_196);
nand U115 (N_115,In_18,In_6);
nand U116 (N_116,In_144,In_119);
nand U117 (N_117,In_171,In_26);
nand U118 (N_118,In_217,In_34);
nor U119 (N_119,In_496,In_456);
nor U120 (N_120,In_134,In_327);
nand U121 (N_121,In_472,In_40);
or U122 (N_122,In_94,In_441);
xnor U123 (N_123,In_140,In_106);
nor U124 (N_124,In_128,In_15);
xnor U125 (N_125,In_5,In_71);
nor U126 (N_126,In_260,In_478);
and U127 (N_127,In_27,In_271);
nor U128 (N_128,In_116,In_243);
nor U129 (N_129,In_224,In_266);
and U130 (N_130,In_127,In_187);
nor U131 (N_131,In_182,In_304);
xnor U132 (N_132,In_377,In_446);
xnor U133 (N_133,In_431,In_281);
or U134 (N_134,In_113,In_296);
nor U135 (N_135,In_82,In_474);
nor U136 (N_136,In_122,In_261);
nor U137 (N_137,In_440,In_139);
and U138 (N_138,In_429,In_305);
and U139 (N_139,In_65,In_104);
xor U140 (N_140,In_287,In_146);
or U141 (N_141,In_11,In_347);
or U142 (N_142,In_231,In_163);
or U143 (N_143,In_389,In_101);
or U144 (N_144,In_397,In_403);
and U145 (N_145,In_141,In_148);
nor U146 (N_146,In_480,In_318);
nor U147 (N_147,In_328,In_154);
nand U148 (N_148,In_210,In_275);
and U149 (N_149,In_482,In_93);
nand U150 (N_150,In_53,In_449);
or U151 (N_151,In_338,In_213);
and U152 (N_152,In_108,In_426);
nor U153 (N_153,In_352,In_42);
nand U154 (N_154,In_365,In_83);
or U155 (N_155,In_244,In_176);
nand U156 (N_156,In_0,In_51);
nand U157 (N_157,In_259,In_384);
xor U158 (N_158,In_393,In_211);
or U159 (N_159,In_405,In_111);
xor U160 (N_160,In_386,In_326);
xnor U161 (N_161,In_312,In_234);
or U162 (N_162,In_165,In_64);
and U163 (N_163,In_413,In_242);
xnor U164 (N_164,In_68,In_300);
or U165 (N_165,In_61,In_276);
nor U166 (N_166,In_214,In_72);
or U167 (N_167,In_201,In_451);
xor U168 (N_168,In_117,In_293);
nor U169 (N_169,In_258,In_427);
or U170 (N_170,In_473,In_7);
and U171 (N_171,In_483,In_142);
xnor U172 (N_172,In_369,In_130);
or U173 (N_173,In_14,In_181);
nor U174 (N_174,In_444,In_168);
and U175 (N_175,In_69,In_269);
or U176 (N_176,In_329,In_230);
xnor U177 (N_177,In_208,In_334);
nor U178 (N_178,In_12,In_132);
nand U179 (N_179,In_493,In_339);
nor U180 (N_180,In_467,In_10);
xnor U181 (N_181,In_48,In_268);
nor U182 (N_182,In_316,In_237);
and U183 (N_183,In_486,In_164);
or U184 (N_184,In_443,In_263);
or U185 (N_185,In_434,In_49);
nor U186 (N_186,In_78,In_324);
or U187 (N_187,In_158,In_417);
or U188 (N_188,In_170,In_306);
nor U189 (N_189,In_206,In_299);
or U190 (N_190,In_332,In_485);
nor U191 (N_191,In_362,In_46);
and U192 (N_192,In_499,In_313);
nand U193 (N_193,In_484,In_98);
xnor U194 (N_194,In_59,In_289);
and U195 (N_195,In_315,In_406);
nand U196 (N_196,In_320,In_407);
or U197 (N_197,In_366,In_207);
or U198 (N_198,In_447,In_220);
nand U199 (N_199,In_30,In_311);
and U200 (N_200,In_487,In_288);
or U201 (N_201,In_161,In_145);
nor U202 (N_202,In_95,In_174);
and U203 (N_203,In_468,In_457);
and U204 (N_204,In_400,In_452);
xor U205 (N_205,In_378,In_370);
xnor U206 (N_206,In_115,In_109);
xnor U207 (N_207,In_322,In_418);
or U208 (N_208,In_151,In_218);
and U209 (N_209,In_123,In_131);
xor U210 (N_210,In_185,In_495);
or U211 (N_211,In_175,In_100);
nor U212 (N_212,In_9,In_238);
nand U213 (N_213,In_463,In_156);
nand U214 (N_214,In_89,In_25);
xnor U215 (N_215,In_193,In_97);
nor U216 (N_216,In_262,In_298);
nor U217 (N_217,In_411,In_194);
and U218 (N_218,In_183,In_219);
or U219 (N_219,In_162,In_382);
nor U220 (N_220,In_310,In_460);
nand U221 (N_221,In_155,In_435);
nor U222 (N_222,In_415,In_477);
and U223 (N_223,In_184,In_291);
or U224 (N_224,In_466,In_152);
nor U225 (N_225,In_160,In_341);
nor U226 (N_226,In_360,In_412);
and U227 (N_227,In_112,In_205);
nand U228 (N_228,In_274,In_19);
nand U229 (N_229,In_239,In_215);
xnor U230 (N_230,In_285,In_43);
xnor U231 (N_231,In_81,In_280);
or U232 (N_232,In_428,In_409);
and U233 (N_233,In_273,In_36);
and U234 (N_234,In_410,In_2);
or U235 (N_235,In_351,In_99);
or U236 (N_236,In_67,In_267);
and U237 (N_237,In_91,In_323);
or U238 (N_238,In_150,In_204);
nand U239 (N_239,In_424,In_87);
nand U240 (N_240,In_52,In_396);
xor U241 (N_241,In_70,In_346);
nand U242 (N_242,In_373,In_33);
nor U243 (N_243,In_344,In_246);
nand U244 (N_244,In_159,In_439);
and U245 (N_245,In_479,In_66);
nand U246 (N_246,In_270,In_120);
xnor U247 (N_247,In_416,In_84);
nand U248 (N_248,In_126,In_179);
nor U249 (N_249,In_192,In_198);
nand U250 (N_250,In_137,In_140);
xor U251 (N_251,In_124,In_137);
or U252 (N_252,In_190,In_388);
xor U253 (N_253,In_65,In_424);
nor U254 (N_254,In_473,In_439);
or U255 (N_255,In_64,In_55);
nand U256 (N_256,In_195,In_115);
nand U257 (N_257,In_127,In_13);
xor U258 (N_258,In_196,In_411);
nor U259 (N_259,In_300,In_474);
or U260 (N_260,In_455,In_348);
nand U261 (N_261,In_486,In_29);
or U262 (N_262,In_482,In_259);
nand U263 (N_263,In_122,In_73);
or U264 (N_264,In_175,In_380);
nand U265 (N_265,In_213,In_180);
and U266 (N_266,In_378,In_429);
xnor U267 (N_267,In_55,In_77);
and U268 (N_268,In_404,In_111);
and U269 (N_269,In_408,In_452);
xor U270 (N_270,In_354,In_232);
nor U271 (N_271,In_402,In_442);
or U272 (N_272,In_19,In_114);
nand U273 (N_273,In_346,In_218);
nand U274 (N_274,In_241,In_257);
or U275 (N_275,In_423,In_425);
xnor U276 (N_276,In_33,In_289);
nand U277 (N_277,In_260,In_367);
xor U278 (N_278,In_449,In_387);
and U279 (N_279,In_387,In_173);
and U280 (N_280,In_83,In_493);
or U281 (N_281,In_210,In_182);
nand U282 (N_282,In_153,In_98);
nand U283 (N_283,In_471,In_47);
or U284 (N_284,In_248,In_11);
nand U285 (N_285,In_419,In_336);
and U286 (N_286,In_464,In_377);
and U287 (N_287,In_308,In_495);
and U288 (N_288,In_395,In_486);
or U289 (N_289,In_106,In_14);
or U290 (N_290,In_99,In_220);
nor U291 (N_291,In_425,In_284);
xnor U292 (N_292,In_198,In_240);
nand U293 (N_293,In_445,In_94);
or U294 (N_294,In_283,In_146);
and U295 (N_295,In_414,In_457);
and U296 (N_296,In_100,In_464);
and U297 (N_297,In_286,In_53);
xor U298 (N_298,In_164,In_188);
xor U299 (N_299,In_372,In_34);
or U300 (N_300,In_384,In_201);
or U301 (N_301,In_454,In_484);
or U302 (N_302,In_201,In_360);
nor U303 (N_303,In_178,In_87);
nand U304 (N_304,In_40,In_313);
or U305 (N_305,In_452,In_395);
xnor U306 (N_306,In_175,In_361);
or U307 (N_307,In_78,In_23);
xnor U308 (N_308,In_135,In_206);
xor U309 (N_309,In_143,In_248);
nor U310 (N_310,In_199,In_289);
xnor U311 (N_311,In_197,In_365);
xnor U312 (N_312,In_149,In_318);
xnor U313 (N_313,In_239,In_46);
nor U314 (N_314,In_315,In_140);
xor U315 (N_315,In_454,In_277);
xnor U316 (N_316,In_272,In_403);
xor U317 (N_317,In_8,In_352);
nand U318 (N_318,In_111,In_309);
xor U319 (N_319,In_248,In_42);
nor U320 (N_320,In_189,In_28);
nor U321 (N_321,In_11,In_318);
nor U322 (N_322,In_327,In_177);
and U323 (N_323,In_440,In_137);
nand U324 (N_324,In_344,In_4);
and U325 (N_325,In_267,In_216);
or U326 (N_326,In_240,In_47);
and U327 (N_327,In_268,In_138);
and U328 (N_328,In_406,In_177);
and U329 (N_329,In_411,In_310);
xnor U330 (N_330,In_415,In_105);
or U331 (N_331,In_186,In_156);
and U332 (N_332,In_486,In_305);
and U333 (N_333,In_420,In_174);
nor U334 (N_334,In_338,In_50);
nand U335 (N_335,In_208,In_155);
xnor U336 (N_336,In_418,In_317);
and U337 (N_337,In_124,In_319);
nor U338 (N_338,In_375,In_421);
xor U339 (N_339,In_110,In_19);
xor U340 (N_340,In_349,In_444);
xnor U341 (N_341,In_66,In_420);
or U342 (N_342,In_59,In_61);
xor U343 (N_343,In_244,In_360);
xnor U344 (N_344,In_405,In_166);
and U345 (N_345,In_91,In_80);
or U346 (N_346,In_280,In_326);
and U347 (N_347,In_175,In_407);
nor U348 (N_348,In_305,In_64);
nor U349 (N_349,In_129,In_366);
or U350 (N_350,In_52,In_158);
and U351 (N_351,In_189,In_394);
or U352 (N_352,In_131,In_486);
nor U353 (N_353,In_209,In_369);
xor U354 (N_354,In_458,In_299);
or U355 (N_355,In_258,In_144);
or U356 (N_356,In_201,In_229);
nand U357 (N_357,In_351,In_84);
or U358 (N_358,In_174,In_138);
or U359 (N_359,In_254,In_243);
nand U360 (N_360,In_121,In_440);
nor U361 (N_361,In_397,In_12);
nand U362 (N_362,In_335,In_470);
nor U363 (N_363,In_191,In_306);
nor U364 (N_364,In_415,In_417);
xnor U365 (N_365,In_218,In_415);
nand U366 (N_366,In_361,In_415);
nor U367 (N_367,In_495,In_195);
or U368 (N_368,In_468,In_34);
or U369 (N_369,In_385,In_388);
or U370 (N_370,In_156,In_26);
nor U371 (N_371,In_407,In_231);
xor U372 (N_372,In_346,In_138);
xor U373 (N_373,In_24,In_433);
and U374 (N_374,In_353,In_206);
or U375 (N_375,In_95,In_331);
and U376 (N_376,In_26,In_110);
or U377 (N_377,In_471,In_312);
nand U378 (N_378,In_474,In_9);
xnor U379 (N_379,In_244,In_296);
and U380 (N_380,In_194,In_187);
and U381 (N_381,In_391,In_272);
or U382 (N_382,In_490,In_190);
nor U383 (N_383,In_152,In_312);
and U384 (N_384,In_110,In_246);
nor U385 (N_385,In_65,In_355);
and U386 (N_386,In_68,In_330);
xnor U387 (N_387,In_384,In_483);
nand U388 (N_388,In_274,In_328);
or U389 (N_389,In_168,In_43);
nand U390 (N_390,In_457,In_462);
nand U391 (N_391,In_42,In_272);
or U392 (N_392,In_168,In_380);
or U393 (N_393,In_138,In_441);
and U394 (N_394,In_94,In_324);
or U395 (N_395,In_31,In_237);
and U396 (N_396,In_306,In_173);
or U397 (N_397,In_51,In_498);
nand U398 (N_398,In_483,In_406);
or U399 (N_399,In_155,In_24);
and U400 (N_400,In_167,In_151);
or U401 (N_401,In_440,In_456);
nand U402 (N_402,In_375,In_252);
or U403 (N_403,In_16,In_237);
xor U404 (N_404,In_450,In_172);
or U405 (N_405,In_146,In_257);
nand U406 (N_406,In_363,In_33);
or U407 (N_407,In_106,In_71);
xor U408 (N_408,In_51,In_312);
and U409 (N_409,In_55,In_325);
nor U410 (N_410,In_396,In_169);
nand U411 (N_411,In_351,In_93);
nor U412 (N_412,In_375,In_176);
nand U413 (N_413,In_85,In_452);
xor U414 (N_414,In_229,In_276);
and U415 (N_415,In_253,In_97);
nor U416 (N_416,In_195,In_314);
and U417 (N_417,In_270,In_327);
or U418 (N_418,In_305,In_108);
xnor U419 (N_419,In_152,In_285);
xor U420 (N_420,In_486,In_111);
xnor U421 (N_421,In_366,In_345);
xnor U422 (N_422,In_363,In_499);
and U423 (N_423,In_488,In_254);
or U424 (N_424,In_409,In_281);
and U425 (N_425,In_25,In_491);
and U426 (N_426,In_121,In_177);
nor U427 (N_427,In_64,In_2);
or U428 (N_428,In_303,In_298);
and U429 (N_429,In_456,In_120);
xor U430 (N_430,In_351,In_378);
and U431 (N_431,In_55,In_265);
nor U432 (N_432,In_370,In_428);
nand U433 (N_433,In_251,In_380);
or U434 (N_434,In_89,In_485);
or U435 (N_435,In_382,In_40);
xor U436 (N_436,In_15,In_132);
nor U437 (N_437,In_246,In_173);
or U438 (N_438,In_273,In_162);
or U439 (N_439,In_468,In_274);
xor U440 (N_440,In_413,In_340);
xor U441 (N_441,In_478,In_19);
nor U442 (N_442,In_338,In_395);
nor U443 (N_443,In_164,In_161);
nor U444 (N_444,In_270,In_28);
or U445 (N_445,In_326,In_359);
nand U446 (N_446,In_282,In_461);
xnor U447 (N_447,In_372,In_64);
or U448 (N_448,In_201,In_442);
nor U449 (N_449,In_150,In_476);
xor U450 (N_450,In_353,In_98);
or U451 (N_451,In_378,In_45);
nor U452 (N_452,In_308,In_458);
or U453 (N_453,In_132,In_473);
nor U454 (N_454,In_30,In_242);
nand U455 (N_455,In_342,In_429);
nand U456 (N_456,In_139,In_74);
or U457 (N_457,In_5,In_308);
or U458 (N_458,In_300,In_497);
nand U459 (N_459,In_281,In_54);
and U460 (N_460,In_117,In_437);
xor U461 (N_461,In_461,In_276);
nand U462 (N_462,In_493,In_205);
or U463 (N_463,In_402,In_195);
or U464 (N_464,In_244,In_378);
xor U465 (N_465,In_221,In_459);
nor U466 (N_466,In_121,In_279);
or U467 (N_467,In_215,In_48);
and U468 (N_468,In_254,In_100);
or U469 (N_469,In_209,In_393);
xnor U470 (N_470,In_410,In_489);
nand U471 (N_471,In_273,In_432);
xor U472 (N_472,In_365,In_305);
xnor U473 (N_473,In_264,In_185);
or U474 (N_474,In_53,In_495);
xnor U475 (N_475,In_322,In_351);
nand U476 (N_476,In_109,In_132);
and U477 (N_477,In_237,In_244);
nand U478 (N_478,In_210,In_172);
nor U479 (N_479,In_334,In_271);
xor U480 (N_480,In_422,In_229);
nand U481 (N_481,In_490,In_495);
or U482 (N_482,In_274,In_488);
or U483 (N_483,In_101,In_357);
or U484 (N_484,In_488,In_280);
or U485 (N_485,In_3,In_169);
nor U486 (N_486,In_22,In_352);
and U487 (N_487,In_317,In_401);
xor U488 (N_488,In_52,In_341);
and U489 (N_489,In_208,In_306);
or U490 (N_490,In_82,In_321);
nor U491 (N_491,In_396,In_170);
xnor U492 (N_492,In_157,In_76);
and U493 (N_493,In_481,In_120);
and U494 (N_494,In_441,In_493);
nor U495 (N_495,In_393,In_49);
and U496 (N_496,In_432,In_96);
and U497 (N_497,In_450,In_231);
nand U498 (N_498,In_473,In_90);
nor U499 (N_499,In_310,In_207);
nor U500 (N_500,In_14,In_494);
xor U501 (N_501,In_245,In_112);
and U502 (N_502,In_366,In_121);
xor U503 (N_503,In_404,In_243);
nor U504 (N_504,In_323,In_475);
nand U505 (N_505,In_176,In_207);
or U506 (N_506,In_249,In_82);
nand U507 (N_507,In_149,In_464);
or U508 (N_508,In_15,In_110);
nand U509 (N_509,In_107,In_53);
or U510 (N_510,In_193,In_269);
or U511 (N_511,In_482,In_231);
xor U512 (N_512,In_122,In_25);
and U513 (N_513,In_47,In_95);
nand U514 (N_514,In_401,In_98);
and U515 (N_515,In_72,In_294);
and U516 (N_516,In_23,In_386);
nand U517 (N_517,In_196,In_62);
and U518 (N_518,In_130,In_463);
nand U519 (N_519,In_419,In_471);
and U520 (N_520,In_178,In_81);
and U521 (N_521,In_162,In_294);
xnor U522 (N_522,In_142,In_162);
and U523 (N_523,In_211,In_249);
and U524 (N_524,In_458,In_103);
nor U525 (N_525,In_121,In_252);
xnor U526 (N_526,In_179,In_22);
nor U527 (N_527,In_97,In_38);
and U528 (N_528,In_409,In_113);
or U529 (N_529,In_429,In_130);
nand U530 (N_530,In_271,In_431);
nand U531 (N_531,In_437,In_308);
or U532 (N_532,In_444,In_67);
nor U533 (N_533,In_214,In_254);
xor U534 (N_534,In_182,In_389);
nor U535 (N_535,In_271,In_28);
nand U536 (N_536,In_382,In_86);
nor U537 (N_537,In_320,In_165);
nand U538 (N_538,In_486,In_258);
or U539 (N_539,In_62,In_246);
nor U540 (N_540,In_64,In_209);
or U541 (N_541,In_262,In_103);
xor U542 (N_542,In_134,In_278);
nor U543 (N_543,In_261,In_147);
xor U544 (N_544,In_26,In_34);
and U545 (N_545,In_432,In_471);
nand U546 (N_546,In_328,In_159);
nand U547 (N_547,In_146,In_73);
nor U548 (N_548,In_125,In_73);
nor U549 (N_549,In_282,In_471);
nand U550 (N_550,In_481,In_218);
nand U551 (N_551,In_342,In_281);
nor U552 (N_552,In_383,In_488);
and U553 (N_553,In_29,In_35);
nand U554 (N_554,In_408,In_497);
nor U555 (N_555,In_110,In_273);
xnor U556 (N_556,In_28,In_111);
nand U557 (N_557,In_312,In_224);
nor U558 (N_558,In_94,In_322);
and U559 (N_559,In_4,In_433);
and U560 (N_560,In_352,In_482);
nor U561 (N_561,In_152,In_157);
or U562 (N_562,In_249,In_42);
nor U563 (N_563,In_188,In_286);
xnor U564 (N_564,In_120,In_11);
xor U565 (N_565,In_366,In_410);
nor U566 (N_566,In_253,In_320);
xnor U567 (N_567,In_64,In_283);
nand U568 (N_568,In_389,In_24);
nand U569 (N_569,In_75,In_329);
nand U570 (N_570,In_249,In_309);
nor U571 (N_571,In_218,In_246);
and U572 (N_572,In_96,In_256);
xor U573 (N_573,In_111,In_202);
xor U574 (N_574,In_499,In_325);
and U575 (N_575,In_142,In_229);
xor U576 (N_576,In_181,In_494);
xnor U577 (N_577,In_207,In_27);
nor U578 (N_578,In_257,In_23);
xnor U579 (N_579,In_41,In_453);
and U580 (N_580,In_182,In_85);
nand U581 (N_581,In_442,In_315);
and U582 (N_582,In_162,In_172);
and U583 (N_583,In_60,In_377);
or U584 (N_584,In_296,In_294);
and U585 (N_585,In_199,In_438);
xor U586 (N_586,In_302,In_206);
nor U587 (N_587,In_247,In_128);
and U588 (N_588,In_84,In_379);
and U589 (N_589,In_303,In_278);
or U590 (N_590,In_249,In_107);
xor U591 (N_591,In_262,In_388);
and U592 (N_592,In_251,In_222);
nor U593 (N_593,In_193,In_425);
nor U594 (N_594,In_83,In_105);
nor U595 (N_595,In_49,In_98);
nand U596 (N_596,In_10,In_37);
xnor U597 (N_597,In_205,In_272);
and U598 (N_598,In_266,In_454);
and U599 (N_599,In_345,In_297);
nand U600 (N_600,N_558,N_510);
or U601 (N_601,N_591,N_341);
nand U602 (N_602,N_163,N_251);
and U603 (N_603,N_226,N_441);
and U604 (N_604,N_314,N_373);
nor U605 (N_605,N_426,N_91);
nand U606 (N_606,N_492,N_130);
xor U607 (N_607,N_168,N_361);
nor U608 (N_608,N_449,N_384);
or U609 (N_609,N_436,N_556);
or U610 (N_610,N_470,N_356);
or U611 (N_611,N_348,N_520);
and U612 (N_612,N_273,N_67);
nor U613 (N_613,N_178,N_458);
and U614 (N_614,N_391,N_491);
xnor U615 (N_615,N_206,N_244);
and U616 (N_616,N_599,N_537);
or U617 (N_617,N_62,N_408);
or U618 (N_618,N_228,N_462);
nor U619 (N_619,N_561,N_197);
nor U620 (N_620,N_464,N_306);
and U621 (N_621,N_380,N_64);
xnor U622 (N_622,N_192,N_574);
xor U623 (N_623,N_302,N_446);
and U624 (N_624,N_499,N_291);
nor U625 (N_625,N_53,N_220);
nor U626 (N_626,N_20,N_75);
nor U627 (N_627,N_587,N_444);
nand U628 (N_628,N_171,N_214);
nand U629 (N_629,N_532,N_198);
xor U630 (N_630,N_9,N_116);
and U631 (N_631,N_478,N_114);
xor U632 (N_632,N_109,N_547);
or U633 (N_633,N_177,N_418);
and U634 (N_634,N_248,N_594);
xnor U635 (N_635,N_593,N_259);
or U636 (N_636,N_503,N_311);
and U637 (N_637,N_488,N_284);
nor U638 (N_638,N_400,N_346);
and U639 (N_639,N_298,N_103);
xnor U640 (N_640,N_497,N_100);
or U641 (N_641,N_385,N_49);
xor U642 (N_642,N_158,N_337);
nor U643 (N_643,N_199,N_12);
and U644 (N_644,N_227,N_598);
and U645 (N_645,N_370,N_122);
nor U646 (N_646,N_76,N_288);
and U647 (N_647,N_552,N_534);
xnor U648 (N_648,N_369,N_50);
nand U649 (N_649,N_434,N_303);
nor U650 (N_650,N_476,N_51);
and U651 (N_651,N_16,N_512);
and U652 (N_652,N_359,N_94);
xor U653 (N_653,N_554,N_580);
or U654 (N_654,N_24,N_431);
or U655 (N_655,N_0,N_107);
nor U656 (N_656,N_527,N_98);
or U657 (N_657,N_521,N_536);
xor U658 (N_658,N_42,N_13);
xnor U659 (N_659,N_252,N_204);
and U660 (N_660,N_422,N_238);
or U661 (N_661,N_209,N_225);
xnor U662 (N_662,N_115,N_48);
nor U663 (N_663,N_516,N_125);
and U664 (N_664,N_166,N_132);
or U665 (N_665,N_597,N_404);
or U666 (N_666,N_23,N_278);
nor U667 (N_667,N_84,N_515);
and U668 (N_668,N_283,N_395);
xnor U669 (N_669,N_567,N_221);
nand U670 (N_670,N_232,N_455);
xnor U671 (N_671,N_445,N_352);
and U672 (N_672,N_242,N_34);
nand U673 (N_673,N_54,N_293);
and U674 (N_674,N_79,N_501);
nand U675 (N_675,N_148,N_172);
and U676 (N_676,N_190,N_454);
xor U677 (N_677,N_36,N_8);
and U678 (N_678,N_301,N_154);
and U679 (N_679,N_41,N_2);
or U680 (N_680,N_280,N_363);
or U681 (N_681,N_43,N_571);
or U682 (N_682,N_263,N_10);
xnor U683 (N_683,N_572,N_200);
xnor U684 (N_684,N_429,N_405);
nand U685 (N_685,N_474,N_270);
and U686 (N_686,N_272,N_72);
and U687 (N_687,N_268,N_297);
nor U688 (N_688,N_469,N_87);
nand U689 (N_689,N_86,N_229);
nand U690 (N_690,N_120,N_504);
nor U691 (N_691,N_265,N_425);
and U692 (N_692,N_165,N_292);
and U693 (N_693,N_279,N_447);
and U694 (N_694,N_397,N_26);
nand U695 (N_695,N_421,N_322);
nand U696 (N_696,N_312,N_456);
nor U697 (N_697,N_457,N_159);
nor U698 (N_698,N_490,N_17);
xor U699 (N_699,N_459,N_411);
and U700 (N_700,N_505,N_546);
nor U701 (N_701,N_553,N_393);
nor U702 (N_702,N_151,N_117);
nand U703 (N_703,N_30,N_285);
nand U704 (N_704,N_290,N_379);
nand U705 (N_705,N_473,N_477);
xnor U706 (N_706,N_60,N_95);
nor U707 (N_707,N_557,N_174);
xnor U708 (N_708,N_568,N_1);
xnor U709 (N_709,N_362,N_465);
xnor U710 (N_710,N_440,N_489);
or U711 (N_711,N_157,N_208);
nor U712 (N_712,N_129,N_354);
nor U713 (N_713,N_245,N_123);
xnor U714 (N_714,N_300,N_155);
nand U715 (N_715,N_482,N_186);
and U716 (N_716,N_216,N_68);
nand U717 (N_717,N_576,N_224);
or U718 (N_718,N_21,N_413);
nand U719 (N_719,N_182,N_328);
and U720 (N_720,N_309,N_203);
nand U721 (N_721,N_383,N_99);
nand U722 (N_722,N_142,N_540);
nor U723 (N_723,N_565,N_78);
xor U724 (N_724,N_506,N_46);
and U725 (N_725,N_551,N_110);
or U726 (N_726,N_342,N_333);
or U727 (N_727,N_202,N_69);
nor U728 (N_728,N_136,N_73);
and U729 (N_729,N_65,N_88);
or U730 (N_730,N_357,N_315);
nor U731 (N_731,N_187,N_524);
xor U732 (N_732,N_555,N_351);
nor U733 (N_733,N_170,N_101);
xor U734 (N_734,N_543,N_570);
and U735 (N_735,N_71,N_294);
or U736 (N_736,N_52,N_105);
nor U737 (N_737,N_525,N_541);
or U738 (N_738,N_326,N_338);
nor U739 (N_739,N_28,N_164);
nor U740 (N_740,N_127,N_276);
nand U741 (N_741,N_485,N_509);
and U742 (N_742,N_40,N_448);
nand U743 (N_743,N_254,N_247);
or U744 (N_744,N_264,N_592);
xnor U745 (N_745,N_266,N_585);
and U746 (N_746,N_223,N_365);
nor U747 (N_747,N_304,N_511);
nand U748 (N_748,N_63,N_234);
xor U749 (N_749,N_37,N_336);
nor U750 (N_750,N_210,N_82);
or U751 (N_751,N_387,N_167);
or U752 (N_752,N_205,N_233);
or U753 (N_753,N_415,N_212);
nor U754 (N_754,N_514,N_286);
and U755 (N_755,N_324,N_250);
or U756 (N_756,N_414,N_193);
nor U757 (N_757,N_6,N_44);
or U758 (N_758,N_584,N_378);
nor U759 (N_759,N_231,N_427);
xnor U760 (N_760,N_409,N_45);
nor U761 (N_761,N_494,N_5);
and U762 (N_762,N_70,N_496);
nor U763 (N_763,N_452,N_329);
nand U764 (N_764,N_310,N_138);
xor U765 (N_765,N_175,N_81);
xnor U766 (N_766,N_194,N_150);
and U767 (N_767,N_360,N_295);
nand U768 (N_768,N_530,N_323);
nand U769 (N_769,N_239,N_305);
nor U770 (N_770,N_230,N_219);
nand U771 (N_771,N_89,N_97);
nand U772 (N_772,N_35,N_108);
nor U773 (N_773,N_519,N_240);
nand U774 (N_774,N_472,N_577);
nand U775 (N_775,N_131,N_569);
and U776 (N_776,N_389,N_267);
and U777 (N_777,N_113,N_358);
nor U778 (N_778,N_334,N_195);
nand U779 (N_779,N_595,N_134);
nand U780 (N_780,N_33,N_140);
and U781 (N_781,N_327,N_162);
nand U782 (N_782,N_590,N_83);
nand U783 (N_783,N_382,N_237);
nor U784 (N_784,N_77,N_102);
xor U785 (N_785,N_392,N_390);
or U786 (N_786,N_588,N_517);
or U787 (N_787,N_374,N_544);
and U788 (N_788,N_161,N_246);
or U789 (N_789,N_14,N_181);
nor U790 (N_790,N_4,N_339);
or U791 (N_791,N_596,N_112);
nor U792 (N_792,N_451,N_15);
and U793 (N_793,N_586,N_169);
nand U794 (N_794,N_11,N_453);
nand U795 (N_795,N_461,N_296);
xnor U796 (N_796,N_345,N_307);
and U797 (N_797,N_367,N_92);
xnor U798 (N_798,N_176,N_319);
nor U799 (N_799,N_443,N_545);
xor U800 (N_800,N_287,N_381);
nand U801 (N_801,N_261,N_529);
and U802 (N_802,N_344,N_222);
xor U803 (N_803,N_406,N_371);
nand U804 (N_804,N_428,N_139);
and U805 (N_805,N_350,N_317);
or U806 (N_806,N_523,N_249);
xnor U807 (N_807,N_217,N_179);
or U808 (N_808,N_468,N_548);
nand U809 (N_809,N_398,N_106);
nor U810 (N_810,N_564,N_236);
and U811 (N_811,N_299,N_111);
nor U812 (N_812,N_213,N_375);
and U813 (N_813,N_423,N_320);
xnor U814 (N_814,N_258,N_364);
nor U815 (N_815,N_59,N_372);
nand U816 (N_816,N_119,N_573);
and U817 (N_817,N_253,N_442);
nand U818 (N_818,N_533,N_47);
nand U819 (N_819,N_18,N_563);
xnor U820 (N_820,N_416,N_522);
nor U821 (N_821,N_57,N_402);
nor U822 (N_822,N_156,N_526);
xnor U823 (N_823,N_347,N_579);
and U824 (N_824,N_463,N_85);
nor U825 (N_825,N_152,N_7);
nor U826 (N_826,N_466,N_211);
xnor U827 (N_827,N_349,N_135);
nor U828 (N_828,N_407,N_316);
or U829 (N_829,N_438,N_196);
nand U830 (N_830,N_321,N_22);
and U831 (N_831,N_386,N_493);
and U832 (N_832,N_332,N_289);
xnor U833 (N_833,N_325,N_61);
xnor U834 (N_834,N_330,N_417);
nand U835 (N_835,N_39,N_589);
xor U836 (N_836,N_483,N_508);
xor U837 (N_837,N_235,N_262);
xor U838 (N_838,N_495,N_126);
nor U839 (N_839,N_366,N_388);
and U840 (N_840,N_394,N_96);
nor U841 (N_841,N_137,N_583);
nor U842 (N_842,N_318,N_58);
or U843 (N_843,N_355,N_104);
xnor U844 (N_844,N_368,N_19);
and U845 (N_845,N_184,N_180);
xnor U846 (N_846,N_343,N_403);
xnor U847 (N_847,N_513,N_188);
and U848 (N_848,N_149,N_582);
nand U849 (N_849,N_260,N_479);
nor U850 (N_850,N_502,N_189);
nand U851 (N_851,N_118,N_562);
and U852 (N_852,N_401,N_218);
nand U853 (N_853,N_215,N_38);
xnor U854 (N_854,N_450,N_183);
and U855 (N_855,N_433,N_141);
nand U856 (N_856,N_420,N_308);
xor U857 (N_857,N_128,N_550);
nor U858 (N_858,N_575,N_331);
or U859 (N_859,N_274,N_549);
and U860 (N_860,N_507,N_437);
nand U861 (N_861,N_281,N_93);
or U862 (N_862,N_145,N_207);
or U863 (N_863,N_256,N_313);
nand U864 (N_864,N_124,N_29);
xor U865 (N_865,N_412,N_335);
nand U866 (N_866,N_255,N_144);
nor U867 (N_867,N_484,N_498);
and U868 (N_868,N_377,N_282);
nand U869 (N_869,N_31,N_143);
nand U870 (N_870,N_340,N_424);
nand U871 (N_871,N_185,N_535);
nor U872 (N_872,N_539,N_578);
and U873 (N_873,N_471,N_3);
nor U874 (N_874,N_410,N_160);
or U875 (N_875,N_32,N_481);
xnor U876 (N_876,N_56,N_475);
xnor U877 (N_877,N_153,N_542);
and U878 (N_878,N_538,N_90);
nand U879 (N_879,N_66,N_500);
nand U880 (N_880,N_419,N_243);
and U881 (N_881,N_133,N_257);
nand U882 (N_882,N_173,N_121);
nor U883 (N_883,N_376,N_432);
or U884 (N_884,N_241,N_269);
or U885 (N_885,N_191,N_25);
xor U886 (N_886,N_467,N_147);
nor U887 (N_887,N_396,N_271);
and U888 (N_888,N_80,N_55);
or U889 (N_889,N_460,N_480);
xnor U890 (N_890,N_435,N_581);
nor U891 (N_891,N_528,N_439);
and U892 (N_892,N_566,N_487);
xor U893 (N_893,N_531,N_399);
nand U894 (N_894,N_518,N_146);
nor U895 (N_895,N_277,N_560);
nand U896 (N_896,N_201,N_27);
or U897 (N_897,N_275,N_353);
or U898 (N_898,N_74,N_486);
nor U899 (N_899,N_559,N_430);
nor U900 (N_900,N_129,N_117);
nor U901 (N_901,N_36,N_358);
xnor U902 (N_902,N_522,N_107);
nand U903 (N_903,N_547,N_598);
xor U904 (N_904,N_469,N_143);
nand U905 (N_905,N_286,N_105);
nand U906 (N_906,N_224,N_470);
xor U907 (N_907,N_496,N_28);
xor U908 (N_908,N_278,N_298);
and U909 (N_909,N_407,N_181);
or U910 (N_910,N_519,N_162);
nor U911 (N_911,N_7,N_251);
xnor U912 (N_912,N_136,N_489);
or U913 (N_913,N_3,N_300);
nand U914 (N_914,N_197,N_168);
xnor U915 (N_915,N_137,N_415);
or U916 (N_916,N_313,N_476);
or U917 (N_917,N_332,N_394);
nor U918 (N_918,N_350,N_61);
or U919 (N_919,N_55,N_50);
nand U920 (N_920,N_40,N_17);
nor U921 (N_921,N_399,N_212);
nand U922 (N_922,N_399,N_374);
or U923 (N_923,N_362,N_378);
nand U924 (N_924,N_210,N_111);
nand U925 (N_925,N_483,N_538);
or U926 (N_926,N_379,N_31);
xnor U927 (N_927,N_453,N_275);
nor U928 (N_928,N_423,N_76);
nor U929 (N_929,N_561,N_196);
nor U930 (N_930,N_430,N_337);
and U931 (N_931,N_186,N_67);
nand U932 (N_932,N_468,N_118);
nand U933 (N_933,N_330,N_338);
xor U934 (N_934,N_568,N_526);
or U935 (N_935,N_320,N_160);
or U936 (N_936,N_594,N_102);
xor U937 (N_937,N_314,N_463);
nand U938 (N_938,N_588,N_29);
xnor U939 (N_939,N_186,N_266);
and U940 (N_940,N_169,N_488);
and U941 (N_941,N_565,N_452);
nor U942 (N_942,N_186,N_398);
nor U943 (N_943,N_342,N_588);
or U944 (N_944,N_326,N_147);
nand U945 (N_945,N_48,N_166);
and U946 (N_946,N_314,N_591);
xnor U947 (N_947,N_506,N_164);
nand U948 (N_948,N_411,N_139);
xnor U949 (N_949,N_343,N_586);
nand U950 (N_950,N_402,N_430);
nor U951 (N_951,N_78,N_589);
nor U952 (N_952,N_19,N_120);
nor U953 (N_953,N_222,N_117);
xor U954 (N_954,N_23,N_144);
nor U955 (N_955,N_140,N_265);
and U956 (N_956,N_272,N_259);
nand U957 (N_957,N_563,N_103);
nor U958 (N_958,N_328,N_86);
and U959 (N_959,N_284,N_579);
nor U960 (N_960,N_528,N_381);
nor U961 (N_961,N_565,N_538);
xor U962 (N_962,N_541,N_536);
or U963 (N_963,N_441,N_83);
nand U964 (N_964,N_349,N_272);
and U965 (N_965,N_121,N_91);
and U966 (N_966,N_341,N_255);
xnor U967 (N_967,N_128,N_355);
and U968 (N_968,N_91,N_133);
xnor U969 (N_969,N_60,N_466);
and U970 (N_970,N_499,N_198);
or U971 (N_971,N_103,N_74);
and U972 (N_972,N_525,N_593);
or U973 (N_973,N_122,N_124);
nor U974 (N_974,N_263,N_115);
or U975 (N_975,N_555,N_334);
xnor U976 (N_976,N_528,N_294);
nand U977 (N_977,N_397,N_448);
nand U978 (N_978,N_225,N_456);
or U979 (N_979,N_325,N_217);
and U980 (N_980,N_437,N_500);
or U981 (N_981,N_57,N_131);
or U982 (N_982,N_512,N_205);
or U983 (N_983,N_546,N_34);
and U984 (N_984,N_45,N_274);
or U985 (N_985,N_125,N_525);
nand U986 (N_986,N_508,N_507);
and U987 (N_987,N_326,N_539);
xor U988 (N_988,N_502,N_43);
xnor U989 (N_989,N_293,N_539);
nor U990 (N_990,N_597,N_113);
nor U991 (N_991,N_375,N_522);
or U992 (N_992,N_361,N_140);
nor U993 (N_993,N_24,N_34);
nor U994 (N_994,N_86,N_238);
or U995 (N_995,N_32,N_312);
nor U996 (N_996,N_373,N_368);
or U997 (N_997,N_478,N_248);
and U998 (N_998,N_79,N_292);
nand U999 (N_999,N_24,N_544);
nor U1000 (N_1000,N_270,N_443);
or U1001 (N_1001,N_51,N_32);
nand U1002 (N_1002,N_35,N_177);
nand U1003 (N_1003,N_13,N_165);
or U1004 (N_1004,N_153,N_523);
xnor U1005 (N_1005,N_351,N_451);
nand U1006 (N_1006,N_589,N_105);
nand U1007 (N_1007,N_158,N_224);
xor U1008 (N_1008,N_330,N_17);
and U1009 (N_1009,N_148,N_210);
nor U1010 (N_1010,N_165,N_87);
xnor U1011 (N_1011,N_182,N_545);
and U1012 (N_1012,N_357,N_594);
xnor U1013 (N_1013,N_103,N_31);
or U1014 (N_1014,N_569,N_396);
xnor U1015 (N_1015,N_257,N_48);
xnor U1016 (N_1016,N_383,N_375);
nand U1017 (N_1017,N_318,N_342);
and U1018 (N_1018,N_53,N_90);
nor U1019 (N_1019,N_279,N_398);
and U1020 (N_1020,N_281,N_508);
xor U1021 (N_1021,N_296,N_530);
nor U1022 (N_1022,N_497,N_281);
xnor U1023 (N_1023,N_212,N_325);
xnor U1024 (N_1024,N_576,N_553);
and U1025 (N_1025,N_25,N_71);
and U1026 (N_1026,N_379,N_70);
nor U1027 (N_1027,N_69,N_492);
and U1028 (N_1028,N_146,N_223);
nand U1029 (N_1029,N_255,N_138);
nand U1030 (N_1030,N_121,N_59);
nor U1031 (N_1031,N_511,N_521);
or U1032 (N_1032,N_332,N_159);
xnor U1033 (N_1033,N_514,N_308);
nand U1034 (N_1034,N_383,N_309);
nand U1035 (N_1035,N_0,N_84);
nor U1036 (N_1036,N_451,N_273);
and U1037 (N_1037,N_259,N_38);
and U1038 (N_1038,N_152,N_154);
xor U1039 (N_1039,N_569,N_326);
xor U1040 (N_1040,N_383,N_270);
xor U1041 (N_1041,N_285,N_374);
xnor U1042 (N_1042,N_472,N_126);
nand U1043 (N_1043,N_377,N_297);
or U1044 (N_1044,N_158,N_504);
nor U1045 (N_1045,N_466,N_308);
xor U1046 (N_1046,N_596,N_501);
xor U1047 (N_1047,N_213,N_24);
xor U1048 (N_1048,N_193,N_87);
or U1049 (N_1049,N_496,N_464);
xnor U1050 (N_1050,N_164,N_270);
and U1051 (N_1051,N_159,N_434);
and U1052 (N_1052,N_440,N_178);
or U1053 (N_1053,N_216,N_453);
nand U1054 (N_1054,N_4,N_254);
nand U1055 (N_1055,N_486,N_372);
nor U1056 (N_1056,N_57,N_525);
and U1057 (N_1057,N_183,N_269);
nor U1058 (N_1058,N_214,N_270);
nand U1059 (N_1059,N_169,N_406);
nand U1060 (N_1060,N_534,N_236);
nor U1061 (N_1061,N_351,N_100);
and U1062 (N_1062,N_557,N_302);
or U1063 (N_1063,N_341,N_479);
nor U1064 (N_1064,N_141,N_414);
nor U1065 (N_1065,N_67,N_193);
and U1066 (N_1066,N_547,N_131);
nand U1067 (N_1067,N_127,N_61);
nand U1068 (N_1068,N_195,N_124);
nor U1069 (N_1069,N_403,N_599);
xnor U1070 (N_1070,N_262,N_284);
or U1071 (N_1071,N_9,N_434);
nor U1072 (N_1072,N_248,N_102);
and U1073 (N_1073,N_426,N_403);
or U1074 (N_1074,N_252,N_545);
or U1075 (N_1075,N_425,N_466);
nand U1076 (N_1076,N_542,N_547);
or U1077 (N_1077,N_485,N_53);
or U1078 (N_1078,N_443,N_1);
or U1079 (N_1079,N_365,N_563);
or U1080 (N_1080,N_588,N_140);
or U1081 (N_1081,N_144,N_465);
xnor U1082 (N_1082,N_39,N_527);
xor U1083 (N_1083,N_394,N_80);
xor U1084 (N_1084,N_187,N_22);
and U1085 (N_1085,N_535,N_152);
and U1086 (N_1086,N_372,N_293);
nand U1087 (N_1087,N_179,N_186);
xnor U1088 (N_1088,N_546,N_213);
nor U1089 (N_1089,N_129,N_46);
nor U1090 (N_1090,N_532,N_372);
or U1091 (N_1091,N_329,N_119);
nand U1092 (N_1092,N_37,N_467);
nand U1093 (N_1093,N_40,N_354);
nor U1094 (N_1094,N_511,N_368);
nand U1095 (N_1095,N_410,N_413);
nand U1096 (N_1096,N_495,N_114);
or U1097 (N_1097,N_406,N_44);
and U1098 (N_1098,N_38,N_39);
and U1099 (N_1099,N_174,N_508);
nand U1100 (N_1100,N_164,N_569);
xnor U1101 (N_1101,N_11,N_570);
or U1102 (N_1102,N_161,N_191);
xnor U1103 (N_1103,N_295,N_452);
nor U1104 (N_1104,N_380,N_76);
xnor U1105 (N_1105,N_541,N_385);
nor U1106 (N_1106,N_596,N_181);
nand U1107 (N_1107,N_333,N_574);
nor U1108 (N_1108,N_502,N_426);
and U1109 (N_1109,N_42,N_547);
or U1110 (N_1110,N_151,N_347);
xnor U1111 (N_1111,N_18,N_535);
xnor U1112 (N_1112,N_230,N_245);
nor U1113 (N_1113,N_198,N_247);
nand U1114 (N_1114,N_330,N_597);
nor U1115 (N_1115,N_484,N_185);
xnor U1116 (N_1116,N_428,N_33);
and U1117 (N_1117,N_523,N_420);
or U1118 (N_1118,N_156,N_486);
xnor U1119 (N_1119,N_211,N_353);
xnor U1120 (N_1120,N_39,N_253);
nand U1121 (N_1121,N_74,N_210);
nor U1122 (N_1122,N_506,N_106);
xnor U1123 (N_1123,N_355,N_588);
nand U1124 (N_1124,N_388,N_457);
xor U1125 (N_1125,N_258,N_145);
nand U1126 (N_1126,N_104,N_221);
and U1127 (N_1127,N_428,N_412);
nand U1128 (N_1128,N_68,N_423);
and U1129 (N_1129,N_335,N_256);
nor U1130 (N_1130,N_227,N_143);
or U1131 (N_1131,N_254,N_474);
nor U1132 (N_1132,N_190,N_262);
nor U1133 (N_1133,N_247,N_517);
and U1134 (N_1134,N_54,N_168);
xnor U1135 (N_1135,N_488,N_94);
nand U1136 (N_1136,N_431,N_333);
or U1137 (N_1137,N_349,N_202);
nor U1138 (N_1138,N_564,N_334);
and U1139 (N_1139,N_53,N_66);
nor U1140 (N_1140,N_212,N_39);
nor U1141 (N_1141,N_121,N_495);
xor U1142 (N_1142,N_72,N_594);
xnor U1143 (N_1143,N_82,N_237);
xor U1144 (N_1144,N_598,N_265);
and U1145 (N_1145,N_64,N_405);
nand U1146 (N_1146,N_446,N_433);
nor U1147 (N_1147,N_591,N_380);
nand U1148 (N_1148,N_246,N_563);
xor U1149 (N_1149,N_64,N_340);
nor U1150 (N_1150,N_282,N_456);
nor U1151 (N_1151,N_446,N_544);
xnor U1152 (N_1152,N_588,N_310);
and U1153 (N_1153,N_543,N_553);
or U1154 (N_1154,N_168,N_8);
nand U1155 (N_1155,N_587,N_250);
nor U1156 (N_1156,N_426,N_47);
and U1157 (N_1157,N_403,N_488);
or U1158 (N_1158,N_203,N_109);
nand U1159 (N_1159,N_110,N_86);
nor U1160 (N_1160,N_202,N_85);
nor U1161 (N_1161,N_0,N_317);
and U1162 (N_1162,N_362,N_369);
nor U1163 (N_1163,N_335,N_279);
or U1164 (N_1164,N_221,N_86);
xor U1165 (N_1165,N_30,N_142);
nand U1166 (N_1166,N_328,N_84);
nand U1167 (N_1167,N_42,N_139);
xnor U1168 (N_1168,N_208,N_49);
nor U1169 (N_1169,N_598,N_189);
and U1170 (N_1170,N_201,N_97);
nand U1171 (N_1171,N_167,N_19);
xnor U1172 (N_1172,N_407,N_473);
nor U1173 (N_1173,N_222,N_230);
and U1174 (N_1174,N_413,N_231);
and U1175 (N_1175,N_380,N_517);
nand U1176 (N_1176,N_59,N_432);
nor U1177 (N_1177,N_7,N_232);
xor U1178 (N_1178,N_287,N_117);
xor U1179 (N_1179,N_103,N_439);
nor U1180 (N_1180,N_116,N_422);
xor U1181 (N_1181,N_483,N_158);
or U1182 (N_1182,N_482,N_489);
or U1183 (N_1183,N_289,N_213);
and U1184 (N_1184,N_227,N_55);
nand U1185 (N_1185,N_214,N_160);
nand U1186 (N_1186,N_80,N_531);
nand U1187 (N_1187,N_248,N_3);
nor U1188 (N_1188,N_566,N_312);
or U1189 (N_1189,N_256,N_226);
nand U1190 (N_1190,N_172,N_405);
nor U1191 (N_1191,N_508,N_411);
and U1192 (N_1192,N_204,N_78);
and U1193 (N_1193,N_419,N_138);
nand U1194 (N_1194,N_7,N_49);
nor U1195 (N_1195,N_182,N_53);
or U1196 (N_1196,N_324,N_288);
and U1197 (N_1197,N_497,N_140);
xor U1198 (N_1198,N_514,N_254);
or U1199 (N_1199,N_32,N_189);
and U1200 (N_1200,N_886,N_987);
or U1201 (N_1201,N_760,N_660);
xnor U1202 (N_1202,N_875,N_1102);
nor U1203 (N_1203,N_611,N_1041);
or U1204 (N_1204,N_787,N_945);
nor U1205 (N_1205,N_967,N_754);
nand U1206 (N_1206,N_642,N_778);
nor U1207 (N_1207,N_1087,N_624);
xnor U1208 (N_1208,N_691,N_688);
nor U1209 (N_1209,N_932,N_1017);
and U1210 (N_1210,N_783,N_654);
and U1211 (N_1211,N_1177,N_813);
or U1212 (N_1212,N_679,N_906);
xnor U1213 (N_1213,N_904,N_990);
nand U1214 (N_1214,N_801,N_1168);
and U1215 (N_1215,N_730,N_795);
xnor U1216 (N_1216,N_829,N_820);
nand U1217 (N_1217,N_1110,N_839);
nor U1218 (N_1218,N_805,N_712);
and U1219 (N_1219,N_616,N_1165);
xnor U1220 (N_1220,N_786,N_713);
nand U1221 (N_1221,N_1016,N_1149);
nand U1222 (N_1222,N_800,N_812);
nand U1223 (N_1223,N_880,N_1069);
nor U1224 (N_1224,N_608,N_1019);
or U1225 (N_1225,N_793,N_975);
nand U1226 (N_1226,N_698,N_1009);
and U1227 (N_1227,N_752,N_872);
and U1228 (N_1228,N_935,N_825);
xnor U1229 (N_1229,N_1072,N_857);
xnor U1230 (N_1230,N_1088,N_741);
nand U1231 (N_1231,N_923,N_1022);
or U1232 (N_1232,N_629,N_956);
or U1233 (N_1233,N_764,N_876);
or U1234 (N_1234,N_621,N_1008);
or U1235 (N_1235,N_613,N_1151);
xnor U1236 (N_1236,N_1095,N_1150);
and U1237 (N_1237,N_1040,N_748);
and U1238 (N_1238,N_1125,N_1006);
and U1239 (N_1239,N_1047,N_1011);
xor U1240 (N_1240,N_732,N_1045);
and U1241 (N_1241,N_1052,N_1014);
or U1242 (N_1242,N_1198,N_1145);
nor U1243 (N_1243,N_803,N_757);
nand U1244 (N_1244,N_668,N_1178);
nand U1245 (N_1245,N_731,N_1174);
nand U1246 (N_1246,N_1156,N_1042);
nor U1247 (N_1247,N_905,N_949);
nand U1248 (N_1248,N_1085,N_1160);
xor U1249 (N_1249,N_742,N_1187);
xor U1250 (N_1250,N_995,N_1070);
nor U1251 (N_1251,N_948,N_677);
nor U1252 (N_1252,N_648,N_1065);
and U1253 (N_1253,N_1073,N_902);
xor U1254 (N_1254,N_1054,N_1028);
and U1255 (N_1255,N_609,N_808);
xor U1256 (N_1256,N_766,N_950);
or U1257 (N_1257,N_1137,N_806);
and U1258 (N_1258,N_1034,N_627);
xnor U1259 (N_1259,N_844,N_958);
nor U1260 (N_1260,N_765,N_969);
and U1261 (N_1261,N_607,N_894);
or U1262 (N_1262,N_964,N_926);
or U1263 (N_1263,N_965,N_650);
or U1264 (N_1264,N_1029,N_637);
nand U1265 (N_1265,N_1184,N_702);
xor U1266 (N_1266,N_780,N_723);
and U1267 (N_1267,N_1051,N_606);
xnor U1268 (N_1268,N_867,N_919);
and U1269 (N_1269,N_604,N_998);
xnor U1270 (N_1270,N_635,N_913);
nor U1271 (N_1271,N_705,N_916);
nor U1272 (N_1272,N_751,N_799);
or U1273 (N_1273,N_1062,N_1119);
or U1274 (N_1274,N_911,N_846);
xor U1275 (N_1275,N_893,N_1079);
or U1276 (N_1276,N_976,N_849);
xnor U1277 (N_1277,N_756,N_1130);
nand U1278 (N_1278,N_737,N_827);
nor U1279 (N_1279,N_1159,N_983);
xor U1280 (N_1280,N_640,N_877);
xnor U1281 (N_1281,N_822,N_678);
and U1282 (N_1282,N_1005,N_670);
or U1283 (N_1283,N_687,N_692);
and U1284 (N_1284,N_796,N_666);
and U1285 (N_1285,N_1092,N_716);
nor U1286 (N_1286,N_667,N_689);
and U1287 (N_1287,N_781,N_1024);
and U1288 (N_1288,N_963,N_866);
or U1289 (N_1289,N_745,N_1173);
or U1290 (N_1290,N_1025,N_665);
or U1291 (N_1291,N_1190,N_1170);
nand U1292 (N_1292,N_854,N_868);
xor U1293 (N_1293,N_1185,N_934);
nand U1294 (N_1294,N_736,N_1060);
nand U1295 (N_1295,N_1131,N_818);
and U1296 (N_1296,N_770,N_978);
nand U1297 (N_1297,N_763,N_651);
xor U1298 (N_1298,N_649,N_862);
nand U1299 (N_1299,N_1192,N_1002);
nor U1300 (N_1300,N_993,N_628);
xnor U1301 (N_1301,N_907,N_643);
or U1302 (N_1302,N_1138,N_882);
or U1303 (N_1303,N_631,N_722);
xor U1304 (N_1304,N_682,N_797);
nand U1305 (N_1305,N_869,N_623);
and U1306 (N_1306,N_1031,N_852);
nand U1307 (N_1307,N_727,N_746);
or U1308 (N_1308,N_1124,N_603);
or U1309 (N_1309,N_618,N_903);
nand U1310 (N_1310,N_632,N_1157);
or U1311 (N_1311,N_938,N_1020);
and U1312 (N_1312,N_755,N_881);
nor U1313 (N_1313,N_1193,N_657);
and U1314 (N_1314,N_1147,N_895);
xor U1315 (N_1315,N_735,N_826);
nor U1316 (N_1316,N_962,N_1012);
xor U1317 (N_1317,N_1115,N_1000);
and U1318 (N_1318,N_762,N_814);
nand U1319 (N_1319,N_817,N_1148);
nor U1320 (N_1320,N_873,N_997);
xnor U1321 (N_1321,N_974,N_1169);
nor U1322 (N_1322,N_870,N_810);
or U1323 (N_1323,N_798,N_714);
xnor U1324 (N_1324,N_848,N_734);
nand U1325 (N_1325,N_1021,N_715);
and U1326 (N_1326,N_675,N_972);
xnor U1327 (N_1327,N_749,N_1143);
and U1328 (N_1328,N_920,N_851);
nor U1329 (N_1329,N_1161,N_874);
or U1330 (N_1330,N_710,N_837);
and U1331 (N_1331,N_1057,N_1037);
and U1332 (N_1332,N_791,N_811);
nand U1333 (N_1333,N_693,N_720);
nand U1334 (N_1334,N_1194,N_1081);
nor U1335 (N_1335,N_1050,N_1077);
xnor U1336 (N_1336,N_685,N_761);
xor U1337 (N_1337,N_733,N_973);
xnor U1338 (N_1338,N_871,N_1126);
nor U1339 (N_1339,N_680,N_992);
or U1340 (N_1340,N_636,N_831);
nand U1341 (N_1341,N_1096,N_991);
nand U1342 (N_1342,N_684,N_909);
nand U1343 (N_1343,N_697,N_729);
xor U1344 (N_1344,N_612,N_1053);
nand U1345 (N_1345,N_1139,N_790);
nand U1346 (N_1346,N_1090,N_999);
nand U1347 (N_1347,N_1015,N_1172);
or U1348 (N_1348,N_901,N_841);
nand U1349 (N_1349,N_985,N_1084);
nor U1350 (N_1350,N_785,N_1082);
nor U1351 (N_1351,N_1108,N_1196);
xor U1352 (N_1352,N_704,N_878);
nand U1353 (N_1353,N_759,N_928);
nand U1354 (N_1354,N_726,N_1046);
xnor U1355 (N_1355,N_840,N_966);
xor U1356 (N_1356,N_833,N_1061);
nand U1357 (N_1357,N_1106,N_674);
xor U1358 (N_1358,N_921,N_937);
and U1359 (N_1359,N_1128,N_695);
xnor U1360 (N_1360,N_1063,N_1167);
and U1361 (N_1361,N_753,N_700);
xnor U1362 (N_1362,N_951,N_1121);
nor U1363 (N_1363,N_625,N_669);
or U1364 (N_1364,N_750,N_955);
and U1365 (N_1365,N_1117,N_673);
nor U1366 (N_1366,N_725,N_979);
xor U1367 (N_1367,N_1109,N_1036);
nand U1368 (N_1368,N_1097,N_931);
xnor U1369 (N_1369,N_896,N_602);
nor U1370 (N_1370,N_619,N_924);
nand U1371 (N_1371,N_672,N_952);
nand U1372 (N_1372,N_816,N_860);
nor U1373 (N_1373,N_626,N_828);
nor U1374 (N_1374,N_696,N_659);
or U1375 (N_1375,N_970,N_912);
nand U1376 (N_1376,N_947,N_789);
or U1377 (N_1377,N_929,N_1166);
or U1378 (N_1378,N_815,N_863);
and U1379 (N_1379,N_996,N_888);
nand U1380 (N_1380,N_1135,N_1094);
and U1381 (N_1381,N_644,N_724);
nand U1382 (N_1382,N_917,N_834);
nor U1383 (N_1383,N_706,N_1064);
or U1384 (N_1384,N_1123,N_1067);
xor U1385 (N_1385,N_823,N_1152);
or U1386 (N_1386,N_933,N_646);
and U1387 (N_1387,N_1195,N_1197);
nor U1388 (N_1388,N_959,N_708);
and U1389 (N_1389,N_1134,N_918);
nor U1390 (N_1390,N_622,N_850);
or U1391 (N_1391,N_676,N_942);
nor U1392 (N_1392,N_1101,N_858);
and U1393 (N_1393,N_819,N_879);
and U1394 (N_1394,N_939,N_1112);
and U1395 (N_1395,N_1033,N_824);
xor U1396 (N_1396,N_639,N_1132);
nor U1397 (N_1397,N_994,N_890);
nand U1398 (N_1398,N_699,N_1154);
and U1399 (N_1399,N_1104,N_686);
or U1400 (N_1400,N_865,N_1066);
nand U1401 (N_1401,N_1181,N_1129);
nor U1402 (N_1402,N_897,N_614);
nor U1403 (N_1403,N_703,N_1027);
nor U1404 (N_1404,N_1179,N_617);
xnor U1405 (N_1405,N_1186,N_1035);
or U1406 (N_1406,N_1155,N_910);
xor U1407 (N_1407,N_601,N_1142);
or U1408 (N_1408,N_804,N_1083);
nor U1409 (N_1409,N_645,N_1001);
nor U1410 (N_1410,N_615,N_855);
nand U1411 (N_1411,N_694,N_1136);
nand U1412 (N_1412,N_743,N_1086);
xnor U1413 (N_1413,N_658,N_1038);
xor U1414 (N_1414,N_662,N_683);
nand U1415 (N_1415,N_1171,N_889);
nor U1416 (N_1416,N_802,N_1032);
or U1417 (N_1417,N_1076,N_1056);
xor U1418 (N_1418,N_767,N_835);
and U1419 (N_1419,N_1175,N_701);
and U1420 (N_1420,N_936,N_977);
and U1421 (N_1421,N_968,N_941);
or U1422 (N_1422,N_794,N_777);
nand U1423 (N_1423,N_1044,N_634);
nor U1424 (N_1424,N_664,N_960);
xnor U1425 (N_1425,N_1144,N_738);
or U1426 (N_1426,N_989,N_986);
nand U1427 (N_1427,N_655,N_864);
xor U1428 (N_1428,N_830,N_1059);
nor U1429 (N_1429,N_930,N_914);
nor U1430 (N_1430,N_899,N_1120);
xnor U1431 (N_1431,N_638,N_856);
nand U1432 (N_1432,N_707,N_1158);
nand U1433 (N_1433,N_744,N_980);
and U1434 (N_1434,N_1043,N_1071);
and U1435 (N_1435,N_940,N_681);
nand U1436 (N_1436,N_663,N_747);
nand U1437 (N_1437,N_1162,N_847);
nor U1438 (N_1438,N_1146,N_656);
nand U1439 (N_1439,N_769,N_845);
nand U1440 (N_1440,N_1113,N_633);
nor U1441 (N_1441,N_984,N_1100);
and U1442 (N_1442,N_1103,N_1183);
and U1443 (N_1443,N_861,N_1030);
or U1444 (N_1444,N_982,N_1080);
nor U1445 (N_1445,N_836,N_1091);
and U1446 (N_1446,N_630,N_946);
nor U1447 (N_1447,N_1068,N_900);
or U1448 (N_1448,N_981,N_1099);
nor U1449 (N_1449,N_792,N_1105);
and U1450 (N_1450,N_1010,N_641);
nand U1451 (N_1451,N_859,N_1004);
or U1452 (N_1452,N_1116,N_1078);
and U1453 (N_1453,N_779,N_1074);
xnor U1454 (N_1454,N_620,N_1180);
xor U1455 (N_1455,N_1003,N_971);
nand U1456 (N_1456,N_719,N_711);
and U1457 (N_1457,N_944,N_647);
xnor U1458 (N_1458,N_1140,N_782);
xnor U1459 (N_1459,N_788,N_961);
nor U1460 (N_1460,N_953,N_1191);
nand U1461 (N_1461,N_922,N_1018);
nand U1462 (N_1462,N_887,N_1127);
xnor U1463 (N_1463,N_775,N_1023);
or U1464 (N_1464,N_1107,N_809);
xnor U1465 (N_1465,N_728,N_1176);
nand U1466 (N_1466,N_1007,N_842);
and U1467 (N_1467,N_1055,N_1049);
and U1468 (N_1468,N_610,N_771);
or U1469 (N_1469,N_1182,N_1058);
nand U1470 (N_1470,N_1153,N_915);
nor U1471 (N_1471,N_773,N_891);
or U1472 (N_1472,N_772,N_1075);
and U1473 (N_1473,N_718,N_838);
and U1474 (N_1474,N_898,N_671);
xor U1475 (N_1475,N_1164,N_1089);
nand U1476 (N_1476,N_885,N_1093);
xor U1477 (N_1477,N_883,N_740);
xor U1478 (N_1478,N_717,N_739);
nor U1479 (N_1479,N_709,N_853);
nor U1480 (N_1480,N_758,N_1189);
nand U1481 (N_1481,N_690,N_943);
and U1482 (N_1482,N_774,N_908);
nor U1483 (N_1483,N_1026,N_843);
or U1484 (N_1484,N_927,N_784);
xnor U1485 (N_1485,N_957,N_1133);
and U1486 (N_1486,N_768,N_1098);
xor U1487 (N_1487,N_721,N_600);
and U1488 (N_1488,N_653,N_988);
nand U1489 (N_1489,N_925,N_807);
and U1490 (N_1490,N_1111,N_1048);
xnor U1491 (N_1491,N_821,N_892);
xor U1492 (N_1492,N_832,N_954);
nand U1493 (N_1493,N_776,N_661);
or U1494 (N_1494,N_1141,N_1114);
or U1495 (N_1495,N_1199,N_1013);
nor U1496 (N_1496,N_1118,N_1039);
nor U1497 (N_1497,N_1163,N_652);
nand U1498 (N_1498,N_884,N_1122);
and U1499 (N_1499,N_605,N_1188);
or U1500 (N_1500,N_938,N_972);
xnor U1501 (N_1501,N_790,N_776);
or U1502 (N_1502,N_1028,N_637);
and U1503 (N_1503,N_984,N_792);
and U1504 (N_1504,N_635,N_1117);
xor U1505 (N_1505,N_708,N_899);
xnor U1506 (N_1506,N_1032,N_881);
or U1507 (N_1507,N_943,N_1119);
xor U1508 (N_1508,N_684,N_783);
nand U1509 (N_1509,N_1053,N_703);
and U1510 (N_1510,N_968,N_969);
and U1511 (N_1511,N_1065,N_1089);
or U1512 (N_1512,N_860,N_937);
nand U1513 (N_1513,N_864,N_627);
xnor U1514 (N_1514,N_963,N_715);
nor U1515 (N_1515,N_997,N_1199);
nor U1516 (N_1516,N_1100,N_1063);
and U1517 (N_1517,N_616,N_1145);
and U1518 (N_1518,N_1047,N_680);
or U1519 (N_1519,N_1093,N_983);
or U1520 (N_1520,N_1078,N_817);
and U1521 (N_1521,N_752,N_1070);
nand U1522 (N_1522,N_1173,N_1055);
nand U1523 (N_1523,N_1118,N_998);
and U1524 (N_1524,N_762,N_872);
and U1525 (N_1525,N_889,N_849);
xnor U1526 (N_1526,N_805,N_819);
nand U1527 (N_1527,N_631,N_821);
or U1528 (N_1528,N_913,N_981);
and U1529 (N_1529,N_874,N_734);
and U1530 (N_1530,N_1098,N_1012);
nor U1531 (N_1531,N_1014,N_948);
xnor U1532 (N_1532,N_615,N_852);
or U1533 (N_1533,N_677,N_899);
nand U1534 (N_1534,N_869,N_1183);
nor U1535 (N_1535,N_1076,N_1156);
xnor U1536 (N_1536,N_990,N_1152);
or U1537 (N_1537,N_933,N_691);
and U1538 (N_1538,N_841,N_665);
and U1539 (N_1539,N_700,N_878);
and U1540 (N_1540,N_827,N_1089);
xnor U1541 (N_1541,N_661,N_987);
and U1542 (N_1542,N_619,N_753);
or U1543 (N_1543,N_1077,N_824);
nand U1544 (N_1544,N_855,N_999);
or U1545 (N_1545,N_1036,N_1001);
or U1546 (N_1546,N_872,N_707);
nor U1547 (N_1547,N_1093,N_812);
nor U1548 (N_1548,N_730,N_769);
nor U1549 (N_1549,N_845,N_903);
nand U1550 (N_1550,N_884,N_1076);
xnor U1551 (N_1551,N_871,N_740);
xor U1552 (N_1552,N_1039,N_618);
and U1553 (N_1553,N_836,N_601);
nor U1554 (N_1554,N_882,N_672);
xnor U1555 (N_1555,N_636,N_644);
and U1556 (N_1556,N_942,N_720);
nand U1557 (N_1557,N_1017,N_693);
and U1558 (N_1558,N_604,N_1086);
nor U1559 (N_1559,N_810,N_1123);
and U1560 (N_1560,N_794,N_1189);
nand U1561 (N_1561,N_796,N_1096);
or U1562 (N_1562,N_1113,N_963);
or U1563 (N_1563,N_719,N_1145);
or U1564 (N_1564,N_634,N_1091);
xor U1565 (N_1565,N_1099,N_1174);
and U1566 (N_1566,N_682,N_1139);
nor U1567 (N_1567,N_791,N_709);
xor U1568 (N_1568,N_1073,N_886);
nand U1569 (N_1569,N_645,N_610);
and U1570 (N_1570,N_991,N_632);
nand U1571 (N_1571,N_950,N_1028);
xnor U1572 (N_1572,N_851,N_760);
and U1573 (N_1573,N_861,N_839);
xor U1574 (N_1574,N_606,N_808);
nor U1575 (N_1575,N_1032,N_702);
xnor U1576 (N_1576,N_687,N_953);
nor U1577 (N_1577,N_627,N_602);
or U1578 (N_1578,N_764,N_966);
nand U1579 (N_1579,N_663,N_1062);
or U1580 (N_1580,N_802,N_990);
and U1581 (N_1581,N_939,N_900);
and U1582 (N_1582,N_1151,N_792);
or U1583 (N_1583,N_1158,N_1159);
or U1584 (N_1584,N_641,N_855);
nand U1585 (N_1585,N_976,N_942);
nand U1586 (N_1586,N_1076,N_655);
and U1587 (N_1587,N_867,N_803);
xnor U1588 (N_1588,N_968,N_862);
or U1589 (N_1589,N_601,N_1169);
or U1590 (N_1590,N_1097,N_833);
xnor U1591 (N_1591,N_644,N_891);
xnor U1592 (N_1592,N_815,N_981);
xor U1593 (N_1593,N_835,N_818);
nor U1594 (N_1594,N_757,N_924);
or U1595 (N_1595,N_655,N_760);
nand U1596 (N_1596,N_849,N_1189);
nor U1597 (N_1597,N_716,N_1041);
xor U1598 (N_1598,N_1058,N_607);
nand U1599 (N_1599,N_612,N_832);
or U1600 (N_1600,N_692,N_711);
or U1601 (N_1601,N_1091,N_684);
nor U1602 (N_1602,N_907,N_1059);
nor U1603 (N_1603,N_731,N_1071);
nand U1604 (N_1604,N_959,N_745);
nand U1605 (N_1605,N_1144,N_1001);
and U1606 (N_1606,N_998,N_610);
or U1607 (N_1607,N_632,N_876);
nor U1608 (N_1608,N_734,N_873);
or U1609 (N_1609,N_1000,N_1198);
nor U1610 (N_1610,N_843,N_780);
and U1611 (N_1611,N_1050,N_890);
xor U1612 (N_1612,N_1142,N_646);
nand U1613 (N_1613,N_761,N_1175);
or U1614 (N_1614,N_1066,N_647);
nand U1615 (N_1615,N_616,N_862);
or U1616 (N_1616,N_758,N_980);
nor U1617 (N_1617,N_1147,N_734);
and U1618 (N_1618,N_860,N_604);
nor U1619 (N_1619,N_1136,N_1152);
or U1620 (N_1620,N_732,N_1114);
nand U1621 (N_1621,N_932,N_985);
and U1622 (N_1622,N_688,N_652);
nor U1623 (N_1623,N_937,N_812);
nor U1624 (N_1624,N_692,N_642);
or U1625 (N_1625,N_720,N_1150);
nor U1626 (N_1626,N_1098,N_745);
or U1627 (N_1627,N_994,N_740);
and U1628 (N_1628,N_1128,N_1065);
nor U1629 (N_1629,N_915,N_730);
nand U1630 (N_1630,N_605,N_826);
xnor U1631 (N_1631,N_1069,N_785);
nand U1632 (N_1632,N_822,N_992);
and U1633 (N_1633,N_835,N_870);
nor U1634 (N_1634,N_1008,N_1012);
xor U1635 (N_1635,N_600,N_881);
and U1636 (N_1636,N_1037,N_1105);
nor U1637 (N_1637,N_842,N_902);
xor U1638 (N_1638,N_640,N_776);
and U1639 (N_1639,N_908,N_988);
and U1640 (N_1640,N_1060,N_982);
or U1641 (N_1641,N_975,N_871);
and U1642 (N_1642,N_958,N_847);
nor U1643 (N_1643,N_1178,N_779);
and U1644 (N_1644,N_654,N_1094);
nand U1645 (N_1645,N_1171,N_1175);
or U1646 (N_1646,N_795,N_934);
or U1647 (N_1647,N_1198,N_723);
xor U1648 (N_1648,N_1117,N_747);
xnor U1649 (N_1649,N_1134,N_760);
or U1650 (N_1650,N_1105,N_958);
and U1651 (N_1651,N_685,N_942);
and U1652 (N_1652,N_1053,N_1136);
nand U1653 (N_1653,N_944,N_1140);
xor U1654 (N_1654,N_1006,N_740);
or U1655 (N_1655,N_996,N_985);
or U1656 (N_1656,N_742,N_843);
or U1657 (N_1657,N_832,N_1135);
xor U1658 (N_1658,N_931,N_1116);
and U1659 (N_1659,N_786,N_860);
nand U1660 (N_1660,N_1109,N_727);
xnor U1661 (N_1661,N_852,N_885);
or U1662 (N_1662,N_628,N_1000);
nor U1663 (N_1663,N_872,N_856);
nor U1664 (N_1664,N_695,N_1187);
xnor U1665 (N_1665,N_876,N_1031);
or U1666 (N_1666,N_894,N_822);
or U1667 (N_1667,N_625,N_760);
and U1668 (N_1668,N_749,N_779);
or U1669 (N_1669,N_1179,N_804);
or U1670 (N_1670,N_1053,N_690);
nand U1671 (N_1671,N_724,N_772);
or U1672 (N_1672,N_965,N_1195);
nand U1673 (N_1673,N_1106,N_1111);
xnor U1674 (N_1674,N_950,N_997);
nor U1675 (N_1675,N_919,N_638);
xnor U1676 (N_1676,N_689,N_872);
or U1677 (N_1677,N_1075,N_892);
xor U1678 (N_1678,N_1160,N_1094);
xnor U1679 (N_1679,N_804,N_1033);
and U1680 (N_1680,N_904,N_940);
xnor U1681 (N_1681,N_779,N_1094);
xnor U1682 (N_1682,N_939,N_1126);
nand U1683 (N_1683,N_1140,N_811);
or U1684 (N_1684,N_1196,N_1192);
and U1685 (N_1685,N_890,N_1002);
nor U1686 (N_1686,N_989,N_1159);
and U1687 (N_1687,N_880,N_725);
or U1688 (N_1688,N_1075,N_1189);
xor U1689 (N_1689,N_1135,N_1040);
nor U1690 (N_1690,N_1157,N_779);
xor U1691 (N_1691,N_640,N_830);
or U1692 (N_1692,N_782,N_1042);
nand U1693 (N_1693,N_1109,N_984);
xnor U1694 (N_1694,N_1088,N_604);
and U1695 (N_1695,N_1164,N_629);
nor U1696 (N_1696,N_1178,N_620);
nor U1697 (N_1697,N_759,N_1166);
or U1698 (N_1698,N_966,N_1008);
and U1699 (N_1699,N_707,N_706);
xor U1700 (N_1700,N_944,N_1189);
and U1701 (N_1701,N_719,N_826);
or U1702 (N_1702,N_739,N_630);
xor U1703 (N_1703,N_703,N_951);
nor U1704 (N_1704,N_1094,N_841);
nor U1705 (N_1705,N_867,N_1022);
xor U1706 (N_1706,N_1152,N_1011);
and U1707 (N_1707,N_987,N_738);
nand U1708 (N_1708,N_935,N_1074);
nand U1709 (N_1709,N_1139,N_1042);
and U1710 (N_1710,N_909,N_856);
nor U1711 (N_1711,N_959,N_1137);
nor U1712 (N_1712,N_1087,N_1131);
or U1713 (N_1713,N_912,N_871);
and U1714 (N_1714,N_604,N_1064);
and U1715 (N_1715,N_874,N_876);
or U1716 (N_1716,N_723,N_690);
nor U1717 (N_1717,N_1022,N_916);
and U1718 (N_1718,N_1156,N_1104);
nor U1719 (N_1719,N_1023,N_1004);
nor U1720 (N_1720,N_1150,N_898);
xnor U1721 (N_1721,N_794,N_1049);
nand U1722 (N_1722,N_671,N_734);
nor U1723 (N_1723,N_925,N_1198);
and U1724 (N_1724,N_1014,N_1170);
and U1725 (N_1725,N_1056,N_639);
xor U1726 (N_1726,N_970,N_678);
or U1727 (N_1727,N_1158,N_665);
and U1728 (N_1728,N_739,N_1011);
and U1729 (N_1729,N_759,N_669);
xor U1730 (N_1730,N_908,N_639);
nor U1731 (N_1731,N_772,N_774);
or U1732 (N_1732,N_806,N_895);
or U1733 (N_1733,N_852,N_637);
and U1734 (N_1734,N_839,N_883);
xor U1735 (N_1735,N_1087,N_917);
nor U1736 (N_1736,N_1038,N_852);
nand U1737 (N_1737,N_669,N_760);
nand U1738 (N_1738,N_1017,N_697);
nand U1739 (N_1739,N_860,N_1144);
nor U1740 (N_1740,N_721,N_765);
and U1741 (N_1741,N_990,N_1026);
nand U1742 (N_1742,N_1087,N_1147);
nand U1743 (N_1743,N_910,N_1109);
nand U1744 (N_1744,N_755,N_981);
xor U1745 (N_1745,N_844,N_803);
nand U1746 (N_1746,N_997,N_809);
nor U1747 (N_1747,N_1029,N_925);
and U1748 (N_1748,N_705,N_600);
nand U1749 (N_1749,N_1094,N_614);
xor U1750 (N_1750,N_700,N_864);
or U1751 (N_1751,N_1103,N_813);
and U1752 (N_1752,N_857,N_958);
or U1753 (N_1753,N_1123,N_1150);
xor U1754 (N_1754,N_924,N_677);
and U1755 (N_1755,N_728,N_839);
or U1756 (N_1756,N_922,N_957);
xnor U1757 (N_1757,N_875,N_615);
nand U1758 (N_1758,N_652,N_1180);
or U1759 (N_1759,N_667,N_713);
nand U1760 (N_1760,N_850,N_895);
nand U1761 (N_1761,N_1157,N_1018);
nor U1762 (N_1762,N_996,N_1193);
xnor U1763 (N_1763,N_840,N_913);
nor U1764 (N_1764,N_669,N_1071);
or U1765 (N_1765,N_1081,N_968);
and U1766 (N_1766,N_1115,N_1195);
nor U1767 (N_1767,N_670,N_636);
or U1768 (N_1768,N_1042,N_858);
or U1769 (N_1769,N_733,N_616);
xor U1770 (N_1770,N_1050,N_903);
nor U1771 (N_1771,N_1058,N_796);
or U1772 (N_1772,N_605,N_1027);
xor U1773 (N_1773,N_756,N_964);
nor U1774 (N_1774,N_1085,N_1019);
xor U1775 (N_1775,N_1117,N_935);
nand U1776 (N_1776,N_790,N_1041);
nand U1777 (N_1777,N_1038,N_936);
or U1778 (N_1778,N_739,N_644);
nor U1779 (N_1779,N_1081,N_821);
nand U1780 (N_1780,N_719,N_1194);
or U1781 (N_1781,N_880,N_1165);
and U1782 (N_1782,N_1136,N_1032);
and U1783 (N_1783,N_778,N_776);
nor U1784 (N_1784,N_693,N_695);
nand U1785 (N_1785,N_949,N_653);
xnor U1786 (N_1786,N_950,N_1159);
or U1787 (N_1787,N_609,N_1024);
xnor U1788 (N_1788,N_632,N_921);
and U1789 (N_1789,N_763,N_675);
xnor U1790 (N_1790,N_867,N_933);
nor U1791 (N_1791,N_1029,N_647);
or U1792 (N_1792,N_1119,N_761);
and U1793 (N_1793,N_867,N_854);
and U1794 (N_1794,N_687,N_600);
nand U1795 (N_1795,N_1057,N_1152);
nor U1796 (N_1796,N_896,N_794);
nand U1797 (N_1797,N_816,N_923);
or U1798 (N_1798,N_647,N_787);
xor U1799 (N_1799,N_654,N_1070);
nor U1800 (N_1800,N_1678,N_1724);
xnor U1801 (N_1801,N_1368,N_1642);
nand U1802 (N_1802,N_1569,N_1329);
nor U1803 (N_1803,N_1531,N_1710);
xor U1804 (N_1804,N_1478,N_1345);
nor U1805 (N_1805,N_1583,N_1592);
xnor U1806 (N_1806,N_1352,N_1558);
xnor U1807 (N_1807,N_1593,N_1759);
nor U1808 (N_1808,N_1357,N_1331);
nand U1809 (N_1809,N_1509,N_1207);
and U1810 (N_1810,N_1714,N_1259);
xnor U1811 (N_1811,N_1280,N_1364);
and U1812 (N_1812,N_1681,N_1372);
xor U1813 (N_1813,N_1279,N_1338);
xnor U1814 (N_1814,N_1321,N_1263);
and U1815 (N_1815,N_1532,N_1718);
and U1816 (N_1816,N_1780,N_1340);
nand U1817 (N_1817,N_1735,N_1218);
and U1818 (N_1818,N_1635,N_1298);
nor U1819 (N_1819,N_1381,N_1536);
nand U1820 (N_1820,N_1533,N_1474);
and U1821 (N_1821,N_1223,N_1779);
xnor U1822 (N_1822,N_1578,N_1265);
xnor U1823 (N_1823,N_1762,N_1416);
and U1824 (N_1824,N_1716,N_1701);
nor U1825 (N_1825,N_1295,N_1395);
nand U1826 (N_1826,N_1247,N_1770);
nor U1827 (N_1827,N_1487,N_1203);
xor U1828 (N_1828,N_1246,N_1616);
and U1829 (N_1829,N_1502,N_1458);
and U1830 (N_1830,N_1495,N_1249);
nand U1831 (N_1831,N_1705,N_1237);
nand U1832 (N_1832,N_1434,N_1758);
and U1833 (N_1833,N_1408,N_1612);
xor U1834 (N_1834,N_1293,N_1524);
nor U1835 (N_1835,N_1589,N_1781);
nor U1836 (N_1836,N_1708,N_1512);
xnor U1837 (N_1837,N_1515,N_1663);
xor U1838 (N_1838,N_1473,N_1647);
and U1839 (N_1839,N_1268,N_1348);
or U1840 (N_1840,N_1244,N_1498);
or U1841 (N_1841,N_1307,N_1335);
and U1842 (N_1842,N_1436,N_1342);
and U1843 (N_1843,N_1383,N_1267);
xnor U1844 (N_1844,N_1205,N_1675);
and U1845 (N_1845,N_1306,N_1665);
nand U1846 (N_1846,N_1517,N_1356);
nor U1847 (N_1847,N_1631,N_1630);
nand U1848 (N_1848,N_1562,N_1564);
and U1849 (N_1849,N_1666,N_1751);
or U1850 (N_1850,N_1305,N_1686);
xnor U1851 (N_1851,N_1354,N_1580);
nor U1852 (N_1852,N_1333,N_1343);
and U1853 (N_1853,N_1645,N_1202);
or U1854 (N_1854,N_1728,N_1755);
nand U1855 (N_1855,N_1513,N_1501);
or U1856 (N_1856,N_1657,N_1411);
nand U1857 (N_1857,N_1455,N_1428);
nand U1858 (N_1858,N_1540,N_1366);
xnor U1859 (N_1859,N_1682,N_1750);
or U1860 (N_1860,N_1370,N_1749);
and U1861 (N_1861,N_1506,N_1559);
xnor U1862 (N_1862,N_1282,N_1667);
nor U1863 (N_1863,N_1433,N_1266);
nand U1864 (N_1864,N_1251,N_1481);
and U1865 (N_1865,N_1378,N_1346);
xor U1866 (N_1866,N_1409,N_1349);
nand U1867 (N_1867,N_1288,N_1521);
and U1868 (N_1868,N_1245,N_1212);
xor U1869 (N_1869,N_1337,N_1427);
or U1870 (N_1870,N_1325,N_1324);
nand U1871 (N_1871,N_1619,N_1507);
nand U1872 (N_1872,N_1339,N_1787);
nand U1873 (N_1873,N_1567,N_1789);
nand U1874 (N_1874,N_1744,N_1304);
nand U1875 (N_1875,N_1351,N_1545);
and U1876 (N_1876,N_1685,N_1404);
or U1877 (N_1877,N_1467,N_1232);
nor U1878 (N_1878,N_1308,N_1275);
nor U1879 (N_1879,N_1233,N_1585);
xor U1880 (N_1880,N_1528,N_1576);
nand U1881 (N_1881,N_1219,N_1615);
or U1882 (N_1882,N_1683,N_1661);
nor U1883 (N_1883,N_1215,N_1632);
xnor U1884 (N_1884,N_1353,N_1200);
and U1885 (N_1885,N_1626,N_1217);
xor U1886 (N_1886,N_1390,N_1622);
and U1887 (N_1887,N_1447,N_1579);
xor U1888 (N_1888,N_1389,N_1426);
nand U1889 (N_1889,N_1542,N_1256);
or U1890 (N_1890,N_1414,N_1387);
xnor U1891 (N_1891,N_1611,N_1550);
or U1892 (N_1892,N_1365,N_1660);
nor U1893 (N_1893,N_1669,N_1281);
nand U1894 (N_1894,N_1407,N_1684);
xor U1895 (N_1895,N_1462,N_1527);
nor U1896 (N_1896,N_1596,N_1651);
and U1897 (N_1897,N_1377,N_1659);
nand U1898 (N_1898,N_1386,N_1729);
or U1899 (N_1899,N_1314,N_1384);
nor U1900 (N_1900,N_1491,N_1733);
and U1901 (N_1901,N_1330,N_1757);
or U1902 (N_1902,N_1373,N_1731);
or U1903 (N_1903,N_1376,N_1312);
nor U1904 (N_1904,N_1690,N_1607);
nor U1905 (N_1905,N_1652,N_1786);
nor U1906 (N_1906,N_1285,N_1327);
xnor U1907 (N_1907,N_1572,N_1556);
nor U1908 (N_1908,N_1764,N_1273);
nand U1909 (N_1909,N_1597,N_1699);
and U1910 (N_1910,N_1523,N_1209);
or U1911 (N_1911,N_1796,N_1225);
nor U1912 (N_1912,N_1760,N_1470);
or U1913 (N_1913,N_1736,N_1719);
nand U1914 (N_1914,N_1336,N_1543);
xor U1915 (N_1915,N_1743,N_1252);
or U1916 (N_1916,N_1319,N_1401);
or U1917 (N_1917,N_1586,N_1697);
or U1918 (N_1918,N_1423,N_1793);
xor U1919 (N_1919,N_1662,N_1700);
and U1920 (N_1920,N_1614,N_1582);
nand U1921 (N_1921,N_1271,N_1405);
xor U1922 (N_1922,N_1425,N_1763);
and U1923 (N_1923,N_1773,N_1276);
xor U1924 (N_1924,N_1466,N_1417);
or U1925 (N_1925,N_1798,N_1403);
nor U1926 (N_1926,N_1790,N_1772);
or U1927 (N_1927,N_1260,N_1571);
or U1928 (N_1928,N_1380,N_1445);
xnor U1929 (N_1929,N_1234,N_1210);
or U1930 (N_1930,N_1537,N_1605);
and U1931 (N_1931,N_1739,N_1713);
xor U1932 (N_1932,N_1486,N_1526);
and U1933 (N_1933,N_1452,N_1374);
nor U1934 (N_1934,N_1519,N_1363);
xnor U1935 (N_1935,N_1516,N_1636);
xnor U1936 (N_1936,N_1476,N_1621);
or U1937 (N_1937,N_1742,N_1732);
xnor U1938 (N_1938,N_1530,N_1283);
or U1939 (N_1939,N_1520,N_1355);
or U1940 (N_1940,N_1482,N_1679);
or U1941 (N_1941,N_1573,N_1323);
and U1942 (N_1942,N_1650,N_1727);
nor U1943 (N_1943,N_1594,N_1471);
nor U1944 (N_1944,N_1264,N_1514);
and U1945 (N_1945,N_1554,N_1654);
and U1946 (N_1946,N_1220,N_1577);
nand U1947 (N_1947,N_1648,N_1320);
xnor U1948 (N_1948,N_1797,N_1463);
or U1949 (N_1949,N_1784,N_1257);
nand U1950 (N_1950,N_1644,N_1453);
and U1951 (N_1951,N_1310,N_1602);
nand U1952 (N_1952,N_1704,N_1670);
nand U1953 (N_1953,N_1769,N_1418);
xor U1954 (N_1954,N_1393,N_1588);
nor U1955 (N_1955,N_1555,N_1284);
xnor U1956 (N_1956,N_1696,N_1688);
xnor U1957 (N_1957,N_1598,N_1634);
or U1958 (N_1958,N_1334,N_1230);
and U1959 (N_1959,N_1775,N_1707);
and U1960 (N_1960,N_1278,N_1689);
xnor U1961 (N_1961,N_1741,N_1546);
xor U1962 (N_1962,N_1613,N_1258);
nor U1963 (N_1963,N_1437,N_1702);
or U1964 (N_1964,N_1449,N_1222);
and U1965 (N_1965,N_1392,N_1723);
nor U1966 (N_1966,N_1698,N_1591);
or U1967 (N_1967,N_1590,N_1618);
or U1968 (N_1968,N_1539,N_1439);
nor U1969 (N_1969,N_1385,N_1254);
nor U1970 (N_1970,N_1347,N_1311);
xnor U1971 (N_1971,N_1413,N_1441);
nor U1972 (N_1972,N_1444,N_1350);
nor U1973 (N_1973,N_1674,N_1238);
nand U1974 (N_1974,N_1479,N_1712);
nand U1975 (N_1975,N_1493,N_1745);
and U1976 (N_1976,N_1406,N_1792);
nor U1977 (N_1977,N_1541,N_1410);
nand U1978 (N_1978,N_1756,N_1313);
nor U1979 (N_1979,N_1766,N_1326);
nand U1980 (N_1980,N_1371,N_1794);
nand U1981 (N_1981,N_1655,N_1277);
or U1982 (N_1982,N_1552,N_1691);
nor U1983 (N_1983,N_1459,N_1231);
xor U1984 (N_1984,N_1344,N_1297);
nor U1985 (N_1985,N_1317,N_1362);
and U1986 (N_1986,N_1668,N_1782);
xnor U1987 (N_1987,N_1302,N_1563);
xnor U1988 (N_1988,N_1315,N_1776);
and U1989 (N_1989,N_1361,N_1269);
and U1990 (N_1990,N_1500,N_1774);
xnor U1991 (N_1991,N_1687,N_1508);
nor U1992 (N_1992,N_1565,N_1431);
xnor U1993 (N_1993,N_1715,N_1777);
and U1994 (N_1994,N_1783,N_1328);
xnor U1995 (N_1995,N_1388,N_1664);
and U1996 (N_1996,N_1641,N_1322);
nand U1997 (N_1997,N_1438,N_1620);
or U1998 (N_1998,N_1496,N_1693);
or U1999 (N_1999,N_1717,N_1640);
xnor U2000 (N_2000,N_1603,N_1609);
xnor U2001 (N_2001,N_1460,N_1560);
and U2002 (N_2002,N_1375,N_1484);
nor U2003 (N_2003,N_1242,N_1213);
nor U2004 (N_2004,N_1360,N_1468);
or U2005 (N_2005,N_1730,N_1791);
xnor U2006 (N_2006,N_1695,N_1456);
xnor U2007 (N_2007,N_1261,N_1457);
xnor U2008 (N_2008,N_1402,N_1461);
or U2009 (N_2009,N_1753,N_1296);
and U2010 (N_2010,N_1379,N_1561);
nand U2011 (N_2011,N_1294,N_1656);
nand U2012 (N_2012,N_1221,N_1442);
xor U2013 (N_2013,N_1653,N_1799);
nor U2014 (N_2014,N_1465,N_1595);
nand U2015 (N_2015,N_1671,N_1291);
or U2016 (N_2016,N_1292,N_1761);
xnor U2017 (N_2017,N_1318,N_1397);
xor U2018 (N_2018,N_1309,N_1240);
nand U2019 (N_2019,N_1446,N_1544);
xor U2020 (N_2020,N_1483,N_1503);
nor U2021 (N_2021,N_1301,N_1469);
nor U2022 (N_2022,N_1584,N_1677);
or U2023 (N_2023,N_1646,N_1680);
nor U2024 (N_2024,N_1420,N_1492);
xor U2025 (N_2025,N_1581,N_1391);
nand U2026 (N_2026,N_1464,N_1511);
xor U2027 (N_2027,N_1568,N_1747);
nand U2028 (N_2028,N_1489,N_1601);
nor U2029 (N_2029,N_1494,N_1649);
nor U2030 (N_2030,N_1250,N_1211);
xor U2031 (N_2031,N_1549,N_1748);
nand U2032 (N_2032,N_1637,N_1208);
and U2033 (N_2033,N_1725,N_1643);
and U2034 (N_2034,N_1658,N_1448);
or U2035 (N_2035,N_1672,N_1606);
nor U2036 (N_2036,N_1538,N_1262);
and U2037 (N_2037,N_1239,N_1499);
xor U2038 (N_2038,N_1272,N_1204);
nand U2039 (N_2039,N_1497,N_1341);
nor U2040 (N_2040,N_1419,N_1216);
xnor U2041 (N_2041,N_1703,N_1477);
nor U2042 (N_2042,N_1504,N_1676);
or U2043 (N_2043,N_1795,N_1765);
nand U2044 (N_2044,N_1505,N_1490);
and U2045 (N_2045,N_1303,N_1399);
nor U2046 (N_2046,N_1746,N_1547);
xor U2047 (N_2047,N_1243,N_1475);
or U2048 (N_2048,N_1299,N_1638);
xor U2049 (N_2049,N_1226,N_1720);
nand U2050 (N_2050,N_1575,N_1422);
nor U2051 (N_2051,N_1412,N_1566);
xnor U2052 (N_2052,N_1400,N_1624);
nor U2053 (N_2053,N_1394,N_1534);
and U2054 (N_2054,N_1270,N_1415);
or U2055 (N_2055,N_1206,N_1548);
xnor U2056 (N_2056,N_1551,N_1435);
nand U2057 (N_2057,N_1286,N_1229);
and U2058 (N_2058,N_1241,N_1553);
or U2059 (N_2059,N_1535,N_1608);
and U2060 (N_2060,N_1274,N_1432);
xor U2061 (N_2061,N_1557,N_1737);
nor U2062 (N_2062,N_1574,N_1740);
nor U2063 (N_2063,N_1767,N_1778);
or U2064 (N_2064,N_1480,N_1639);
nand U2065 (N_2065,N_1625,N_1692);
and U2066 (N_2066,N_1424,N_1711);
or U2067 (N_2067,N_1398,N_1332);
nor U2068 (N_2068,N_1617,N_1529);
nor U2069 (N_2069,N_1785,N_1610);
or U2070 (N_2070,N_1600,N_1673);
or U2071 (N_2071,N_1771,N_1706);
or U2072 (N_2072,N_1367,N_1253);
nand U2073 (N_2073,N_1485,N_1599);
or U2074 (N_2074,N_1768,N_1227);
nor U2075 (N_2075,N_1726,N_1451);
or U2076 (N_2076,N_1722,N_1358);
or U2077 (N_2077,N_1228,N_1510);
xnor U2078 (N_2078,N_1248,N_1396);
and U2079 (N_2079,N_1623,N_1628);
and U2080 (N_2080,N_1709,N_1359);
or U2081 (N_2081,N_1214,N_1235);
nand U2082 (N_2082,N_1738,N_1450);
nor U2083 (N_2083,N_1201,N_1627);
xor U2084 (N_2084,N_1604,N_1316);
xor U2085 (N_2085,N_1488,N_1570);
nand U2086 (N_2086,N_1525,N_1224);
or U2087 (N_2087,N_1522,N_1289);
and U2088 (N_2088,N_1788,N_1382);
nand U2089 (N_2089,N_1287,N_1290);
nor U2090 (N_2090,N_1629,N_1754);
nand U2091 (N_2091,N_1429,N_1472);
nor U2092 (N_2092,N_1633,N_1430);
nand U2093 (N_2093,N_1454,N_1421);
or U2094 (N_2094,N_1369,N_1752);
or U2095 (N_2095,N_1694,N_1734);
and U2096 (N_2096,N_1300,N_1721);
and U2097 (N_2097,N_1255,N_1443);
nor U2098 (N_2098,N_1587,N_1236);
or U2099 (N_2099,N_1440,N_1518);
nand U2100 (N_2100,N_1614,N_1260);
and U2101 (N_2101,N_1799,N_1636);
or U2102 (N_2102,N_1215,N_1523);
and U2103 (N_2103,N_1495,N_1550);
xor U2104 (N_2104,N_1600,N_1308);
nand U2105 (N_2105,N_1790,N_1498);
nor U2106 (N_2106,N_1628,N_1640);
or U2107 (N_2107,N_1334,N_1760);
nor U2108 (N_2108,N_1657,N_1740);
nand U2109 (N_2109,N_1386,N_1630);
nor U2110 (N_2110,N_1780,N_1426);
and U2111 (N_2111,N_1740,N_1230);
or U2112 (N_2112,N_1467,N_1769);
and U2113 (N_2113,N_1689,N_1407);
nand U2114 (N_2114,N_1268,N_1673);
xor U2115 (N_2115,N_1564,N_1753);
and U2116 (N_2116,N_1673,N_1625);
or U2117 (N_2117,N_1643,N_1469);
nand U2118 (N_2118,N_1254,N_1455);
nor U2119 (N_2119,N_1490,N_1704);
or U2120 (N_2120,N_1432,N_1414);
nor U2121 (N_2121,N_1495,N_1316);
nor U2122 (N_2122,N_1337,N_1767);
nand U2123 (N_2123,N_1526,N_1243);
xnor U2124 (N_2124,N_1329,N_1797);
and U2125 (N_2125,N_1662,N_1568);
nor U2126 (N_2126,N_1330,N_1503);
nor U2127 (N_2127,N_1578,N_1499);
nand U2128 (N_2128,N_1236,N_1362);
xnor U2129 (N_2129,N_1549,N_1229);
nor U2130 (N_2130,N_1749,N_1750);
nor U2131 (N_2131,N_1495,N_1768);
nand U2132 (N_2132,N_1589,N_1479);
nand U2133 (N_2133,N_1709,N_1365);
xnor U2134 (N_2134,N_1412,N_1387);
or U2135 (N_2135,N_1348,N_1415);
nand U2136 (N_2136,N_1472,N_1702);
or U2137 (N_2137,N_1340,N_1481);
or U2138 (N_2138,N_1385,N_1541);
and U2139 (N_2139,N_1794,N_1679);
xor U2140 (N_2140,N_1589,N_1749);
and U2141 (N_2141,N_1765,N_1658);
and U2142 (N_2142,N_1747,N_1461);
nor U2143 (N_2143,N_1568,N_1401);
xor U2144 (N_2144,N_1511,N_1288);
nand U2145 (N_2145,N_1238,N_1551);
and U2146 (N_2146,N_1404,N_1576);
nand U2147 (N_2147,N_1727,N_1235);
nand U2148 (N_2148,N_1695,N_1462);
and U2149 (N_2149,N_1712,N_1271);
or U2150 (N_2150,N_1515,N_1332);
nor U2151 (N_2151,N_1572,N_1410);
nor U2152 (N_2152,N_1459,N_1740);
xor U2153 (N_2153,N_1579,N_1548);
nor U2154 (N_2154,N_1785,N_1241);
and U2155 (N_2155,N_1227,N_1601);
nor U2156 (N_2156,N_1534,N_1366);
nor U2157 (N_2157,N_1291,N_1512);
and U2158 (N_2158,N_1692,N_1216);
or U2159 (N_2159,N_1257,N_1394);
and U2160 (N_2160,N_1418,N_1797);
and U2161 (N_2161,N_1737,N_1380);
nor U2162 (N_2162,N_1248,N_1240);
nand U2163 (N_2163,N_1241,N_1359);
xor U2164 (N_2164,N_1767,N_1672);
or U2165 (N_2165,N_1688,N_1360);
xnor U2166 (N_2166,N_1522,N_1797);
and U2167 (N_2167,N_1248,N_1381);
or U2168 (N_2168,N_1642,N_1573);
and U2169 (N_2169,N_1787,N_1597);
and U2170 (N_2170,N_1788,N_1689);
xor U2171 (N_2171,N_1346,N_1714);
nor U2172 (N_2172,N_1597,N_1773);
and U2173 (N_2173,N_1745,N_1534);
nor U2174 (N_2174,N_1672,N_1299);
or U2175 (N_2175,N_1648,N_1300);
xor U2176 (N_2176,N_1209,N_1743);
and U2177 (N_2177,N_1244,N_1249);
nand U2178 (N_2178,N_1245,N_1559);
nand U2179 (N_2179,N_1506,N_1741);
xor U2180 (N_2180,N_1264,N_1780);
xnor U2181 (N_2181,N_1514,N_1561);
nor U2182 (N_2182,N_1752,N_1566);
xnor U2183 (N_2183,N_1297,N_1754);
xor U2184 (N_2184,N_1747,N_1663);
or U2185 (N_2185,N_1679,N_1556);
or U2186 (N_2186,N_1563,N_1715);
and U2187 (N_2187,N_1227,N_1210);
nand U2188 (N_2188,N_1408,N_1592);
and U2189 (N_2189,N_1598,N_1772);
nand U2190 (N_2190,N_1212,N_1464);
and U2191 (N_2191,N_1258,N_1750);
and U2192 (N_2192,N_1338,N_1251);
or U2193 (N_2193,N_1659,N_1796);
nand U2194 (N_2194,N_1315,N_1565);
or U2195 (N_2195,N_1486,N_1266);
nand U2196 (N_2196,N_1575,N_1636);
nor U2197 (N_2197,N_1363,N_1305);
or U2198 (N_2198,N_1757,N_1779);
or U2199 (N_2199,N_1460,N_1753);
and U2200 (N_2200,N_1372,N_1649);
or U2201 (N_2201,N_1548,N_1200);
or U2202 (N_2202,N_1294,N_1339);
and U2203 (N_2203,N_1682,N_1684);
nand U2204 (N_2204,N_1633,N_1795);
nor U2205 (N_2205,N_1795,N_1460);
xnor U2206 (N_2206,N_1713,N_1711);
and U2207 (N_2207,N_1460,N_1515);
nor U2208 (N_2208,N_1514,N_1695);
nor U2209 (N_2209,N_1211,N_1336);
or U2210 (N_2210,N_1492,N_1436);
xor U2211 (N_2211,N_1496,N_1609);
and U2212 (N_2212,N_1413,N_1705);
or U2213 (N_2213,N_1483,N_1487);
xnor U2214 (N_2214,N_1329,N_1619);
nor U2215 (N_2215,N_1553,N_1504);
nor U2216 (N_2216,N_1751,N_1425);
or U2217 (N_2217,N_1522,N_1496);
or U2218 (N_2218,N_1234,N_1268);
nand U2219 (N_2219,N_1357,N_1229);
or U2220 (N_2220,N_1709,N_1786);
nor U2221 (N_2221,N_1599,N_1790);
nor U2222 (N_2222,N_1772,N_1721);
or U2223 (N_2223,N_1373,N_1521);
or U2224 (N_2224,N_1628,N_1519);
nor U2225 (N_2225,N_1456,N_1659);
and U2226 (N_2226,N_1739,N_1768);
xor U2227 (N_2227,N_1334,N_1555);
xnor U2228 (N_2228,N_1615,N_1353);
and U2229 (N_2229,N_1258,N_1703);
xnor U2230 (N_2230,N_1609,N_1656);
xor U2231 (N_2231,N_1683,N_1676);
nand U2232 (N_2232,N_1377,N_1635);
nor U2233 (N_2233,N_1525,N_1240);
xnor U2234 (N_2234,N_1226,N_1271);
nor U2235 (N_2235,N_1495,N_1514);
xor U2236 (N_2236,N_1261,N_1688);
nor U2237 (N_2237,N_1556,N_1445);
nand U2238 (N_2238,N_1334,N_1614);
or U2239 (N_2239,N_1536,N_1732);
nand U2240 (N_2240,N_1268,N_1434);
xnor U2241 (N_2241,N_1263,N_1547);
and U2242 (N_2242,N_1467,N_1341);
or U2243 (N_2243,N_1241,N_1366);
nor U2244 (N_2244,N_1206,N_1525);
xnor U2245 (N_2245,N_1404,N_1659);
xnor U2246 (N_2246,N_1233,N_1692);
and U2247 (N_2247,N_1679,N_1786);
nor U2248 (N_2248,N_1551,N_1316);
and U2249 (N_2249,N_1248,N_1390);
or U2250 (N_2250,N_1271,N_1475);
nor U2251 (N_2251,N_1509,N_1465);
nor U2252 (N_2252,N_1520,N_1770);
and U2253 (N_2253,N_1200,N_1313);
and U2254 (N_2254,N_1388,N_1589);
xnor U2255 (N_2255,N_1708,N_1455);
xor U2256 (N_2256,N_1269,N_1587);
nor U2257 (N_2257,N_1449,N_1746);
nor U2258 (N_2258,N_1492,N_1269);
nor U2259 (N_2259,N_1623,N_1385);
xnor U2260 (N_2260,N_1720,N_1668);
nand U2261 (N_2261,N_1494,N_1531);
nand U2262 (N_2262,N_1590,N_1558);
nand U2263 (N_2263,N_1230,N_1207);
and U2264 (N_2264,N_1671,N_1276);
nand U2265 (N_2265,N_1551,N_1670);
nand U2266 (N_2266,N_1452,N_1233);
nand U2267 (N_2267,N_1269,N_1212);
nor U2268 (N_2268,N_1596,N_1550);
or U2269 (N_2269,N_1650,N_1718);
or U2270 (N_2270,N_1666,N_1694);
xor U2271 (N_2271,N_1377,N_1778);
or U2272 (N_2272,N_1258,N_1213);
and U2273 (N_2273,N_1275,N_1566);
nor U2274 (N_2274,N_1399,N_1771);
nor U2275 (N_2275,N_1202,N_1725);
nand U2276 (N_2276,N_1666,N_1577);
nand U2277 (N_2277,N_1793,N_1638);
nand U2278 (N_2278,N_1246,N_1772);
xnor U2279 (N_2279,N_1311,N_1475);
or U2280 (N_2280,N_1706,N_1752);
nor U2281 (N_2281,N_1567,N_1606);
nor U2282 (N_2282,N_1387,N_1224);
nand U2283 (N_2283,N_1237,N_1551);
xor U2284 (N_2284,N_1472,N_1519);
nor U2285 (N_2285,N_1278,N_1380);
xor U2286 (N_2286,N_1469,N_1603);
and U2287 (N_2287,N_1577,N_1610);
nor U2288 (N_2288,N_1227,N_1794);
nor U2289 (N_2289,N_1765,N_1215);
and U2290 (N_2290,N_1269,N_1677);
nor U2291 (N_2291,N_1523,N_1394);
xor U2292 (N_2292,N_1423,N_1743);
nand U2293 (N_2293,N_1675,N_1417);
and U2294 (N_2294,N_1676,N_1266);
xor U2295 (N_2295,N_1518,N_1247);
xnor U2296 (N_2296,N_1548,N_1518);
nor U2297 (N_2297,N_1473,N_1656);
xor U2298 (N_2298,N_1523,N_1535);
or U2299 (N_2299,N_1473,N_1243);
xnor U2300 (N_2300,N_1427,N_1598);
xnor U2301 (N_2301,N_1629,N_1494);
xor U2302 (N_2302,N_1286,N_1493);
nand U2303 (N_2303,N_1218,N_1606);
or U2304 (N_2304,N_1508,N_1710);
or U2305 (N_2305,N_1448,N_1370);
and U2306 (N_2306,N_1234,N_1237);
nor U2307 (N_2307,N_1382,N_1325);
nand U2308 (N_2308,N_1322,N_1476);
xnor U2309 (N_2309,N_1317,N_1216);
nor U2310 (N_2310,N_1656,N_1747);
nand U2311 (N_2311,N_1774,N_1400);
xor U2312 (N_2312,N_1283,N_1613);
and U2313 (N_2313,N_1293,N_1549);
nor U2314 (N_2314,N_1586,N_1733);
and U2315 (N_2315,N_1640,N_1544);
or U2316 (N_2316,N_1686,N_1438);
nand U2317 (N_2317,N_1680,N_1409);
nand U2318 (N_2318,N_1300,N_1316);
and U2319 (N_2319,N_1592,N_1780);
and U2320 (N_2320,N_1364,N_1519);
and U2321 (N_2321,N_1306,N_1553);
xor U2322 (N_2322,N_1719,N_1624);
xor U2323 (N_2323,N_1543,N_1350);
nor U2324 (N_2324,N_1764,N_1531);
or U2325 (N_2325,N_1230,N_1404);
or U2326 (N_2326,N_1455,N_1290);
nor U2327 (N_2327,N_1466,N_1418);
nand U2328 (N_2328,N_1782,N_1578);
and U2329 (N_2329,N_1347,N_1721);
xnor U2330 (N_2330,N_1439,N_1797);
nand U2331 (N_2331,N_1701,N_1734);
xnor U2332 (N_2332,N_1700,N_1435);
nand U2333 (N_2333,N_1422,N_1782);
and U2334 (N_2334,N_1639,N_1503);
or U2335 (N_2335,N_1654,N_1384);
or U2336 (N_2336,N_1620,N_1719);
or U2337 (N_2337,N_1595,N_1546);
and U2338 (N_2338,N_1718,N_1592);
or U2339 (N_2339,N_1280,N_1325);
and U2340 (N_2340,N_1509,N_1776);
nor U2341 (N_2341,N_1606,N_1474);
nor U2342 (N_2342,N_1299,N_1523);
nand U2343 (N_2343,N_1628,N_1260);
and U2344 (N_2344,N_1209,N_1734);
nand U2345 (N_2345,N_1793,N_1424);
or U2346 (N_2346,N_1685,N_1607);
or U2347 (N_2347,N_1535,N_1452);
or U2348 (N_2348,N_1422,N_1463);
nand U2349 (N_2349,N_1439,N_1720);
or U2350 (N_2350,N_1252,N_1662);
nor U2351 (N_2351,N_1607,N_1494);
nand U2352 (N_2352,N_1310,N_1468);
nor U2353 (N_2353,N_1389,N_1371);
nand U2354 (N_2354,N_1674,N_1611);
nor U2355 (N_2355,N_1561,N_1554);
and U2356 (N_2356,N_1235,N_1510);
nand U2357 (N_2357,N_1799,N_1500);
nand U2358 (N_2358,N_1531,N_1321);
or U2359 (N_2359,N_1477,N_1210);
or U2360 (N_2360,N_1230,N_1675);
xor U2361 (N_2361,N_1236,N_1303);
or U2362 (N_2362,N_1315,N_1353);
nand U2363 (N_2363,N_1250,N_1334);
and U2364 (N_2364,N_1405,N_1706);
xor U2365 (N_2365,N_1583,N_1763);
or U2366 (N_2366,N_1794,N_1653);
nor U2367 (N_2367,N_1461,N_1559);
nand U2368 (N_2368,N_1511,N_1325);
xor U2369 (N_2369,N_1481,N_1657);
nand U2370 (N_2370,N_1459,N_1585);
nor U2371 (N_2371,N_1334,N_1653);
nand U2372 (N_2372,N_1727,N_1344);
nor U2373 (N_2373,N_1222,N_1553);
and U2374 (N_2374,N_1379,N_1611);
and U2375 (N_2375,N_1487,N_1221);
nand U2376 (N_2376,N_1784,N_1506);
xnor U2377 (N_2377,N_1431,N_1542);
nand U2378 (N_2378,N_1571,N_1749);
nor U2379 (N_2379,N_1538,N_1599);
nand U2380 (N_2380,N_1673,N_1709);
or U2381 (N_2381,N_1554,N_1693);
nand U2382 (N_2382,N_1275,N_1449);
nand U2383 (N_2383,N_1253,N_1498);
and U2384 (N_2384,N_1620,N_1549);
or U2385 (N_2385,N_1559,N_1253);
and U2386 (N_2386,N_1651,N_1390);
nor U2387 (N_2387,N_1790,N_1719);
nand U2388 (N_2388,N_1360,N_1479);
or U2389 (N_2389,N_1651,N_1732);
nand U2390 (N_2390,N_1687,N_1499);
xor U2391 (N_2391,N_1453,N_1324);
nand U2392 (N_2392,N_1659,N_1409);
xnor U2393 (N_2393,N_1254,N_1552);
xor U2394 (N_2394,N_1498,N_1415);
or U2395 (N_2395,N_1732,N_1274);
and U2396 (N_2396,N_1529,N_1320);
and U2397 (N_2397,N_1772,N_1628);
nor U2398 (N_2398,N_1603,N_1624);
nor U2399 (N_2399,N_1773,N_1769);
and U2400 (N_2400,N_2114,N_2205);
nand U2401 (N_2401,N_1829,N_1883);
or U2402 (N_2402,N_1890,N_2283);
xnor U2403 (N_2403,N_1935,N_2008);
or U2404 (N_2404,N_1851,N_1916);
and U2405 (N_2405,N_2204,N_1995);
xor U2406 (N_2406,N_2234,N_2392);
nand U2407 (N_2407,N_2179,N_2316);
nand U2408 (N_2408,N_2369,N_1957);
or U2409 (N_2409,N_2365,N_2351);
nor U2410 (N_2410,N_1948,N_1819);
and U2411 (N_2411,N_2166,N_2130);
nor U2412 (N_2412,N_2184,N_1894);
nor U2413 (N_2413,N_2198,N_1955);
and U2414 (N_2414,N_2226,N_2339);
or U2415 (N_2415,N_2359,N_2071);
xor U2416 (N_2416,N_2138,N_2066);
nor U2417 (N_2417,N_2153,N_1941);
xor U2418 (N_2418,N_1860,N_1994);
or U2419 (N_2419,N_1858,N_1892);
nor U2420 (N_2420,N_1977,N_2218);
and U2421 (N_2421,N_1901,N_2037);
nor U2422 (N_2422,N_1964,N_2187);
or U2423 (N_2423,N_2010,N_2251);
xnor U2424 (N_2424,N_2046,N_2113);
and U2425 (N_2425,N_2096,N_1850);
or U2426 (N_2426,N_2201,N_1874);
xor U2427 (N_2427,N_1867,N_1853);
nand U2428 (N_2428,N_2284,N_2348);
xnor U2429 (N_2429,N_2196,N_2274);
nand U2430 (N_2430,N_1872,N_1818);
nand U2431 (N_2431,N_1975,N_2346);
xor U2432 (N_2432,N_1893,N_2292);
or U2433 (N_2433,N_2299,N_2028);
or U2434 (N_2434,N_2014,N_2297);
nor U2435 (N_2435,N_2344,N_1820);
and U2436 (N_2436,N_1800,N_2220);
and U2437 (N_2437,N_1871,N_2132);
and U2438 (N_2438,N_2151,N_2026);
and U2439 (N_2439,N_2105,N_1811);
or U2440 (N_2440,N_2330,N_2280);
nand U2441 (N_2441,N_2327,N_2051);
and U2442 (N_2442,N_1914,N_2202);
xnor U2443 (N_2443,N_2325,N_2161);
or U2444 (N_2444,N_1880,N_1943);
or U2445 (N_2445,N_2362,N_1884);
or U2446 (N_2446,N_1988,N_2143);
or U2447 (N_2447,N_2265,N_2216);
nand U2448 (N_2448,N_1990,N_2210);
xnor U2449 (N_2449,N_1832,N_2070);
nor U2450 (N_2450,N_1925,N_2188);
and U2451 (N_2451,N_1920,N_2065);
xor U2452 (N_2452,N_1963,N_2322);
nor U2453 (N_2453,N_2200,N_2199);
and U2454 (N_2454,N_1993,N_2318);
nor U2455 (N_2455,N_2170,N_2399);
xor U2456 (N_2456,N_2156,N_1813);
xnor U2457 (N_2457,N_1970,N_1812);
or U2458 (N_2458,N_1959,N_2129);
nor U2459 (N_2459,N_2023,N_2389);
nor U2460 (N_2460,N_2367,N_2063);
xor U2461 (N_2461,N_1909,N_2334);
nor U2462 (N_2462,N_2194,N_1998);
nor U2463 (N_2463,N_2239,N_1848);
and U2464 (N_2464,N_2385,N_2183);
nor U2465 (N_2465,N_2233,N_1846);
and U2466 (N_2466,N_1942,N_2064);
xnor U2467 (N_2467,N_1862,N_2128);
xor U2468 (N_2468,N_1999,N_2139);
nand U2469 (N_2469,N_2288,N_1900);
or U2470 (N_2470,N_2090,N_2147);
and U2471 (N_2471,N_2285,N_1849);
and U2472 (N_2472,N_1953,N_2341);
and U2473 (N_2473,N_2397,N_1857);
nand U2474 (N_2474,N_1961,N_1912);
nor U2475 (N_2475,N_2276,N_2058);
nor U2476 (N_2476,N_1917,N_2068);
or U2477 (N_2477,N_2387,N_2350);
nand U2478 (N_2478,N_1947,N_1974);
xnor U2479 (N_2479,N_2300,N_2035);
nand U2480 (N_2480,N_1972,N_2012);
nand U2481 (N_2481,N_1810,N_1958);
or U2482 (N_2482,N_2015,N_2106);
nand U2483 (N_2483,N_1952,N_2287);
or U2484 (N_2484,N_2141,N_1861);
nand U2485 (N_2485,N_1944,N_1840);
or U2486 (N_2486,N_2353,N_1907);
nand U2487 (N_2487,N_2236,N_1989);
nor U2488 (N_2488,N_1919,N_2003);
nand U2489 (N_2489,N_2272,N_1991);
or U2490 (N_2490,N_2006,N_2031);
and U2491 (N_2491,N_2270,N_1875);
or U2492 (N_2492,N_2343,N_2078);
or U2493 (N_2493,N_1842,N_1814);
nand U2494 (N_2494,N_1928,N_2331);
nor U2495 (N_2495,N_2213,N_1804);
nor U2496 (N_2496,N_2264,N_1802);
and U2497 (N_2497,N_2395,N_2286);
xnor U2498 (N_2498,N_2328,N_1946);
nor U2499 (N_2499,N_2137,N_2177);
nand U2500 (N_2500,N_1815,N_2145);
or U2501 (N_2501,N_2085,N_1915);
and U2502 (N_2502,N_2025,N_2326);
or U2503 (N_2503,N_2221,N_2335);
nand U2504 (N_2504,N_2057,N_1807);
and U2505 (N_2505,N_2380,N_2033);
xor U2506 (N_2506,N_1831,N_2004);
or U2507 (N_2507,N_2281,N_2157);
and U2508 (N_2508,N_2340,N_2257);
nor U2509 (N_2509,N_2089,N_2371);
xor U2510 (N_2510,N_2102,N_1803);
and U2511 (N_2511,N_2142,N_2056);
nand U2512 (N_2512,N_1929,N_2342);
nor U2513 (N_2513,N_2376,N_2247);
or U2514 (N_2514,N_2171,N_2036);
or U2515 (N_2515,N_2323,N_1835);
and U2516 (N_2516,N_1801,N_2394);
and U2517 (N_2517,N_2396,N_1971);
nand U2518 (N_2518,N_1859,N_2225);
nand U2519 (N_2519,N_1841,N_2393);
or U2520 (N_2520,N_1967,N_2192);
nor U2521 (N_2521,N_2048,N_2030);
xor U2522 (N_2522,N_1969,N_2088);
or U2523 (N_2523,N_2047,N_1904);
nor U2524 (N_2524,N_1825,N_1992);
or U2525 (N_2525,N_2214,N_2172);
xor U2526 (N_2526,N_2178,N_1954);
or U2527 (N_2527,N_2013,N_2290);
xnor U2528 (N_2528,N_2313,N_2258);
and U2529 (N_2529,N_2277,N_2358);
and U2530 (N_2530,N_1997,N_2146);
and U2531 (N_2531,N_1878,N_2310);
or U2532 (N_2532,N_2373,N_1809);
xnor U2533 (N_2533,N_1996,N_2241);
and U2534 (N_2534,N_2246,N_2303);
and U2535 (N_2535,N_1923,N_1838);
nor U2536 (N_2536,N_1927,N_2163);
xor U2537 (N_2537,N_1933,N_2232);
nor U2538 (N_2538,N_2268,N_2377);
xnor U2539 (N_2539,N_2317,N_2080);
or U2540 (N_2540,N_2061,N_2195);
nand U2541 (N_2541,N_2098,N_2049);
xor U2542 (N_2542,N_2298,N_1905);
and U2543 (N_2543,N_2381,N_1956);
or U2544 (N_2544,N_1965,N_2185);
or U2545 (N_2545,N_2231,N_2109);
or U2546 (N_2546,N_2165,N_2275);
xor U2547 (N_2547,N_2055,N_2269);
xnor U2548 (N_2548,N_2228,N_2144);
and U2549 (N_2549,N_2116,N_1827);
nor U2550 (N_2550,N_1937,N_2079);
or U2551 (N_2551,N_2017,N_2301);
xnor U2552 (N_2552,N_2248,N_2242);
nor U2553 (N_2553,N_2197,N_2100);
nand U2554 (N_2554,N_1940,N_2117);
nor U2555 (N_2555,N_1833,N_2095);
or U2556 (N_2556,N_2315,N_1903);
xnor U2557 (N_2557,N_2243,N_1865);
or U2558 (N_2558,N_2319,N_2094);
nor U2559 (N_2559,N_2181,N_2000);
nor U2560 (N_2560,N_2398,N_2122);
xnor U2561 (N_2561,N_1830,N_2019);
and U2562 (N_2562,N_2186,N_2108);
or U2563 (N_2563,N_2075,N_2304);
nand U2564 (N_2564,N_1966,N_2308);
nor U2565 (N_2565,N_2238,N_2230);
nor U2566 (N_2566,N_2160,N_1910);
and U2567 (N_2567,N_1864,N_2133);
or U2568 (N_2568,N_1985,N_2249);
xnor U2569 (N_2569,N_2045,N_2329);
and U2570 (N_2570,N_1962,N_2262);
xnor U2571 (N_2571,N_1844,N_1918);
nor U2572 (N_2572,N_2180,N_2305);
nand U2573 (N_2573,N_1945,N_2021);
nand U2574 (N_2574,N_2345,N_2361);
xnor U2575 (N_2575,N_1895,N_2193);
nor U2576 (N_2576,N_2386,N_1922);
and U2577 (N_2577,N_1806,N_1866);
and U2578 (N_2578,N_2282,N_2278);
or U2579 (N_2579,N_2034,N_2307);
xnor U2580 (N_2580,N_1837,N_1817);
xnor U2581 (N_2581,N_2223,N_2357);
or U2582 (N_2582,N_2084,N_1879);
xor U2583 (N_2583,N_2158,N_2054);
and U2584 (N_2584,N_2254,N_2067);
and U2585 (N_2585,N_1856,N_2235);
and U2586 (N_2586,N_2311,N_2149);
or U2587 (N_2587,N_2115,N_2148);
xnor U2588 (N_2588,N_1854,N_1979);
nor U2589 (N_2589,N_1987,N_2125);
nor U2590 (N_2590,N_1887,N_2208);
nor U2591 (N_2591,N_2383,N_2333);
or U2592 (N_2592,N_2041,N_2364);
xnor U2593 (N_2593,N_2119,N_1881);
or U2594 (N_2594,N_2124,N_1869);
and U2595 (N_2595,N_1852,N_1845);
or U2596 (N_2596,N_2349,N_2120);
xnor U2597 (N_2597,N_2127,N_2244);
nand U2598 (N_2598,N_2289,N_1821);
xnor U2599 (N_2599,N_2022,N_2378);
or U2600 (N_2600,N_2002,N_2296);
xnor U2601 (N_2601,N_2168,N_2255);
nand U2602 (N_2602,N_2382,N_2118);
xnor U2603 (N_2603,N_1843,N_2103);
xor U2604 (N_2604,N_2217,N_2306);
and U2605 (N_2605,N_2169,N_2206);
xor U2606 (N_2606,N_1897,N_1888);
nand U2607 (N_2607,N_2082,N_2294);
and U2608 (N_2608,N_2073,N_2167);
xor U2609 (N_2609,N_1896,N_2352);
xnor U2610 (N_2610,N_1938,N_2229);
nor U2611 (N_2611,N_1873,N_2101);
nor U2612 (N_2612,N_2263,N_2111);
and U2613 (N_2613,N_1886,N_1902);
nand U2614 (N_2614,N_2044,N_1911);
nand U2615 (N_2615,N_2293,N_2043);
xor U2616 (N_2616,N_2279,N_2107);
or U2617 (N_2617,N_2093,N_2099);
xor U2618 (N_2618,N_2302,N_1839);
xnor U2619 (N_2619,N_2052,N_2375);
and U2620 (N_2620,N_2029,N_2011);
and U2621 (N_2621,N_1876,N_2134);
nor U2622 (N_2622,N_2074,N_2391);
or U2623 (N_2623,N_2032,N_2211);
nand U2624 (N_2624,N_1870,N_2092);
nor U2625 (N_2625,N_2266,N_2072);
xor U2626 (N_2626,N_2087,N_2131);
nand U2627 (N_2627,N_2240,N_2291);
nor U2628 (N_2628,N_2347,N_2175);
and U2629 (N_2629,N_2091,N_1921);
or U2630 (N_2630,N_2374,N_2354);
xor U2631 (N_2631,N_2182,N_2212);
nand U2632 (N_2632,N_2069,N_2273);
nor U2633 (N_2633,N_1868,N_2271);
nor U2634 (N_2634,N_1924,N_1816);
and U2635 (N_2635,N_1949,N_2162);
or U2636 (N_2636,N_2059,N_2038);
nand U2637 (N_2637,N_2321,N_1824);
xor U2638 (N_2638,N_1968,N_2159);
or U2639 (N_2639,N_2336,N_1877);
nor U2640 (N_2640,N_2366,N_2007);
nand U2641 (N_2641,N_1882,N_2126);
and U2642 (N_2642,N_2173,N_2190);
or U2643 (N_2643,N_2388,N_2356);
and U2644 (N_2644,N_1855,N_2152);
xnor U2645 (N_2645,N_2155,N_2267);
or U2646 (N_2646,N_1808,N_1932);
nand U2647 (N_2647,N_1934,N_2136);
or U2648 (N_2648,N_2123,N_2215);
nand U2649 (N_2649,N_2135,N_2027);
xor U2650 (N_2650,N_2001,N_2042);
and U2651 (N_2651,N_2081,N_2189);
nand U2652 (N_2652,N_2252,N_2250);
and U2653 (N_2653,N_2140,N_2039);
nor U2654 (N_2654,N_2363,N_1828);
nor U2655 (N_2655,N_2370,N_2053);
or U2656 (N_2656,N_1978,N_1847);
nand U2657 (N_2657,N_1986,N_2261);
nand U2658 (N_2658,N_2309,N_2076);
and U2659 (N_2659,N_1930,N_2368);
nor U2660 (N_2660,N_1976,N_1891);
nor U2661 (N_2661,N_2384,N_2050);
nor U2662 (N_2662,N_2355,N_1951);
xor U2663 (N_2663,N_2314,N_1899);
xnor U2664 (N_2664,N_1980,N_2176);
and U2665 (N_2665,N_1984,N_2222);
nand U2666 (N_2666,N_1950,N_1908);
nand U2667 (N_2667,N_2372,N_2040);
nor U2668 (N_2668,N_2083,N_1931);
xor U2669 (N_2669,N_1936,N_1885);
or U2670 (N_2670,N_2338,N_2203);
nand U2671 (N_2671,N_2062,N_2256);
and U2672 (N_2672,N_1939,N_1889);
nand U2673 (N_2673,N_2312,N_2150);
nor U2674 (N_2674,N_1863,N_2324);
or U2675 (N_2675,N_2104,N_2295);
nor U2676 (N_2676,N_2320,N_2360);
or U2677 (N_2677,N_2110,N_2260);
nand U2678 (N_2678,N_2020,N_2086);
and U2679 (N_2679,N_2154,N_1805);
xnor U2680 (N_2680,N_1982,N_1926);
nor U2681 (N_2681,N_2253,N_2077);
and U2682 (N_2682,N_2112,N_2207);
and U2683 (N_2683,N_1983,N_2191);
nand U2684 (N_2684,N_2237,N_1823);
and U2685 (N_2685,N_2245,N_2024);
nand U2686 (N_2686,N_1973,N_2121);
nand U2687 (N_2687,N_1960,N_2097);
xor U2688 (N_2688,N_2259,N_2005);
nor U2689 (N_2689,N_2174,N_1913);
nand U2690 (N_2690,N_2219,N_1981);
or U2691 (N_2691,N_2224,N_2337);
nor U2692 (N_2692,N_2227,N_2060);
nand U2693 (N_2693,N_2332,N_2009);
and U2694 (N_2694,N_2016,N_2164);
nor U2695 (N_2695,N_1822,N_2018);
nand U2696 (N_2696,N_2390,N_1836);
and U2697 (N_2697,N_1906,N_1898);
nand U2698 (N_2698,N_1826,N_2379);
xnor U2699 (N_2699,N_2209,N_1834);
xor U2700 (N_2700,N_2174,N_2273);
and U2701 (N_2701,N_1832,N_1842);
and U2702 (N_2702,N_1932,N_2378);
nor U2703 (N_2703,N_2077,N_1807);
xnor U2704 (N_2704,N_2366,N_2340);
nand U2705 (N_2705,N_2305,N_2250);
and U2706 (N_2706,N_2306,N_2396);
and U2707 (N_2707,N_2023,N_1879);
and U2708 (N_2708,N_2270,N_2244);
and U2709 (N_2709,N_2194,N_1872);
or U2710 (N_2710,N_1903,N_2319);
and U2711 (N_2711,N_2127,N_1944);
or U2712 (N_2712,N_2011,N_2229);
and U2713 (N_2713,N_1804,N_1991);
nand U2714 (N_2714,N_2283,N_2308);
and U2715 (N_2715,N_2012,N_1889);
xnor U2716 (N_2716,N_2119,N_2081);
and U2717 (N_2717,N_2353,N_1972);
xnor U2718 (N_2718,N_2234,N_2332);
and U2719 (N_2719,N_1803,N_2224);
or U2720 (N_2720,N_1995,N_2117);
or U2721 (N_2721,N_2138,N_2025);
nand U2722 (N_2722,N_1853,N_2109);
nand U2723 (N_2723,N_2313,N_1889);
nand U2724 (N_2724,N_2151,N_2203);
nand U2725 (N_2725,N_1998,N_1949);
nand U2726 (N_2726,N_1951,N_2032);
nand U2727 (N_2727,N_2089,N_2335);
nor U2728 (N_2728,N_2130,N_2216);
nor U2729 (N_2729,N_2195,N_2279);
xor U2730 (N_2730,N_2228,N_2093);
nand U2731 (N_2731,N_1882,N_2338);
nand U2732 (N_2732,N_2361,N_2151);
or U2733 (N_2733,N_2225,N_2271);
xor U2734 (N_2734,N_2357,N_2363);
and U2735 (N_2735,N_2186,N_2318);
or U2736 (N_2736,N_2072,N_1928);
nand U2737 (N_2737,N_2180,N_2163);
nand U2738 (N_2738,N_1929,N_2318);
nor U2739 (N_2739,N_2127,N_2051);
xor U2740 (N_2740,N_1829,N_1857);
and U2741 (N_2741,N_2002,N_2134);
nor U2742 (N_2742,N_2335,N_1909);
xor U2743 (N_2743,N_2303,N_1927);
and U2744 (N_2744,N_2165,N_2221);
and U2745 (N_2745,N_1913,N_1802);
nand U2746 (N_2746,N_1968,N_2394);
nand U2747 (N_2747,N_2227,N_1889);
and U2748 (N_2748,N_2177,N_1986);
nor U2749 (N_2749,N_1964,N_2379);
xor U2750 (N_2750,N_1817,N_2053);
nand U2751 (N_2751,N_2185,N_1930);
nor U2752 (N_2752,N_1823,N_1834);
nor U2753 (N_2753,N_2010,N_2269);
and U2754 (N_2754,N_2191,N_2269);
or U2755 (N_2755,N_1873,N_2154);
or U2756 (N_2756,N_1821,N_2002);
nand U2757 (N_2757,N_2350,N_2001);
nor U2758 (N_2758,N_2075,N_1857);
and U2759 (N_2759,N_1845,N_2308);
nor U2760 (N_2760,N_2308,N_1987);
or U2761 (N_2761,N_2303,N_2182);
nand U2762 (N_2762,N_2309,N_1822);
nand U2763 (N_2763,N_2359,N_1887);
nand U2764 (N_2764,N_1984,N_2127);
and U2765 (N_2765,N_2178,N_1863);
nand U2766 (N_2766,N_1927,N_2267);
nand U2767 (N_2767,N_2217,N_1949);
nor U2768 (N_2768,N_1954,N_2162);
xnor U2769 (N_2769,N_2147,N_2272);
and U2770 (N_2770,N_2113,N_1979);
and U2771 (N_2771,N_2247,N_1816);
nand U2772 (N_2772,N_2045,N_2062);
or U2773 (N_2773,N_2303,N_2116);
and U2774 (N_2774,N_2183,N_2064);
nor U2775 (N_2775,N_2394,N_1845);
xnor U2776 (N_2776,N_2144,N_2333);
and U2777 (N_2777,N_2090,N_2121);
xnor U2778 (N_2778,N_2385,N_2203);
xor U2779 (N_2779,N_2088,N_2333);
nand U2780 (N_2780,N_1909,N_2204);
nor U2781 (N_2781,N_1913,N_2142);
nor U2782 (N_2782,N_1914,N_2222);
nor U2783 (N_2783,N_2018,N_1880);
nor U2784 (N_2784,N_2183,N_2318);
xor U2785 (N_2785,N_1993,N_2354);
nor U2786 (N_2786,N_2371,N_2116);
or U2787 (N_2787,N_2162,N_1956);
or U2788 (N_2788,N_2347,N_1953);
and U2789 (N_2789,N_1980,N_2354);
or U2790 (N_2790,N_1958,N_2272);
nor U2791 (N_2791,N_1845,N_2286);
nor U2792 (N_2792,N_2367,N_2336);
and U2793 (N_2793,N_2251,N_2192);
nor U2794 (N_2794,N_1837,N_1847);
nand U2795 (N_2795,N_2177,N_2220);
or U2796 (N_2796,N_2111,N_2081);
or U2797 (N_2797,N_1880,N_2044);
nor U2798 (N_2798,N_2108,N_2148);
xnor U2799 (N_2799,N_2128,N_2075);
nor U2800 (N_2800,N_2298,N_2128);
xor U2801 (N_2801,N_2247,N_2262);
nand U2802 (N_2802,N_2343,N_1906);
or U2803 (N_2803,N_1868,N_2336);
or U2804 (N_2804,N_2140,N_2329);
xor U2805 (N_2805,N_1872,N_2102);
nor U2806 (N_2806,N_1927,N_2244);
nand U2807 (N_2807,N_2098,N_2034);
or U2808 (N_2808,N_2052,N_2224);
nand U2809 (N_2809,N_2257,N_1817);
or U2810 (N_2810,N_1953,N_1995);
or U2811 (N_2811,N_2267,N_2184);
nand U2812 (N_2812,N_1907,N_2397);
nand U2813 (N_2813,N_2224,N_1925);
nor U2814 (N_2814,N_2200,N_2296);
nand U2815 (N_2815,N_2386,N_2342);
or U2816 (N_2816,N_2357,N_1899);
nand U2817 (N_2817,N_1924,N_1856);
or U2818 (N_2818,N_2188,N_2046);
and U2819 (N_2819,N_1960,N_2030);
nor U2820 (N_2820,N_2187,N_2372);
and U2821 (N_2821,N_2335,N_2219);
xor U2822 (N_2822,N_1912,N_2346);
nand U2823 (N_2823,N_1973,N_1963);
nand U2824 (N_2824,N_2338,N_1839);
and U2825 (N_2825,N_1878,N_1846);
or U2826 (N_2826,N_1930,N_2374);
nand U2827 (N_2827,N_2109,N_2383);
and U2828 (N_2828,N_2029,N_2054);
nor U2829 (N_2829,N_2357,N_2347);
and U2830 (N_2830,N_2364,N_2234);
nand U2831 (N_2831,N_1921,N_2312);
nand U2832 (N_2832,N_1901,N_1949);
nand U2833 (N_2833,N_1956,N_1859);
or U2834 (N_2834,N_2065,N_1979);
nor U2835 (N_2835,N_2253,N_2232);
xor U2836 (N_2836,N_2383,N_2170);
nand U2837 (N_2837,N_2275,N_2131);
and U2838 (N_2838,N_1971,N_2060);
or U2839 (N_2839,N_2091,N_2141);
xnor U2840 (N_2840,N_2228,N_2140);
or U2841 (N_2841,N_2288,N_2202);
or U2842 (N_2842,N_2066,N_2324);
nor U2843 (N_2843,N_2260,N_1927);
nand U2844 (N_2844,N_2367,N_2033);
xnor U2845 (N_2845,N_2308,N_2264);
xnor U2846 (N_2846,N_2374,N_1891);
and U2847 (N_2847,N_1902,N_2124);
xnor U2848 (N_2848,N_2049,N_2052);
nor U2849 (N_2849,N_2069,N_2110);
nand U2850 (N_2850,N_1960,N_1961);
or U2851 (N_2851,N_2382,N_1843);
nand U2852 (N_2852,N_2297,N_1963);
or U2853 (N_2853,N_1921,N_1948);
nor U2854 (N_2854,N_1913,N_1880);
or U2855 (N_2855,N_2170,N_2148);
and U2856 (N_2856,N_2327,N_1816);
nand U2857 (N_2857,N_1856,N_2081);
nand U2858 (N_2858,N_1804,N_2246);
and U2859 (N_2859,N_2363,N_1892);
nand U2860 (N_2860,N_2178,N_2219);
nand U2861 (N_2861,N_2009,N_2354);
xor U2862 (N_2862,N_2306,N_2169);
xnor U2863 (N_2863,N_2353,N_2321);
and U2864 (N_2864,N_2294,N_2211);
and U2865 (N_2865,N_1965,N_1914);
and U2866 (N_2866,N_1901,N_2091);
xor U2867 (N_2867,N_1919,N_1982);
nand U2868 (N_2868,N_2060,N_1827);
xor U2869 (N_2869,N_2065,N_1927);
nor U2870 (N_2870,N_2083,N_2039);
nor U2871 (N_2871,N_2053,N_1943);
xor U2872 (N_2872,N_1828,N_2186);
xnor U2873 (N_2873,N_1843,N_2192);
or U2874 (N_2874,N_1897,N_2248);
nand U2875 (N_2875,N_1923,N_2188);
nor U2876 (N_2876,N_1980,N_2287);
nand U2877 (N_2877,N_2166,N_2202);
and U2878 (N_2878,N_1943,N_1933);
or U2879 (N_2879,N_1912,N_2064);
xnor U2880 (N_2880,N_2194,N_2289);
or U2881 (N_2881,N_2351,N_2045);
nand U2882 (N_2882,N_1860,N_2000);
xor U2883 (N_2883,N_2349,N_1903);
nor U2884 (N_2884,N_2007,N_2176);
xnor U2885 (N_2885,N_2293,N_2276);
nor U2886 (N_2886,N_1966,N_2275);
nor U2887 (N_2887,N_2180,N_1874);
nor U2888 (N_2888,N_1950,N_1840);
xor U2889 (N_2889,N_2164,N_2028);
nand U2890 (N_2890,N_2073,N_2219);
or U2891 (N_2891,N_2120,N_2311);
nor U2892 (N_2892,N_2355,N_1928);
or U2893 (N_2893,N_2268,N_1806);
nor U2894 (N_2894,N_1837,N_2317);
nor U2895 (N_2895,N_2181,N_2011);
nand U2896 (N_2896,N_2204,N_2144);
nor U2897 (N_2897,N_1974,N_2056);
nor U2898 (N_2898,N_2342,N_2378);
or U2899 (N_2899,N_2276,N_2095);
nor U2900 (N_2900,N_2195,N_1830);
nor U2901 (N_2901,N_1927,N_2208);
nor U2902 (N_2902,N_1850,N_1843);
nor U2903 (N_2903,N_1916,N_2176);
xnor U2904 (N_2904,N_2399,N_2228);
xnor U2905 (N_2905,N_2163,N_1995);
nand U2906 (N_2906,N_2161,N_2297);
nand U2907 (N_2907,N_2155,N_1973);
xor U2908 (N_2908,N_1906,N_2268);
nor U2909 (N_2909,N_2195,N_2077);
and U2910 (N_2910,N_2123,N_1874);
xnor U2911 (N_2911,N_2114,N_2159);
or U2912 (N_2912,N_1854,N_2366);
or U2913 (N_2913,N_2307,N_2144);
and U2914 (N_2914,N_2061,N_1862);
and U2915 (N_2915,N_2276,N_2202);
xnor U2916 (N_2916,N_2390,N_1928);
and U2917 (N_2917,N_1805,N_2157);
nor U2918 (N_2918,N_2076,N_2186);
nand U2919 (N_2919,N_2076,N_1867);
xnor U2920 (N_2920,N_2213,N_2183);
and U2921 (N_2921,N_2099,N_2344);
or U2922 (N_2922,N_2387,N_2277);
xor U2923 (N_2923,N_2331,N_1902);
nand U2924 (N_2924,N_2073,N_2106);
nor U2925 (N_2925,N_2018,N_2001);
xor U2926 (N_2926,N_2062,N_2373);
or U2927 (N_2927,N_2277,N_1812);
and U2928 (N_2928,N_2219,N_1845);
xnor U2929 (N_2929,N_2223,N_2334);
or U2930 (N_2930,N_1836,N_2238);
or U2931 (N_2931,N_1813,N_1893);
nor U2932 (N_2932,N_2203,N_1903);
xnor U2933 (N_2933,N_2255,N_2263);
or U2934 (N_2934,N_1815,N_1920);
nand U2935 (N_2935,N_2133,N_2254);
and U2936 (N_2936,N_1859,N_2247);
xor U2937 (N_2937,N_1857,N_1885);
nor U2938 (N_2938,N_2133,N_1913);
nor U2939 (N_2939,N_1876,N_2247);
or U2940 (N_2940,N_2379,N_2108);
nand U2941 (N_2941,N_2262,N_1957);
nand U2942 (N_2942,N_1972,N_1814);
nand U2943 (N_2943,N_2177,N_1971);
nand U2944 (N_2944,N_1936,N_2372);
and U2945 (N_2945,N_1873,N_2325);
nand U2946 (N_2946,N_1939,N_2177);
and U2947 (N_2947,N_2175,N_2253);
or U2948 (N_2948,N_1884,N_2283);
or U2949 (N_2949,N_2263,N_1998);
nand U2950 (N_2950,N_2101,N_2027);
xor U2951 (N_2951,N_2295,N_2238);
xnor U2952 (N_2952,N_2353,N_1930);
nand U2953 (N_2953,N_2369,N_2334);
nor U2954 (N_2954,N_2081,N_2030);
xor U2955 (N_2955,N_2189,N_2230);
xor U2956 (N_2956,N_2271,N_2038);
xor U2957 (N_2957,N_1982,N_2375);
or U2958 (N_2958,N_2073,N_2186);
xnor U2959 (N_2959,N_1936,N_2319);
or U2960 (N_2960,N_2255,N_1836);
xnor U2961 (N_2961,N_2330,N_1854);
xnor U2962 (N_2962,N_2007,N_1839);
and U2963 (N_2963,N_2102,N_2141);
and U2964 (N_2964,N_2138,N_2059);
or U2965 (N_2965,N_1855,N_2264);
or U2966 (N_2966,N_2090,N_2075);
nor U2967 (N_2967,N_2170,N_2058);
nor U2968 (N_2968,N_1895,N_2155);
nand U2969 (N_2969,N_2270,N_2250);
or U2970 (N_2970,N_2399,N_2392);
xor U2971 (N_2971,N_2103,N_2217);
or U2972 (N_2972,N_2075,N_2367);
and U2973 (N_2973,N_1878,N_2301);
or U2974 (N_2974,N_2378,N_2231);
and U2975 (N_2975,N_2010,N_1949);
xnor U2976 (N_2976,N_1839,N_2023);
and U2977 (N_2977,N_1966,N_1994);
xnor U2978 (N_2978,N_2300,N_1855);
and U2979 (N_2979,N_2266,N_2276);
nand U2980 (N_2980,N_2243,N_2150);
and U2981 (N_2981,N_2136,N_1953);
xor U2982 (N_2982,N_2002,N_2174);
nor U2983 (N_2983,N_2002,N_1970);
nand U2984 (N_2984,N_2174,N_2023);
xor U2985 (N_2985,N_2260,N_1901);
xnor U2986 (N_2986,N_2380,N_1946);
and U2987 (N_2987,N_2173,N_2271);
xor U2988 (N_2988,N_2047,N_2097);
and U2989 (N_2989,N_2221,N_1875);
or U2990 (N_2990,N_2126,N_2221);
or U2991 (N_2991,N_1886,N_1821);
nand U2992 (N_2992,N_2353,N_1896);
nor U2993 (N_2993,N_1815,N_2299);
nor U2994 (N_2994,N_1916,N_2036);
and U2995 (N_2995,N_2377,N_1956);
nand U2996 (N_2996,N_1890,N_2116);
xor U2997 (N_2997,N_2191,N_1893);
nand U2998 (N_2998,N_1950,N_2217);
nand U2999 (N_2999,N_2175,N_2374);
and UO_0 (O_0,N_2476,N_2739);
nand UO_1 (O_1,N_2964,N_2929);
nor UO_2 (O_2,N_2803,N_2994);
xor UO_3 (O_3,N_2794,N_2896);
nor UO_4 (O_4,N_2636,N_2804);
xnor UO_5 (O_5,N_2858,N_2546);
nor UO_6 (O_6,N_2903,N_2710);
or UO_7 (O_7,N_2860,N_2509);
xor UO_8 (O_8,N_2721,N_2902);
and UO_9 (O_9,N_2652,N_2642);
nand UO_10 (O_10,N_2879,N_2907);
and UO_11 (O_11,N_2746,N_2419);
nand UO_12 (O_12,N_2665,N_2944);
nand UO_13 (O_13,N_2745,N_2431);
nor UO_14 (O_14,N_2924,N_2428);
nand UO_15 (O_15,N_2468,N_2751);
nand UO_16 (O_16,N_2409,N_2748);
nor UO_17 (O_17,N_2969,N_2884);
xnor UO_18 (O_18,N_2706,N_2436);
nand UO_19 (O_19,N_2893,N_2894);
or UO_20 (O_20,N_2523,N_2805);
xor UO_21 (O_21,N_2811,N_2559);
nand UO_22 (O_22,N_2480,N_2566);
xor UO_23 (O_23,N_2795,N_2998);
xor UO_24 (O_24,N_2897,N_2533);
nor UO_25 (O_25,N_2977,N_2458);
nand UO_26 (O_26,N_2440,N_2908);
xor UO_27 (O_27,N_2762,N_2914);
xor UO_28 (O_28,N_2404,N_2779);
or UO_29 (O_29,N_2420,N_2841);
and UO_30 (O_30,N_2500,N_2617);
nor UO_31 (O_31,N_2493,N_2402);
nor UO_32 (O_32,N_2590,N_2542);
xor UO_33 (O_33,N_2560,N_2750);
xor UO_34 (O_34,N_2901,N_2687);
or UO_35 (O_35,N_2938,N_2427);
and UO_36 (O_36,N_2928,N_2505);
or UO_37 (O_37,N_2723,N_2892);
xnor UO_38 (O_38,N_2796,N_2904);
xor UO_39 (O_39,N_2960,N_2640);
nor UO_40 (O_40,N_2953,N_2962);
nand UO_41 (O_41,N_2465,N_2780);
nor UO_42 (O_42,N_2595,N_2774);
nand UO_43 (O_43,N_2426,N_2555);
or UO_44 (O_44,N_2806,N_2678);
nor UO_45 (O_45,N_2781,N_2684);
or UO_46 (O_46,N_2733,N_2987);
nor UO_47 (O_47,N_2663,N_2722);
nor UO_48 (O_48,N_2838,N_2947);
xnor UO_49 (O_49,N_2561,N_2618);
xor UO_50 (O_50,N_2454,N_2418);
nor UO_51 (O_51,N_2443,N_2726);
nor UO_52 (O_52,N_2868,N_2708);
xnor UO_53 (O_53,N_2818,N_2905);
and UO_54 (O_54,N_2898,N_2686);
xnor UO_55 (O_55,N_2830,N_2582);
xnor UO_56 (O_56,N_2408,N_2629);
nand UO_57 (O_57,N_2494,N_2876);
nor UO_58 (O_58,N_2516,N_2588);
and UO_59 (O_59,N_2850,N_2675);
and UO_60 (O_60,N_2571,N_2909);
and UO_61 (O_61,N_2943,N_2683);
nor UO_62 (O_62,N_2615,N_2452);
xor UO_63 (O_63,N_2627,N_2954);
or UO_64 (O_64,N_2711,N_2548);
xnor UO_65 (O_65,N_2633,N_2719);
and UO_66 (O_66,N_2579,N_2670);
xnor UO_67 (O_67,N_2882,N_2713);
nand UO_68 (O_68,N_2718,N_2671);
nor UO_69 (O_69,N_2421,N_2931);
or UO_70 (O_70,N_2643,N_2935);
and UO_71 (O_71,N_2410,N_2932);
nor UO_72 (O_72,N_2478,N_2600);
xor UO_73 (O_73,N_2502,N_2715);
and UO_74 (O_74,N_2470,N_2535);
and UO_75 (O_75,N_2517,N_2575);
or UO_76 (O_76,N_2587,N_2817);
xor UO_77 (O_77,N_2814,N_2842);
nand UO_78 (O_78,N_2870,N_2689);
or UO_79 (O_79,N_2758,N_2699);
xnor UO_80 (O_80,N_2867,N_2741);
nor UO_81 (O_81,N_2784,N_2596);
nand UO_82 (O_82,N_2793,N_2639);
and UO_83 (O_83,N_2651,N_2936);
nor UO_84 (O_84,N_2414,N_2716);
and UO_85 (O_85,N_2899,N_2637);
or UO_86 (O_86,N_2744,N_2520);
nand UO_87 (O_87,N_2433,N_2484);
and UO_88 (O_88,N_2623,N_2564);
and UO_89 (O_89,N_2845,N_2531);
or UO_90 (O_90,N_2926,N_2536);
and UO_91 (O_91,N_2967,N_2720);
nand UO_92 (O_92,N_2910,N_2401);
nand UO_93 (O_93,N_2406,N_2598);
nor UO_94 (O_94,N_2562,N_2752);
and UO_95 (O_95,N_2812,N_2423);
and UO_96 (O_96,N_2990,N_2819);
or UO_97 (O_97,N_2768,N_2906);
and UO_98 (O_98,N_2513,N_2757);
nand UO_99 (O_99,N_2847,N_2585);
nor UO_100 (O_100,N_2444,N_2974);
xor UO_101 (O_101,N_2527,N_2833);
or UO_102 (O_102,N_2995,N_2705);
or UO_103 (O_103,N_2547,N_2690);
nand UO_104 (O_104,N_2735,N_2952);
and UO_105 (O_105,N_2603,N_2495);
and UO_106 (O_106,N_2552,N_2473);
and UO_107 (O_107,N_2696,N_2597);
and UO_108 (O_108,N_2619,N_2791);
or UO_109 (O_109,N_2655,N_2872);
nor UO_110 (O_110,N_2407,N_2518);
nand UO_111 (O_111,N_2790,N_2773);
and UO_112 (O_112,N_2631,N_2415);
and UO_113 (O_113,N_2992,N_2761);
nand UO_114 (O_114,N_2949,N_2709);
nor UO_115 (O_115,N_2688,N_2921);
or UO_116 (O_116,N_2883,N_2797);
or UO_117 (O_117,N_2770,N_2424);
nand UO_118 (O_118,N_2743,N_2783);
nor UO_119 (O_119,N_2612,N_2856);
xor UO_120 (O_120,N_2788,N_2417);
or UO_121 (O_121,N_2490,N_2422);
nor UO_122 (O_122,N_2455,N_2767);
xor UO_123 (O_123,N_2601,N_2591);
nor UO_124 (O_124,N_2725,N_2625);
xnor UO_125 (O_125,N_2732,N_2568);
nor UO_126 (O_126,N_2835,N_2738);
xor UO_127 (O_127,N_2873,N_2650);
and UO_128 (O_128,N_2832,N_2963);
nand UO_129 (O_129,N_2462,N_2945);
nand UO_130 (O_130,N_2869,N_2874);
and UO_131 (O_131,N_2460,N_2890);
xor UO_132 (O_132,N_2975,N_2809);
and UO_133 (O_133,N_2772,N_2888);
nand UO_134 (O_134,N_2979,N_2859);
xor UO_135 (O_135,N_2742,N_2474);
xnor UO_136 (O_136,N_2503,N_2672);
or UO_137 (O_137,N_2605,N_2983);
and UO_138 (O_138,N_2815,N_2464);
or UO_139 (O_139,N_2463,N_2438);
nand UO_140 (O_140,N_2567,N_2729);
nor UO_141 (O_141,N_2666,N_2577);
xnor UO_142 (O_142,N_2753,N_2545);
nor UO_143 (O_143,N_2430,N_2965);
and UO_144 (O_144,N_2429,N_2578);
xnor UO_145 (O_145,N_2829,N_2680);
nand UO_146 (O_146,N_2487,N_2456);
and UO_147 (O_147,N_2861,N_2707);
nor UO_148 (O_148,N_2581,N_2446);
or UO_149 (O_149,N_2466,N_2717);
nand UO_150 (O_150,N_2556,N_2912);
nand UO_151 (O_151,N_2628,N_2886);
or UO_152 (O_152,N_2692,N_2471);
or UO_153 (O_153,N_2824,N_2828);
xnor UO_154 (O_154,N_2712,N_2816);
nand UO_155 (O_155,N_2498,N_2755);
or UO_156 (O_156,N_2855,N_2827);
or UO_157 (O_157,N_2594,N_2918);
and UO_158 (O_158,N_2551,N_2731);
nand UO_159 (O_159,N_2934,N_2925);
nand UO_160 (O_160,N_2413,N_2988);
nand UO_161 (O_161,N_2632,N_2878);
or UO_162 (O_162,N_2543,N_2403);
nor UO_163 (O_163,N_2800,N_2854);
or UO_164 (O_164,N_2961,N_2572);
and UO_165 (O_165,N_2769,N_2785);
nand UO_166 (O_166,N_2787,N_2837);
xnor UO_167 (O_167,N_2621,N_2823);
or UO_168 (O_168,N_2849,N_2626);
and UO_169 (O_169,N_2589,N_2702);
and UO_170 (O_170,N_2584,N_2442);
nand UO_171 (O_171,N_2537,N_2563);
xor UO_172 (O_172,N_2756,N_2865);
nand UO_173 (O_173,N_2461,N_2459);
nand UO_174 (O_174,N_2662,N_2411);
or UO_175 (O_175,N_2948,N_2540);
or UO_176 (O_176,N_2959,N_2432);
nor UO_177 (O_177,N_2613,N_2911);
nand UO_178 (O_178,N_2654,N_2647);
xnor UO_179 (O_179,N_2864,N_2951);
xnor UO_180 (O_180,N_2851,N_2986);
xnor UO_181 (O_181,N_2942,N_2734);
nand UO_182 (O_182,N_2558,N_2553);
nand UO_183 (O_183,N_2669,N_2507);
xor UO_184 (O_184,N_2481,N_2622);
nand UO_185 (O_185,N_2754,N_2514);
nor UO_186 (O_186,N_2808,N_2610);
or UO_187 (O_187,N_2641,N_2919);
and UO_188 (O_188,N_2497,N_2747);
nand UO_189 (O_189,N_2766,N_2810);
or UO_190 (O_190,N_2698,N_2950);
nand UO_191 (O_191,N_2853,N_2638);
and UO_192 (O_192,N_2989,N_2664);
or UO_193 (O_193,N_2501,N_2997);
and UO_194 (O_194,N_2616,N_2656);
nand UO_195 (O_195,N_2544,N_2852);
nor UO_196 (O_196,N_2940,N_2844);
and UO_197 (O_197,N_2957,N_2915);
nand UO_198 (O_198,N_2922,N_2450);
xnor UO_199 (O_199,N_2441,N_2661);
xor UO_200 (O_200,N_2447,N_2880);
and UO_201 (O_201,N_2697,N_2649);
nand UO_202 (O_202,N_2453,N_2539);
and UO_203 (O_203,N_2993,N_2802);
xnor UO_204 (O_204,N_2982,N_2524);
nand UO_205 (O_205,N_2831,N_2614);
nor UO_206 (O_206,N_2703,N_2435);
nor UO_207 (O_207,N_2472,N_2635);
nor UO_208 (O_208,N_2515,N_2510);
nand UO_209 (O_209,N_2630,N_2887);
nor UO_210 (O_210,N_2857,N_2846);
nor UO_211 (O_211,N_2512,N_2530);
and UO_212 (O_212,N_2984,N_2607);
and UO_213 (O_213,N_2765,N_2620);
nor UO_214 (O_214,N_2674,N_2866);
and UO_215 (O_215,N_2681,N_2848);
and UO_216 (O_216,N_2956,N_2927);
xor UO_217 (O_217,N_2682,N_2400);
and UO_218 (O_218,N_2467,N_2593);
and UO_219 (O_219,N_2759,N_2599);
xnor UO_220 (O_220,N_2881,N_2968);
nor UO_221 (O_221,N_2506,N_2714);
xnor UO_222 (O_222,N_2786,N_2668);
and UO_223 (O_223,N_2840,N_2519);
xor UO_224 (O_224,N_2492,N_2801);
or UO_225 (O_225,N_2653,N_2798);
and UO_226 (O_226,N_2775,N_2491);
nor UO_227 (O_227,N_2972,N_2538);
nand UO_228 (O_228,N_2736,N_2966);
xor UO_229 (O_229,N_2475,N_2891);
or UO_230 (O_230,N_2836,N_2822);
nand UO_231 (O_231,N_2496,N_2526);
nor UO_232 (O_232,N_2807,N_2659);
nor UO_233 (O_233,N_2958,N_2937);
and UO_234 (O_234,N_2602,N_2978);
nand UO_235 (O_235,N_2673,N_2624);
and UO_236 (O_236,N_2933,N_2724);
nor UO_237 (O_237,N_2991,N_2694);
or UO_238 (O_238,N_2416,N_2508);
and UO_239 (O_239,N_2477,N_2955);
xor UO_240 (O_240,N_2917,N_2875);
nand UO_241 (O_241,N_2693,N_2946);
nand UO_242 (O_242,N_2405,N_2486);
and UO_243 (O_243,N_2685,N_2550);
nor UO_244 (O_244,N_2980,N_2541);
or UO_245 (O_245,N_2691,N_2499);
or UO_246 (O_246,N_2425,N_2843);
and UO_247 (O_247,N_2820,N_2437);
nor UO_248 (O_248,N_2985,N_2789);
nor UO_249 (O_249,N_2608,N_2760);
nand UO_250 (O_250,N_2549,N_2728);
nor UO_251 (O_251,N_2439,N_2970);
nand UO_252 (O_252,N_2451,N_2586);
nor UO_253 (O_253,N_2634,N_2877);
nand UO_254 (O_254,N_2448,N_2569);
xnor UO_255 (O_255,N_2782,N_2996);
and UO_256 (O_256,N_2862,N_2825);
nor UO_257 (O_257,N_2565,N_2525);
xor UO_258 (O_258,N_2604,N_2580);
and UO_259 (O_259,N_2973,N_2763);
and UO_260 (O_260,N_2749,N_2667);
xor UO_261 (O_261,N_2792,N_2930);
nor UO_262 (O_262,N_2971,N_2813);
or UO_263 (O_263,N_2863,N_2777);
and UO_264 (O_264,N_2557,N_2412);
or UO_265 (O_265,N_2457,N_2695);
and UO_266 (O_266,N_2704,N_2727);
xor UO_267 (O_267,N_2923,N_2449);
xor UO_268 (O_268,N_2871,N_2889);
nand UO_269 (O_269,N_2445,N_2981);
xnor UO_270 (O_270,N_2916,N_2677);
xnor UO_271 (O_271,N_2488,N_2469);
nand UO_272 (O_272,N_2576,N_2839);
xnor UO_273 (O_273,N_2489,N_2485);
nor UO_274 (O_274,N_2737,N_2657);
nor UO_275 (O_275,N_2939,N_2999);
xor UO_276 (O_276,N_2764,N_2554);
xor UO_277 (O_277,N_2821,N_2611);
or UO_278 (O_278,N_2776,N_2976);
nand UO_279 (O_279,N_2529,N_2482);
and UO_280 (O_280,N_2895,N_2532);
or UO_281 (O_281,N_2730,N_2522);
xnor UO_282 (O_282,N_2913,N_2504);
nand UO_283 (O_283,N_2479,N_2574);
nand UO_284 (O_284,N_2676,N_2606);
xor UO_285 (O_285,N_2570,N_2646);
nand UO_286 (O_286,N_2679,N_2573);
nand UO_287 (O_287,N_2592,N_2583);
and UO_288 (O_288,N_2700,N_2778);
and UO_289 (O_289,N_2660,N_2920);
xnor UO_290 (O_290,N_2528,N_2900);
nand UO_291 (O_291,N_2511,N_2644);
nand UO_292 (O_292,N_2483,N_2740);
or UO_293 (O_293,N_2534,N_2645);
nor UO_294 (O_294,N_2434,N_2771);
and UO_295 (O_295,N_2658,N_2826);
xnor UO_296 (O_296,N_2799,N_2941);
nand UO_297 (O_297,N_2609,N_2885);
xnor UO_298 (O_298,N_2648,N_2701);
xnor UO_299 (O_299,N_2834,N_2521);
nor UO_300 (O_300,N_2466,N_2607);
nand UO_301 (O_301,N_2934,N_2433);
or UO_302 (O_302,N_2592,N_2503);
nand UO_303 (O_303,N_2558,N_2596);
nor UO_304 (O_304,N_2696,N_2738);
nand UO_305 (O_305,N_2505,N_2675);
or UO_306 (O_306,N_2570,N_2790);
nand UO_307 (O_307,N_2701,N_2946);
nand UO_308 (O_308,N_2726,N_2429);
or UO_309 (O_309,N_2943,N_2681);
xnor UO_310 (O_310,N_2974,N_2926);
and UO_311 (O_311,N_2608,N_2457);
nand UO_312 (O_312,N_2956,N_2545);
nand UO_313 (O_313,N_2801,N_2915);
and UO_314 (O_314,N_2948,N_2901);
and UO_315 (O_315,N_2924,N_2868);
nor UO_316 (O_316,N_2623,N_2578);
nand UO_317 (O_317,N_2923,N_2876);
nand UO_318 (O_318,N_2996,N_2421);
nor UO_319 (O_319,N_2834,N_2714);
and UO_320 (O_320,N_2570,N_2814);
nand UO_321 (O_321,N_2659,N_2622);
xor UO_322 (O_322,N_2840,N_2911);
nand UO_323 (O_323,N_2779,N_2895);
xor UO_324 (O_324,N_2599,N_2979);
xnor UO_325 (O_325,N_2844,N_2484);
and UO_326 (O_326,N_2652,N_2855);
or UO_327 (O_327,N_2599,N_2885);
or UO_328 (O_328,N_2608,N_2789);
or UO_329 (O_329,N_2732,N_2961);
or UO_330 (O_330,N_2981,N_2812);
nor UO_331 (O_331,N_2982,N_2953);
xnor UO_332 (O_332,N_2696,N_2635);
or UO_333 (O_333,N_2536,N_2553);
xor UO_334 (O_334,N_2537,N_2647);
xnor UO_335 (O_335,N_2768,N_2908);
nor UO_336 (O_336,N_2928,N_2624);
nand UO_337 (O_337,N_2604,N_2462);
xor UO_338 (O_338,N_2689,N_2765);
nor UO_339 (O_339,N_2600,N_2617);
xnor UO_340 (O_340,N_2978,N_2559);
or UO_341 (O_341,N_2815,N_2589);
nand UO_342 (O_342,N_2754,N_2489);
and UO_343 (O_343,N_2538,N_2963);
and UO_344 (O_344,N_2429,N_2706);
nor UO_345 (O_345,N_2611,N_2796);
and UO_346 (O_346,N_2566,N_2733);
xnor UO_347 (O_347,N_2765,N_2407);
xor UO_348 (O_348,N_2822,N_2706);
xor UO_349 (O_349,N_2789,N_2826);
nor UO_350 (O_350,N_2420,N_2515);
and UO_351 (O_351,N_2522,N_2844);
xnor UO_352 (O_352,N_2409,N_2430);
nand UO_353 (O_353,N_2594,N_2870);
and UO_354 (O_354,N_2943,N_2576);
nor UO_355 (O_355,N_2583,N_2608);
or UO_356 (O_356,N_2643,N_2464);
xor UO_357 (O_357,N_2555,N_2453);
xor UO_358 (O_358,N_2980,N_2738);
nor UO_359 (O_359,N_2821,N_2628);
and UO_360 (O_360,N_2950,N_2597);
nand UO_361 (O_361,N_2826,N_2889);
nor UO_362 (O_362,N_2722,N_2960);
and UO_363 (O_363,N_2604,N_2735);
and UO_364 (O_364,N_2946,N_2511);
nor UO_365 (O_365,N_2943,N_2735);
and UO_366 (O_366,N_2648,N_2966);
xor UO_367 (O_367,N_2741,N_2476);
nor UO_368 (O_368,N_2884,N_2982);
and UO_369 (O_369,N_2863,N_2613);
and UO_370 (O_370,N_2624,N_2783);
xor UO_371 (O_371,N_2460,N_2794);
nand UO_372 (O_372,N_2995,N_2653);
nor UO_373 (O_373,N_2743,N_2652);
nand UO_374 (O_374,N_2843,N_2520);
xor UO_375 (O_375,N_2981,N_2525);
nand UO_376 (O_376,N_2461,N_2934);
and UO_377 (O_377,N_2802,N_2443);
or UO_378 (O_378,N_2589,N_2462);
nor UO_379 (O_379,N_2642,N_2428);
nor UO_380 (O_380,N_2941,N_2648);
xnor UO_381 (O_381,N_2599,N_2415);
xor UO_382 (O_382,N_2755,N_2818);
or UO_383 (O_383,N_2580,N_2948);
nand UO_384 (O_384,N_2631,N_2747);
and UO_385 (O_385,N_2478,N_2759);
nand UO_386 (O_386,N_2898,N_2699);
nand UO_387 (O_387,N_2632,N_2985);
nand UO_388 (O_388,N_2995,N_2475);
or UO_389 (O_389,N_2986,N_2935);
xor UO_390 (O_390,N_2527,N_2733);
or UO_391 (O_391,N_2402,N_2936);
xor UO_392 (O_392,N_2977,N_2747);
nand UO_393 (O_393,N_2865,N_2937);
or UO_394 (O_394,N_2792,N_2447);
nand UO_395 (O_395,N_2887,N_2614);
nand UO_396 (O_396,N_2900,N_2744);
nand UO_397 (O_397,N_2576,N_2910);
nand UO_398 (O_398,N_2597,N_2946);
and UO_399 (O_399,N_2854,N_2964);
nor UO_400 (O_400,N_2496,N_2998);
xnor UO_401 (O_401,N_2565,N_2974);
and UO_402 (O_402,N_2708,N_2926);
or UO_403 (O_403,N_2513,N_2519);
and UO_404 (O_404,N_2552,N_2612);
nor UO_405 (O_405,N_2446,N_2688);
or UO_406 (O_406,N_2873,N_2879);
or UO_407 (O_407,N_2675,N_2840);
and UO_408 (O_408,N_2959,N_2748);
and UO_409 (O_409,N_2471,N_2957);
xnor UO_410 (O_410,N_2530,N_2864);
xnor UO_411 (O_411,N_2824,N_2654);
and UO_412 (O_412,N_2474,N_2866);
nor UO_413 (O_413,N_2618,N_2773);
nor UO_414 (O_414,N_2764,N_2753);
and UO_415 (O_415,N_2900,N_2690);
xor UO_416 (O_416,N_2752,N_2815);
nand UO_417 (O_417,N_2840,N_2958);
nand UO_418 (O_418,N_2730,N_2587);
xnor UO_419 (O_419,N_2886,N_2865);
nor UO_420 (O_420,N_2476,N_2733);
nand UO_421 (O_421,N_2773,N_2706);
or UO_422 (O_422,N_2443,N_2842);
nand UO_423 (O_423,N_2812,N_2898);
nor UO_424 (O_424,N_2865,N_2769);
or UO_425 (O_425,N_2957,N_2580);
xnor UO_426 (O_426,N_2443,N_2487);
nor UO_427 (O_427,N_2863,N_2951);
or UO_428 (O_428,N_2905,N_2558);
xor UO_429 (O_429,N_2686,N_2431);
nor UO_430 (O_430,N_2624,N_2681);
or UO_431 (O_431,N_2884,N_2805);
nor UO_432 (O_432,N_2708,N_2949);
or UO_433 (O_433,N_2688,N_2624);
nand UO_434 (O_434,N_2817,N_2762);
xor UO_435 (O_435,N_2846,N_2559);
or UO_436 (O_436,N_2594,N_2887);
xnor UO_437 (O_437,N_2865,N_2950);
nand UO_438 (O_438,N_2903,N_2528);
nand UO_439 (O_439,N_2478,N_2589);
or UO_440 (O_440,N_2485,N_2558);
or UO_441 (O_441,N_2637,N_2875);
and UO_442 (O_442,N_2415,N_2427);
nor UO_443 (O_443,N_2864,N_2790);
and UO_444 (O_444,N_2753,N_2466);
nor UO_445 (O_445,N_2993,N_2688);
xnor UO_446 (O_446,N_2984,N_2905);
nand UO_447 (O_447,N_2616,N_2770);
nand UO_448 (O_448,N_2466,N_2925);
nor UO_449 (O_449,N_2752,N_2578);
nor UO_450 (O_450,N_2646,N_2713);
or UO_451 (O_451,N_2710,N_2802);
nor UO_452 (O_452,N_2736,N_2699);
nand UO_453 (O_453,N_2772,N_2992);
nor UO_454 (O_454,N_2503,N_2720);
or UO_455 (O_455,N_2588,N_2700);
and UO_456 (O_456,N_2569,N_2708);
nand UO_457 (O_457,N_2464,N_2842);
nor UO_458 (O_458,N_2500,N_2885);
or UO_459 (O_459,N_2744,N_2979);
or UO_460 (O_460,N_2796,N_2404);
nor UO_461 (O_461,N_2653,N_2427);
nand UO_462 (O_462,N_2489,N_2568);
or UO_463 (O_463,N_2519,N_2421);
nand UO_464 (O_464,N_2932,N_2619);
xnor UO_465 (O_465,N_2744,N_2569);
xor UO_466 (O_466,N_2465,N_2969);
xnor UO_467 (O_467,N_2864,N_2603);
nor UO_468 (O_468,N_2963,N_2745);
nor UO_469 (O_469,N_2901,N_2588);
nor UO_470 (O_470,N_2640,N_2478);
or UO_471 (O_471,N_2586,N_2471);
nand UO_472 (O_472,N_2976,N_2703);
or UO_473 (O_473,N_2623,N_2705);
xor UO_474 (O_474,N_2644,N_2645);
and UO_475 (O_475,N_2944,N_2534);
and UO_476 (O_476,N_2686,N_2827);
nand UO_477 (O_477,N_2461,N_2607);
nand UO_478 (O_478,N_2831,N_2575);
and UO_479 (O_479,N_2446,N_2815);
and UO_480 (O_480,N_2853,N_2701);
nor UO_481 (O_481,N_2511,N_2523);
xnor UO_482 (O_482,N_2965,N_2970);
or UO_483 (O_483,N_2673,N_2757);
or UO_484 (O_484,N_2528,N_2464);
xor UO_485 (O_485,N_2508,N_2438);
or UO_486 (O_486,N_2628,N_2616);
nor UO_487 (O_487,N_2724,N_2557);
and UO_488 (O_488,N_2404,N_2467);
xnor UO_489 (O_489,N_2539,N_2626);
nand UO_490 (O_490,N_2946,N_2569);
xor UO_491 (O_491,N_2920,N_2550);
and UO_492 (O_492,N_2949,N_2774);
or UO_493 (O_493,N_2849,N_2941);
xnor UO_494 (O_494,N_2620,N_2417);
xor UO_495 (O_495,N_2818,N_2569);
nand UO_496 (O_496,N_2884,N_2484);
nor UO_497 (O_497,N_2580,N_2491);
nand UO_498 (O_498,N_2691,N_2403);
nand UO_499 (O_499,N_2957,N_2917);
endmodule