module basic_1000_10000_1500_50_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
and U0 (N_0,In_670,In_483);
xnor U1 (N_1,In_639,In_431);
or U2 (N_2,In_692,In_360);
nand U3 (N_3,In_420,In_939);
and U4 (N_4,In_791,In_212);
nand U5 (N_5,In_895,In_123);
xor U6 (N_6,In_761,In_259);
and U7 (N_7,In_814,In_587);
or U8 (N_8,In_163,In_345);
and U9 (N_9,In_595,In_580);
xnor U10 (N_10,In_645,In_975);
nor U11 (N_11,In_144,In_781);
nand U12 (N_12,In_347,In_170);
nand U13 (N_13,In_450,In_547);
nand U14 (N_14,In_344,In_885);
or U15 (N_15,In_97,In_999);
xnor U16 (N_16,In_55,In_494);
nand U17 (N_17,In_278,In_500);
nor U18 (N_18,In_63,In_575);
xnor U19 (N_19,In_216,In_410);
nor U20 (N_20,In_658,In_510);
xor U21 (N_21,In_441,In_870);
and U22 (N_22,In_274,In_523);
or U23 (N_23,In_768,In_798);
nor U24 (N_24,In_774,In_140);
and U25 (N_25,In_795,In_377);
and U26 (N_26,In_88,In_730);
or U27 (N_27,In_907,In_892);
nand U28 (N_28,In_602,In_74);
xor U29 (N_29,In_598,In_363);
nand U30 (N_30,In_825,In_970);
nor U31 (N_31,In_766,In_669);
xor U32 (N_32,In_506,In_303);
nand U33 (N_33,In_818,In_644);
nor U34 (N_34,In_316,In_596);
nor U35 (N_35,In_79,In_529);
nor U36 (N_36,In_401,In_439);
nor U37 (N_37,In_414,In_810);
xor U38 (N_38,In_426,In_495);
xnor U39 (N_39,In_754,In_972);
xor U40 (N_40,In_926,In_748);
xor U41 (N_41,In_49,In_464);
xnor U42 (N_42,In_826,In_807);
xor U43 (N_43,In_951,In_735);
nor U44 (N_44,In_704,In_663);
and U45 (N_45,In_337,In_332);
nor U46 (N_46,In_200,In_508);
and U47 (N_47,In_260,In_214);
nor U48 (N_48,In_513,In_722);
xnor U49 (N_49,In_91,In_531);
nor U50 (N_50,In_582,In_412);
nand U51 (N_51,In_484,In_434);
xnor U52 (N_52,In_243,In_908);
nor U53 (N_53,In_89,In_779);
or U54 (N_54,In_323,In_339);
and U55 (N_55,In_697,In_737);
or U56 (N_56,In_119,In_935);
or U57 (N_57,In_720,In_78);
nand U58 (N_58,In_925,In_35);
or U59 (N_59,In_906,In_958);
or U60 (N_60,In_364,In_640);
and U61 (N_61,In_492,In_609);
xnor U62 (N_62,In_237,In_10);
or U63 (N_63,In_399,In_176);
nand U64 (N_64,In_920,In_558);
xnor U65 (N_65,In_728,In_762);
and U66 (N_66,In_330,In_246);
xor U67 (N_67,In_563,In_184);
nand U68 (N_68,In_812,In_108);
and U69 (N_69,In_477,In_352);
and U70 (N_70,In_808,In_594);
or U71 (N_71,In_665,In_425);
xor U72 (N_72,In_777,In_631);
nand U73 (N_73,In_372,In_806);
xor U74 (N_74,In_819,In_677);
or U75 (N_75,In_309,In_950);
xor U76 (N_76,In_385,In_158);
nand U77 (N_77,In_11,In_784);
xor U78 (N_78,In_226,In_980);
or U79 (N_79,In_407,In_853);
xor U80 (N_80,In_541,In_205);
nand U81 (N_81,In_866,In_509);
nand U82 (N_82,In_874,In_817);
nand U83 (N_83,In_206,In_955);
xnor U84 (N_84,In_707,In_335);
nand U85 (N_85,In_408,In_979);
xnor U86 (N_86,In_277,In_124);
and U87 (N_87,In_307,In_788);
xnor U88 (N_88,In_954,In_799);
or U89 (N_89,In_914,In_72);
nand U90 (N_90,In_963,In_695);
and U91 (N_91,In_183,In_660);
or U92 (N_92,In_288,In_753);
and U93 (N_93,In_440,In_394);
and U94 (N_94,In_376,In_462);
nor U95 (N_95,In_305,In_13);
and U96 (N_96,In_579,In_395);
xor U97 (N_97,In_387,In_952);
nor U98 (N_98,In_890,In_336);
nand U99 (N_99,In_936,In_151);
or U100 (N_100,In_396,In_931);
xor U101 (N_101,In_685,In_282);
nor U102 (N_102,In_624,In_995);
nand U103 (N_103,In_867,In_365);
and U104 (N_104,In_153,In_900);
nor U105 (N_105,In_776,In_630);
nand U106 (N_106,In_789,In_195);
and U107 (N_107,In_542,In_133);
and U108 (N_108,In_850,In_836);
nor U109 (N_109,In_493,In_422);
nand U110 (N_110,In_338,In_256);
xnor U111 (N_111,In_66,In_27);
or U112 (N_112,In_327,In_266);
nand U113 (N_113,In_985,In_75);
nor U114 (N_114,In_272,In_374);
nor U115 (N_115,In_267,In_934);
nor U116 (N_116,In_815,In_947);
or U117 (N_117,In_570,In_486);
nor U118 (N_118,In_326,In_354);
nor U119 (N_119,In_681,In_647);
nand U120 (N_120,In_472,In_627);
and U121 (N_121,In_312,In_99);
nand U122 (N_122,In_504,In_898);
and U123 (N_123,In_94,In_592);
or U124 (N_124,In_359,In_161);
nand U125 (N_125,In_743,In_904);
or U126 (N_126,In_865,In_745);
and U127 (N_127,In_383,In_240);
nor U128 (N_128,In_899,In_751);
nor U129 (N_129,In_71,In_933);
and U130 (N_130,In_527,In_519);
nand U131 (N_131,In_992,In_51);
or U132 (N_132,In_969,In_576);
xnor U133 (N_133,In_386,In_785);
and U134 (N_134,In_971,In_371);
xor U135 (N_135,In_569,In_370);
xnor U136 (N_136,In_3,In_889);
xor U137 (N_137,In_60,In_820);
or U138 (N_138,In_511,In_832);
xnor U139 (N_139,In_18,In_912);
or U140 (N_140,In_600,In_923);
and U141 (N_141,In_471,In_869);
and U142 (N_142,In_112,In_943);
xor U143 (N_143,In_538,In_404);
nand U144 (N_144,In_118,In_586);
nand U145 (N_145,In_432,In_479);
and U146 (N_146,In_960,In_251);
or U147 (N_147,In_796,In_875);
and U148 (N_148,In_845,In_20);
nor U149 (N_149,In_651,In_147);
nand U150 (N_150,In_505,In_136);
xor U151 (N_151,In_227,In_622);
nand U152 (N_152,In_460,In_905);
xnor U153 (N_153,In_829,In_553);
xor U154 (N_154,In_549,In_961);
nand U155 (N_155,In_679,In_86);
and U156 (N_156,In_182,In_626);
xor U157 (N_157,In_167,In_192);
xnor U158 (N_158,In_621,In_185);
xnor U159 (N_159,In_202,In_56);
nand U160 (N_160,In_449,In_366);
xnor U161 (N_161,In_612,In_536);
xnor U162 (N_162,In_328,In_314);
xnor U163 (N_163,In_655,In_224);
or U164 (N_164,In_684,In_320);
or U165 (N_165,In_716,In_887);
nand U166 (N_166,In_358,In_524);
nor U167 (N_167,In_275,In_667);
xnor U168 (N_168,In_263,In_593);
and U169 (N_169,In_638,In_48);
xor U170 (N_170,In_919,In_427);
nand U171 (N_171,In_962,In_714);
or U172 (N_172,In_646,In_423);
and U173 (N_173,In_773,In_26);
nand U174 (N_174,In_910,In_641);
nor U175 (N_175,In_252,In_245);
and U176 (N_176,In_672,In_848);
and U177 (N_177,In_85,In_46);
nand U178 (N_178,In_417,In_98);
and U179 (N_179,In_203,In_283);
and U180 (N_180,In_52,In_73);
or U181 (N_181,In_67,In_886);
nor U182 (N_182,In_828,In_141);
and U183 (N_183,In_659,In_107);
nand U184 (N_184,In_114,In_827);
nor U185 (N_185,In_254,In_105);
nand U186 (N_186,In_437,In_948);
nand U187 (N_187,In_528,In_909);
nor U188 (N_188,In_126,In_121);
xnor U189 (N_189,In_556,In_871);
or U190 (N_190,In_403,In_732);
nand U191 (N_191,In_800,In_555);
and U192 (N_192,In_792,In_381);
and U193 (N_193,In_380,In_740);
nand U194 (N_194,In_37,In_30);
and U195 (N_195,In_9,In_652);
xor U196 (N_196,In_468,In_991);
nor U197 (N_197,In_194,In_451);
nor U198 (N_198,In_131,In_548);
or U199 (N_199,In_498,In_125);
nand U200 (N_200,N_95,In_973);
or U201 (N_201,In_430,N_42);
and U202 (N_202,In_325,In_847);
nor U203 (N_203,In_415,N_185);
xor U204 (N_204,In_574,In_564);
nand U205 (N_205,In_215,In_689);
nor U206 (N_206,In_682,N_92);
or U207 (N_207,In_22,In_193);
xor U208 (N_208,In_362,In_544);
xor U209 (N_209,In_250,N_189);
nor U210 (N_210,In_628,In_858);
and U211 (N_211,In_674,In_937);
nor U212 (N_212,N_51,In_990);
nand U213 (N_213,N_15,In_379);
xnor U214 (N_214,In_255,N_53);
xnor U215 (N_215,In_308,In_533);
xnor U216 (N_216,In_321,In_608);
nand U217 (N_217,In_113,In_264);
nor U218 (N_218,In_149,In_470);
nand U219 (N_219,N_49,In_546);
nor U220 (N_220,N_199,N_182);
nand U221 (N_221,N_3,In_616);
nor U222 (N_222,In_213,In_45);
nor U223 (N_223,In_518,In_726);
or U224 (N_224,In_552,In_270);
and U225 (N_225,In_285,In_474);
xor U226 (N_226,N_2,N_83);
nand U227 (N_227,In_770,In_597);
and U228 (N_228,In_881,In_96);
or U229 (N_229,In_128,In_302);
nand U230 (N_230,In_838,In_953);
xnor U231 (N_231,In_225,In_258);
nand U232 (N_232,N_160,N_75);
nand U233 (N_233,In_443,In_614);
nor U234 (N_234,In_287,In_775);
nand U235 (N_235,In_356,In_668);
nor U236 (N_236,In_711,In_210);
nor U237 (N_237,In_653,In_868);
xor U238 (N_238,N_113,N_134);
and U239 (N_239,In_606,In_562);
nor U240 (N_240,N_73,In_599);
and U241 (N_241,N_107,In_944);
nand U242 (N_242,In_452,In_150);
and U243 (N_243,N_180,In_666);
nand U244 (N_244,In_53,N_24);
nand U245 (N_245,In_680,In_839);
nand U246 (N_246,In_965,In_301);
and U247 (N_247,In_877,In_299);
or U248 (N_248,In_19,In_173);
nor U249 (N_249,In_34,In_70);
nand U250 (N_250,In_521,N_5);
nand U251 (N_251,N_71,In_291);
nor U252 (N_252,In_346,In_411);
nor U253 (N_253,In_87,In_69);
nand U254 (N_254,In_981,In_28);
nand U255 (N_255,N_89,In_949);
and U256 (N_256,In_130,N_150);
xnor U257 (N_257,In_139,N_123);
nor U258 (N_258,In_296,N_63);
nor U259 (N_259,In_987,In_604);
xor U260 (N_260,In_901,N_157);
or U261 (N_261,N_80,In_485);
nand U262 (N_262,In_110,In_801);
nor U263 (N_263,In_248,N_23);
or U264 (N_264,In_769,N_4);
nor U265 (N_265,In_989,In_433);
xnor U266 (N_266,In_578,In_710);
nor U267 (N_267,N_34,N_163);
xor U268 (N_268,In_135,In_294);
nand U269 (N_269,N_179,In_54);
xor U270 (N_270,In_932,In_234);
and U271 (N_271,In_794,In_476);
and U272 (N_272,In_457,In_535);
nand U273 (N_273,N_18,N_8);
nand U274 (N_274,N_28,In_349);
and U275 (N_275,N_40,In_77);
xor U276 (N_276,In_165,N_198);
xnor U277 (N_277,N_176,In_664);
nand U278 (N_278,In_883,N_84);
xnor U279 (N_279,In_530,N_25);
xor U280 (N_280,N_152,In_725);
nor U281 (N_281,N_41,In_632);
nand U282 (N_282,N_138,In_473);
xor U283 (N_283,In_893,N_132);
xnor U284 (N_284,In_879,In_539);
and U285 (N_285,N_170,In_465);
or U286 (N_286,N_70,N_22);
nand U287 (N_287,In_560,In_189);
nor U288 (N_288,In_872,In_755);
and U289 (N_289,N_60,In_29);
nand U290 (N_290,In_805,N_145);
and U291 (N_291,N_35,In_221);
or U292 (N_292,In_127,In_100);
nor U293 (N_293,In_611,N_135);
or U294 (N_294,N_79,In_787);
nor U295 (N_295,In_284,In_843);
and U296 (N_296,In_489,In_902);
nor U297 (N_297,In_715,N_76);
nor U298 (N_298,N_52,In_12);
nand U299 (N_299,N_20,In_341);
xnor U300 (N_300,N_57,In_279);
and U301 (N_301,N_21,N_78);
or U302 (N_302,In_863,In_691);
nor U303 (N_303,N_111,In_233);
nor U304 (N_304,In_453,In_581);
nand U305 (N_305,In_261,In_102);
or U306 (N_306,N_55,In_104);
nand U307 (N_307,In_24,In_831);
and U308 (N_308,In_392,N_9);
nand U309 (N_309,In_613,In_650);
xnor U310 (N_310,In_375,N_32);
xor U311 (N_311,N_47,In_945);
or U312 (N_312,In_116,In_873);
nand U313 (N_313,In_16,In_913);
and U314 (N_314,In_583,In_610);
or U315 (N_315,N_124,N_12);
and U316 (N_316,In_705,In_706);
xor U317 (N_317,In_601,In_840);
xor U318 (N_318,In_537,In_315);
and U319 (N_319,N_184,In_44);
or U320 (N_320,In_760,In_859);
nand U321 (N_321,N_64,In_146);
nand U322 (N_322,In_703,In_218);
nor U323 (N_323,In_334,In_230);
xor U324 (N_324,N_167,In_64);
or U325 (N_325,In_717,N_102);
and U326 (N_326,In_353,N_119);
nor U327 (N_327,In_171,In_76);
or U328 (N_328,In_854,In_635);
xnor U329 (N_329,In_607,In_180);
nand U330 (N_330,In_57,N_10);
xnor U331 (N_331,In_696,In_928);
nor U332 (N_332,In_813,In_676);
and U333 (N_333,In_648,In_993);
or U334 (N_334,In_700,N_117);
nand U335 (N_335,In_573,In_475);
or U336 (N_336,N_98,In_134);
nor U337 (N_337,In_804,In_497);
and U338 (N_338,In_92,N_99);
or U339 (N_339,N_1,In_577);
or U340 (N_340,N_105,N_48);
or U341 (N_341,In_469,In_772);
nor U342 (N_342,N_178,In_724);
nand U343 (N_343,In_741,In_852);
nand U344 (N_344,In_0,In_657);
or U345 (N_345,In_391,In_388);
xor U346 (N_346,N_122,In_154);
and U347 (N_347,In_502,In_997);
nor U348 (N_348,In_585,In_257);
or U349 (N_349,In_297,N_81);
and U350 (N_350,In_84,In_368);
nand U351 (N_351,N_130,N_149);
nor U352 (N_352,In_752,In_393);
nor U353 (N_353,In_117,In_629);
xnor U354 (N_354,In_445,In_447);
xor U355 (N_355,In_824,In_33);
and U356 (N_356,In_765,In_461);
nor U357 (N_357,N_6,In_983);
xor U358 (N_358,N_120,In_809);
and U359 (N_359,N_27,In_367);
or U360 (N_360,In_713,In_930);
nand U361 (N_361,In_851,N_31);
nand U362 (N_362,N_59,In_93);
nor U363 (N_363,In_351,In_342);
nand U364 (N_364,In_155,N_197);
and U365 (N_365,In_187,In_208);
nor U366 (N_366,N_114,N_118);
and U367 (N_367,In_178,In_217);
and U368 (N_368,N_103,N_65);
nand U369 (N_369,N_39,N_86);
nor U370 (N_370,In_802,In_159);
nand U371 (N_371,In_499,In_842);
or U372 (N_372,In_736,In_406);
nand U373 (N_373,In_688,In_554);
nor U374 (N_374,In_615,In_317);
and U375 (N_375,In_290,In_348);
xor U376 (N_376,N_194,In_623);
nand U377 (N_377,In_324,N_147);
and U378 (N_378,N_133,In_940);
nor U379 (N_379,In_557,N_116);
or U380 (N_380,In_702,In_888);
nor U381 (N_381,In_516,In_120);
nor U382 (N_382,N_154,N_126);
xor U383 (N_383,N_156,N_0);
and U384 (N_384,In_490,N_19);
nor U385 (N_385,In_238,In_157);
and U386 (N_386,In_409,In_172);
and U387 (N_387,In_634,In_145);
and U388 (N_388,In_390,N_85);
nor U389 (N_389,In_982,In_80);
nand U390 (N_390,In_496,In_115);
nand U391 (N_391,In_956,In_164);
or U392 (N_392,N_87,N_45);
nor U393 (N_393,In_750,In_924);
or U394 (N_394,In_739,In_276);
nand U395 (N_395,In_397,In_855);
nand U396 (N_396,In_378,In_491);
and U397 (N_397,In_239,N_74);
nor U398 (N_398,In_487,In_236);
nor U399 (N_399,In_211,N_166);
nand U400 (N_400,N_36,In_786);
nor U401 (N_401,In_429,N_273);
nand U402 (N_402,In_673,N_140);
xnor U403 (N_403,N_283,N_205);
or U404 (N_404,In_894,N_317);
or U405 (N_405,N_357,In_7);
and U406 (N_406,N_272,In_103);
or U407 (N_407,N_131,N_177);
nor U408 (N_408,N_327,N_293);
and U409 (N_409,In_822,N_262);
and U410 (N_410,In_265,N_322);
nor U411 (N_411,N_191,In_122);
nor U412 (N_412,N_175,N_223);
or U413 (N_413,In_137,In_976);
nor U414 (N_414,In_444,N_244);
xor U415 (N_415,N_13,In_82);
nor U416 (N_416,In_729,N_373);
xnor U417 (N_417,In_559,N_336);
nor U418 (N_418,N_255,In_821);
nor U419 (N_419,N_304,N_329);
xor U420 (N_420,In_32,N_286);
and U421 (N_421,N_210,N_266);
nor U422 (N_422,N_326,N_82);
nand U423 (N_423,In_222,N_356);
and U424 (N_424,N_50,N_338);
or U425 (N_425,In_333,In_620);
xnor U426 (N_426,In_816,In_382);
or U427 (N_427,N_234,N_246);
and U428 (N_428,N_67,In_229);
nand U429 (N_429,In_389,In_946);
and U430 (N_430,N_37,N_390);
and U431 (N_431,N_161,In_860);
xor U432 (N_432,In_844,N_69);
and U433 (N_433,In_835,N_324);
or U434 (N_434,In_778,N_248);
xnor U435 (N_435,N_112,In_58);
xor U436 (N_436,In_271,In_803);
or U437 (N_437,N_270,N_162);
xor U438 (N_438,In_738,In_719);
xnor U439 (N_439,N_249,In_269);
nand U440 (N_440,In_938,In_177);
nor U441 (N_441,In_293,N_305);
xor U442 (N_442,In_156,N_364);
or U443 (N_443,In_253,In_633);
and U444 (N_444,In_618,In_384);
and U445 (N_445,N_261,In_857);
or U446 (N_446,In_793,N_200);
or U447 (N_447,In_718,In_884);
nand U448 (N_448,N_44,In_590);
nand U449 (N_449,In_683,N_97);
or U450 (N_450,N_275,In_514);
nor U451 (N_451,N_33,N_106);
or U452 (N_452,In_169,In_918);
nor U453 (N_453,N_344,In_191);
or U454 (N_454,In_687,N_245);
or U455 (N_455,In_693,In_543);
nand U456 (N_456,In_757,N_104);
xnor U457 (N_457,N_362,In_61);
and U458 (N_458,N_220,In_780);
and U459 (N_459,N_88,In_31);
xnor U460 (N_460,In_463,N_377);
nor U461 (N_461,In_988,In_603);
nand U462 (N_462,In_168,N_386);
and U463 (N_463,In_994,In_571);
and U464 (N_464,N_168,In_219);
xnor U465 (N_465,N_351,N_314);
xor U466 (N_466,In_38,N_127);
nor U467 (N_467,In_458,N_54);
nand U468 (N_468,N_339,N_94);
or U469 (N_469,N_153,N_229);
xnor U470 (N_470,In_132,In_481);
nand U471 (N_471,N_396,In_17);
nor U472 (N_472,In_747,N_316);
xor U473 (N_473,In_428,In_550);
nand U474 (N_474,In_534,In_617);
nand U475 (N_475,In_727,N_312);
nand U476 (N_476,In_111,In_152);
or U477 (N_477,N_350,N_331);
xor U478 (N_478,In_295,In_767);
nand U479 (N_479,N_340,In_734);
xnor U480 (N_480,N_212,N_253);
nand U481 (N_481,In_488,N_165);
nand U482 (N_482,N_366,N_91);
or U483 (N_483,N_181,In_897);
nor U484 (N_484,N_379,In_723);
nand U485 (N_485,N_241,In_281);
nor U486 (N_486,N_195,In_273);
or U487 (N_487,In_978,N_142);
xor U488 (N_488,In_520,N_292);
and U489 (N_489,N_393,N_43);
and U490 (N_490,N_267,In_39);
or U491 (N_491,In_964,N_265);
xnor U492 (N_492,In_916,N_343);
or U493 (N_493,In_361,N_361);
or U494 (N_494,In_694,N_269);
or U495 (N_495,In_977,In_249);
nand U496 (N_496,In_442,N_230);
and U497 (N_497,N_321,N_298);
and U498 (N_498,N_371,In_849);
xnor U499 (N_499,N_375,N_17);
nor U500 (N_500,In_690,N_125);
and U501 (N_501,N_93,In_742);
or U502 (N_502,N_225,In_968);
nand U503 (N_503,In_166,In_41);
nor U504 (N_504,N_56,N_137);
nor U505 (N_505,In_966,In_568);
xnor U506 (N_506,N_66,In_231);
nand U507 (N_507,In_179,In_223);
xnor U508 (N_508,In_456,N_381);
and U509 (N_509,In_701,In_232);
and U510 (N_510,In_996,In_306);
or U511 (N_511,N_192,N_228);
xor U512 (N_512,N_345,In_605);
and U513 (N_513,N_100,In_446);
or U514 (N_514,In_405,In_861);
and U515 (N_515,N_395,N_346);
nor U516 (N_516,N_258,In_517);
nand U517 (N_517,In_129,N_313);
or U518 (N_518,In_42,N_164);
xnor U519 (N_519,N_257,In_619);
or U520 (N_520,In_424,In_731);
and U521 (N_521,In_589,N_146);
and U522 (N_522,N_202,In_478);
nand U523 (N_523,In_322,N_334);
and U524 (N_524,In_186,In_25);
nand U525 (N_525,N_303,In_400);
or U526 (N_526,In_526,In_959);
nor U527 (N_527,In_565,N_29);
nor U528 (N_528,In_101,N_151);
nand U529 (N_529,N_369,In_331);
xnor U530 (N_530,N_264,In_59);
xor U531 (N_531,In_242,N_193);
or U532 (N_532,In_833,N_239);
nor U533 (N_533,N_333,In_856);
or U534 (N_534,N_306,In_209);
nor U535 (N_535,In_2,In_4);
nand U536 (N_536,In_797,N_310);
or U537 (N_537,N_284,N_235);
and U538 (N_538,N_358,N_206);
nor U539 (N_539,N_354,In_656);
nand U540 (N_540,N_378,In_174);
nand U541 (N_541,N_335,In_15);
nand U542 (N_542,In_418,In_878);
and U543 (N_543,In_196,In_65);
and U544 (N_544,N_288,N_121);
or U545 (N_545,N_308,N_171);
xnor U546 (N_546,N_388,N_46);
xnor U547 (N_547,In_204,In_318);
nand U548 (N_548,N_325,In_106);
nor U549 (N_549,N_300,In_709);
or U550 (N_550,In_876,In_435);
xor U551 (N_551,In_142,In_764);
or U552 (N_552,N_311,N_77);
nor U553 (N_553,In_198,N_204);
or U554 (N_554,In_448,In_190);
or U555 (N_555,N_224,In_501);
and U556 (N_556,In_220,N_183);
nor U557 (N_557,In_942,In_984);
nor U558 (N_558,N_216,N_238);
nor U559 (N_559,N_360,N_309);
nand U560 (N_560,N_348,N_332);
nand U561 (N_561,N_211,In_83);
xor U562 (N_562,In_675,N_172);
or U563 (N_563,In_834,In_746);
xor U564 (N_564,N_277,N_190);
and U565 (N_565,N_382,N_318);
or U566 (N_566,In_419,In_572);
xnor U567 (N_567,In_525,In_864);
nor U568 (N_568,In_915,In_891);
nor U569 (N_569,N_222,N_374);
xnor U570 (N_570,In_642,In_591);
and U571 (N_571,N_256,N_233);
and U572 (N_572,In_712,N_218);
nand U573 (N_573,In_749,In_625);
xnor U574 (N_574,N_330,N_363);
nand U575 (N_575,N_368,N_282);
or U576 (N_576,N_278,In_758);
and U577 (N_577,N_353,In_503);
or U578 (N_578,In_671,In_319);
or U579 (N_579,N_144,In_343);
xor U580 (N_580,In_522,In_466);
nand U581 (N_581,In_438,In_247);
xor U582 (N_582,In_36,In_532);
or U583 (N_583,In_512,N_389);
nor U584 (N_584,N_250,N_294);
xnor U585 (N_585,In_421,In_304);
xnor U586 (N_586,In_823,N_7);
or U587 (N_587,N_274,N_342);
nand U588 (N_588,N_271,N_268);
and U589 (N_589,N_217,N_207);
and U590 (N_590,N_139,N_260);
and U591 (N_591,In_841,N_196);
or U592 (N_592,In_698,N_61);
or U593 (N_593,N_108,In_357);
and U594 (N_594,In_148,In_921);
and U595 (N_595,In_903,In_298);
nor U596 (N_596,N_380,N_188);
or U597 (N_597,N_319,In_416);
and U598 (N_598,N_68,In_300);
and U599 (N_599,N_352,In_998);
nor U600 (N_600,In_340,N_129);
xnor U601 (N_601,In_160,N_397);
nor U602 (N_602,N_444,N_553);
nand U603 (N_603,N_451,N_297);
nor U604 (N_604,N_480,N_280);
or U605 (N_605,N_291,N_489);
or U606 (N_606,N_315,N_428);
nand U607 (N_607,In_733,In_350);
xnor U608 (N_608,N_497,In_23);
and U609 (N_609,In_459,N_506);
and U610 (N_610,N_158,In_90);
and U611 (N_611,N_526,N_96);
nand U612 (N_612,N_221,N_495);
and U613 (N_613,N_472,In_480);
or U614 (N_614,In_207,In_310);
xnor U615 (N_615,N_337,N_458);
nor U616 (N_616,In_637,N_551);
and U617 (N_617,N_599,N_493);
or U618 (N_618,N_488,N_565);
and U619 (N_619,N_413,N_473);
nand U620 (N_620,In_515,In_654);
or U621 (N_621,N_450,N_541);
nor U622 (N_622,N_571,N_301);
nor U623 (N_623,N_62,N_550);
xor U624 (N_624,N_383,N_583);
nor U625 (N_625,N_355,In_882);
or U626 (N_626,In_109,N_446);
xnor U627 (N_627,N_14,N_285);
xor U628 (N_628,In_846,N_400);
nor U629 (N_629,N_498,N_136);
nor U630 (N_630,In_896,N_543);
or U631 (N_631,N_209,In_436);
and U632 (N_632,In_68,N_510);
or U633 (N_633,In_369,N_432);
xnor U634 (N_634,In_95,N_401);
nand U635 (N_635,N_307,In_6);
nor U636 (N_636,In_643,N_569);
nand U637 (N_637,N_479,N_579);
nor U638 (N_638,In_790,In_373);
nand U639 (N_639,In_143,N_592);
or U640 (N_640,N_582,N_567);
nand U641 (N_641,N_213,N_540);
xor U642 (N_642,In_50,N_449);
nand U643 (N_643,N_110,In_175);
or U644 (N_644,In_311,In_540);
or U645 (N_645,In_40,N_546);
nor U646 (N_646,N_232,N_148);
xnor U647 (N_647,N_555,In_922);
or U648 (N_648,N_482,N_16);
nand U649 (N_649,N_394,N_290);
or U650 (N_650,N_445,N_527);
or U651 (N_651,N_584,N_387);
nor U652 (N_652,N_219,N_243);
nand U653 (N_653,N_538,N_585);
or U654 (N_654,N_578,N_418);
nand U655 (N_655,N_591,In_228);
nor U656 (N_656,N_548,N_143);
or U657 (N_657,N_507,N_514);
nand U658 (N_658,N_468,N_58);
nand U659 (N_659,N_545,In_241);
nor U660 (N_660,N_399,N_328);
nand U661 (N_661,N_38,N_226);
or U662 (N_662,In_1,N_347);
or U663 (N_663,In_782,In_662);
or U664 (N_664,N_486,In_235);
and U665 (N_665,N_431,N_452);
or U666 (N_666,N_470,N_577);
and U667 (N_667,In_262,In_957);
and U668 (N_668,In_551,N_558);
or U669 (N_669,N_483,In_636);
and U670 (N_670,N_423,In_811);
or U671 (N_671,N_173,N_242);
nor U672 (N_672,In_986,N_586);
and U673 (N_673,N_559,N_438);
and U674 (N_674,In_268,In_917);
or U675 (N_675,N_518,N_574);
xnor U676 (N_676,N_414,N_484);
and U677 (N_677,N_570,In_967);
nand U678 (N_678,N_478,N_251);
nand U679 (N_679,N_494,In_880);
and U680 (N_680,N_508,N_159);
and U681 (N_681,N_323,N_560);
and U682 (N_682,N_513,N_115);
or U683 (N_683,N_422,N_461);
xnor U684 (N_684,N_512,N_341);
xor U685 (N_685,N_441,N_392);
nand U686 (N_686,N_215,N_491);
nor U687 (N_687,N_534,In_566);
and U688 (N_688,N_365,N_406);
nand U689 (N_689,N_421,N_552);
nor U690 (N_690,N_572,N_522);
xnor U691 (N_691,N_227,In_455);
xnor U692 (N_692,N_367,N_240);
nand U693 (N_693,N_516,N_174);
or U694 (N_694,N_463,N_403);
nand U695 (N_695,N_155,In_62);
xnor U696 (N_696,N_128,In_783);
nand U697 (N_697,N_503,N_504);
nor U698 (N_698,N_520,In_561);
nor U699 (N_699,N_30,N_169);
nor U700 (N_700,In_911,N_448);
and U701 (N_701,N_459,In_402);
or U702 (N_702,In_649,N_420);
and U703 (N_703,N_443,In_862);
and U704 (N_704,N_402,In_81);
nor U705 (N_705,N_425,In_313);
or U706 (N_706,N_434,N_384);
or U707 (N_707,N_295,N_568);
and U708 (N_708,N_237,N_433);
or U709 (N_709,N_440,N_528);
xnor U710 (N_710,N_524,In_188);
xor U711 (N_711,N_519,N_517);
nand U712 (N_712,N_281,N_372);
or U713 (N_713,In_927,N_385);
nand U714 (N_714,In_280,N_593);
nor U715 (N_715,N_536,N_462);
or U716 (N_716,N_455,N_515);
nor U717 (N_717,In_181,N_410);
nand U718 (N_718,N_587,In_584);
nor U719 (N_719,N_466,N_496);
or U720 (N_720,In_244,N_460);
or U721 (N_721,N_287,N_561);
nor U722 (N_722,N_557,In_398);
or U723 (N_723,N_535,In_355);
nor U724 (N_724,In_5,N_487);
or U725 (N_725,N_581,N_547);
xnor U726 (N_726,N_259,N_407);
nor U727 (N_727,N_415,N_302);
xor U728 (N_728,N_236,N_456);
xnor U729 (N_729,In_482,N_511);
and U730 (N_730,N_475,In_47);
nor U731 (N_731,In_289,N_404);
xnor U732 (N_732,In_138,N_26);
and U733 (N_733,In_199,N_398);
or U734 (N_734,N_549,N_201);
xnor U735 (N_735,N_454,N_598);
or U736 (N_736,N_109,N_469);
nand U737 (N_737,N_539,N_501);
xnor U738 (N_738,N_186,N_72);
and U739 (N_739,N_525,N_474);
xnor U740 (N_740,N_521,N_101);
nor U741 (N_741,In_686,N_203);
nor U742 (N_742,N_376,In_699);
or U743 (N_743,N_476,In_837);
nor U744 (N_744,N_263,N_437);
and U745 (N_745,N_537,N_533);
or U746 (N_746,N_416,N_542);
xor U747 (N_747,N_187,In_197);
or U748 (N_748,N_435,In_467);
and U749 (N_749,N_573,In_756);
or U750 (N_750,N_439,N_349);
and U751 (N_751,In_329,N_417);
nand U752 (N_752,In_830,N_141);
xnor U753 (N_753,N_477,In_974);
xor U754 (N_754,N_453,N_566);
or U755 (N_755,N_530,In_21);
xnor U756 (N_756,N_502,N_485);
xnor U757 (N_757,N_464,N_481);
nor U758 (N_758,N_231,N_424);
and U759 (N_759,N_247,In_771);
and U760 (N_760,N_505,In_286);
xnor U761 (N_761,N_252,N_457);
xor U762 (N_762,In_413,N_597);
xor U763 (N_763,N_411,N_465);
xnor U764 (N_764,N_499,N_289);
nand U765 (N_765,N_563,N_429);
xor U766 (N_766,N_588,N_430);
xor U767 (N_767,N_580,N_447);
nand U768 (N_768,N_419,N_442);
or U769 (N_769,N_509,In_744);
xnor U770 (N_770,In_941,In_507);
nand U771 (N_771,In_292,N_500);
nand U772 (N_772,N_595,N_436);
nand U773 (N_773,N_299,N_589);
or U774 (N_774,N_427,In_8);
nor U775 (N_775,In_759,N_214);
or U776 (N_776,N_11,N_467);
nand U777 (N_777,N_562,N_391);
nand U778 (N_778,In_929,In_162);
and U779 (N_779,In_454,In_567);
nand U780 (N_780,In_14,N_370);
nor U781 (N_781,N_208,In_721);
or U782 (N_782,N_492,In_545);
nand U783 (N_783,N_409,N_320);
nor U784 (N_784,N_529,N_490);
nand U785 (N_785,N_296,In_43);
nand U786 (N_786,N_564,N_576);
or U787 (N_787,N_523,N_531);
and U788 (N_788,In_661,N_575);
nor U789 (N_789,N_544,N_426);
xnor U790 (N_790,N_408,N_405);
nand U791 (N_791,N_594,N_532);
nor U792 (N_792,In_588,N_590);
nor U793 (N_793,In_678,N_412);
xnor U794 (N_794,N_596,N_554);
xor U795 (N_795,N_556,In_708);
xor U796 (N_796,N_279,N_359);
or U797 (N_797,In_763,N_276);
xnor U798 (N_798,N_471,N_90);
and U799 (N_799,In_201,N_254);
xnor U800 (N_800,N_615,N_651);
or U801 (N_801,N_756,N_650);
nand U802 (N_802,N_764,N_772);
nand U803 (N_803,N_728,N_675);
xnor U804 (N_804,N_660,N_681);
and U805 (N_805,N_750,N_731);
nor U806 (N_806,N_741,N_623);
nand U807 (N_807,N_722,N_672);
xor U808 (N_808,N_739,N_685);
nor U809 (N_809,N_788,N_669);
nor U810 (N_810,N_676,N_605);
or U811 (N_811,N_686,N_677);
or U812 (N_812,N_698,N_704);
and U813 (N_813,N_618,N_687);
or U814 (N_814,N_769,N_740);
or U815 (N_815,N_743,N_600);
or U816 (N_816,N_707,N_665);
or U817 (N_817,N_785,N_789);
nor U818 (N_818,N_748,N_620);
xnor U819 (N_819,N_710,N_774);
nand U820 (N_820,N_631,N_648);
and U821 (N_821,N_634,N_638);
nand U822 (N_822,N_683,N_787);
xnor U823 (N_823,N_642,N_610);
nand U824 (N_824,N_694,N_799);
nor U825 (N_825,N_747,N_689);
xnor U826 (N_826,N_757,N_752);
or U827 (N_827,N_790,N_652);
and U828 (N_828,N_655,N_705);
and U829 (N_829,N_716,N_626);
xnor U830 (N_830,N_663,N_637);
xnor U831 (N_831,N_745,N_732);
xnor U832 (N_832,N_627,N_635);
xnor U833 (N_833,N_649,N_770);
or U834 (N_834,N_733,N_612);
or U835 (N_835,N_622,N_690);
and U836 (N_836,N_718,N_738);
xnor U837 (N_837,N_670,N_727);
nand U838 (N_838,N_614,N_751);
nor U839 (N_839,N_673,N_749);
xor U840 (N_840,N_761,N_656);
nand U841 (N_841,N_674,N_645);
and U842 (N_842,N_602,N_702);
and U843 (N_843,N_763,N_601);
or U844 (N_844,N_606,N_712);
nand U845 (N_845,N_619,N_767);
nand U846 (N_846,N_793,N_742);
nand U847 (N_847,N_782,N_682);
and U848 (N_848,N_736,N_717);
xor U849 (N_849,N_695,N_706);
xor U850 (N_850,N_617,N_697);
and U851 (N_851,N_709,N_730);
nor U852 (N_852,N_778,N_791);
nand U853 (N_853,N_781,N_758);
nand U854 (N_854,N_629,N_678);
and U855 (N_855,N_680,N_762);
xnor U856 (N_856,N_714,N_766);
xor U857 (N_857,N_688,N_644);
nand U858 (N_858,N_625,N_621);
and U859 (N_859,N_724,N_607);
or U860 (N_860,N_628,N_630);
nor U861 (N_861,N_720,N_658);
nand U862 (N_862,N_613,N_603);
xnor U863 (N_863,N_735,N_792);
nand U864 (N_864,N_616,N_693);
nor U865 (N_865,N_771,N_783);
and U866 (N_866,N_715,N_759);
or U867 (N_867,N_633,N_608);
and U868 (N_868,N_624,N_657);
and U869 (N_869,N_796,N_713);
xor U870 (N_870,N_641,N_725);
or U871 (N_871,N_640,N_780);
xor U872 (N_872,N_646,N_737);
or U873 (N_873,N_773,N_662);
xnor U874 (N_874,N_684,N_696);
or U875 (N_875,N_755,N_643);
or U876 (N_876,N_779,N_711);
nand U877 (N_877,N_671,N_719);
nand U878 (N_878,N_632,N_786);
and U879 (N_879,N_667,N_726);
nor U880 (N_880,N_775,N_691);
nand U881 (N_881,N_794,N_760);
or U882 (N_882,N_765,N_744);
nand U883 (N_883,N_679,N_708);
xnor U884 (N_884,N_664,N_703);
xnor U885 (N_885,N_639,N_699);
nand U886 (N_886,N_795,N_701);
xor U887 (N_887,N_797,N_700);
nand U888 (N_888,N_661,N_668);
xor U889 (N_889,N_768,N_721);
nor U890 (N_890,N_776,N_729);
or U891 (N_891,N_798,N_609);
nand U892 (N_892,N_666,N_746);
xor U893 (N_893,N_647,N_604);
and U894 (N_894,N_734,N_611);
nand U895 (N_895,N_784,N_692);
and U896 (N_896,N_636,N_723);
nand U897 (N_897,N_753,N_777);
nand U898 (N_898,N_754,N_654);
and U899 (N_899,N_659,N_653);
xor U900 (N_900,N_672,N_766);
nor U901 (N_901,N_756,N_703);
and U902 (N_902,N_649,N_793);
or U903 (N_903,N_736,N_786);
nor U904 (N_904,N_686,N_664);
nor U905 (N_905,N_658,N_647);
nand U906 (N_906,N_719,N_723);
or U907 (N_907,N_718,N_600);
nor U908 (N_908,N_613,N_617);
nand U909 (N_909,N_769,N_794);
and U910 (N_910,N_787,N_755);
and U911 (N_911,N_651,N_669);
nor U912 (N_912,N_668,N_798);
nand U913 (N_913,N_718,N_766);
and U914 (N_914,N_753,N_754);
or U915 (N_915,N_736,N_749);
or U916 (N_916,N_788,N_786);
or U917 (N_917,N_631,N_601);
and U918 (N_918,N_790,N_646);
nand U919 (N_919,N_627,N_659);
xor U920 (N_920,N_651,N_677);
or U921 (N_921,N_641,N_674);
nor U922 (N_922,N_696,N_708);
nor U923 (N_923,N_652,N_695);
or U924 (N_924,N_724,N_774);
and U925 (N_925,N_644,N_620);
xnor U926 (N_926,N_732,N_644);
nor U927 (N_927,N_609,N_787);
and U928 (N_928,N_693,N_725);
and U929 (N_929,N_732,N_695);
nand U930 (N_930,N_708,N_785);
or U931 (N_931,N_747,N_600);
nor U932 (N_932,N_647,N_761);
or U933 (N_933,N_777,N_652);
nand U934 (N_934,N_721,N_690);
and U935 (N_935,N_761,N_643);
nand U936 (N_936,N_786,N_757);
and U937 (N_937,N_652,N_680);
or U938 (N_938,N_647,N_733);
xnor U939 (N_939,N_749,N_773);
and U940 (N_940,N_602,N_669);
or U941 (N_941,N_683,N_700);
and U942 (N_942,N_612,N_646);
or U943 (N_943,N_675,N_620);
and U944 (N_944,N_668,N_677);
or U945 (N_945,N_622,N_605);
and U946 (N_946,N_645,N_683);
xor U947 (N_947,N_664,N_741);
nor U948 (N_948,N_646,N_721);
or U949 (N_949,N_682,N_616);
and U950 (N_950,N_756,N_723);
xnor U951 (N_951,N_687,N_741);
xnor U952 (N_952,N_661,N_680);
or U953 (N_953,N_642,N_627);
nor U954 (N_954,N_725,N_755);
nor U955 (N_955,N_786,N_707);
nor U956 (N_956,N_613,N_760);
or U957 (N_957,N_677,N_796);
nand U958 (N_958,N_744,N_712);
nand U959 (N_959,N_670,N_750);
nand U960 (N_960,N_695,N_694);
and U961 (N_961,N_771,N_799);
and U962 (N_962,N_607,N_720);
and U963 (N_963,N_637,N_755);
xor U964 (N_964,N_624,N_718);
and U965 (N_965,N_634,N_684);
nand U966 (N_966,N_619,N_620);
nor U967 (N_967,N_741,N_681);
xor U968 (N_968,N_613,N_639);
nor U969 (N_969,N_725,N_738);
xnor U970 (N_970,N_766,N_757);
xnor U971 (N_971,N_601,N_771);
nor U972 (N_972,N_640,N_797);
xor U973 (N_973,N_621,N_658);
or U974 (N_974,N_781,N_650);
nand U975 (N_975,N_773,N_729);
or U976 (N_976,N_709,N_636);
nor U977 (N_977,N_737,N_666);
nand U978 (N_978,N_772,N_605);
nand U979 (N_979,N_688,N_759);
or U980 (N_980,N_722,N_795);
and U981 (N_981,N_797,N_722);
and U982 (N_982,N_659,N_797);
or U983 (N_983,N_714,N_660);
or U984 (N_984,N_612,N_759);
and U985 (N_985,N_737,N_701);
or U986 (N_986,N_692,N_670);
nor U987 (N_987,N_794,N_765);
nand U988 (N_988,N_765,N_672);
or U989 (N_989,N_789,N_702);
nand U990 (N_990,N_631,N_779);
nand U991 (N_991,N_626,N_641);
or U992 (N_992,N_645,N_601);
nand U993 (N_993,N_733,N_625);
or U994 (N_994,N_791,N_681);
nand U995 (N_995,N_648,N_776);
nand U996 (N_996,N_672,N_756);
or U997 (N_997,N_798,N_610);
or U998 (N_998,N_613,N_662);
nor U999 (N_999,N_716,N_672);
nor U1000 (N_1000,N_861,N_954);
xnor U1001 (N_1001,N_947,N_935);
or U1002 (N_1002,N_996,N_851);
nand U1003 (N_1003,N_847,N_856);
and U1004 (N_1004,N_900,N_911);
xnor U1005 (N_1005,N_960,N_898);
and U1006 (N_1006,N_916,N_872);
xor U1007 (N_1007,N_836,N_945);
or U1008 (N_1008,N_992,N_824);
nand U1009 (N_1009,N_814,N_907);
xor U1010 (N_1010,N_942,N_949);
nand U1011 (N_1011,N_906,N_970);
and U1012 (N_1012,N_983,N_905);
xnor U1013 (N_1013,N_815,N_967);
or U1014 (N_1014,N_821,N_839);
nor U1015 (N_1015,N_908,N_976);
xnor U1016 (N_1016,N_914,N_820);
or U1017 (N_1017,N_936,N_832);
or U1018 (N_1018,N_912,N_998);
nand U1019 (N_1019,N_931,N_854);
xor U1020 (N_1020,N_822,N_893);
nor U1021 (N_1021,N_875,N_878);
or U1022 (N_1022,N_818,N_962);
or U1023 (N_1023,N_895,N_807);
nor U1024 (N_1024,N_899,N_830);
xor U1025 (N_1025,N_800,N_950);
and U1026 (N_1026,N_913,N_987);
xnor U1027 (N_1027,N_886,N_981);
or U1028 (N_1028,N_866,N_903);
xnor U1029 (N_1029,N_940,N_871);
nand U1030 (N_1030,N_964,N_852);
or U1031 (N_1031,N_892,N_829);
and U1032 (N_1032,N_953,N_811);
xor U1033 (N_1033,N_986,N_877);
nor U1034 (N_1034,N_926,N_923);
nor U1035 (N_1035,N_833,N_834);
nor U1036 (N_1036,N_828,N_928);
xnor U1037 (N_1037,N_890,N_885);
xnor U1038 (N_1038,N_805,N_946);
and U1039 (N_1039,N_952,N_816);
and U1040 (N_1040,N_819,N_944);
nand U1041 (N_1041,N_880,N_846);
nand U1042 (N_1042,N_802,N_867);
and U1043 (N_1043,N_922,N_969);
xor U1044 (N_1044,N_984,N_997);
nand U1045 (N_1045,N_989,N_827);
nand U1046 (N_1046,N_844,N_803);
nand U1047 (N_1047,N_873,N_904);
nand U1048 (N_1048,N_897,N_990);
nor U1049 (N_1049,N_881,N_848);
or U1050 (N_1050,N_993,N_838);
nor U1051 (N_1051,N_974,N_801);
or U1052 (N_1052,N_850,N_980);
or U1053 (N_1053,N_939,N_902);
or U1054 (N_1054,N_894,N_868);
xnor U1055 (N_1055,N_841,N_973);
nand U1056 (N_1056,N_963,N_959);
nor U1057 (N_1057,N_910,N_994);
and U1058 (N_1058,N_978,N_977);
or U1059 (N_1059,N_930,N_991);
or U1060 (N_1060,N_941,N_859);
nand U1061 (N_1061,N_896,N_917);
nor U1062 (N_1062,N_937,N_876);
or U1063 (N_1063,N_812,N_882);
nor U1064 (N_1064,N_862,N_938);
xor U1065 (N_1065,N_849,N_813);
xnor U1066 (N_1066,N_835,N_879);
or U1067 (N_1067,N_810,N_888);
nor U1068 (N_1068,N_891,N_804);
and U1069 (N_1069,N_837,N_918);
nor U1070 (N_1070,N_808,N_982);
nand U1071 (N_1071,N_975,N_934);
nand U1072 (N_1072,N_979,N_853);
or U1073 (N_1073,N_831,N_965);
xor U1074 (N_1074,N_921,N_925);
or U1075 (N_1075,N_948,N_855);
or U1076 (N_1076,N_889,N_865);
nand U1077 (N_1077,N_927,N_809);
nor U1078 (N_1078,N_901,N_863);
nand U1079 (N_1079,N_870,N_966);
nand U1080 (N_1080,N_806,N_817);
nor U1081 (N_1081,N_845,N_929);
or U1082 (N_1082,N_972,N_864);
or U1083 (N_1083,N_924,N_826);
and U1084 (N_1084,N_857,N_909);
and U1085 (N_1085,N_956,N_843);
nand U1086 (N_1086,N_825,N_957);
xor U1087 (N_1087,N_883,N_919);
or U1088 (N_1088,N_823,N_932);
xor U1089 (N_1089,N_869,N_955);
and U1090 (N_1090,N_915,N_858);
nand U1091 (N_1091,N_968,N_999);
and U1092 (N_1092,N_943,N_933);
nand U1093 (N_1093,N_988,N_958);
nand U1094 (N_1094,N_884,N_840);
or U1095 (N_1095,N_874,N_887);
nand U1096 (N_1096,N_951,N_971);
nor U1097 (N_1097,N_860,N_920);
xor U1098 (N_1098,N_985,N_995);
nor U1099 (N_1099,N_961,N_842);
or U1100 (N_1100,N_926,N_837);
or U1101 (N_1101,N_989,N_801);
and U1102 (N_1102,N_959,N_896);
or U1103 (N_1103,N_946,N_907);
xor U1104 (N_1104,N_973,N_871);
xnor U1105 (N_1105,N_908,N_964);
xor U1106 (N_1106,N_939,N_852);
xor U1107 (N_1107,N_834,N_967);
xor U1108 (N_1108,N_817,N_971);
nor U1109 (N_1109,N_983,N_841);
nor U1110 (N_1110,N_931,N_858);
nand U1111 (N_1111,N_886,N_957);
nand U1112 (N_1112,N_837,N_943);
nand U1113 (N_1113,N_893,N_990);
nor U1114 (N_1114,N_983,N_847);
nor U1115 (N_1115,N_811,N_976);
nor U1116 (N_1116,N_891,N_964);
xnor U1117 (N_1117,N_820,N_867);
xor U1118 (N_1118,N_904,N_870);
nand U1119 (N_1119,N_923,N_800);
and U1120 (N_1120,N_949,N_847);
and U1121 (N_1121,N_831,N_918);
nand U1122 (N_1122,N_986,N_961);
xor U1123 (N_1123,N_899,N_832);
or U1124 (N_1124,N_932,N_945);
xor U1125 (N_1125,N_883,N_822);
xor U1126 (N_1126,N_828,N_941);
xnor U1127 (N_1127,N_824,N_867);
nand U1128 (N_1128,N_920,N_809);
nor U1129 (N_1129,N_810,N_927);
xor U1130 (N_1130,N_956,N_995);
and U1131 (N_1131,N_804,N_926);
and U1132 (N_1132,N_898,N_867);
or U1133 (N_1133,N_892,N_964);
nand U1134 (N_1134,N_925,N_868);
or U1135 (N_1135,N_948,N_866);
and U1136 (N_1136,N_971,N_886);
xnor U1137 (N_1137,N_947,N_809);
or U1138 (N_1138,N_953,N_822);
nor U1139 (N_1139,N_942,N_977);
nand U1140 (N_1140,N_972,N_842);
or U1141 (N_1141,N_880,N_819);
xnor U1142 (N_1142,N_858,N_933);
or U1143 (N_1143,N_924,N_926);
or U1144 (N_1144,N_907,N_929);
and U1145 (N_1145,N_973,N_923);
or U1146 (N_1146,N_975,N_994);
and U1147 (N_1147,N_840,N_864);
xor U1148 (N_1148,N_951,N_867);
and U1149 (N_1149,N_810,N_997);
and U1150 (N_1150,N_822,N_986);
nand U1151 (N_1151,N_845,N_850);
nor U1152 (N_1152,N_971,N_890);
nor U1153 (N_1153,N_812,N_904);
or U1154 (N_1154,N_824,N_990);
nand U1155 (N_1155,N_803,N_863);
or U1156 (N_1156,N_864,N_956);
or U1157 (N_1157,N_859,N_825);
nor U1158 (N_1158,N_825,N_853);
nor U1159 (N_1159,N_989,N_926);
xor U1160 (N_1160,N_853,N_945);
nand U1161 (N_1161,N_808,N_810);
xor U1162 (N_1162,N_808,N_888);
xnor U1163 (N_1163,N_834,N_897);
and U1164 (N_1164,N_975,N_866);
nor U1165 (N_1165,N_886,N_906);
or U1166 (N_1166,N_958,N_951);
nor U1167 (N_1167,N_837,N_802);
xnor U1168 (N_1168,N_980,N_935);
or U1169 (N_1169,N_942,N_855);
and U1170 (N_1170,N_860,N_847);
nand U1171 (N_1171,N_942,N_921);
nor U1172 (N_1172,N_820,N_864);
and U1173 (N_1173,N_920,N_894);
nor U1174 (N_1174,N_987,N_819);
nand U1175 (N_1175,N_834,N_974);
and U1176 (N_1176,N_974,N_975);
and U1177 (N_1177,N_966,N_812);
xor U1178 (N_1178,N_844,N_985);
xnor U1179 (N_1179,N_838,N_885);
nor U1180 (N_1180,N_820,N_940);
nor U1181 (N_1181,N_904,N_938);
nor U1182 (N_1182,N_994,N_942);
xor U1183 (N_1183,N_850,N_807);
xnor U1184 (N_1184,N_834,N_839);
and U1185 (N_1185,N_965,N_829);
nand U1186 (N_1186,N_907,N_950);
nand U1187 (N_1187,N_817,N_946);
nand U1188 (N_1188,N_995,N_849);
or U1189 (N_1189,N_968,N_947);
and U1190 (N_1190,N_922,N_879);
xnor U1191 (N_1191,N_860,N_816);
xnor U1192 (N_1192,N_898,N_984);
nand U1193 (N_1193,N_838,N_908);
or U1194 (N_1194,N_998,N_856);
nor U1195 (N_1195,N_883,N_860);
nand U1196 (N_1196,N_934,N_973);
xnor U1197 (N_1197,N_993,N_803);
and U1198 (N_1198,N_890,N_824);
nand U1199 (N_1199,N_897,N_995);
or U1200 (N_1200,N_1037,N_1079);
xnor U1201 (N_1201,N_1194,N_1035);
nor U1202 (N_1202,N_1113,N_1030);
or U1203 (N_1203,N_1098,N_1123);
nor U1204 (N_1204,N_1154,N_1043);
or U1205 (N_1205,N_1017,N_1041);
nand U1206 (N_1206,N_1054,N_1001);
and U1207 (N_1207,N_1197,N_1146);
nor U1208 (N_1208,N_1062,N_1010);
and U1209 (N_1209,N_1080,N_1163);
or U1210 (N_1210,N_1169,N_1187);
xor U1211 (N_1211,N_1150,N_1122);
nor U1212 (N_1212,N_1024,N_1021);
xnor U1213 (N_1213,N_1152,N_1031);
xnor U1214 (N_1214,N_1020,N_1053);
nand U1215 (N_1215,N_1137,N_1044);
xnor U1216 (N_1216,N_1107,N_1090);
or U1217 (N_1217,N_1072,N_1014);
nand U1218 (N_1218,N_1160,N_1029);
nor U1219 (N_1219,N_1015,N_1129);
and U1220 (N_1220,N_1130,N_1166);
nor U1221 (N_1221,N_1089,N_1140);
nand U1222 (N_1222,N_1019,N_1084);
xor U1223 (N_1223,N_1048,N_1064);
xor U1224 (N_1224,N_1077,N_1082);
or U1225 (N_1225,N_1003,N_1094);
nand U1226 (N_1226,N_1157,N_1008);
nand U1227 (N_1227,N_1110,N_1022);
or U1228 (N_1228,N_1143,N_1078);
xor U1229 (N_1229,N_1056,N_1153);
nand U1230 (N_1230,N_1161,N_1081);
xor U1231 (N_1231,N_1092,N_1033);
and U1232 (N_1232,N_1145,N_1174);
or U1233 (N_1233,N_1005,N_1059);
nand U1234 (N_1234,N_1147,N_1112);
nor U1235 (N_1235,N_1032,N_1095);
nor U1236 (N_1236,N_1004,N_1002);
xnor U1237 (N_1237,N_1135,N_1100);
nand U1238 (N_1238,N_1189,N_1007);
nor U1239 (N_1239,N_1118,N_1139);
or U1240 (N_1240,N_1119,N_1061);
and U1241 (N_1241,N_1088,N_1047);
xnor U1242 (N_1242,N_1184,N_1182);
nor U1243 (N_1243,N_1192,N_1038);
xor U1244 (N_1244,N_1199,N_1124);
nand U1245 (N_1245,N_1051,N_1013);
nand U1246 (N_1246,N_1085,N_1126);
xnor U1247 (N_1247,N_1173,N_1067);
xnor U1248 (N_1248,N_1065,N_1068);
xor U1249 (N_1249,N_1018,N_1138);
and U1250 (N_1250,N_1128,N_1193);
or U1251 (N_1251,N_1009,N_1191);
and U1252 (N_1252,N_1083,N_1093);
nand U1253 (N_1253,N_1060,N_1023);
nand U1254 (N_1254,N_1097,N_1196);
nand U1255 (N_1255,N_1141,N_1116);
nand U1256 (N_1256,N_1016,N_1034);
xnor U1257 (N_1257,N_1120,N_1149);
or U1258 (N_1258,N_1000,N_1050);
or U1259 (N_1259,N_1167,N_1087);
xnor U1260 (N_1260,N_1177,N_1052);
xor U1261 (N_1261,N_1086,N_1103);
nor U1262 (N_1262,N_1102,N_1106);
xnor U1263 (N_1263,N_1104,N_1162);
or U1264 (N_1264,N_1076,N_1108);
or U1265 (N_1265,N_1171,N_1172);
nand U1266 (N_1266,N_1028,N_1091);
nor U1267 (N_1267,N_1131,N_1027);
nor U1268 (N_1268,N_1170,N_1069);
xnor U1269 (N_1269,N_1178,N_1144);
xor U1270 (N_1270,N_1063,N_1114);
nand U1271 (N_1271,N_1148,N_1115);
nand U1272 (N_1272,N_1159,N_1151);
nor U1273 (N_1273,N_1164,N_1190);
nor U1274 (N_1274,N_1179,N_1168);
and U1275 (N_1275,N_1071,N_1165);
nor U1276 (N_1276,N_1183,N_1176);
and U1277 (N_1277,N_1111,N_1055);
nor U1278 (N_1278,N_1026,N_1073);
nand U1279 (N_1279,N_1136,N_1006);
nand U1280 (N_1280,N_1158,N_1133);
nand U1281 (N_1281,N_1117,N_1175);
nand U1282 (N_1282,N_1127,N_1036);
nor U1283 (N_1283,N_1185,N_1075);
nor U1284 (N_1284,N_1046,N_1180);
nor U1285 (N_1285,N_1045,N_1101);
or U1286 (N_1286,N_1070,N_1121);
nor U1287 (N_1287,N_1039,N_1109);
nand U1288 (N_1288,N_1096,N_1074);
nor U1289 (N_1289,N_1132,N_1186);
nand U1290 (N_1290,N_1011,N_1134);
nor U1291 (N_1291,N_1156,N_1049);
or U1292 (N_1292,N_1195,N_1066);
and U1293 (N_1293,N_1057,N_1040);
xor U1294 (N_1294,N_1198,N_1042);
xor U1295 (N_1295,N_1125,N_1181);
or U1296 (N_1296,N_1188,N_1105);
or U1297 (N_1297,N_1025,N_1099);
nand U1298 (N_1298,N_1012,N_1142);
nand U1299 (N_1299,N_1155,N_1058);
nor U1300 (N_1300,N_1006,N_1120);
and U1301 (N_1301,N_1094,N_1195);
xnor U1302 (N_1302,N_1166,N_1139);
xor U1303 (N_1303,N_1127,N_1031);
nor U1304 (N_1304,N_1053,N_1144);
and U1305 (N_1305,N_1134,N_1067);
or U1306 (N_1306,N_1112,N_1150);
xnor U1307 (N_1307,N_1042,N_1199);
nor U1308 (N_1308,N_1152,N_1095);
xor U1309 (N_1309,N_1105,N_1046);
or U1310 (N_1310,N_1087,N_1088);
nand U1311 (N_1311,N_1064,N_1123);
or U1312 (N_1312,N_1040,N_1046);
or U1313 (N_1313,N_1069,N_1116);
nand U1314 (N_1314,N_1007,N_1061);
or U1315 (N_1315,N_1155,N_1119);
nand U1316 (N_1316,N_1161,N_1061);
and U1317 (N_1317,N_1008,N_1018);
xor U1318 (N_1318,N_1067,N_1068);
or U1319 (N_1319,N_1106,N_1138);
and U1320 (N_1320,N_1032,N_1119);
or U1321 (N_1321,N_1122,N_1072);
or U1322 (N_1322,N_1113,N_1036);
nand U1323 (N_1323,N_1192,N_1186);
nor U1324 (N_1324,N_1124,N_1181);
and U1325 (N_1325,N_1075,N_1007);
nor U1326 (N_1326,N_1067,N_1116);
nor U1327 (N_1327,N_1165,N_1155);
and U1328 (N_1328,N_1068,N_1003);
or U1329 (N_1329,N_1155,N_1174);
and U1330 (N_1330,N_1185,N_1196);
and U1331 (N_1331,N_1016,N_1074);
nor U1332 (N_1332,N_1160,N_1175);
xor U1333 (N_1333,N_1185,N_1146);
nand U1334 (N_1334,N_1131,N_1118);
nor U1335 (N_1335,N_1159,N_1025);
or U1336 (N_1336,N_1075,N_1022);
nor U1337 (N_1337,N_1042,N_1183);
nor U1338 (N_1338,N_1086,N_1104);
xor U1339 (N_1339,N_1049,N_1099);
and U1340 (N_1340,N_1125,N_1069);
nor U1341 (N_1341,N_1113,N_1086);
nor U1342 (N_1342,N_1070,N_1057);
nand U1343 (N_1343,N_1184,N_1141);
nand U1344 (N_1344,N_1182,N_1033);
xor U1345 (N_1345,N_1036,N_1117);
nor U1346 (N_1346,N_1144,N_1049);
xor U1347 (N_1347,N_1134,N_1145);
and U1348 (N_1348,N_1174,N_1062);
nor U1349 (N_1349,N_1191,N_1173);
nand U1350 (N_1350,N_1118,N_1193);
xnor U1351 (N_1351,N_1020,N_1089);
nor U1352 (N_1352,N_1028,N_1163);
xor U1353 (N_1353,N_1198,N_1196);
or U1354 (N_1354,N_1086,N_1026);
or U1355 (N_1355,N_1147,N_1052);
nor U1356 (N_1356,N_1052,N_1078);
nor U1357 (N_1357,N_1189,N_1103);
or U1358 (N_1358,N_1042,N_1149);
nor U1359 (N_1359,N_1082,N_1033);
xnor U1360 (N_1360,N_1068,N_1055);
and U1361 (N_1361,N_1038,N_1040);
nand U1362 (N_1362,N_1181,N_1008);
nand U1363 (N_1363,N_1193,N_1063);
xnor U1364 (N_1364,N_1097,N_1104);
or U1365 (N_1365,N_1085,N_1003);
nor U1366 (N_1366,N_1164,N_1046);
nor U1367 (N_1367,N_1154,N_1117);
or U1368 (N_1368,N_1154,N_1175);
or U1369 (N_1369,N_1151,N_1133);
nand U1370 (N_1370,N_1151,N_1130);
xnor U1371 (N_1371,N_1115,N_1091);
xnor U1372 (N_1372,N_1066,N_1002);
and U1373 (N_1373,N_1104,N_1106);
nor U1374 (N_1374,N_1009,N_1061);
xnor U1375 (N_1375,N_1057,N_1197);
and U1376 (N_1376,N_1024,N_1116);
or U1377 (N_1377,N_1022,N_1025);
nor U1378 (N_1378,N_1072,N_1153);
or U1379 (N_1379,N_1139,N_1018);
nand U1380 (N_1380,N_1139,N_1049);
xnor U1381 (N_1381,N_1140,N_1047);
xor U1382 (N_1382,N_1100,N_1134);
nor U1383 (N_1383,N_1029,N_1134);
or U1384 (N_1384,N_1076,N_1042);
xnor U1385 (N_1385,N_1151,N_1040);
xnor U1386 (N_1386,N_1039,N_1185);
xor U1387 (N_1387,N_1150,N_1027);
nand U1388 (N_1388,N_1087,N_1016);
nor U1389 (N_1389,N_1011,N_1151);
or U1390 (N_1390,N_1146,N_1014);
xor U1391 (N_1391,N_1111,N_1174);
nand U1392 (N_1392,N_1070,N_1044);
nand U1393 (N_1393,N_1049,N_1178);
xor U1394 (N_1394,N_1057,N_1051);
xor U1395 (N_1395,N_1173,N_1023);
xnor U1396 (N_1396,N_1148,N_1175);
and U1397 (N_1397,N_1190,N_1187);
nor U1398 (N_1398,N_1129,N_1190);
and U1399 (N_1399,N_1125,N_1117);
or U1400 (N_1400,N_1321,N_1209);
nor U1401 (N_1401,N_1381,N_1390);
and U1402 (N_1402,N_1374,N_1322);
nor U1403 (N_1403,N_1278,N_1287);
or U1404 (N_1404,N_1257,N_1235);
and U1405 (N_1405,N_1254,N_1228);
nor U1406 (N_1406,N_1326,N_1301);
and U1407 (N_1407,N_1219,N_1217);
xor U1408 (N_1408,N_1268,N_1393);
xor U1409 (N_1409,N_1259,N_1271);
and U1410 (N_1410,N_1221,N_1345);
and U1411 (N_1411,N_1351,N_1303);
nor U1412 (N_1412,N_1281,N_1330);
and U1413 (N_1413,N_1250,N_1230);
and U1414 (N_1414,N_1289,N_1391);
nor U1415 (N_1415,N_1332,N_1333);
and U1416 (N_1416,N_1372,N_1280);
or U1417 (N_1417,N_1223,N_1261);
or U1418 (N_1418,N_1357,N_1324);
and U1419 (N_1419,N_1376,N_1350);
and U1420 (N_1420,N_1310,N_1383);
xnor U1421 (N_1421,N_1343,N_1234);
or U1422 (N_1422,N_1279,N_1236);
or U1423 (N_1423,N_1312,N_1215);
xnor U1424 (N_1424,N_1202,N_1258);
or U1425 (N_1425,N_1243,N_1389);
nand U1426 (N_1426,N_1212,N_1360);
and U1427 (N_1427,N_1249,N_1238);
or U1428 (N_1428,N_1331,N_1262);
or U1429 (N_1429,N_1328,N_1292);
or U1430 (N_1430,N_1361,N_1348);
and U1431 (N_1431,N_1338,N_1335);
nor U1432 (N_1432,N_1384,N_1283);
xor U1433 (N_1433,N_1399,N_1340);
nand U1434 (N_1434,N_1255,N_1210);
nor U1435 (N_1435,N_1318,N_1339);
nor U1436 (N_1436,N_1298,N_1222);
and U1437 (N_1437,N_1285,N_1233);
or U1438 (N_1438,N_1251,N_1371);
and U1439 (N_1439,N_1225,N_1355);
nand U1440 (N_1440,N_1398,N_1378);
nor U1441 (N_1441,N_1375,N_1267);
nand U1442 (N_1442,N_1241,N_1311);
or U1443 (N_1443,N_1307,N_1299);
or U1444 (N_1444,N_1213,N_1203);
nor U1445 (N_1445,N_1227,N_1308);
nand U1446 (N_1446,N_1309,N_1353);
nand U1447 (N_1447,N_1247,N_1356);
xor U1448 (N_1448,N_1269,N_1366);
and U1449 (N_1449,N_1265,N_1349);
nor U1450 (N_1450,N_1276,N_1242);
or U1451 (N_1451,N_1362,N_1205);
or U1452 (N_1452,N_1337,N_1245);
xor U1453 (N_1453,N_1346,N_1231);
and U1454 (N_1454,N_1296,N_1305);
nor U1455 (N_1455,N_1368,N_1320);
and U1456 (N_1456,N_1237,N_1282);
nor U1457 (N_1457,N_1352,N_1358);
xnor U1458 (N_1458,N_1388,N_1341);
or U1459 (N_1459,N_1288,N_1380);
or U1460 (N_1460,N_1314,N_1291);
or U1461 (N_1461,N_1273,N_1373);
nor U1462 (N_1462,N_1260,N_1379);
nor U1463 (N_1463,N_1240,N_1208);
or U1464 (N_1464,N_1300,N_1207);
or U1465 (N_1465,N_1263,N_1377);
nand U1466 (N_1466,N_1329,N_1214);
nor U1467 (N_1467,N_1369,N_1274);
nand U1468 (N_1468,N_1218,N_1284);
or U1469 (N_1469,N_1295,N_1396);
and U1470 (N_1470,N_1232,N_1253);
and U1471 (N_1471,N_1275,N_1395);
and U1472 (N_1472,N_1270,N_1370);
nand U1473 (N_1473,N_1319,N_1290);
nand U1474 (N_1474,N_1293,N_1385);
nor U1475 (N_1475,N_1327,N_1264);
or U1476 (N_1476,N_1323,N_1204);
nor U1477 (N_1477,N_1397,N_1317);
xor U1478 (N_1478,N_1313,N_1387);
xor U1479 (N_1479,N_1315,N_1316);
or U1480 (N_1480,N_1256,N_1342);
and U1481 (N_1481,N_1304,N_1392);
nand U1482 (N_1482,N_1252,N_1359);
xnor U1483 (N_1483,N_1277,N_1266);
nor U1484 (N_1484,N_1325,N_1229);
nor U1485 (N_1485,N_1347,N_1365);
nand U1486 (N_1486,N_1200,N_1226);
or U1487 (N_1487,N_1364,N_1246);
and U1488 (N_1488,N_1367,N_1239);
nand U1489 (N_1489,N_1363,N_1272);
or U1490 (N_1490,N_1297,N_1220);
nor U1491 (N_1491,N_1382,N_1206);
and U1492 (N_1492,N_1394,N_1344);
or U1493 (N_1493,N_1354,N_1336);
nor U1494 (N_1494,N_1211,N_1216);
and U1495 (N_1495,N_1244,N_1334);
nand U1496 (N_1496,N_1302,N_1294);
or U1497 (N_1497,N_1386,N_1286);
xnor U1498 (N_1498,N_1224,N_1248);
xor U1499 (N_1499,N_1306,N_1201);
xor U1500 (N_1500,N_1315,N_1323);
or U1501 (N_1501,N_1350,N_1285);
nor U1502 (N_1502,N_1270,N_1342);
nor U1503 (N_1503,N_1206,N_1288);
or U1504 (N_1504,N_1328,N_1304);
nor U1505 (N_1505,N_1248,N_1261);
or U1506 (N_1506,N_1300,N_1353);
and U1507 (N_1507,N_1264,N_1247);
nand U1508 (N_1508,N_1287,N_1312);
or U1509 (N_1509,N_1367,N_1221);
or U1510 (N_1510,N_1399,N_1386);
nand U1511 (N_1511,N_1229,N_1231);
and U1512 (N_1512,N_1275,N_1238);
nand U1513 (N_1513,N_1286,N_1293);
nand U1514 (N_1514,N_1291,N_1254);
nor U1515 (N_1515,N_1259,N_1388);
and U1516 (N_1516,N_1271,N_1261);
or U1517 (N_1517,N_1391,N_1203);
nor U1518 (N_1518,N_1282,N_1300);
and U1519 (N_1519,N_1373,N_1307);
nor U1520 (N_1520,N_1374,N_1376);
nor U1521 (N_1521,N_1240,N_1383);
and U1522 (N_1522,N_1397,N_1325);
xnor U1523 (N_1523,N_1238,N_1288);
and U1524 (N_1524,N_1222,N_1257);
xnor U1525 (N_1525,N_1351,N_1346);
or U1526 (N_1526,N_1331,N_1285);
xor U1527 (N_1527,N_1345,N_1211);
or U1528 (N_1528,N_1245,N_1278);
xor U1529 (N_1529,N_1248,N_1242);
and U1530 (N_1530,N_1390,N_1321);
nand U1531 (N_1531,N_1206,N_1337);
and U1532 (N_1532,N_1267,N_1327);
and U1533 (N_1533,N_1366,N_1309);
nor U1534 (N_1534,N_1244,N_1363);
nand U1535 (N_1535,N_1348,N_1357);
or U1536 (N_1536,N_1397,N_1281);
xnor U1537 (N_1537,N_1225,N_1370);
xor U1538 (N_1538,N_1332,N_1279);
or U1539 (N_1539,N_1297,N_1284);
nor U1540 (N_1540,N_1291,N_1353);
and U1541 (N_1541,N_1282,N_1362);
or U1542 (N_1542,N_1316,N_1218);
nand U1543 (N_1543,N_1253,N_1357);
or U1544 (N_1544,N_1311,N_1278);
nor U1545 (N_1545,N_1397,N_1349);
nor U1546 (N_1546,N_1226,N_1242);
and U1547 (N_1547,N_1258,N_1273);
xor U1548 (N_1548,N_1313,N_1352);
and U1549 (N_1549,N_1364,N_1260);
or U1550 (N_1550,N_1389,N_1370);
and U1551 (N_1551,N_1234,N_1373);
nand U1552 (N_1552,N_1219,N_1379);
nor U1553 (N_1553,N_1365,N_1300);
or U1554 (N_1554,N_1276,N_1283);
nand U1555 (N_1555,N_1372,N_1234);
nand U1556 (N_1556,N_1376,N_1371);
and U1557 (N_1557,N_1281,N_1221);
nand U1558 (N_1558,N_1222,N_1368);
nor U1559 (N_1559,N_1372,N_1248);
nor U1560 (N_1560,N_1379,N_1394);
nor U1561 (N_1561,N_1378,N_1292);
nor U1562 (N_1562,N_1210,N_1205);
nand U1563 (N_1563,N_1233,N_1216);
xnor U1564 (N_1564,N_1291,N_1247);
or U1565 (N_1565,N_1335,N_1336);
nor U1566 (N_1566,N_1333,N_1393);
nor U1567 (N_1567,N_1394,N_1368);
nor U1568 (N_1568,N_1291,N_1211);
nand U1569 (N_1569,N_1382,N_1298);
or U1570 (N_1570,N_1250,N_1350);
nor U1571 (N_1571,N_1287,N_1208);
nor U1572 (N_1572,N_1383,N_1366);
and U1573 (N_1573,N_1355,N_1219);
or U1574 (N_1574,N_1295,N_1323);
nor U1575 (N_1575,N_1306,N_1324);
and U1576 (N_1576,N_1391,N_1340);
nand U1577 (N_1577,N_1242,N_1348);
and U1578 (N_1578,N_1338,N_1385);
nand U1579 (N_1579,N_1389,N_1339);
nand U1580 (N_1580,N_1311,N_1379);
nor U1581 (N_1581,N_1319,N_1229);
xnor U1582 (N_1582,N_1337,N_1251);
nand U1583 (N_1583,N_1212,N_1248);
and U1584 (N_1584,N_1376,N_1373);
xnor U1585 (N_1585,N_1238,N_1236);
nand U1586 (N_1586,N_1243,N_1328);
xor U1587 (N_1587,N_1263,N_1343);
nand U1588 (N_1588,N_1239,N_1270);
or U1589 (N_1589,N_1240,N_1328);
and U1590 (N_1590,N_1327,N_1359);
nand U1591 (N_1591,N_1352,N_1217);
nand U1592 (N_1592,N_1384,N_1320);
and U1593 (N_1593,N_1268,N_1398);
nand U1594 (N_1594,N_1347,N_1226);
nor U1595 (N_1595,N_1383,N_1382);
xnor U1596 (N_1596,N_1261,N_1329);
nor U1597 (N_1597,N_1215,N_1367);
nand U1598 (N_1598,N_1321,N_1362);
nor U1599 (N_1599,N_1281,N_1384);
nand U1600 (N_1600,N_1434,N_1555);
nand U1601 (N_1601,N_1535,N_1483);
nor U1602 (N_1602,N_1580,N_1497);
and U1603 (N_1603,N_1442,N_1542);
nor U1604 (N_1604,N_1563,N_1577);
nand U1605 (N_1605,N_1583,N_1566);
and U1606 (N_1606,N_1456,N_1436);
xnor U1607 (N_1607,N_1430,N_1552);
nand U1608 (N_1608,N_1545,N_1559);
or U1609 (N_1609,N_1575,N_1443);
nand U1610 (N_1610,N_1576,N_1549);
nor U1611 (N_1611,N_1496,N_1570);
or U1612 (N_1612,N_1546,N_1595);
and U1613 (N_1613,N_1447,N_1529);
xor U1614 (N_1614,N_1551,N_1424);
or U1615 (N_1615,N_1517,N_1428);
nor U1616 (N_1616,N_1467,N_1544);
nor U1617 (N_1617,N_1416,N_1597);
xor U1618 (N_1618,N_1413,N_1573);
nand U1619 (N_1619,N_1564,N_1585);
xnor U1620 (N_1620,N_1525,N_1533);
xor U1621 (N_1621,N_1536,N_1418);
or U1622 (N_1622,N_1522,N_1485);
and U1623 (N_1623,N_1515,N_1490);
and U1624 (N_1624,N_1593,N_1579);
or U1625 (N_1625,N_1403,N_1561);
nor U1626 (N_1626,N_1598,N_1444);
xnor U1627 (N_1627,N_1588,N_1574);
or U1628 (N_1628,N_1537,N_1468);
and U1629 (N_1629,N_1402,N_1568);
nor U1630 (N_1630,N_1586,N_1590);
xor U1631 (N_1631,N_1569,N_1441);
nand U1632 (N_1632,N_1550,N_1565);
and U1633 (N_1633,N_1412,N_1404);
or U1634 (N_1634,N_1464,N_1477);
nand U1635 (N_1635,N_1431,N_1465);
and U1636 (N_1636,N_1526,N_1448);
nor U1637 (N_1637,N_1459,N_1511);
or U1638 (N_1638,N_1400,N_1591);
nor U1639 (N_1639,N_1524,N_1445);
nand U1640 (N_1640,N_1407,N_1421);
or U1641 (N_1641,N_1452,N_1541);
and U1642 (N_1642,N_1401,N_1491);
nand U1643 (N_1643,N_1474,N_1503);
nand U1644 (N_1644,N_1499,N_1506);
or U1645 (N_1645,N_1558,N_1548);
nor U1646 (N_1646,N_1417,N_1420);
or U1647 (N_1647,N_1440,N_1534);
nand U1648 (N_1648,N_1543,N_1571);
nand U1649 (N_1649,N_1433,N_1501);
nor U1650 (N_1650,N_1406,N_1481);
xor U1651 (N_1651,N_1446,N_1556);
xor U1652 (N_1652,N_1553,N_1594);
nor U1653 (N_1653,N_1419,N_1581);
or U1654 (N_1654,N_1495,N_1449);
nand U1655 (N_1655,N_1560,N_1531);
nand U1656 (N_1656,N_1518,N_1427);
nor U1657 (N_1657,N_1508,N_1502);
xnor U1658 (N_1658,N_1482,N_1516);
xor U1659 (N_1659,N_1457,N_1409);
nor U1660 (N_1660,N_1587,N_1513);
xor U1661 (N_1661,N_1514,N_1423);
and U1662 (N_1662,N_1547,N_1469);
nor U1663 (N_1663,N_1429,N_1500);
xnor U1664 (N_1664,N_1472,N_1486);
xor U1665 (N_1665,N_1596,N_1432);
xor U1666 (N_1666,N_1435,N_1478);
nand U1667 (N_1667,N_1425,N_1422);
nand U1668 (N_1668,N_1487,N_1527);
or U1669 (N_1669,N_1453,N_1538);
or U1670 (N_1670,N_1461,N_1521);
xnor U1671 (N_1671,N_1540,N_1466);
nor U1672 (N_1672,N_1523,N_1528);
or U1673 (N_1673,N_1498,N_1492);
nand U1674 (N_1674,N_1584,N_1557);
nand U1675 (N_1675,N_1562,N_1480);
nand U1676 (N_1676,N_1450,N_1494);
nor U1677 (N_1677,N_1414,N_1475);
nor U1678 (N_1678,N_1572,N_1473);
xor U1679 (N_1679,N_1520,N_1519);
xor U1680 (N_1680,N_1512,N_1439);
and U1681 (N_1681,N_1451,N_1504);
and U1682 (N_1682,N_1426,N_1470);
or U1683 (N_1683,N_1455,N_1463);
nor U1684 (N_1684,N_1493,N_1589);
nand U1685 (N_1685,N_1437,N_1484);
nor U1686 (N_1686,N_1460,N_1510);
nor U1687 (N_1687,N_1471,N_1410);
xnor U1688 (N_1688,N_1462,N_1582);
nor U1689 (N_1689,N_1599,N_1539);
nand U1690 (N_1690,N_1505,N_1592);
or U1691 (N_1691,N_1509,N_1438);
nor U1692 (N_1692,N_1479,N_1507);
or U1693 (N_1693,N_1567,N_1411);
xor U1694 (N_1694,N_1408,N_1554);
nor U1695 (N_1695,N_1530,N_1476);
xnor U1696 (N_1696,N_1454,N_1532);
nor U1697 (N_1697,N_1488,N_1415);
xor U1698 (N_1698,N_1405,N_1489);
or U1699 (N_1699,N_1458,N_1578);
nor U1700 (N_1700,N_1541,N_1544);
xnor U1701 (N_1701,N_1541,N_1487);
nand U1702 (N_1702,N_1508,N_1589);
xor U1703 (N_1703,N_1561,N_1520);
or U1704 (N_1704,N_1461,N_1493);
nand U1705 (N_1705,N_1437,N_1514);
or U1706 (N_1706,N_1459,N_1540);
nor U1707 (N_1707,N_1537,N_1585);
or U1708 (N_1708,N_1597,N_1529);
and U1709 (N_1709,N_1597,N_1558);
xor U1710 (N_1710,N_1520,N_1442);
and U1711 (N_1711,N_1539,N_1522);
nand U1712 (N_1712,N_1478,N_1429);
nor U1713 (N_1713,N_1554,N_1468);
nand U1714 (N_1714,N_1471,N_1445);
or U1715 (N_1715,N_1415,N_1407);
xor U1716 (N_1716,N_1428,N_1544);
or U1717 (N_1717,N_1406,N_1540);
and U1718 (N_1718,N_1499,N_1593);
and U1719 (N_1719,N_1599,N_1463);
nor U1720 (N_1720,N_1516,N_1500);
nor U1721 (N_1721,N_1519,N_1412);
or U1722 (N_1722,N_1480,N_1447);
nand U1723 (N_1723,N_1581,N_1575);
and U1724 (N_1724,N_1553,N_1469);
nand U1725 (N_1725,N_1406,N_1500);
or U1726 (N_1726,N_1526,N_1566);
nand U1727 (N_1727,N_1422,N_1428);
or U1728 (N_1728,N_1448,N_1518);
xnor U1729 (N_1729,N_1527,N_1500);
nand U1730 (N_1730,N_1500,N_1440);
xor U1731 (N_1731,N_1453,N_1413);
nand U1732 (N_1732,N_1400,N_1559);
or U1733 (N_1733,N_1566,N_1571);
nand U1734 (N_1734,N_1508,N_1559);
and U1735 (N_1735,N_1422,N_1470);
or U1736 (N_1736,N_1504,N_1484);
and U1737 (N_1737,N_1570,N_1518);
nor U1738 (N_1738,N_1493,N_1430);
nor U1739 (N_1739,N_1544,N_1439);
or U1740 (N_1740,N_1530,N_1434);
nor U1741 (N_1741,N_1546,N_1469);
nand U1742 (N_1742,N_1451,N_1440);
nor U1743 (N_1743,N_1448,N_1528);
or U1744 (N_1744,N_1492,N_1530);
or U1745 (N_1745,N_1568,N_1433);
nor U1746 (N_1746,N_1554,N_1534);
nor U1747 (N_1747,N_1429,N_1417);
xor U1748 (N_1748,N_1594,N_1557);
nor U1749 (N_1749,N_1596,N_1550);
and U1750 (N_1750,N_1513,N_1404);
and U1751 (N_1751,N_1455,N_1445);
xor U1752 (N_1752,N_1476,N_1451);
nor U1753 (N_1753,N_1413,N_1548);
or U1754 (N_1754,N_1405,N_1515);
and U1755 (N_1755,N_1509,N_1517);
and U1756 (N_1756,N_1475,N_1471);
and U1757 (N_1757,N_1484,N_1428);
nor U1758 (N_1758,N_1557,N_1445);
nand U1759 (N_1759,N_1433,N_1444);
nor U1760 (N_1760,N_1545,N_1494);
xnor U1761 (N_1761,N_1531,N_1426);
xnor U1762 (N_1762,N_1562,N_1425);
or U1763 (N_1763,N_1465,N_1505);
nor U1764 (N_1764,N_1475,N_1587);
and U1765 (N_1765,N_1539,N_1446);
xnor U1766 (N_1766,N_1466,N_1553);
or U1767 (N_1767,N_1454,N_1428);
or U1768 (N_1768,N_1419,N_1597);
and U1769 (N_1769,N_1481,N_1430);
nor U1770 (N_1770,N_1419,N_1438);
xor U1771 (N_1771,N_1417,N_1451);
nand U1772 (N_1772,N_1422,N_1552);
xnor U1773 (N_1773,N_1527,N_1426);
xor U1774 (N_1774,N_1580,N_1532);
xor U1775 (N_1775,N_1583,N_1508);
xnor U1776 (N_1776,N_1441,N_1494);
and U1777 (N_1777,N_1451,N_1516);
nand U1778 (N_1778,N_1484,N_1479);
nand U1779 (N_1779,N_1563,N_1402);
or U1780 (N_1780,N_1535,N_1401);
nand U1781 (N_1781,N_1594,N_1461);
nand U1782 (N_1782,N_1548,N_1490);
and U1783 (N_1783,N_1588,N_1448);
and U1784 (N_1784,N_1534,N_1502);
nor U1785 (N_1785,N_1556,N_1519);
nand U1786 (N_1786,N_1449,N_1440);
nor U1787 (N_1787,N_1588,N_1554);
nand U1788 (N_1788,N_1528,N_1571);
or U1789 (N_1789,N_1533,N_1408);
nand U1790 (N_1790,N_1525,N_1518);
nor U1791 (N_1791,N_1503,N_1446);
and U1792 (N_1792,N_1531,N_1498);
and U1793 (N_1793,N_1480,N_1530);
nor U1794 (N_1794,N_1501,N_1429);
nor U1795 (N_1795,N_1578,N_1521);
nand U1796 (N_1796,N_1413,N_1472);
and U1797 (N_1797,N_1467,N_1421);
nor U1798 (N_1798,N_1438,N_1401);
nor U1799 (N_1799,N_1551,N_1483);
nor U1800 (N_1800,N_1635,N_1640);
nor U1801 (N_1801,N_1776,N_1716);
nor U1802 (N_1802,N_1792,N_1661);
xnor U1803 (N_1803,N_1689,N_1780);
xnor U1804 (N_1804,N_1646,N_1624);
and U1805 (N_1805,N_1673,N_1739);
nand U1806 (N_1806,N_1772,N_1628);
or U1807 (N_1807,N_1731,N_1629);
nor U1808 (N_1808,N_1724,N_1741);
xor U1809 (N_1809,N_1777,N_1759);
nand U1810 (N_1810,N_1799,N_1773);
nand U1811 (N_1811,N_1730,N_1649);
or U1812 (N_1812,N_1729,N_1656);
xnor U1813 (N_1813,N_1658,N_1634);
nand U1814 (N_1814,N_1708,N_1665);
nand U1815 (N_1815,N_1625,N_1722);
nor U1816 (N_1816,N_1756,N_1745);
or U1817 (N_1817,N_1618,N_1668);
or U1818 (N_1818,N_1647,N_1762);
nand U1819 (N_1819,N_1788,N_1636);
nor U1820 (N_1820,N_1648,N_1601);
or U1821 (N_1821,N_1727,N_1717);
and U1822 (N_1822,N_1767,N_1642);
and U1823 (N_1823,N_1796,N_1753);
and U1824 (N_1824,N_1736,N_1734);
xor U1825 (N_1825,N_1627,N_1686);
nor U1826 (N_1826,N_1652,N_1651);
nor U1827 (N_1827,N_1698,N_1757);
xor U1828 (N_1828,N_1755,N_1691);
nand U1829 (N_1829,N_1603,N_1763);
xor U1830 (N_1830,N_1700,N_1781);
or U1831 (N_1831,N_1630,N_1619);
xor U1832 (N_1832,N_1703,N_1768);
nor U1833 (N_1833,N_1742,N_1679);
nand U1834 (N_1834,N_1637,N_1670);
xor U1835 (N_1835,N_1687,N_1733);
nand U1836 (N_1836,N_1682,N_1662);
and U1837 (N_1837,N_1790,N_1655);
and U1838 (N_1838,N_1617,N_1611);
xnor U1839 (N_1839,N_1709,N_1723);
and U1840 (N_1840,N_1675,N_1654);
xnor U1841 (N_1841,N_1795,N_1732);
nor U1842 (N_1842,N_1650,N_1692);
or U1843 (N_1843,N_1684,N_1794);
or U1844 (N_1844,N_1664,N_1787);
nor U1845 (N_1845,N_1643,N_1713);
nand U1846 (N_1846,N_1688,N_1631);
and U1847 (N_1847,N_1743,N_1786);
nand U1848 (N_1848,N_1605,N_1669);
nand U1849 (N_1849,N_1750,N_1632);
xnor U1850 (N_1850,N_1707,N_1602);
nand U1851 (N_1851,N_1798,N_1633);
and U1852 (N_1852,N_1746,N_1663);
or U1853 (N_1853,N_1667,N_1789);
or U1854 (N_1854,N_1770,N_1740);
nor U1855 (N_1855,N_1641,N_1769);
xnor U1856 (N_1856,N_1657,N_1712);
and U1857 (N_1857,N_1749,N_1711);
nor U1858 (N_1858,N_1725,N_1674);
or U1859 (N_1859,N_1685,N_1678);
nor U1860 (N_1860,N_1613,N_1760);
or U1861 (N_1861,N_1761,N_1620);
xor U1862 (N_1862,N_1666,N_1683);
xnor U1863 (N_1863,N_1728,N_1639);
nor U1864 (N_1864,N_1653,N_1719);
or U1865 (N_1865,N_1748,N_1735);
or U1866 (N_1866,N_1701,N_1775);
xor U1867 (N_1867,N_1737,N_1785);
xor U1868 (N_1868,N_1609,N_1720);
and U1869 (N_1869,N_1695,N_1784);
and U1870 (N_1870,N_1771,N_1751);
xor U1871 (N_1871,N_1680,N_1704);
nor U1872 (N_1872,N_1793,N_1797);
nand U1873 (N_1873,N_1774,N_1766);
nand U1874 (N_1874,N_1677,N_1612);
xor U1875 (N_1875,N_1659,N_1660);
nand U1876 (N_1876,N_1623,N_1606);
and U1877 (N_1877,N_1778,N_1783);
or U1878 (N_1878,N_1718,N_1693);
and U1879 (N_1879,N_1738,N_1616);
nand U1880 (N_1880,N_1715,N_1690);
xnor U1881 (N_1881,N_1604,N_1644);
or U1882 (N_1882,N_1754,N_1779);
nand U1883 (N_1883,N_1607,N_1621);
nor U1884 (N_1884,N_1744,N_1600);
nand U1885 (N_1885,N_1764,N_1638);
or U1886 (N_1886,N_1615,N_1752);
xnor U1887 (N_1887,N_1671,N_1681);
nand U1888 (N_1888,N_1714,N_1696);
or U1889 (N_1889,N_1702,N_1608);
nand U1890 (N_1890,N_1676,N_1694);
nand U1891 (N_1891,N_1705,N_1726);
or U1892 (N_1892,N_1710,N_1645);
xor U1893 (N_1893,N_1610,N_1699);
nor U1894 (N_1894,N_1614,N_1721);
nor U1895 (N_1895,N_1758,N_1706);
xnor U1896 (N_1896,N_1672,N_1626);
xor U1897 (N_1897,N_1622,N_1697);
nor U1898 (N_1898,N_1791,N_1782);
xnor U1899 (N_1899,N_1747,N_1765);
nor U1900 (N_1900,N_1691,N_1784);
or U1901 (N_1901,N_1737,N_1752);
or U1902 (N_1902,N_1644,N_1647);
xnor U1903 (N_1903,N_1615,N_1621);
and U1904 (N_1904,N_1788,N_1675);
xor U1905 (N_1905,N_1625,N_1788);
or U1906 (N_1906,N_1734,N_1751);
and U1907 (N_1907,N_1667,N_1609);
or U1908 (N_1908,N_1742,N_1635);
and U1909 (N_1909,N_1601,N_1624);
and U1910 (N_1910,N_1794,N_1679);
or U1911 (N_1911,N_1773,N_1762);
and U1912 (N_1912,N_1625,N_1633);
nor U1913 (N_1913,N_1667,N_1652);
xor U1914 (N_1914,N_1637,N_1720);
nand U1915 (N_1915,N_1770,N_1783);
nor U1916 (N_1916,N_1681,N_1633);
or U1917 (N_1917,N_1607,N_1698);
xnor U1918 (N_1918,N_1789,N_1747);
and U1919 (N_1919,N_1779,N_1690);
nor U1920 (N_1920,N_1756,N_1685);
or U1921 (N_1921,N_1610,N_1705);
nor U1922 (N_1922,N_1777,N_1667);
or U1923 (N_1923,N_1676,N_1780);
xor U1924 (N_1924,N_1791,N_1795);
nand U1925 (N_1925,N_1722,N_1705);
and U1926 (N_1926,N_1771,N_1769);
xor U1927 (N_1927,N_1671,N_1629);
or U1928 (N_1928,N_1635,N_1669);
nor U1929 (N_1929,N_1611,N_1747);
or U1930 (N_1930,N_1644,N_1610);
nand U1931 (N_1931,N_1700,N_1763);
nor U1932 (N_1932,N_1772,N_1731);
nor U1933 (N_1933,N_1756,N_1785);
or U1934 (N_1934,N_1759,N_1652);
nor U1935 (N_1935,N_1789,N_1678);
xnor U1936 (N_1936,N_1656,N_1783);
or U1937 (N_1937,N_1703,N_1731);
nand U1938 (N_1938,N_1784,N_1767);
xor U1939 (N_1939,N_1613,N_1666);
nor U1940 (N_1940,N_1724,N_1789);
xnor U1941 (N_1941,N_1614,N_1687);
or U1942 (N_1942,N_1700,N_1786);
nand U1943 (N_1943,N_1672,N_1636);
nand U1944 (N_1944,N_1644,N_1633);
or U1945 (N_1945,N_1602,N_1755);
xor U1946 (N_1946,N_1776,N_1783);
nand U1947 (N_1947,N_1792,N_1622);
nor U1948 (N_1948,N_1741,N_1644);
and U1949 (N_1949,N_1798,N_1789);
nor U1950 (N_1950,N_1748,N_1704);
and U1951 (N_1951,N_1769,N_1698);
or U1952 (N_1952,N_1765,N_1783);
nand U1953 (N_1953,N_1651,N_1793);
or U1954 (N_1954,N_1739,N_1775);
and U1955 (N_1955,N_1621,N_1602);
xor U1956 (N_1956,N_1610,N_1782);
or U1957 (N_1957,N_1729,N_1720);
xnor U1958 (N_1958,N_1633,N_1791);
nor U1959 (N_1959,N_1633,N_1789);
xnor U1960 (N_1960,N_1627,N_1737);
nand U1961 (N_1961,N_1691,N_1792);
and U1962 (N_1962,N_1608,N_1631);
xor U1963 (N_1963,N_1749,N_1779);
and U1964 (N_1964,N_1601,N_1606);
nand U1965 (N_1965,N_1698,N_1743);
or U1966 (N_1966,N_1629,N_1770);
or U1967 (N_1967,N_1722,N_1752);
nand U1968 (N_1968,N_1705,N_1661);
and U1969 (N_1969,N_1667,N_1712);
nor U1970 (N_1970,N_1716,N_1707);
nor U1971 (N_1971,N_1618,N_1621);
nand U1972 (N_1972,N_1650,N_1764);
and U1973 (N_1973,N_1783,N_1608);
or U1974 (N_1974,N_1680,N_1742);
nor U1975 (N_1975,N_1712,N_1672);
and U1976 (N_1976,N_1670,N_1742);
nand U1977 (N_1977,N_1747,N_1771);
and U1978 (N_1978,N_1682,N_1685);
nor U1979 (N_1979,N_1719,N_1794);
xor U1980 (N_1980,N_1733,N_1703);
and U1981 (N_1981,N_1682,N_1749);
or U1982 (N_1982,N_1691,N_1667);
xor U1983 (N_1983,N_1759,N_1757);
and U1984 (N_1984,N_1736,N_1752);
or U1985 (N_1985,N_1730,N_1737);
xor U1986 (N_1986,N_1689,N_1695);
or U1987 (N_1987,N_1621,N_1776);
nor U1988 (N_1988,N_1605,N_1661);
nand U1989 (N_1989,N_1601,N_1789);
or U1990 (N_1990,N_1688,N_1718);
nand U1991 (N_1991,N_1736,N_1697);
nor U1992 (N_1992,N_1735,N_1645);
xnor U1993 (N_1993,N_1676,N_1759);
or U1994 (N_1994,N_1792,N_1755);
and U1995 (N_1995,N_1646,N_1612);
and U1996 (N_1996,N_1654,N_1692);
xor U1997 (N_1997,N_1708,N_1694);
nand U1998 (N_1998,N_1725,N_1798);
nand U1999 (N_1999,N_1755,N_1760);
xnor U2000 (N_2000,N_1925,N_1891);
xnor U2001 (N_2001,N_1804,N_1887);
nor U2002 (N_2002,N_1823,N_1868);
nor U2003 (N_2003,N_1927,N_1986);
or U2004 (N_2004,N_1808,N_1842);
or U2005 (N_2005,N_1846,N_1806);
nor U2006 (N_2006,N_1888,N_1910);
nor U2007 (N_2007,N_1947,N_1997);
nand U2008 (N_2008,N_1968,N_1926);
xnor U2009 (N_2009,N_1861,N_1839);
xnor U2010 (N_2010,N_1973,N_1885);
xnor U2011 (N_2011,N_1875,N_1800);
nand U2012 (N_2012,N_1884,N_1976);
or U2013 (N_2013,N_1834,N_1992);
or U2014 (N_2014,N_1890,N_1825);
nand U2015 (N_2015,N_1993,N_1984);
nand U2016 (N_2016,N_1841,N_1961);
nor U2017 (N_2017,N_1813,N_1911);
and U2018 (N_2018,N_1867,N_1994);
and U2019 (N_2019,N_1991,N_1971);
nor U2020 (N_2020,N_1960,N_1955);
or U2021 (N_2021,N_1957,N_1965);
or U2022 (N_2022,N_1900,N_1939);
nor U2023 (N_2023,N_1801,N_1873);
and U2024 (N_2024,N_1810,N_1920);
xnor U2025 (N_2025,N_1824,N_1978);
nor U2026 (N_2026,N_1905,N_1933);
xor U2027 (N_2027,N_1835,N_1959);
and U2028 (N_2028,N_1909,N_1871);
and U2029 (N_2029,N_1901,N_1859);
nand U2030 (N_2030,N_1892,N_1923);
and U2031 (N_2031,N_1822,N_1903);
and U2032 (N_2032,N_1934,N_1860);
nor U2033 (N_2033,N_1815,N_1880);
and U2034 (N_2034,N_1844,N_1914);
nor U2035 (N_2035,N_1847,N_1811);
nor U2036 (N_2036,N_1995,N_1958);
nand U2037 (N_2037,N_1938,N_1848);
nor U2038 (N_2038,N_1896,N_1814);
xnor U2039 (N_2039,N_1831,N_1952);
or U2040 (N_2040,N_1948,N_1819);
nand U2041 (N_2041,N_1970,N_1951);
xnor U2042 (N_2042,N_1937,N_1881);
or U2043 (N_2043,N_1982,N_1866);
xnor U2044 (N_2044,N_1953,N_1969);
nor U2045 (N_2045,N_1912,N_1865);
or U2046 (N_2046,N_1830,N_1803);
or U2047 (N_2047,N_1963,N_1941);
and U2048 (N_2048,N_1907,N_1893);
and U2049 (N_2049,N_1820,N_1832);
or U2050 (N_2050,N_1836,N_1878);
nand U2051 (N_2051,N_1977,N_1802);
and U2052 (N_2052,N_1990,N_1829);
nor U2053 (N_2053,N_1929,N_1996);
xor U2054 (N_2054,N_1989,N_1854);
nand U2055 (N_2055,N_1877,N_1974);
nor U2056 (N_2056,N_1809,N_1833);
xnor U2057 (N_2057,N_1928,N_1998);
or U2058 (N_2058,N_1899,N_1858);
and U2059 (N_2059,N_1906,N_1882);
and U2060 (N_2060,N_1883,N_1975);
and U2061 (N_2061,N_1856,N_1898);
or U2062 (N_2062,N_1950,N_1840);
xor U2063 (N_2063,N_1853,N_1897);
or U2064 (N_2064,N_1837,N_1843);
or U2065 (N_2065,N_1943,N_1855);
nand U2066 (N_2066,N_1827,N_1935);
nand U2067 (N_2067,N_1944,N_1894);
or U2068 (N_2068,N_1918,N_1966);
nand U2069 (N_2069,N_1904,N_1886);
xnor U2070 (N_2070,N_1869,N_1852);
or U2071 (N_2071,N_1850,N_1936);
and U2072 (N_2072,N_1828,N_1964);
or U2073 (N_2073,N_1930,N_1940);
nand U2074 (N_2074,N_1816,N_1879);
and U2075 (N_2075,N_1863,N_1956);
nor U2076 (N_2076,N_1916,N_1987);
and U2077 (N_2077,N_1949,N_1919);
and U2078 (N_2078,N_1895,N_1979);
or U2079 (N_2079,N_1932,N_1999);
xnor U2080 (N_2080,N_1838,N_1981);
and U2081 (N_2081,N_1972,N_1849);
or U2082 (N_2082,N_1805,N_1983);
or U2083 (N_2083,N_1845,N_1988);
xor U2084 (N_2084,N_1922,N_1921);
nand U2085 (N_2085,N_1872,N_1913);
xor U2086 (N_2086,N_1985,N_1851);
nand U2087 (N_2087,N_1807,N_1946);
nand U2088 (N_2088,N_1931,N_1942);
nor U2089 (N_2089,N_1812,N_1915);
or U2090 (N_2090,N_1817,N_1967);
and U2091 (N_2091,N_1876,N_1954);
and U2092 (N_2092,N_1821,N_1902);
or U2093 (N_2093,N_1874,N_1818);
or U2094 (N_2094,N_1980,N_1917);
nor U2095 (N_2095,N_1862,N_1962);
and U2096 (N_2096,N_1924,N_1908);
nor U2097 (N_2097,N_1945,N_1870);
and U2098 (N_2098,N_1889,N_1864);
nor U2099 (N_2099,N_1857,N_1826);
or U2100 (N_2100,N_1856,N_1808);
nand U2101 (N_2101,N_1985,N_1923);
and U2102 (N_2102,N_1964,N_1875);
and U2103 (N_2103,N_1865,N_1805);
xnor U2104 (N_2104,N_1892,N_1877);
xnor U2105 (N_2105,N_1984,N_1998);
or U2106 (N_2106,N_1875,N_1851);
nand U2107 (N_2107,N_1832,N_1804);
or U2108 (N_2108,N_1982,N_1910);
nand U2109 (N_2109,N_1800,N_1921);
and U2110 (N_2110,N_1828,N_1853);
and U2111 (N_2111,N_1817,N_1829);
nor U2112 (N_2112,N_1917,N_1894);
nand U2113 (N_2113,N_1839,N_1931);
xnor U2114 (N_2114,N_1908,N_1894);
xor U2115 (N_2115,N_1939,N_1858);
nor U2116 (N_2116,N_1872,N_1917);
or U2117 (N_2117,N_1974,N_1906);
nor U2118 (N_2118,N_1905,N_1892);
xor U2119 (N_2119,N_1861,N_1909);
nor U2120 (N_2120,N_1936,N_1885);
and U2121 (N_2121,N_1840,N_1829);
xnor U2122 (N_2122,N_1805,N_1929);
or U2123 (N_2123,N_1841,N_1922);
nor U2124 (N_2124,N_1886,N_1948);
nand U2125 (N_2125,N_1908,N_1826);
or U2126 (N_2126,N_1861,N_1825);
and U2127 (N_2127,N_1944,N_1979);
xor U2128 (N_2128,N_1923,N_1801);
xnor U2129 (N_2129,N_1886,N_1847);
and U2130 (N_2130,N_1924,N_1877);
nor U2131 (N_2131,N_1930,N_1927);
nor U2132 (N_2132,N_1831,N_1900);
nor U2133 (N_2133,N_1812,N_1986);
nor U2134 (N_2134,N_1870,N_1979);
or U2135 (N_2135,N_1898,N_1921);
xor U2136 (N_2136,N_1872,N_1989);
xnor U2137 (N_2137,N_1962,N_1931);
nand U2138 (N_2138,N_1965,N_1937);
nor U2139 (N_2139,N_1962,N_1941);
nor U2140 (N_2140,N_1940,N_1883);
or U2141 (N_2141,N_1889,N_1833);
or U2142 (N_2142,N_1917,N_1979);
nor U2143 (N_2143,N_1953,N_1842);
nand U2144 (N_2144,N_1836,N_1843);
or U2145 (N_2145,N_1883,N_1938);
nand U2146 (N_2146,N_1909,N_1841);
or U2147 (N_2147,N_1955,N_1901);
nor U2148 (N_2148,N_1816,N_1897);
or U2149 (N_2149,N_1839,N_1943);
or U2150 (N_2150,N_1835,N_1875);
and U2151 (N_2151,N_1887,N_1889);
nor U2152 (N_2152,N_1916,N_1883);
or U2153 (N_2153,N_1867,N_1989);
or U2154 (N_2154,N_1812,N_1894);
xnor U2155 (N_2155,N_1891,N_1841);
xor U2156 (N_2156,N_1860,N_1932);
or U2157 (N_2157,N_1824,N_1927);
nand U2158 (N_2158,N_1859,N_1829);
xor U2159 (N_2159,N_1814,N_1873);
or U2160 (N_2160,N_1999,N_1841);
nand U2161 (N_2161,N_1850,N_1861);
and U2162 (N_2162,N_1998,N_1839);
nand U2163 (N_2163,N_1961,N_1900);
and U2164 (N_2164,N_1946,N_1948);
nor U2165 (N_2165,N_1847,N_1915);
or U2166 (N_2166,N_1824,N_1955);
and U2167 (N_2167,N_1892,N_1876);
xnor U2168 (N_2168,N_1859,N_1969);
xor U2169 (N_2169,N_1923,N_1878);
nor U2170 (N_2170,N_1914,N_1818);
nand U2171 (N_2171,N_1902,N_1908);
or U2172 (N_2172,N_1900,N_1816);
or U2173 (N_2173,N_1926,N_1853);
or U2174 (N_2174,N_1964,N_1935);
nand U2175 (N_2175,N_1826,N_1815);
nand U2176 (N_2176,N_1872,N_1919);
and U2177 (N_2177,N_1863,N_1936);
nand U2178 (N_2178,N_1822,N_1821);
or U2179 (N_2179,N_1912,N_1893);
or U2180 (N_2180,N_1944,N_1856);
and U2181 (N_2181,N_1960,N_1852);
or U2182 (N_2182,N_1882,N_1974);
nand U2183 (N_2183,N_1911,N_1926);
nand U2184 (N_2184,N_1987,N_1851);
nor U2185 (N_2185,N_1874,N_1872);
or U2186 (N_2186,N_1850,N_1927);
nand U2187 (N_2187,N_1920,N_1981);
and U2188 (N_2188,N_1921,N_1976);
nor U2189 (N_2189,N_1872,N_1964);
and U2190 (N_2190,N_1947,N_1940);
nand U2191 (N_2191,N_1882,N_1950);
or U2192 (N_2192,N_1888,N_1847);
xor U2193 (N_2193,N_1861,N_1920);
nor U2194 (N_2194,N_1897,N_1834);
nor U2195 (N_2195,N_1940,N_1819);
and U2196 (N_2196,N_1955,N_1848);
and U2197 (N_2197,N_1879,N_1825);
or U2198 (N_2198,N_1890,N_1823);
nand U2199 (N_2199,N_1873,N_1946);
nand U2200 (N_2200,N_2095,N_2142);
xnor U2201 (N_2201,N_2131,N_2091);
xor U2202 (N_2202,N_2030,N_2073);
xor U2203 (N_2203,N_2161,N_2099);
xor U2204 (N_2204,N_2184,N_2017);
nand U2205 (N_2205,N_2005,N_2086);
nand U2206 (N_2206,N_2188,N_2033);
and U2207 (N_2207,N_2066,N_2122);
xor U2208 (N_2208,N_2021,N_2039);
and U2209 (N_2209,N_2117,N_2082);
nand U2210 (N_2210,N_2153,N_2135);
nand U2211 (N_2211,N_2182,N_2047);
nand U2212 (N_2212,N_2156,N_2138);
or U2213 (N_2213,N_2111,N_2072);
or U2214 (N_2214,N_2051,N_2195);
xor U2215 (N_2215,N_2025,N_2013);
xnor U2216 (N_2216,N_2026,N_2133);
or U2217 (N_2217,N_2015,N_2067);
xnor U2218 (N_2218,N_2046,N_2063);
and U2219 (N_2219,N_2132,N_2007);
or U2220 (N_2220,N_2010,N_2089);
xnor U2221 (N_2221,N_2198,N_2029);
nor U2222 (N_2222,N_2110,N_2183);
nand U2223 (N_2223,N_2085,N_2125);
and U2224 (N_2224,N_2147,N_2162);
nor U2225 (N_2225,N_2056,N_2155);
or U2226 (N_2226,N_2105,N_2020);
nor U2227 (N_2227,N_2001,N_2052);
nand U2228 (N_2228,N_2000,N_2027);
or U2229 (N_2229,N_2103,N_2093);
xor U2230 (N_2230,N_2045,N_2194);
nand U2231 (N_2231,N_2060,N_2121);
or U2232 (N_2232,N_2053,N_2149);
xor U2233 (N_2233,N_2024,N_2168);
or U2234 (N_2234,N_2163,N_2065);
xor U2235 (N_2235,N_2115,N_2080);
nor U2236 (N_2236,N_2128,N_2075);
or U2237 (N_2237,N_2187,N_2057);
and U2238 (N_2238,N_2108,N_2196);
or U2239 (N_2239,N_2169,N_2035);
and U2240 (N_2240,N_2130,N_2112);
and U2241 (N_2241,N_2151,N_2160);
and U2242 (N_2242,N_2102,N_2127);
or U2243 (N_2243,N_2094,N_2174);
nor U2244 (N_2244,N_2074,N_2144);
nor U2245 (N_2245,N_2158,N_2088);
nand U2246 (N_2246,N_2172,N_2018);
nand U2247 (N_2247,N_2043,N_2034);
xnor U2248 (N_2248,N_2146,N_2055);
or U2249 (N_2249,N_2143,N_2070);
or U2250 (N_2250,N_2054,N_2123);
xnor U2251 (N_2251,N_2019,N_2077);
or U2252 (N_2252,N_2129,N_2036);
or U2253 (N_2253,N_2136,N_2186);
xnor U2254 (N_2254,N_2031,N_2148);
and U2255 (N_2255,N_2199,N_2120);
nor U2256 (N_2256,N_2006,N_2061);
xnor U2257 (N_2257,N_2109,N_2170);
nor U2258 (N_2258,N_2141,N_2139);
nand U2259 (N_2259,N_2197,N_2038);
nand U2260 (N_2260,N_2119,N_2049);
and U2261 (N_2261,N_2078,N_2040);
and U2262 (N_2262,N_2171,N_2193);
xnor U2263 (N_2263,N_2176,N_2076);
xor U2264 (N_2264,N_2069,N_2003);
xor U2265 (N_2265,N_2137,N_2087);
xnor U2266 (N_2266,N_2037,N_2106);
nor U2267 (N_2267,N_2028,N_2081);
or U2268 (N_2268,N_2175,N_2008);
nand U2269 (N_2269,N_2107,N_2180);
nand U2270 (N_2270,N_2097,N_2068);
nand U2271 (N_2271,N_2181,N_2071);
xnor U2272 (N_2272,N_2002,N_2165);
xnor U2273 (N_2273,N_2090,N_2004);
xnor U2274 (N_2274,N_2032,N_2022);
and U2275 (N_2275,N_2014,N_2145);
xor U2276 (N_2276,N_2118,N_2041);
nand U2277 (N_2277,N_2126,N_2092);
nor U2278 (N_2278,N_2101,N_2079);
and U2279 (N_2279,N_2050,N_2059);
nor U2280 (N_2280,N_2084,N_2179);
and U2281 (N_2281,N_2134,N_2116);
xor U2282 (N_2282,N_2100,N_2058);
xor U2283 (N_2283,N_2009,N_2113);
or U2284 (N_2284,N_2178,N_2152);
nor U2285 (N_2285,N_2167,N_2062);
xor U2286 (N_2286,N_2157,N_2154);
xnor U2287 (N_2287,N_2159,N_2011);
nor U2288 (N_2288,N_2048,N_2083);
and U2289 (N_2289,N_2189,N_2185);
nand U2290 (N_2290,N_2012,N_2173);
and U2291 (N_2291,N_2150,N_2192);
and U2292 (N_2292,N_2140,N_2098);
and U2293 (N_2293,N_2166,N_2114);
and U2294 (N_2294,N_2124,N_2016);
or U2295 (N_2295,N_2104,N_2064);
nand U2296 (N_2296,N_2096,N_2164);
nand U2297 (N_2297,N_2042,N_2191);
and U2298 (N_2298,N_2190,N_2044);
nor U2299 (N_2299,N_2023,N_2177);
xor U2300 (N_2300,N_2062,N_2086);
nand U2301 (N_2301,N_2044,N_2182);
nor U2302 (N_2302,N_2098,N_2029);
nand U2303 (N_2303,N_2005,N_2019);
nor U2304 (N_2304,N_2188,N_2192);
or U2305 (N_2305,N_2122,N_2011);
nand U2306 (N_2306,N_2095,N_2155);
nor U2307 (N_2307,N_2106,N_2019);
xnor U2308 (N_2308,N_2097,N_2063);
nor U2309 (N_2309,N_2028,N_2003);
nor U2310 (N_2310,N_2048,N_2149);
xor U2311 (N_2311,N_2009,N_2199);
and U2312 (N_2312,N_2048,N_2194);
or U2313 (N_2313,N_2091,N_2129);
or U2314 (N_2314,N_2124,N_2020);
nand U2315 (N_2315,N_2158,N_2182);
and U2316 (N_2316,N_2100,N_2175);
nand U2317 (N_2317,N_2050,N_2149);
and U2318 (N_2318,N_2104,N_2048);
or U2319 (N_2319,N_2150,N_2113);
nand U2320 (N_2320,N_2076,N_2018);
xor U2321 (N_2321,N_2061,N_2192);
xnor U2322 (N_2322,N_2039,N_2195);
nor U2323 (N_2323,N_2068,N_2168);
nor U2324 (N_2324,N_2038,N_2012);
nand U2325 (N_2325,N_2016,N_2184);
nand U2326 (N_2326,N_2065,N_2153);
xnor U2327 (N_2327,N_2195,N_2182);
xor U2328 (N_2328,N_2010,N_2188);
xor U2329 (N_2329,N_2110,N_2187);
and U2330 (N_2330,N_2016,N_2104);
nand U2331 (N_2331,N_2117,N_2172);
and U2332 (N_2332,N_2011,N_2074);
nor U2333 (N_2333,N_2063,N_2133);
or U2334 (N_2334,N_2029,N_2100);
nand U2335 (N_2335,N_2083,N_2105);
or U2336 (N_2336,N_2032,N_2092);
xor U2337 (N_2337,N_2198,N_2146);
xnor U2338 (N_2338,N_2115,N_2107);
xor U2339 (N_2339,N_2097,N_2077);
and U2340 (N_2340,N_2132,N_2020);
nor U2341 (N_2341,N_2171,N_2199);
nand U2342 (N_2342,N_2126,N_2000);
and U2343 (N_2343,N_2086,N_2145);
and U2344 (N_2344,N_2089,N_2066);
or U2345 (N_2345,N_2095,N_2164);
or U2346 (N_2346,N_2079,N_2085);
and U2347 (N_2347,N_2068,N_2140);
and U2348 (N_2348,N_2097,N_2176);
and U2349 (N_2349,N_2111,N_2069);
nor U2350 (N_2350,N_2019,N_2063);
xor U2351 (N_2351,N_2073,N_2176);
nor U2352 (N_2352,N_2006,N_2148);
xor U2353 (N_2353,N_2150,N_2078);
and U2354 (N_2354,N_2019,N_2008);
nand U2355 (N_2355,N_2162,N_2180);
xnor U2356 (N_2356,N_2196,N_2174);
nand U2357 (N_2357,N_2118,N_2107);
and U2358 (N_2358,N_2142,N_2139);
or U2359 (N_2359,N_2146,N_2186);
or U2360 (N_2360,N_2030,N_2141);
or U2361 (N_2361,N_2031,N_2083);
and U2362 (N_2362,N_2111,N_2164);
and U2363 (N_2363,N_2114,N_2027);
and U2364 (N_2364,N_2194,N_2046);
or U2365 (N_2365,N_2100,N_2030);
xnor U2366 (N_2366,N_2069,N_2178);
xor U2367 (N_2367,N_2068,N_2130);
nand U2368 (N_2368,N_2025,N_2135);
nor U2369 (N_2369,N_2107,N_2061);
or U2370 (N_2370,N_2101,N_2134);
nor U2371 (N_2371,N_2051,N_2136);
nand U2372 (N_2372,N_2119,N_2095);
or U2373 (N_2373,N_2102,N_2075);
nor U2374 (N_2374,N_2023,N_2196);
nand U2375 (N_2375,N_2140,N_2096);
xnor U2376 (N_2376,N_2095,N_2029);
nor U2377 (N_2377,N_2159,N_2079);
nand U2378 (N_2378,N_2016,N_2059);
xnor U2379 (N_2379,N_2145,N_2098);
nand U2380 (N_2380,N_2039,N_2100);
and U2381 (N_2381,N_2109,N_2037);
or U2382 (N_2382,N_2034,N_2102);
and U2383 (N_2383,N_2055,N_2189);
and U2384 (N_2384,N_2179,N_2010);
or U2385 (N_2385,N_2068,N_2116);
and U2386 (N_2386,N_2007,N_2045);
xnor U2387 (N_2387,N_2043,N_2115);
xor U2388 (N_2388,N_2057,N_2109);
nor U2389 (N_2389,N_2186,N_2110);
and U2390 (N_2390,N_2134,N_2129);
nand U2391 (N_2391,N_2003,N_2159);
and U2392 (N_2392,N_2149,N_2068);
xnor U2393 (N_2393,N_2132,N_2088);
xnor U2394 (N_2394,N_2055,N_2184);
and U2395 (N_2395,N_2099,N_2139);
or U2396 (N_2396,N_2161,N_2091);
xor U2397 (N_2397,N_2148,N_2074);
or U2398 (N_2398,N_2186,N_2098);
xor U2399 (N_2399,N_2193,N_2091);
nor U2400 (N_2400,N_2367,N_2230);
nand U2401 (N_2401,N_2347,N_2275);
xnor U2402 (N_2402,N_2332,N_2344);
or U2403 (N_2403,N_2290,N_2269);
or U2404 (N_2404,N_2286,N_2353);
nor U2405 (N_2405,N_2390,N_2358);
and U2406 (N_2406,N_2341,N_2233);
or U2407 (N_2407,N_2261,N_2243);
and U2408 (N_2408,N_2387,N_2299);
xnor U2409 (N_2409,N_2293,N_2316);
and U2410 (N_2410,N_2352,N_2291);
or U2411 (N_2411,N_2399,N_2264);
xor U2412 (N_2412,N_2278,N_2396);
nand U2413 (N_2413,N_2246,N_2305);
nor U2414 (N_2414,N_2254,N_2378);
nor U2415 (N_2415,N_2223,N_2279);
and U2416 (N_2416,N_2220,N_2251);
or U2417 (N_2417,N_2273,N_2292);
nand U2418 (N_2418,N_2391,N_2248);
xor U2419 (N_2419,N_2232,N_2274);
or U2420 (N_2420,N_2311,N_2349);
xor U2421 (N_2421,N_2270,N_2322);
nand U2422 (N_2422,N_2304,N_2371);
nor U2423 (N_2423,N_2268,N_2308);
xnor U2424 (N_2424,N_2361,N_2395);
nand U2425 (N_2425,N_2375,N_2242);
or U2426 (N_2426,N_2366,N_2345);
xor U2427 (N_2427,N_2348,N_2235);
and U2428 (N_2428,N_2386,N_2217);
nor U2429 (N_2429,N_2372,N_2388);
nor U2430 (N_2430,N_2309,N_2272);
nor U2431 (N_2431,N_2257,N_2357);
nor U2432 (N_2432,N_2227,N_2351);
and U2433 (N_2433,N_2258,N_2222);
nor U2434 (N_2434,N_2221,N_2207);
or U2435 (N_2435,N_2295,N_2382);
nand U2436 (N_2436,N_2225,N_2389);
nor U2437 (N_2437,N_2283,N_2383);
and U2438 (N_2438,N_2379,N_2393);
xor U2439 (N_2439,N_2206,N_2398);
nand U2440 (N_2440,N_2296,N_2219);
nor U2441 (N_2441,N_2317,N_2284);
or U2442 (N_2442,N_2218,N_2256);
and U2443 (N_2443,N_2280,N_2330);
xnor U2444 (N_2444,N_2370,N_2333);
nand U2445 (N_2445,N_2315,N_2381);
and U2446 (N_2446,N_2300,N_2240);
and U2447 (N_2447,N_2241,N_2238);
nand U2448 (N_2448,N_2329,N_2320);
nor U2449 (N_2449,N_2343,N_2369);
and U2450 (N_2450,N_2239,N_2252);
or U2451 (N_2451,N_2356,N_2323);
or U2452 (N_2452,N_2355,N_2208);
or U2453 (N_2453,N_2302,N_2215);
and U2454 (N_2454,N_2392,N_2314);
nor U2455 (N_2455,N_2237,N_2331);
nand U2456 (N_2456,N_2262,N_2337);
nor U2457 (N_2457,N_2271,N_2362);
and U2458 (N_2458,N_2212,N_2339);
xnor U2459 (N_2459,N_2267,N_2321);
xnor U2460 (N_2460,N_2319,N_2397);
and U2461 (N_2461,N_2282,N_2294);
nor U2462 (N_2462,N_2211,N_2368);
or U2463 (N_2463,N_2354,N_2377);
or U2464 (N_2464,N_2335,N_2203);
nor U2465 (N_2465,N_2340,N_2298);
nor U2466 (N_2466,N_2385,N_2285);
nand U2467 (N_2467,N_2204,N_2245);
or U2468 (N_2468,N_2205,N_2216);
nand U2469 (N_2469,N_2338,N_2310);
or U2470 (N_2470,N_2301,N_2249);
nand U2471 (N_2471,N_2328,N_2229);
nor U2472 (N_2472,N_2281,N_2307);
nand U2473 (N_2473,N_2394,N_2259);
xor U2474 (N_2474,N_2214,N_2365);
nand U2475 (N_2475,N_2376,N_2231);
nand U2476 (N_2476,N_2226,N_2334);
xor U2477 (N_2477,N_2255,N_2250);
nor U2478 (N_2478,N_2313,N_2209);
or U2479 (N_2479,N_2236,N_2303);
or U2480 (N_2480,N_2234,N_2363);
and U2481 (N_2481,N_2200,N_2380);
and U2482 (N_2482,N_2260,N_2350);
nor U2483 (N_2483,N_2228,N_2210);
and U2484 (N_2484,N_2364,N_2224);
or U2485 (N_2485,N_2244,N_2201);
nand U2486 (N_2486,N_2326,N_2247);
nor U2487 (N_2487,N_2276,N_2287);
nand U2488 (N_2488,N_2374,N_2277);
or U2489 (N_2489,N_2266,N_2312);
and U2490 (N_2490,N_2346,N_2289);
and U2491 (N_2491,N_2306,N_2373);
and U2492 (N_2492,N_2342,N_2297);
nand U2493 (N_2493,N_2359,N_2318);
and U2494 (N_2494,N_2325,N_2324);
xor U2495 (N_2495,N_2253,N_2360);
and U2496 (N_2496,N_2288,N_2336);
or U2497 (N_2497,N_2263,N_2202);
or U2498 (N_2498,N_2384,N_2327);
xnor U2499 (N_2499,N_2213,N_2265);
nor U2500 (N_2500,N_2397,N_2331);
and U2501 (N_2501,N_2257,N_2332);
or U2502 (N_2502,N_2253,N_2237);
nor U2503 (N_2503,N_2300,N_2278);
xnor U2504 (N_2504,N_2304,N_2250);
nor U2505 (N_2505,N_2241,N_2246);
nor U2506 (N_2506,N_2353,N_2241);
xor U2507 (N_2507,N_2240,N_2332);
xnor U2508 (N_2508,N_2374,N_2322);
nor U2509 (N_2509,N_2245,N_2341);
or U2510 (N_2510,N_2385,N_2387);
and U2511 (N_2511,N_2272,N_2248);
nor U2512 (N_2512,N_2358,N_2311);
and U2513 (N_2513,N_2320,N_2336);
nand U2514 (N_2514,N_2333,N_2369);
nand U2515 (N_2515,N_2369,N_2367);
xnor U2516 (N_2516,N_2255,N_2231);
nor U2517 (N_2517,N_2230,N_2312);
nand U2518 (N_2518,N_2245,N_2238);
and U2519 (N_2519,N_2363,N_2347);
xnor U2520 (N_2520,N_2220,N_2371);
nand U2521 (N_2521,N_2219,N_2376);
nand U2522 (N_2522,N_2250,N_2267);
nand U2523 (N_2523,N_2328,N_2290);
and U2524 (N_2524,N_2382,N_2320);
or U2525 (N_2525,N_2288,N_2367);
nand U2526 (N_2526,N_2307,N_2232);
or U2527 (N_2527,N_2298,N_2229);
nor U2528 (N_2528,N_2267,N_2377);
nor U2529 (N_2529,N_2226,N_2261);
and U2530 (N_2530,N_2387,N_2341);
or U2531 (N_2531,N_2299,N_2328);
nand U2532 (N_2532,N_2305,N_2263);
nor U2533 (N_2533,N_2380,N_2379);
and U2534 (N_2534,N_2209,N_2278);
nand U2535 (N_2535,N_2232,N_2316);
xor U2536 (N_2536,N_2304,N_2224);
and U2537 (N_2537,N_2243,N_2217);
xnor U2538 (N_2538,N_2287,N_2291);
or U2539 (N_2539,N_2239,N_2284);
or U2540 (N_2540,N_2211,N_2294);
and U2541 (N_2541,N_2388,N_2343);
or U2542 (N_2542,N_2218,N_2233);
and U2543 (N_2543,N_2371,N_2232);
and U2544 (N_2544,N_2386,N_2334);
nand U2545 (N_2545,N_2329,N_2250);
and U2546 (N_2546,N_2206,N_2393);
nand U2547 (N_2547,N_2374,N_2237);
xnor U2548 (N_2548,N_2243,N_2245);
xnor U2549 (N_2549,N_2265,N_2388);
or U2550 (N_2550,N_2227,N_2341);
or U2551 (N_2551,N_2393,N_2219);
or U2552 (N_2552,N_2382,N_2245);
xnor U2553 (N_2553,N_2364,N_2374);
nand U2554 (N_2554,N_2391,N_2277);
or U2555 (N_2555,N_2386,N_2206);
xor U2556 (N_2556,N_2280,N_2245);
nor U2557 (N_2557,N_2330,N_2364);
nor U2558 (N_2558,N_2397,N_2327);
or U2559 (N_2559,N_2369,N_2388);
nor U2560 (N_2560,N_2208,N_2250);
nor U2561 (N_2561,N_2372,N_2240);
and U2562 (N_2562,N_2232,N_2309);
xnor U2563 (N_2563,N_2348,N_2379);
nor U2564 (N_2564,N_2201,N_2203);
or U2565 (N_2565,N_2229,N_2297);
and U2566 (N_2566,N_2370,N_2353);
or U2567 (N_2567,N_2249,N_2211);
nand U2568 (N_2568,N_2272,N_2364);
or U2569 (N_2569,N_2337,N_2291);
nand U2570 (N_2570,N_2254,N_2313);
and U2571 (N_2571,N_2258,N_2262);
or U2572 (N_2572,N_2279,N_2258);
nand U2573 (N_2573,N_2208,N_2262);
or U2574 (N_2574,N_2315,N_2365);
or U2575 (N_2575,N_2353,N_2343);
and U2576 (N_2576,N_2236,N_2313);
xnor U2577 (N_2577,N_2262,N_2279);
nor U2578 (N_2578,N_2385,N_2212);
nand U2579 (N_2579,N_2258,N_2371);
or U2580 (N_2580,N_2222,N_2219);
xor U2581 (N_2581,N_2389,N_2379);
xnor U2582 (N_2582,N_2344,N_2372);
or U2583 (N_2583,N_2380,N_2396);
and U2584 (N_2584,N_2238,N_2326);
nor U2585 (N_2585,N_2283,N_2366);
or U2586 (N_2586,N_2373,N_2368);
xnor U2587 (N_2587,N_2298,N_2315);
or U2588 (N_2588,N_2266,N_2337);
and U2589 (N_2589,N_2327,N_2202);
and U2590 (N_2590,N_2237,N_2292);
and U2591 (N_2591,N_2225,N_2320);
or U2592 (N_2592,N_2222,N_2318);
xor U2593 (N_2593,N_2228,N_2298);
or U2594 (N_2594,N_2271,N_2227);
nor U2595 (N_2595,N_2334,N_2347);
nor U2596 (N_2596,N_2254,N_2374);
or U2597 (N_2597,N_2305,N_2361);
xnor U2598 (N_2598,N_2378,N_2263);
nand U2599 (N_2599,N_2345,N_2298);
nor U2600 (N_2600,N_2497,N_2522);
or U2601 (N_2601,N_2583,N_2424);
and U2602 (N_2602,N_2501,N_2564);
and U2603 (N_2603,N_2426,N_2535);
and U2604 (N_2604,N_2495,N_2428);
and U2605 (N_2605,N_2556,N_2576);
nor U2606 (N_2606,N_2536,N_2460);
or U2607 (N_2607,N_2485,N_2479);
or U2608 (N_2608,N_2409,N_2591);
nand U2609 (N_2609,N_2567,N_2587);
and U2610 (N_2610,N_2417,N_2425);
xor U2611 (N_2611,N_2450,N_2527);
nand U2612 (N_2612,N_2571,N_2403);
xor U2613 (N_2613,N_2490,N_2470);
xor U2614 (N_2614,N_2506,N_2480);
or U2615 (N_2615,N_2528,N_2447);
or U2616 (N_2616,N_2590,N_2458);
xnor U2617 (N_2617,N_2513,N_2469);
nand U2618 (N_2618,N_2541,N_2456);
or U2619 (N_2619,N_2415,N_2560);
xor U2620 (N_2620,N_2549,N_2525);
and U2621 (N_2621,N_2510,N_2435);
xnor U2622 (N_2622,N_2486,N_2595);
xnor U2623 (N_2623,N_2419,N_2451);
nor U2624 (N_2624,N_2531,N_2410);
or U2625 (N_2625,N_2499,N_2588);
or U2626 (N_2626,N_2577,N_2464);
or U2627 (N_2627,N_2534,N_2558);
nand U2628 (N_2628,N_2579,N_2401);
nor U2629 (N_2629,N_2438,N_2526);
or U2630 (N_2630,N_2551,N_2493);
xnor U2631 (N_2631,N_2584,N_2599);
nor U2632 (N_2632,N_2533,N_2483);
or U2633 (N_2633,N_2563,N_2440);
and U2634 (N_2634,N_2462,N_2429);
xnor U2635 (N_2635,N_2406,N_2530);
xor U2636 (N_2636,N_2523,N_2433);
and U2637 (N_2637,N_2412,N_2474);
xnor U2638 (N_2638,N_2413,N_2521);
nor U2639 (N_2639,N_2565,N_2572);
nand U2640 (N_2640,N_2466,N_2511);
xor U2641 (N_2641,N_2407,N_2524);
nand U2642 (N_2642,N_2594,N_2484);
and U2643 (N_2643,N_2503,N_2494);
xnor U2644 (N_2644,N_2538,N_2573);
nand U2645 (N_2645,N_2442,N_2491);
and U2646 (N_2646,N_2508,N_2507);
or U2647 (N_2647,N_2422,N_2547);
nor U2648 (N_2648,N_2540,N_2418);
or U2649 (N_2649,N_2585,N_2596);
or U2650 (N_2650,N_2487,N_2504);
xnor U2651 (N_2651,N_2553,N_2539);
nand U2652 (N_2652,N_2416,N_2457);
nand U2653 (N_2653,N_2562,N_2488);
xnor U2654 (N_2654,N_2465,N_2537);
nand U2655 (N_2655,N_2581,N_2446);
nor U2656 (N_2656,N_2402,N_2554);
or U2657 (N_2657,N_2498,N_2453);
nor U2658 (N_2658,N_2569,N_2589);
nor U2659 (N_2659,N_2592,N_2548);
and U2660 (N_2660,N_2542,N_2439);
or U2661 (N_2661,N_2582,N_2550);
nor U2662 (N_2662,N_2546,N_2408);
and U2663 (N_2663,N_2586,N_2515);
nor U2664 (N_2664,N_2545,N_2505);
xor U2665 (N_2665,N_2459,N_2471);
nand U2666 (N_2666,N_2489,N_2405);
nor U2667 (N_2667,N_2432,N_2492);
and U2668 (N_2668,N_2452,N_2502);
nand U2669 (N_2669,N_2404,N_2544);
and U2670 (N_2670,N_2520,N_2518);
or U2671 (N_2671,N_2580,N_2454);
and U2672 (N_2672,N_2436,N_2512);
and U2673 (N_2673,N_2461,N_2420);
nor U2674 (N_2674,N_2444,N_2568);
nand U2675 (N_2675,N_2500,N_2434);
xnor U2676 (N_2676,N_2443,N_2597);
nand U2677 (N_2677,N_2445,N_2449);
and U2678 (N_2678,N_2421,N_2575);
or U2679 (N_2679,N_2463,N_2437);
and U2680 (N_2680,N_2482,N_2543);
and U2681 (N_2681,N_2557,N_2578);
nor U2682 (N_2682,N_2517,N_2561);
xor U2683 (N_2683,N_2411,N_2555);
xor U2684 (N_2684,N_2552,N_2481);
nand U2685 (N_2685,N_2593,N_2472);
nor U2686 (N_2686,N_2414,N_2598);
nor U2687 (N_2687,N_2532,N_2467);
or U2688 (N_2688,N_2427,N_2559);
or U2689 (N_2689,N_2529,N_2476);
xor U2690 (N_2690,N_2574,N_2566);
xor U2691 (N_2691,N_2478,N_2519);
or U2692 (N_2692,N_2431,N_2448);
nor U2693 (N_2693,N_2570,N_2496);
or U2694 (N_2694,N_2475,N_2477);
nand U2695 (N_2695,N_2400,N_2441);
and U2696 (N_2696,N_2509,N_2423);
nand U2697 (N_2697,N_2516,N_2473);
nor U2698 (N_2698,N_2514,N_2455);
nand U2699 (N_2699,N_2468,N_2430);
and U2700 (N_2700,N_2408,N_2523);
and U2701 (N_2701,N_2585,N_2441);
xnor U2702 (N_2702,N_2559,N_2537);
nor U2703 (N_2703,N_2439,N_2504);
nand U2704 (N_2704,N_2541,N_2539);
or U2705 (N_2705,N_2565,N_2411);
and U2706 (N_2706,N_2587,N_2464);
nor U2707 (N_2707,N_2466,N_2468);
nor U2708 (N_2708,N_2554,N_2595);
or U2709 (N_2709,N_2432,N_2418);
or U2710 (N_2710,N_2455,N_2520);
and U2711 (N_2711,N_2592,N_2529);
or U2712 (N_2712,N_2517,N_2580);
xnor U2713 (N_2713,N_2430,N_2562);
nand U2714 (N_2714,N_2540,N_2443);
xnor U2715 (N_2715,N_2519,N_2556);
xnor U2716 (N_2716,N_2477,N_2551);
nand U2717 (N_2717,N_2511,N_2588);
xor U2718 (N_2718,N_2545,N_2580);
xor U2719 (N_2719,N_2401,N_2420);
nor U2720 (N_2720,N_2510,N_2489);
nor U2721 (N_2721,N_2492,N_2509);
and U2722 (N_2722,N_2439,N_2584);
xnor U2723 (N_2723,N_2431,N_2566);
nand U2724 (N_2724,N_2520,N_2474);
or U2725 (N_2725,N_2596,N_2520);
or U2726 (N_2726,N_2457,N_2515);
nor U2727 (N_2727,N_2569,N_2542);
xnor U2728 (N_2728,N_2545,N_2471);
or U2729 (N_2729,N_2562,N_2409);
and U2730 (N_2730,N_2408,N_2545);
xnor U2731 (N_2731,N_2593,N_2449);
nor U2732 (N_2732,N_2475,N_2501);
and U2733 (N_2733,N_2421,N_2564);
xnor U2734 (N_2734,N_2580,N_2436);
nor U2735 (N_2735,N_2502,N_2468);
nor U2736 (N_2736,N_2433,N_2444);
xor U2737 (N_2737,N_2453,N_2452);
and U2738 (N_2738,N_2561,N_2453);
nor U2739 (N_2739,N_2503,N_2518);
or U2740 (N_2740,N_2486,N_2516);
nor U2741 (N_2741,N_2535,N_2456);
xnor U2742 (N_2742,N_2557,N_2426);
xor U2743 (N_2743,N_2459,N_2499);
xnor U2744 (N_2744,N_2556,N_2456);
nand U2745 (N_2745,N_2511,N_2450);
nor U2746 (N_2746,N_2496,N_2572);
xor U2747 (N_2747,N_2443,N_2428);
or U2748 (N_2748,N_2545,N_2508);
nand U2749 (N_2749,N_2541,N_2414);
or U2750 (N_2750,N_2487,N_2597);
nand U2751 (N_2751,N_2465,N_2402);
and U2752 (N_2752,N_2461,N_2515);
xor U2753 (N_2753,N_2555,N_2561);
and U2754 (N_2754,N_2441,N_2524);
or U2755 (N_2755,N_2439,N_2451);
xor U2756 (N_2756,N_2419,N_2410);
xor U2757 (N_2757,N_2444,N_2555);
xnor U2758 (N_2758,N_2484,N_2570);
nor U2759 (N_2759,N_2568,N_2427);
xor U2760 (N_2760,N_2402,N_2577);
nand U2761 (N_2761,N_2480,N_2516);
or U2762 (N_2762,N_2490,N_2452);
nor U2763 (N_2763,N_2594,N_2465);
and U2764 (N_2764,N_2478,N_2527);
xnor U2765 (N_2765,N_2488,N_2518);
xor U2766 (N_2766,N_2432,N_2489);
or U2767 (N_2767,N_2515,N_2578);
or U2768 (N_2768,N_2480,N_2434);
nor U2769 (N_2769,N_2512,N_2401);
and U2770 (N_2770,N_2486,N_2547);
and U2771 (N_2771,N_2411,N_2448);
and U2772 (N_2772,N_2450,N_2483);
nand U2773 (N_2773,N_2409,N_2518);
nand U2774 (N_2774,N_2598,N_2503);
nor U2775 (N_2775,N_2521,N_2538);
or U2776 (N_2776,N_2403,N_2492);
xnor U2777 (N_2777,N_2494,N_2509);
xor U2778 (N_2778,N_2503,N_2400);
nor U2779 (N_2779,N_2594,N_2496);
xor U2780 (N_2780,N_2504,N_2575);
xnor U2781 (N_2781,N_2571,N_2498);
nand U2782 (N_2782,N_2437,N_2595);
or U2783 (N_2783,N_2490,N_2440);
xnor U2784 (N_2784,N_2482,N_2573);
nand U2785 (N_2785,N_2591,N_2505);
or U2786 (N_2786,N_2482,N_2440);
xor U2787 (N_2787,N_2503,N_2455);
or U2788 (N_2788,N_2572,N_2552);
xor U2789 (N_2789,N_2525,N_2474);
or U2790 (N_2790,N_2407,N_2440);
xnor U2791 (N_2791,N_2515,N_2435);
nand U2792 (N_2792,N_2422,N_2556);
nor U2793 (N_2793,N_2480,N_2592);
nand U2794 (N_2794,N_2470,N_2461);
or U2795 (N_2795,N_2426,N_2580);
xnor U2796 (N_2796,N_2565,N_2418);
nor U2797 (N_2797,N_2483,N_2493);
nand U2798 (N_2798,N_2499,N_2470);
nor U2799 (N_2799,N_2589,N_2490);
or U2800 (N_2800,N_2618,N_2722);
nand U2801 (N_2801,N_2600,N_2657);
nor U2802 (N_2802,N_2675,N_2682);
or U2803 (N_2803,N_2785,N_2711);
and U2804 (N_2804,N_2670,N_2760);
nand U2805 (N_2805,N_2639,N_2614);
xnor U2806 (N_2806,N_2681,N_2655);
nor U2807 (N_2807,N_2635,N_2611);
nor U2808 (N_2808,N_2633,N_2658);
or U2809 (N_2809,N_2673,N_2691);
and U2810 (N_2810,N_2780,N_2629);
nand U2811 (N_2811,N_2708,N_2634);
nand U2812 (N_2812,N_2701,N_2688);
nand U2813 (N_2813,N_2703,N_2757);
nand U2814 (N_2814,N_2797,N_2799);
nor U2815 (N_2815,N_2695,N_2648);
nand U2816 (N_2816,N_2781,N_2713);
xnor U2817 (N_2817,N_2630,N_2684);
or U2818 (N_2818,N_2735,N_2687);
xor U2819 (N_2819,N_2741,N_2724);
and U2820 (N_2820,N_2668,N_2750);
nor U2821 (N_2821,N_2712,N_2734);
xnor U2822 (N_2822,N_2602,N_2621);
nand U2823 (N_2823,N_2709,N_2715);
and U2824 (N_2824,N_2693,N_2702);
nor U2825 (N_2825,N_2637,N_2774);
nor U2826 (N_2826,N_2676,N_2680);
nand U2827 (N_2827,N_2798,N_2727);
or U2828 (N_2828,N_2766,N_2686);
xor U2829 (N_2829,N_2651,N_2689);
nand U2830 (N_2830,N_2776,N_2656);
nor U2831 (N_2831,N_2731,N_2640);
or U2832 (N_2832,N_2671,N_2754);
or U2833 (N_2833,N_2758,N_2787);
xnor U2834 (N_2834,N_2728,N_2643);
nand U2835 (N_2835,N_2669,N_2793);
or U2836 (N_2836,N_2733,N_2784);
nand U2837 (N_2837,N_2765,N_2606);
nor U2838 (N_2838,N_2775,N_2654);
nand U2839 (N_2839,N_2645,N_2672);
nor U2840 (N_2840,N_2663,N_2738);
nor U2841 (N_2841,N_2753,N_2725);
nand U2842 (N_2842,N_2789,N_2755);
nor U2843 (N_2843,N_2644,N_2739);
and U2844 (N_2844,N_2652,N_2636);
xor U2845 (N_2845,N_2726,N_2772);
xnor U2846 (N_2846,N_2748,N_2716);
nand U2847 (N_2847,N_2768,N_2770);
or U2848 (N_2848,N_2622,N_2746);
xor U2849 (N_2849,N_2761,N_2619);
nand U2850 (N_2850,N_2665,N_2647);
xor U2851 (N_2851,N_2661,N_2704);
xor U2852 (N_2852,N_2719,N_2723);
xnor U2853 (N_2853,N_2698,N_2777);
nor U2854 (N_2854,N_2613,N_2626);
xnor U2855 (N_2855,N_2762,N_2745);
xor U2856 (N_2856,N_2683,N_2678);
and U2857 (N_2857,N_2783,N_2740);
nand U2858 (N_2858,N_2617,N_2718);
nand U2859 (N_2859,N_2778,N_2685);
and U2860 (N_2860,N_2749,N_2608);
and U2861 (N_2861,N_2792,N_2660);
or U2862 (N_2862,N_2664,N_2641);
and U2863 (N_2863,N_2756,N_2769);
nand U2864 (N_2864,N_2659,N_2742);
nor U2865 (N_2865,N_2690,N_2627);
nor U2866 (N_2866,N_2620,N_2791);
and U2867 (N_2867,N_2638,N_2767);
or U2868 (N_2868,N_2794,N_2603);
nor U2869 (N_2869,N_2623,N_2625);
and U2870 (N_2870,N_2632,N_2649);
nor U2871 (N_2871,N_2662,N_2612);
xor U2872 (N_2872,N_2679,N_2697);
nand U2873 (N_2873,N_2710,N_2700);
xor U2874 (N_2874,N_2752,N_2790);
nor U2875 (N_2875,N_2786,N_2714);
or U2876 (N_2876,N_2694,N_2759);
xnor U2877 (N_2877,N_2705,N_2604);
xnor U2878 (N_2878,N_2751,N_2607);
or U2879 (N_2879,N_2707,N_2601);
nand U2880 (N_2880,N_2667,N_2696);
or U2881 (N_2881,N_2699,N_2610);
xor U2882 (N_2882,N_2732,N_2646);
nor U2883 (N_2883,N_2642,N_2795);
xnor U2884 (N_2884,N_2788,N_2773);
or U2885 (N_2885,N_2628,N_2706);
xor U2886 (N_2886,N_2782,N_2779);
nor U2887 (N_2887,N_2650,N_2737);
nor U2888 (N_2888,N_2631,N_2616);
nand U2889 (N_2889,N_2692,N_2674);
and U2890 (N_2890,N_2771,N_2729);
and U2891 (N_2891,N_2721,N_2666);
xor U2892 (N_2892,N_2796,N_2609);
nor U2893 (N_2893,N_2677,N_2717);
or U2894 (N_2894,N_2605,N_2736);
nand U2895 (N_2895,N_2653,N_2744);
xnor U2896 (N_2896,N_2763,N_2730);
xnor U2897 (N_2897,N_2747,N_2624);
or U2898 (N_2898,N_2743,N_2615);
nor U2899 (N_2899,N_2764,N_2720);
or U2900 (N_2900,N_2775,N_2753);
nor U2901 (N_2901,N_2750,N_2688);
xnor U2902 (N_2902,N_2624,N_2696);
nand U2903 (N_2903,N_2740,N_2717);
nand U2904 (N_2904,N_2725,N_2727);
xor U2905 (N_2905,N_2646,N_2692);
and U2906 (N_2906,N_2632,N_2761);
or U2907 (N_2907,N_2760,N_2663);
nand U2908 (N_2908,N_2728,N_2630);
xor U2909 (N_2909,N_2680,N_2776);
or U2910 (N_2910,N_2688,N_2780);
nand U2911 (N_2911,N_2735,N_2790);
nand U2912 (N_2912,N_2600,N_2620);
nor U2913 (N_2913,N_2759,N_2715);
and U2914 (N_2914,N_2648,N_2767);
nor U2915 (N_2915,N_2631,N_2713);
nand U2916 (N_2916,N_2753,N_2632);
and U2917 (N_2917,N_2674,N_2650);
nor U2918 (N_2918,N_2747,N_2648);
xor U2919 (N_2919,N_2604,N_2725);
nand U2920 (N_2920,N_2605,N_2600);
nor U2921 (N_2921,N_2610,N_2689);
and U2922 (N_2922,N_2747,N_2742);
nand U2923 (N_2923,N_2689,N_2620);
nor U2924 (N_2924,N_2739,N_2612);
and U2925 (N_2925,N_2640,N_2752);
or U2926 (N_2926,N_2677,N_2604);
or U2927 (N_2927,N_2791,N_2792);
and U2928 (N_2928,N_2637,N_2750);
nor U2929 (N_2929,N_2763,N_2792);
and U2930 (N_2930,N_2770,N_2671);
nand U2931 (N_2931,N_2668,N_2628);
and U2932 (N_2932,N_2757,N_2797);
or U2933 (N_2933,N_2791,N_2780);
or U2934 (N_2934,N_2714,N_2739);
and U2935 (N_2935,N_2696,N_2645);
and U2936 (N_2936,N_2707,N_2768);
and U2937 (N_2937,N_2764,N_2609);
and U2938 (N_2938,N_2753,N_2675);
nor U2939 (N_2939,N_2723,N_2620);
and U2940 (N_2940,N_2655,N_2743);
or U2941 (N_2941,N_2780,N_2700);
and U2942 (N_2942,N_2645,N_2735);
nand U2943 (N_2943,N_2681,N_2685);
xor U2944 (N_2944,N_2643,N_2754);
nand U2945 (N_2945,N_2781,N_2797);
nor U2946 (N_2946,N_2768,N_2674);
nor U2947 (N_2947,N_2794,N_2795);
or U2948 (N_2948,N_2784,N_2715);
nand U2949 (N_2949,N_2776,N_2780);
nor U2950 (N_2950,N_2604,N_2643);
xnor U2951 (N_2951,N_2711,N_2615);
or U2952 (N_2952,N_2790,N_2721);
xor U2953 (N_2953,N_2603,N_2724);
and U2954 (N_2954,N_2726,N_2632);
and U2955 (N_2955,N_2758,N_2669);
nor U2956 (N_2956,N_2774,N_2770);
or U2957 (N_2957,N_2763,N_2696);
nand U2958 (N_2958,N_2673,N_2729);
or U2959 (N_2959,N_2632,N_2777);
nand U2960 (N_2960,N_2603,N_2715);
xnor U2961 (N_2961,N_2664,N_2723);
or U2962 (N_2962,N_2689,N_2648);
nand U2963 (N_2963,N_2634,N_2693);
and U2964 (N_2964,N_2704,N_2646);
nand U2965 (N_2965,N_2658,N_2716);
or U2966 (N_2966,N_2631,N_2768);
xnor U2967 (N_2967,N_2744,N_2640);
xor U2968 (N_2968,N_2605,N_2701);
and U2969 (N_2969,N_2742,N_2662);
nor U2970 (N_2970,N_2625,N_2779);
and U2971 (N_2971,N_2715,N_2687);
nand U2972 (N_2972,N_2726,N_2654);
nand U2973 (N_2973,N_2798,N_2678);
or U2974 (N_2974,N_2602,N_2723);
and U2975 (N_2975,N_2623,N_2749);
and U2976 (N_2976,N_2751,N_2700);
or U2977 (N_2977,N_2691,N_2614);
nor U2978 (N_2978,N_2749,N_2719);
nand U2979 (N_2979,N_2634,N_2689);
or U2980 (N_2980,N_2625,N_2691);
or U2981 (N_2981,N_2618,N_2757);
nor U2982 (N_2982,N_2748,N_2774);
or U2983 (N_2983,N_2786,N_2611);
xnor U2984 (N_2984,N_2748,N_2750);
and U2985 (N_2985,N_2732,N_2631);
and U2986 (N_2986,N_2627,N_2797);
xor U2987 (N_2987,N_2796,N_2693);
or U2988 (N_2988,N_2684,N_2601);
and U2989 (N_2989,N_2680,N_2782);
nand U2990 (N_2990,N_2690,N_2676);
or U2991 (N_2991,N_2691,N_2768);
and U2992 (N_2992,N_2637,N_2706);
xor U2993 (N_2993,N_2724,N_2710);
xor U2994 (N_2994,N_2615,N_2706);
xor U2995 (N_2995,N_2791,N_2631);
or U2996 (N_2996,N_2759,N_2628);
xnor U2997 (N_2997,N_2621,N_2738);
xor U2998 (N_2998,N_2761,N_2661);
xor U2999 (N_2999,N_2790,N_2617);
and U3000 (N_3000,N_2859,N_2810);
and U3001 (N_3001,N_2881,N_2818);
nand U3002 (N_3002,N_2895,N_2920);
nand U3003 (N_3003,N_2955,N_2876);
nand U3004 (N_3004,N_2970,N_2861);
nand U3005 (N_3005,N_2957,N_2851);
nor U3006 (N_3006,N_2935,N_2854);
xor U3007 (N_3007,N_2944,N_2879);
nor U3008 (N_3008,N_2963,N_2969);
xnor U3009 (N_3009,N_2889,N_2880);
nand U3010 (N_3010,N_2839,N_2902);
xor U3011 (N_3011,N_2996,N_2960);
nor U3012 (N_3012,N_2932,N_2847);
or U3013 (N_3013,N_2968,N_2974);
or U3014 (N_3014,N_2983,N_2891);
or U3015 (N_3015,N_2800,N_2894);
nand U3016 (N_3016,N_2988,N_2997);
nand U3017 (N_3017,N_2975,N_2841);
or U3018 (N_3018,N_2871,N_2952);
nand U3019 (N_3019,N_2834,N_2831);
xnor U3020 (N_3020,N_2925,N_2865);
or U3021 (N_3021,N_2921,N_2907);
xnor U3022 (N_3022,N_2931,N_2805);
xnor U3023 (N_3023,N_2803,N_2977);
and U3024 (N_3024,N_2840,N_2954);
nand U3025 (N_3025,N_2832,N_2890);
or U3026 (N_3026,N_2965,N_2812);
xor U3027 (N_3027,N_2905,N_2922);
nand U3028 (N_3028,N_2815,N_2824);
xor U3029 (N_3029,N_2914,N_2936);
and U3030 (N_3030,N_2823,N_2971);
and U3031 (N_3031,N_2978,N_2918);
or U3032 (N_3032,N_2924,N_2848);
nand U3033 (N_3033,N_2951,N_2884);
or U3034 (N_3034,N_2862,N_2982);
and U3035 (N_3035,N_2844,N_2911);
and U3036 (N_3036,N_2950,N_2868);
nor U3037 (N_3037,N_2899,N_2850);
xnor U3038 (N_3038,N_2984,N_2942);
nor U3039 (N_3039,N_2973,N_2806);
nand U3040 (N_3040,N_2961,N_2927);
or U3041 (N_3041,N_2985,N_2819);
xnor U3042 (N_3042,N_2945,N_2908);
or U3043 (N_3043,N_2825,N_2919);
nor U3044 (N_3044,N_2822,N_2993);
nand U3045 (N_3045,N_2943,N_2915);
xor U3046 (N_3046,N_2941,N_2937);
xnor U3047 (N_3047,N_2949,N_2864);
nand U3048 (N_3048,N_2897,N_2933);
and U3049 (N_3049,N_2808,N_2833);
nor U3050 (N_3050,N_2888,N_2853);
and U3051 (N_3051,N_2910,N_2928);
or U3052 (N_3052,N_2959,N_2877);
xnor U3053 (N_3053,N_2867,N_2893);
nor U3054 (N_3054,N_2998,N_2842);
and U3055 (N_3055,N_2878,N_2896);
nor U3056 (N_3056,N_2870,N_2820);
xor U3057 (N_3057,N_2912,N_2938);
xnor U3058 (N_3058,N_2830,N_2883);
nand U3059 (N_3059,N_2916,N_2992);
nor U3060 (N_3060,N_2845,N_2873);
nor U3061 (N_3061,N_2940,N_2999);
nand U3062 (N_3062,N_2885,N_2837);
and U3063 (N_3063,N_2906,N_2947);
and U3064 (N_3064,N_2962,N_2882);
nor U3065 (N_3065,N_2892,N_2826);
xor U3066 (N_3066,N_2811,N_2934);
nor U3067 (N_3067,N_2948,N_2856);
xor U3068 (N_3068,N_2804,N_2900);
nor U3069 (N_3069,N_2858,N_2855);
or U3070 (N_3070,N_2958,N_2835);
and U3071 (N_3071,N_2953,N_2964);
or U3072 (N_3072,N_2986,N_2980);
xor U3073 (N_3073,N_2989,N_2990);
nor U3074 (N_3074,N_2976,N_2981);
xnor U3075 (N_3075,N_2813,N_2994);
or U3076 (N_3076,N_2860,N_2817);
or U3077 (N_3077,N_2901,N_2909);
xor U3078 (N_3078,N_2887,N_2903);
xnor U3079 (N_3079,N_2874,N_2821);
xor U3080 (N_3080,N_2966,N_2849);
nand U3081 (N_3081,N_2816,N_2946);
xor U3082 (N_3082,N_2913,N_2898);
nand U3083 (N_3083,N_2995,N_2869);
or U3084 (N_3084,N_2875,N_2972);
xor U3085 (N_3085,N_2939,N_2809);
nor U3086 (N_3086,N_2863,N_2843);
nor U3087 (N_3087,N_2987,N_2886);
nand U3088 (N_3088,N_2991,N_2866);
nand U3089 (N_3089,N_2838,N_2967);
xor U3090 (N_3090,N_2829,N_2917);
nor U3091 (N_3091,N_2814,N_2852);
nand U3092 (N_3092,N_2930,N_2828);
xor U3093 (N_3093,N_2956,N_2979);
nand U3094 (N_3094,N_2904,N_2801);
and U3095 (N_3095,N_2807,N_2923);
or U3096 (N_3096,N_2827,N_2926);
or U3097 (N_3097,N_2802,N_2857);
and U3098 (N_3098,N_2836,N_2872);
or U3099 (N_3099,N_2846,N_2929);
and U3100 (N_3100,N_2844,N_2813);
and U3101 (N_3101,N_2816,N_2834);
and U3102 (N_3102,N_2823,N_2934);
nor U3103 (N_3103,N_2898,N_2915);
nand U3104 (N_3104,N_2932,N_2824);
xnor U3105 (N_3105,N_2801,N_2873);
nand U3106 (N_3106,N_2829,N_2897);
nand U3107 (N_3107,N_2918,N_2909);
and U3108 (N_3108,N_2940,N_2820);
and U3109 (N_3109,N_2878,N_2884);
nor U3110 (N_3110,N_2965,N_2933);
or U3111 (N_3111,N_2894,N_2823);
nor U3112 (N_3112,N_2949,N_2997);
nor U3113 (N_3113,N_2969,N_2946);
nor U3114 (N_3114,N_2911,N_2821);
or U3115 (N_3115,N_2806,N_2928);
xnor U3116 (N_3116,N_2939,N_2933);
and U3117 (N_3117,N_2925,N_2944);
xor U3118 (N_3118,N_2817,N_2954);
or U3119 (N_3119,N_2838,N_2828);
nor U3120 (N_3120,N_2971,N_2949);
nor U3121 (N_3121,N_2818,N_2931);
nor U3122 (N_3122,N_2937,N_2814);
nor U3123 (N_3123,N_2988,N_2976);
xor U3124 (N_3124,N_2821,N_2814);
nand U3125 (N_3125,N_2827,N_2882);
and U3126 (N_3126,N_2838,N_2943);
or U3127 (N_3127,N_2861,N_2961);
or U3128 (N_3128,N_2928,N_2927);
nand U3129 (N_3129,N_2871,N_2972);
xor U3130 (N_3130,N_2886,N_2935);
xnor U3131 (N_3131,N_2877,N_2918);
or U3132 (N_3132,N_2880,N_2926);
xor U3133 (N_3133,N_2869,N_2864);
and U3134 (N_3134,N_2882,N_2917);
nor U3135 (N_3135,N_2924,N_2863);
and U3136 (N_3136,N_2843,N_2866);
and U3137 (N_3137,N_2967,N_2946);
nor U3138 (N_3138,N_2937,N_2834);
nand U3139 (N_3139,N_2940,N_2857);
and U3140 (N_3140,N_2854,N_2887);
nor U3141 (N_3141,N_2872,N_2972);
and U3142 (N_3142,N_2986,N_2924);
or U3143 (N_3143,N_2974,N_2907);
nor U3144 (N_3144,N_2872,N_2813);
nand U3145 (N_3145,N_2907,N_2813);
nand U3146 (N_3146,N_2922,N_2887);
or U3147 (N_3147,N_2885,N_2882);
and U3148 (N_3148,N_2935,N_2859);
xnor U3149 (N_3149,N_2886,N_2927);
or U3150 (N_3150,N_2839,N_2942);
and U3151 (N_3151,N_2890,N_2967);
and U3152 (N_3152,N_2831,N_2960);
nor U3153 (N_3153,N_2951,N_2970);
and U3154 (N_3154,N_2825,N_2953);
nand U3155 (N_3155,N_2916,N_2963);
xnor U3156 (N_3156,N_2867,N_2953);
nor U3157 (N_3157,N_2931,N_2903);
nor U3158 (N_3158,N_2918,N_2964);
xnor U3159 (N_3159,N_2809,N_2838);
or U3160 (N_3160,N_2928,N_2897);
xor U3161 (N_3161,N_2853,N_2993);
xor U3162 (N_3162,N_2999,N_2824);
nor U3163 (N_3163,N_2861,N_2925);
or U3164 (N_3164,N_2884,N_2979);
nor U3165 (N_3165,N_2901,N_2958);
or U3166 (N_3166,N_2912,N_2874);
or U3167 (N_3167,N_2867,N_2878);
xor U3168 (N_3168,N_2985,N_2835);
and U3169 (N_3169,N_2908,N_2874);
nand U3170 (N_3170,N_2889,N_2956);
nand U3171 (N_3171,N_2864,N_2835);
nor U3172 (N_3172,N_2913,N_2935);
xnor U3173 (N_3173,N_2982,N_2998);
xor U3174 (N_3174,N_2953,N_2905);
xor U3175 (N_3175,N_2879,N_2802);
nand U3176 (N_3176,N_2894,N_2918);
xnor U3177 (N_3177,N_2806,N_2877);
nor U3178 (N_3178,N_2909,N_2818);
or U3179 (N_3179,N_2802,N_2903);
or U3180 (N_3180,N_2816,N_2928);
nand U3181 (N_3181,N_2960,N_2906);
nor U3182 (N_3182,N_2997,N_2903);
and U3183 (N_3183,N_2844,N_2990);
nand U3184 (N_3184,N_2874,N_2964);
or U3185 (N_3185,N_2879,N_2969);
nor U3186 (N_3186,N_2826,N_2919);
nor U3187 (N_3187,N_2854,N_2893);
nor U3188 (N_3188,N_2994,N_2872);
nor U3189 (N_3189,N_2924,N_2903);
nor U3190 (N_3190,N_2834,N_2846);
or U3191 (N_3191,N_2891,N_2997);
or U3192 (N_3192,N_2809,N_2901);
xor U3193 (N_3193,N_2987,N_2811);
nor U3194 (N_3194,N_2943,N_2997);
nand U3195 (N_3195,N_2860,N_2808);
and U3196 (N_3196,N_2984,N_2870);
nor U3197 (N_3197,N_2931,N_2921);
nor U3198 (N_3198,N_2918,N_2896);
or U3199 (N_3199,N_2933,N_2898);
nor U3200 (N_3200,N_3110,N_3079);
nor U3201 (N_3201,N_3044,N_3074);
and U3202 (N_3202,N_3071,N_3050);
and U3203 (N_3203,N_3017,N_3016);
xnor U3204 (N_3204,N_3081,N_3197);
or U3205 (N_3205,N_3148,N_3164);
and U3206 (N_3206,N_3166,N_3128);
and U3207 (N_3207,N_3008,N_3045);
nor U3208 (N_3208,N_3133,N_3112);
and U3209 (N_3209,N_3199,N_3023);
and U3210 (N_3210,N_3090,N_3073);
xnor U3211 (N_3211,N_3134,N_3139);
and U3212 (N_3212,N_3012,N_3018);
and U3213 (N_3213,N_3025,N_3123);
nor U3214 (N_3214,N_3150,N_3097);
nor U3215 (N_3215,N_3154,N_3000);
and U3216 (N_3216,N_3046,N_3092);
xor U3217 (N_3217,N_3184,N_3019);
nor U3218 (N_3218,N_3195,N_3068);
or U3219 (N_3219,N_3189,N_3135);
xnor U3220 (N_3220,N_3014,N_3055);
nor U3221 (N_3221,N_3083,N_3084);
xor U3222 (N_3222,N_3161,N_3137);
nand U3223 (N_3223,N_3069,N_3052);
nor U3224 (N_3224,N_3051,N_3030);
xnor U3225 (N_3225,N_3113,N_3144);
nand U3226 (N_3226,N_3102,N_3104);
and U3227 (N_3227,N_3086,N_3140);
xnor U3228 (N_3228,N_3165,N_3136);
and U3229 (N_3229,N_3060,N_3070);
nand U3230 (N_3230,N_3032,N_3168);
nor U3231 (N_3231,N_3117,N_3151);
and U3232 (N_3232,N_3067,N_3088);
and U3233 (N_3233,N_3066,N_3033);
nor U3234 (N_3234,N_3127,N_3196);
xnor U3235 (N_3235,N_3167,N_3076);
xnor U3236 (N_3236,N_3173,N_3095);
xnor U3237 (N_3237,N_3034,N_3130);
or U3238 (N_3238,N_3115,N_3147);
and U3239 (N_3239,N_3036,N_3190);
and U3240 (N_3240,N_3027,N_3180);
and U3241 (N_3241,N_3061,N_3149);
or U3242 (N_3242,N_3049,N_3091);
and U3243 (N_3243,N_3125,N_3120);
or U3244 (N_3244,N_3035,N_3058);
nand U3245 (N_3245,N_3116,N_3080);
nor U3246 (N_3246,N_3157,N_3109);
xnor U3247 (N_3247,N_3169,N_3163);
nor U3248 (N_3248,N_3111,N_3022);
or U3249 (N_3249,N_3077,N_3142);
xnor U3250 (N_3250,N_3087,N_3059);
or U3251 (N_3251,N_3155,N_3124);
nor U3252 (N_3252,N_3182,N_3170);
or U3253 (N_3253,N_3054,N_3024);
xnor U3254 (N_3254,N_3099,N_3179);
nor U3255 (N_3255,N_3089,N_3021);
nand U3256 (N_3256,N_3174,N_3181);
xor U3257 (N_3257,N_3192,N_3031);
xor U3258 (N_3258,N_3043,N_3108);
nor U3259 (N_3259,N_3094,N_3039);
nor U3260 (N_3260,N_3141,N_3193);
nand U3261 (N_3261,N_3082,N_3187);
nand U3262 (N_3262,N_3106,N_3006);
or U3263 (N_3263,N_3093,N_3114);
nand U3264 (N_3264,N_3075,N_3153);
and U3265 (N_3265,N_3065,N_3096);
or U3266 (N_3266,N_3064,N_3177);
nor U3267 (N_3267,N_3146,N_3162);
nand U3268 (N_3268,N_3013,N_3103);
xor U3269 (N_3269,N_3194,N_3085);
nor U3270 (N_3270,N_3029,N_3053);
nor U3271 (N_3271,N_3118,N_3158);
nor U3272 (N_3272,N_3001,N_3188);
nor U3273 (N_3273,N_3152,N_3056);
nand U3274 (N_3274,N_3172,N_3105);
nand U3275 (N_3275,N_3185,N_3107);
nand U3276 (N_3276,N_3156,N_3057);
xor U3277 (N_3277,N_3011,N_3119);
nor U3278 (N_3278,N_3122,N_3191);
nor U3279 (N_3279,N_3132,N_3159);
and U3280 (N_3280,N_3131,N_3005);
nand U3281 (N_3281,N_3042,N_3048);
xor U3282 (N_3282,N_3072,N_3004);
nor U3283 (N_3283,N_3186,N_3121);
nor U3284 (N_3284,N_3143,N_3198);
nand U3285 (N_3285,N_3098,N_3078);
xnor U3286 (N_3286,N_3040,N_3028);
nand U3287 (N_3287,N_3007,N_3002);
xor U3288 (N_3288,N_3175,N_3183);
xor U3289 (N_3289,N_3101,N_3063);
nand U3290 (N_3290,N_3038,N_3126);
xnor U3291 (N_3291,N_3026,N_3176);
xor U3292 (N_3292,N_3009,N_3145);
xnor U3293 (N_3293,N_3062,N_3178);
and U3294 (N_3294,N_3020,N_3160);
xor U3295 (N_3295,N_3047,N_3041);
or U3296 (N_3296,N_3037,N_3171);
and U3297 (N_3297,N_3015,N_3138);
nand U3298 (N_3298,N_3003,N_3129);
and U3299 (N_3299,N_3010,N_3100);
nand U3300 (N_3300,N_3102,N_3179);
nor U3301 (N_3301,N_3179,N_3156);
or U3302 (N_3302,N_3171,N_3156);
and U3303 (N_3303,N_3089,N_3172);
nand U3304 (N_3304,N_3027,N_3144);
and U3305 (N_3305,N_3162,N_3113);
nand U3306 (N_3306,N_3180,N_3039);
nor U3307 (N_3307,N_3162,N_3063);
nand U3308 (N_3308,N_3089,N_3114);
nand U3309 (N_3309,N_3014,N_3021);
nand U3310 (N_3310,N_3177,N_3101);
nand U3311 (N_3311,N_3191,N_3139);
and U3312 (N_3312,N_3051,N_3102);
nor U3313 (N_3313,N_3182,N_3037);
and U3314 (N_3314,N_3185,N_3124);
nand U3315 (N_3315,N_3075,N_3026);
or U3316 (N_3316,N_3007,N_3094);
or U3317 (N_3317,N_3159,N_3047);
or U3318 (N_3318,N_3024,N_3050);
and U3319 (N_3319,N_3107,N_3183);
nand U3320 (N_3320,N_3104,N_3032);
nor U3321 (N_3321,N_3173,N_3042);
nor U3322 (N_3322,N_3169,N_3136);
and U3323 (N_3323,N_3014,N_3009);
nor U3324 (N_3324,N_3132,N_3145);
nor U3325 (N_3325,N_3161,N_3071);
nor U3326 (N_3326,N_3027,N_3145);
xor U3327 (N_3327,N_3107,N_3192);
and U3328 (N_3328,N_3196,N_3141);
nor U3329 (N_3329,N_3094,N_3067);
nor U3330 (N_3330,N_3009,N_3198);
or U3331 (N_3331,N_3008,N_3005);
or U3332 (N_3332,N_3038,N_3089);
xnor U3333 (N_3333,N_3073,N_3018);
xnor U3334 (N_3334,N_3104,N_3108);
or U3335 (N_3335,N_3059,N_3018);
nor U3336 (N_3336,N_3191,N_3076);
nor U3337 (N_3337,N_3160,N_3014);
and U3338 (N_3338,N_3016,N_3091);
xor U3339 (N_3339,N_3147,N_3189);
nand U3340 (N_3340,N_3144,N_3066);
or U3341 (N_3341,N_3073,N_3194);
and U3342 (N_3342,N_3035,N_3016);
xnor U3343 (N_3343,N_3103,N_3045);
xor U3344 (N_3344,N_3144,N_3112);
nand U3345 (N_3345,N_3091,N_3134);
or U3346 (N_3346,N_3054,N_3038);
nand U3347 (N_3347,N_3041,N_3018);
nand U3348 (N_3348,N_3084,N_3111);
nor U3349 (N_3349,N_3167,N_3024);
nand U3350 (N_3350,N_3127,N_3058);
nand U3351 (N_3351,N_3013,N_3094);
or U3352 (N_3352,N_3049,N_3071);
or U3353 (N_3353,N_3123,N_3164);
nor U3354 (N_3354,N_3192,N_3054);
xor U3355 (N_3355,N_3141,N_3024);
nor U3356 (N_3356,N_3142,N_3155);
or U3357 (N_3357,N_3073,N_3136);
or U3358 (N_3358,N_3137,N_3022);
nand U3359 (N_3359,N_3129,N_3124);
nand U3360 (N_3360,N_3045,N_3163);
nand U3361 (N_3361,N_3041,N_3078);
or U3362 (N_3362,N_3145,N_3125);
and U3363 (N_3363,N_3067,N_3151);
nand U3364 (N_3364,N_3012,N_3056);
nor U3365 (N_3365,N_3176,N_3061);
xnor U3366 (N_3366,N_3162,N_3084);
xnor U3367 (N_3367,N_3190,N_3010);
nand U3368 (N_3368,N_3184,N_3146);
nor U3369 (N_3369,N_3000,N_3006);
nand U3370 (N_3370,N_3067,N_3189);
xnor U3371 (N_3371,N_3142,N_3124);
xor U3372 (N_3372,N_3101,N_3038);
xor U3373 (N_3373,N_3199,N_3160);
and U3374 (N_3374,N_3087,N_3039);
xnor U3375 (N_3375,N_3151,N_3060);
xnor U3376 (N_3376,N_3177,N_3117);
nand U3377 (N_3377,N_3105,N_3157);
and U3378 (N_3378,N_3092,N_3182);
xor U3379 (N_3379,N_3118,N_3159);
and U3380 (N_3380,N_3015,N_3043);
nand U3381 (N_3381,N_3075,N_3080);
or U3382 (N_3382,N_3007,N_3167);
nand U3383 (N_3383,N_3044,N_3147);
xor U3384 (N_3384,N_3107,N_3113);
nand U3385 (N_3385,N_3176,N_3072);
nor U3386 (N_3386,N_3133,N_3044);
and U3387 (N_3387,N_3090,N_3153);
or U3388 (N_3388,N_3045,N_3019);
xor U3389 (N_3389,N_3083,N_3010);
nor U3390 (N_3390,N_3152,N_3109);
and U3391 (N_3391,N_3048,N_3166);
nor U3392 (N_3392,N_3018,N_3049);
nand U3393 (N_3393,N_3092,N_3031);
xnor U3394 (N_3394,N_3162,N_3137);
or U3395 (N_3395,N_3010,N_3113);
nor U3396 (N_3396,N_3092,N_3109);
xnor U3397 (N_3397,N_3012,N_3045);
and U3398 (N_3398,N_3134,N_3191);
nand U3399 (N_3399,N_3134,N_3051);
nor U3400 (N_3400,N_3372,N_3296);
nor U3401 (N_3401,N_3232,N_3281);
nand U3402 (N_3402,N_3378,N_3270);
nand U3403 (N_3403,N_3261,N_3208);
or U3404 (N_3404,N_3236,N_3304);
or U3405 (N_3405,N_3279,N_3379);
xor U3406 (N_3406,N_3395,N_3399);
and U3407 (N_3407,N_3329,N_3201);
xnor U3408 (N_3408,N_3357,N_3323);
xor U3409 (N_3409,N_3374,N_3202);
xor U3410 (N_3410,N_3312,N_3210);
nor U3411 (N_3411,N_3269,N_3308);
or U3412 (N_3412,N_3334,N_3206);
nand U3413 (N_3413,N_3211,N_3346);
or U3414 (N_3414,N_3386,N_3360);
nor U3415 (N_3415,N_3366,N_3248);
xor U3416 (N_3416,N_3291,N_3226);
nor U3417 (N_3417,N_3337,N_3348);
or U3418 (N_3418,N_3364,N_3382);
xnor U3419 (N_3419,N_3282,N_3349);
xor U3420 (N_3420,N_3305,N_3396);
nor U3421 (N_3421,N_3328,N_3369);
or U3422 (N_3422,N_3246,N_3322);
xor U3423 (N_3423,N_3274,N_3362);
or U3424 (N_3424,N_3326,N_3275);
nand U3425 (N_3425,N_3242,N_3373);
nor U3426 (N_3426,N_3223,N_3300);
nand U3427 (N_3427,N_3393,N_3286);
xor U3428 (N_3428,N_3257,N_3339);
and U3429 (N_3429,N_3341,N_3367);
nand U3430 (N_3430,N_3229,N_3289);
xnor U3431 (N_3431,N_3335,N_3214);
nor U3432 (N_3432,N_3240,N_3319);
nand U3433 (N_3433,N_3390,N_3306);
nand U3434 (N_3434,N_3253,N_3301);
xor U3435 (N_3435,N_3219,N_3247);
nand U3436 (N_3436,N_3287,N_3207);
nand U3437 (N_3437,N_3254,N_3200);
nand U3438 (N_3438,N_3255,N_3344);
and U3439 (N_3439,N_3316,N_3384);
or U3440 (N_3440,N_3381,N_3385);
nor U3441 (N_3441,N_3302,N_3325);
or U3442 (N_3442,N_3377,N_3350);
or U3443 (N_3443,N_3224,N_3262);
or U3444 (N_3444,N_3342,N_3370);
nand U3445 (N_3445,N_3288,N_3318);
or U3446 (N_3446,N_3388,N_3237);
or U3447 (N_3447,N_3265,N_3297);
nor U3448 (N_3448,N_3230,N_3313);
and U3449 (N_3449,N_3345,N_3397);
and U3450 (N_3450,N_3298,N_3215);
xnor U3451 (N_3451,N_3303,N_3234);
or U3452 (N_3452,N_3243,N_3310);
or U3453 (N_3453,N_3205,N_3389);
or U3454 (N_3454,N_3365,N_3343);
or U3455 (N_3455,N_3225,N_3320);
and U3456 (N_3456,N_3266,N_3212);
nand U3457 (N_3457,N_3327,N_3241);
or U3458 (N_3458,N_3259,N_3256);
and U3459 (N_3459,N_3317,N_3260);
or U3460 (N_3460,N_3292,N_3250);
nor U3461 (N_3461,N_3368,N_3371);
nand U3462 (N_3462,N_3204,N_3267);
and U3463 (N_3463,N_3280,N_3272);
nand U3464 (N_3464,N_3330,N_3340);
and U3465 (N_3465,N_3263,N_3347);
xnor U3466 (N_3466,N_3264,N_3391);
nor U3467 (N_3467,N_3249,N_3353);
nor U3468 (N_3468,N_3203,N_3380);
and U3469 (N_3469,N_3358,N_3392);
xnor U3470 (N_3470,N_3231,N_3359);
and U3471 (N_3471,N_3299,N_3277);
or U3472 (N_3472,N_3216,N_3273);
or U3473 (N_3473,N_3354,N_3235);
and U3474 (N_3474,N_3307,N_3228);
nor U3475 (N_3475,N_3375,N_3239);
or U3476 (N_3476,N_3258,N_3361);
or U3477 (N_3477,N_3271,N_3251);
and U3478 (N_3478,N_3387,N_3295);
nand U3479 (N_3479,N_3338,N_3233);
xor U3480 (N_3480,N_3209,N_3221);
or U3481 (N_3481,N_3278,N_3363);
or U3482 (N_3482,N_3398,N_3331);
xor U3483 (N_3483,N_3268,N_3227);
nor U3484 (N_3484,N_3293,N_3315);
nand U3485 (N_3485,N_3238,N_3218);
xnor U3486 (N_3486,N_3321,N_3314);
or U3487 (N_3487,N_3352,N_3332);
and U3488 (N_3488,N_3351,N_3285);
or U3489 (N_3489,N_3356,N_3333);
and U3490 (N_3490,N_3213,N_3294);
xor U3491 (N_3491,N_3244,N_3222);
xor U3492 (N_3492,N_3220,N_3284);
xor U3493 (N_3493,N_3355,N_3290);
nand U3494 (N_3494,N_3276,N_3394);
nand U3495 (N_3495,N_3383,N_3245);
or U3496 (N_3496,N_3252,N_3336);
nand U3497 (N_3497,N_3376,N_3309);
or U3498 (N_3498,N_3283,N_3324);
nand U3499 (N_3499,N_3311,N_3217);
or U3500 (N_3500,N_3248,N_3280);
nor U3501 (N_3501,N_3291,N_3380);
xnor U3502 (N_3502,N_3252,N_3334);
xnor U3503 (N_3503,N_3214,N_3396);
and U3504 (N_3504,N_3307,N_3365);
nand U3505 (N_3505,N_3309,N_3224);
and U3506 (N_3506,N_3213,N_3207);
nor U3507 (N_3507,N_3381,N_3294);
nor U3508 (N_3508,N_3315,N_3292);
nand U3509 (N_3509,N_3211,N_3286);
or U3510 (N_3510,N_3391,N_3269);
or U3511 (N_3511,N_3371,N_3272);
xor U3512 (N_3512,N_3309,N_3348);
or U3513 (N_3513,N_3375,N_3230);
xnor U3514 (N_3514,N_3312,N_3387);
or U3515 (N_3515,N_3351,N_3335);
and U3516 (N_3516,N_3399,N_3286);
nand U3517 (N_3517,N_3258,N_3233);
and U3518 (N_3518,N_3373,N_3233);
or U3519 (N_3519,N_3278,N_3315);
or U3520 (N_3520,N_3209,N_3333);
nand U3521 (N_3521,N_3358,N_3258);
nor U3522 (N_3522,N_3262,N_3259);
or U3523 (N_3523,N_3292,N_3313);
nor U3524 (N_3524,N_3276,N_3329);
and U3525 (N_3525,N_3301,N_3263);
xor U3526 (N_3526,N_3267,N_3237);
xor U3527 (N_3527,N_3275,N_3376);
or U3528 (N_3528,N_3284,N_3358);
or U3529 (N_3529,N_3396,N_3223);
nand U3530 (N_3530,N_3361,N_3295);
nor U3531 (N_3531,N_3323,N_3244);
nor U3532 (N_3532,N_3228,N_3299);
and U3533 (N_3533,N_3285,N_3316);
xor U3534 (N_3534,N_3323,N_3314);
or U3535 (N_3535,N_3291,N_3300);
and U3536 (N_3536,N_3272,N_3221);
nand U3537 (N_3537,N_3292,N_3289);
nor U3538 (N_3538,N_3215,N_3269);
and U3539 (N_3539,N_3205,N_3249);
and U3540 (N_3540,N_3301,N_3300);
or U3541 (N_3541,N_3201,N_3374);
and U3542 (N_3542,N_3203,N_3331);
nand U3543 (N_3543,N_3214,N_3227);
or U3544 (N_3544,N_3265,N_3353);
nor U3545 (N_3545,N_3310,N_3273);
xnor U3546 (N_3546,N_3253,N_3349);
or U3547 (N_3547,N_3292,N_3245);
nor U3548 (N_3548,N_3296,N_3297);
xor U3549 (N_3549,N_3264,N_3387);
xor U3550 (N_3550,N_3286,N_3361);
and U3551 (N_3551,N_3270,N_3234);
nor U3552 (N_3552,N_3364,N_3308);
or U3553 (N_3553,N_3228,N_3296);
nand U3554 (N_3554,N_3323,N_3317);
and U3555 (N_3555,N_3356,N_3338);
or U3556 (N_3556,N_3300,N_3306);
nand U3557 (N_3557,N_3395,N_3359);
or U3558 (N_3558,N_3203,N_3251);
nor U3559 (N_3559,N_3295,N_3298);
and U3560 (N_3560,N_3331,N_3309);
nand U3561 (N_3561,N_3211,N_3397);
or U3562 (N_3562,N_3375,N_3234);
nor U3563 (N_3563,N_3204,N_3202);
nand U3564 (N_3564,N_3298,N_3330);
nor U3565 (N_3565,N_3383,N_3392);
nand U3566 (N_3566,N_3398,N_3308);
xnor U3567 (N_3567,N_3215,N_3332);
or U3568 (N_3568,N_3201,N_3207);
or U3569 (N_3569,N_3260,N_3368);
and U3570 (N_3570,N_3399,N_3269);
xor U3571 (N_3571,N_3359,N_3385);
nor U3572 (N_3572,N_3289,N_3253);
nand U3573 (N_3573,N_3296,N_3232);
nor U3574 (N_3574,N_3240,N_3339);
and U3575 (N_3575,N_3250,N_3242);
and U3576 (N_3576,N_3305,N_3235);
xnor U3577 (N_3577,N_3266,N_3267);
nand U3578 (N_3578,N_3275,N_3290);
nand U3579 (N_3579,N_3379,N_3370);
and U3580 (N_3580,N_3253,N_3311);
nand U3581 (N_3581,N_3267,N_3351);
nor U3582 (N_3582,N_3271,N_3218);
nand U3583 (N_3583,N_3326,N_3377);
nand U3584 (N_3584,N_3252,N_3384);
or U3585 (N_3585,N_3267,N_3321);
xor U3586 (N_3586,N_3208,N_3321);
xor U3587 (N_3587,N_3284,N_3294);
or U3588 (N_3588,N_3266,N_3352);
xnor U3589 (N_3589,N_3343,N_3218);
nor U3590 (N_3590,N_3289,N_3203);
or U3591 (N_3591,N_3291,N_3267);
xnor U3592 (N_3592,N_3278,N_3376);
nand U3593 (N_3593,N_3390,N_3284);
or U3594 (N_3594,N_3363,N_3376);
nand U3595 (N_3595,N_3272,N_3301);
or U3596 (N_3596,N_3316,N_3271);
nor U3597 (N_3597,N_3213,N_3399);
xnor U3598 (N_3598,N_3240,N_3362);
and U3599 (N_3599,N_3255,N_3222);
nor U3600 (N_3600,N_3550,N_3448);
xor U3601 (N_3601,N_3595,N_3446);
nor U3602 (N_3602,N_3419,N_3513);
or U3603 (N_3603,N_3503,N_3599);
or U3604 (N_3604,N_3456,N_3575);
xor U3605 (N_3605,N_3413,N_3571);
nand U3606 (N_3606,N_3515,N_3493);
and U3607 (N_3607,N_3400,N_3527);
and U3608 (N_3608,N_3423,N_3586);
and U3609 (N_3609,N_3472,N_3468);
and U3610 (N_3610,N_3487,N_3430);
nand U3611 (N_3611,N_3505,N_3582);
nand U3612 (N_3612,N_3558,N_3577);
nor U3613 (N_3613,N_3408,N_3551);
nand U3614 (N_3614,N_3526,N_3480);
xor U3615 (N_3615,N_3498,N_3414);
nor U3616 (N_3616,N_3581,N_3520);
nor U3617 (N_3617,N_3445,N_3422);
xor U3618 (N_3618,N_3579,N_3417);
and U3619 (N_3619,N_3510,N_3507);
nand U3620 (N_3620,N_3403,N_3421);
nand U3621 (N_3621,N_3454,N_3467);
nand U3622 (N_3622,N_3411,N_3434);
nor U3623 (N_3623,N_3464,N_3452);
nor U3624 (N_3624,N_3590,N_3585);
nor U3625 (N_3625,N_3587,N_3431);
xnor U3626 (N_3626,N_3509,N_3502);
or U3627 (N_3627,N_3405,N_3516);
and U3628 (N_3628,N_3524,N_3598);
or U3629 (N_3629,N_3447,N_3404);
xnor U3630 (N_3630,N_3457,N_3596);
nor U3631 (N_3631,N_3436,N_3549);
xnor U3632 (N_3632,N_3574,N_3496);
nor U3633 (N_3633,N_3425,N_3578);
xor U3634 (N_3634,N_3450,N_3478);
xnor U3635 (N_3635,N_3542,N_3583);
or U3636 (N_3636,N_3554,N_3449);
nor U3637 (N_3637,N_3569,N_3566);
xnor U3638 (N_3638,N_3429,N_3428);
nor U3639 (N_3639,N_3512,N_3466);
and U3640 (N_3640,N_3552,N_3471);
nand U3641 (N_3641,N_3415,N_3420);
nor U3642 (N_3642,N_3592,N_3492);
nor U3643 (N_3643,N_3412,N_3458);
nor U3644 (N_3644,N_3546,N_3557);
nor U3645 (N_3645,N_3489,N_3561);
and U3646 (N_3646,N_3435,N_3494);
nand U3647 (N_3647,N_3532,N_3555);
xnor U3648 (N_3648,N_3534,N_3538);
and U3649 (N_3649,N_3451,N_3591);
nor U3650 (N_3650,N_3495,N_3588);
nor U3651 (N_3651,N_3402,N_3461);
or U3652 (N_3652,N_3539,N_3463);
xnor U3653 (N_3653,N_3475,N_3562);
and U3654 (N_3654,N_3584,N_3432);
nand U3655 (N_3655,N_3409,N_3514);
xnor U3656 (N_3656,N_3479,N_3427);
and U3657 (N_3657,N_3486,N_3517);
and U3658 (N_3658,N_3518,N_3544);
xor U3659 (N_3659,N_3568,N_3519);
or U3660 (N_3660,N_3504,N_3441);
nand U3661 (N_3661,N_3491,N_3473);
or U3662 (N_3662,N_3401,N_3482);
xnor U3663 (N_3663,N_3597,N_3444);
nand U3664 (N_3664,N_3476,N_3416);
nor U3665 (N_3665,N_3418,N_3469);
and U3666 (N_3666,N_3594,N_3501);
nand U3667 (N_3667,N_3474,N_3490);
and U3668 (N_3668,N_3465,N_3572);
and U3669 (N_3669,N_3523,N_3543);
xnor U3670 (N_3670,N_3508,N_3439);
and U3671 (N_3671,N_3533,N_3442);
or U3672 (N_3672,N_3426,N_3548);
or U3673 (N_3673,N_3455,N_3570);
and U3674 (N_3674,N_3481,N_3470);
and U3675 (N_3675,N_3499,N_3545);
nor U3676 (N_3676,N_3460,N_3531);
nor U3677 (N_3677,N_3540,N_3410);
xnor U3678 (N_3678,N_3440,N_3593);
and U3679 (N_3679,N_3556,N_3528);
xnor U3680 (N_3680,N_3563,N_3564);
xor U3681 (N_3681,N_3536,N_3530);
and U3682 (N_3682,N_3406,N_3559);
xor U3683 (N_3683,N_3553,N_3547);
nor U3684 (N_3684,N_3541,N_3459);
or U3685 (N_3685,N_3477,N_3453);
xor U3686 (N_3686,N_3497,N_3511);
nand U3687 (N_3687,N_3506,N_3443);
and U3688 (N_3688,N_3424,N_3407);
nor U3689 (N_3689,N_3580,N_3485);
or U3690 (N_3690,N_3483,N_3484);
nor U3691 (N_3691,N_3500,N_3438);
nor U3692 (N_3692,N_3535,N_3488);
xnor U3693 (N_3693,N_3537,N_3576);
nand U3694 (N_3694,N_3589,N_3522);
and U3695 (N_3695,N_3565,N_3529);
nor U3696 (N_3696,N_3433,N_3462);
or U3697 (N_3697,N_3573,N_3560);
and U3698 (N_3698,N_3521,N_3567);
and U3699 (N_3699,N_3437,N_3525);
nand U3700 (N_3700,N_3471,N_3400);
nand U3701 (N_3701,N_3588,N_3548);
or U3702 (N_3702,N_3519,N_3432);
and U3703 (N_3703,N_3552,N_3405);
nand U3704 (N_3704,N_3475,N_3435);
nor U3705 (N_3705,N_3567,N_3598);
nand U3706 (N_3706,N_3591,N_3404);
xnor U3707 (N_3707,N_3555,N_3473);
nand U3708 (N_3708,N_3502,N_3585);
and U3709 (N_3709,N_3595,N_3578);
and U3710 (N_3710,N_3536,N_3433);
and U3711 (N_3711,N_3418,N_3552);
or U3712 (N_3712,N_3580,N_3411);
nand U3713 (N_3713,N_3560,N_3511);
xor U3714 (N_3714,N_3529,N_3430);
nand U3715 (N_3715,N_3575,N_3578);
nor U3716 (N_3716,N_3557,N_3422);
or U3717 (N_3717,N_3524,N_3574);
or U3718 (N_3718,N_3495,N_3581);
or U3719 (N_3719,N_3411,N_3417);
nand U3720 (N_3720,N_3475,N_3511);
or U3721 (N_3721,N_3404,N_3516);
or U3722 (N_3722,N_3563,N_3546);
and U3723 (N_3723,N_3413,N_3463);
xor U3724 (N_3724,N_3482,N_3568);
or U3725 (N_3725,N_3487,N_3488);
nor U3726 (N_3726,N_3516,N_3418);
nand U3727 (N_3727,N_3574,N_3545);
and U3728 (N_3728,N_3458,N_3466);
nand U3729 (N_3729,N_3582,N_3590);
nand U3730 (N_3730,N_3495,N_3596);
nand U3731 (N_3731,N_3425,N_3527);
xnor U3732 (N_3732,N_3522,N_3537);
nand U3733 (N_3733,N_3426,N_3419);
nand U3734 (N_3734,N_3524,N_3597);
or U3735 (N_3735,N_3535,N_3528);
and U3736 (N_3736,N_3560,N_3440);
xnor U3737 (N_3737,N_3517,N_3518);
nand U3738 (N_3738,N_3597,N_3453);
or U3739 (N_3739,N_3466,N_3522);
or U3740 (N_3740,N_3512,N_3553);
xnor U3741 (N_3741,N_3507,N_3460);
xnor U3742 (N_3742,N_3456,N_3589);
xor U3743 (N_3743,N_3442,N_3494);
and U3744 (N_3744,N_3422,N_3484);
and U3745 (N_3745,N_3431,N_3439);
and U3746 (N_3746,N_3595,N_3541);
or U3747 (N_3747,N_3577,N_3565);
nand U3748 (N_3748,N_3591,N_3523);
nand U3749 (N_3749,N_3445,N_3433);
nor U3750 (N_3750,N_3415,N_3525);
and U3751 (N_3751,N_3513,N_3484);
nand U3752 (N_3752,N_3415,N_3566);
xor U3753 (N_3753,N_3599,N_3520);
and U3754 (N_3754,N_3518,N_3478);
and U3755 (N_3755,N_3431,N_3542);
nand U3756 (N_3756,N_3594,N_3516);
and U3757 (N_3757,N_3563,N_3557);
nor U3758 (N_3758,N_3463,N_3455);
nor U3759 (N_3759,N_3463,N_3490);
or U3760 (N_3760,N_3541,N_3475);
or U3761 (N_3761,N_3548,N_3488);
xor U3762 (N_3762,N_3580,N_3450);
nand U3763 (N_3763,N_3501,N_3416);
xnor U3764 (N_3764,N_3428,N_3406);
nor U3765 (N_3765,N_3569,N_3592);
or U3766 (N_3766,N_3565,N_3549);
xor U3767 (N_3767,N_3578,N_3533);
or U3768 (N_3768,N_3499,N_3523);
xnor U3769 (N_3769,N_3434,N_3465);
nor U3770 (N_3770,N_3492,N_3449);
or U3771 (N_3771,N_3554,N_3532);
and U3772 (N_3772,N_3471,N_3548);
nor U3773 (N_3773,N_3509,N_3416);
or U3774 (N_3774,N_3530,N_3513);
nor U3775 (N_3775,N_3583,N_3564);
and U3776 (N_3776,N_3566,N_3585);
or U3777 (N_3777,N_3418,N_3490);
xor U3778 (N_3778,N_3562,N_3409);
and U3779 (N_3779,N_3511,N_3575);
nor U3780 (N_3780,N_3483,N_3589);
and U3781 (N_3781,N_3584,N_3443);
or U3782 (N_3782,N_3446,N_3503);
xor U3783 (N_3783,N_3503,N_3423);
nand U3784 (N_3784,N_3518,N_3490);
nor U3785 (N_3785,N_3557,N_3574);
or U3786 (N_3786,N_3421,N_3413);
xnor U3787 (N_3787,N_3599,N_3578);
nand U3788 (N_3788,N_3574,N_3589);
nor U3789 (N_3789,N_3577,N_3520);
nand U3790 (N_3790,N_3559,N_3439);
nand U3791 (N_3791,N_3497,N_3499);
and U3792 (N_3792,N_3531,N_3407);
and U3793 (N_3793,N_3483,N_3585);
and U3794 (N_3794,N_3506,N_3541);
or U3795 (N_3795,N_3494,N_3554);
nor U3796 (N_3796,N_3475,N_3473);
and U3797 (N_3797,N_3574,N_3521);
and U3798 (N_3798,N_3407,N_3449);
xor U3799 (N_3799,N_3402,N_3408);
nand U3800 (N_3800,N_3601,N_3680);
nand U3801 (N_3801,N_3742,N_3702);
nor U3802 (N_3802,N_3765,N_3770);
nand U3803 (N_3803,N_3689,N_3690);
and U3804 (N_3804,N_3713,N_3648);
or U3805 (N_3805,N_3766,N_3686);
nand U3806 (N_3806,N_3757,N_3753);
or U3807 (N_3807,N_3692,N_3738);
nand U3808 (N_3808,N_3710,N_3661);
or U3809 (N_3809,N_3636,N_3656);
xnor U3810 (N_3810,N_3730,N_3647);
and U3811 (N_3811,N_3662,N_3634);
and U3812 (N_3812,N_3653,N_3696);
nand U3813 (N_3813,N_3651,N_3794);
xnor U3814 (N_3814,N_3673,N_3688);
nand U3815 (N_3815,N_3625,N_3623);
nand U3816 (N_3816,N_3719,N_3685);
nand U3817 (N_3817,N_3695,N_3758);
xnor U3818 (N_3818,N_3600,N_3632);
xnor U3819 (N_3819,N_3748,N_3678);
and U3820 (N_3820,N_3641,N_3752);
and U3821 (N_3821,N_3618,N_3698);
xor U3822 (N_3822,N_3603,N_3644);
nor U3823 (N_3823,N_3646,N_3792);
nand U3824 (N_3824,N_3797,N_3654);
nand U3825 (N_3825,N_3631,N_3649);
nand U3826 (N_3826,N_3708,N_3782);
and U3827 (N_3827,N_3699,N_3683);
nand U3828 (N_3828,N_3774,N_3739);
xor U3829 (N_3829,N_3743,N_3779);
nor U3830 (N_3830,N_3672,N_3640);
or U3831 (N_3831,N_3660,N_3731);
and U3832 (N_3832,N_3781,N_3620);
and U3833 (N_3833,N_3612,N_3628);
and U3834 (N_3834,N_3705,N_3772);
xnor U3835 (N_3835,N_3700,N_3609);
and U3836 (N_3836,N_3747,N_3762);
and U3837 (N_3837,N_3670,N_3751);
nor U3838 (N_3838,N_3605,N_3643);
nand U3839 (N_3839,N_3773,N_3621);
xor U3840 (N_3840,N_3733,N_3724);
nand U3841 (N_3841,N_3629,N_3637);
or U3842 (N_3842,N_3740,N_3764);
nand U3843 (N_3843,N_3606,N_3741);
or U3844 (N_3844,N_3712,N_3754);
xnor U3845 (N_3845,N_3761,N_3615);
and U3846 (N_3846,N_3775,N_3703);
and U3847 (N_3847,N_3791,N_3729);
nor U3848 (N_3848,N_3626,N_3674);
and U3849 (N_3849,N_3617,N_3650);
nor U3850 (N_3850,N_3767,N_3777);
or U3851 (N_3851,N_3796,N_3602);
or U3852 (N_3852,N_3614,N_3732);
nand U3853 (N_3853,N_3768,N_3746);
or U3854 (N_3854,N_3611,N_3671);
and U3855 (N_3855,N_3677,N_3760);
xor U3856 (N_3856,N_3622,N_3720);
nand U3857 (N_3857,N_3610,N_3667);
and U3858 (N_3858,N_3635,N_3736);
or U3859 (N_3859,N_3693,N_3676);
xnor U3860 (N_3860,N_3776,N_3607);
or U3861 (N_3861,N_3639,N_3769);
and U3862 (N_3862,N_3709,N_3799);
and U3863 (N_3863,N_3645,N_3734);
xnor U3864 (N_3864,N_3784,N_3726);
or U3865 (N_3865,N_3727,N_3679);
and U3866 (N_3866,N_3663,N_3745);
xor U3867 (N_3867,N_3707,N_3613);
nor U3868 (N_3868,N_3658,N_3785);
nand U3869 (N_3869,N_3638,N_3735);
nor U3870 (N_3870,N_3681,N_3722);
nor U3871 (N_3871,N_3659,N_3737);
and U3872 (N_3872,N_3789,N_3771);
xor U3873 (N_3873,N_3608,N_3721);
xor U3874 (N_3874,N_3604,N_3701);
xnor U3875 (N_3875,N_3763,N_3728);
and U3876 (N_3876,N_3711,N_3675);
xnor U3877 (N_3877,N_3697,N_3642);
xnor U3878 (N_3878,N_3669,N_3795);
nand U3879 (N_3879,N_3714,N_3691);
or U3880 (N_3880,N_3715,N_3633);
nor U3881 (N_3881,N_3788,N_3790);
nand U3882 (N_3882,N_3744,N_3725);
nand U3883 (N_3883,N_3787,N_3793);
nand U3884 (N_3884,N_3717,N_3780);
and U3885 (N_3885,N_3723,N_3657);
xnor U3886 (N_3886,N_3666,N_3627);
nand U3887 (N_3887,N_3665,N_3759);
and U3888 (N_3888,N_3664,N_3687);
nand U3889 (N_3889,N_3652,N_3786);
and U3890 (N_3890,N_3655,N_3756);
nor U3891 (N_3891,N_3718,N_3694);
xor U3892 (N_3892,N_3619,N_3750);
and U3893 (N_3893,N_3716,N_3684);
xor U3894 (N_3894,N_3682,N_3668);
nor U3895 (N_3895,N_3624,N_3706);
or U3896 (N_3896,N_3798,N_3783);
and U3897 (N_3897,N_3778,N_3749);
and U3898 (N_3898,N_3630,N_3755);
and U3899 (N_3899,N_3704,N_3616);
or U3900 (N_3900,N_3737,N_3731);
nand U3901 (N_3901,N_3797,N_3685);
nand U3902 (N_3902,N_3784,N_3735);
nand U3903 (N_3903,N_3789,N_3707);
and U3904 (N_3904,N_3601,N_3671);
nor U3905 (N_3905,N_3688,N_3757);
or U3906 (N_3906,N_3687,N_3765);
and U3907 (N_3907,N_3607,N_3613);
nor U3908 (N_3908,N_3700,N_3635);
xor U3909 (N_3909,N_3677,N_3792);
or U3910 (N_3910,N_3603,N_3637);
and U3911 (N_3911,N_3752,N_3724);
xor U3912 (N_3912,N_3732,N_3755);
nor U3913 (N_3913,N_3630,N_3611);
and U3914 (N_3914,N_3663,N_3708);
or U3915 (N_3915,N_3742,N_3672);
xnor U3916 (N_3916,N_3692,N_3623);
nand U3917 (N_3917,N_3712,N_3761);
nand U3918 (N_3918,N_3644,N_3771);
and U3919 (N_3919,N_3649,N_3785);
xnor U3920 (N_3920,N_3734,N_3767);
xnor U3921 (N_3921,N_3775,N_3797);
or U3922 (N_3922,N_3717,N_3671);
and U3923 (N_3923,N_3632,N_3791);
nand U3924 (N_3924,N_3616,N_3690);
or U3925 (N_3925,N_3617,N_3668);
nand U3926 (N_3926,N_3620,N_3683);
xor U3927 (N_3927,N_3661,N_3796);
nor U3928 (N_3928,N_3680,N_3735);
nor U3929 (N_3929,N_3637,N_3616);
and U3930 (N_3930,N_3719,N_3636);
and U3931 (N_3931,N_3760,N_3749);
nand U3932 (N_3932,N_3619,N_3656);
xnor U3933 (N_3933,N_3629,N_3679);
nor U3934 (N_3934,N_3656,N_3684);
and U3935 (N_3935,N_3787,N_3769);
and U3936 (N_3936,N_3601,N_3733);
nand U3937 (N_3937,N_3660,N_3785);
xor U3938 (N_3938,N_3616,N_3670);
xor U3939 (N_3939,N_3685,N_3698);
and U3940 (N_3940,N_3669,N_3653);
nand U3941 (N_3941,N_3707,N_3690);
nand U3942 (N_3942,N_3705,N_3608);
nand U3943 (N_3943,N_3622,N_3675);
and U3944 (N_3944,N_3716,N_3786);
nor U3945 (N_3945,N_3661,N_3684);
nor U3946 (N_3946,N_3706,N_3788);
nor U3947 (N_3947,N_3678,N_3696);
xnor U3948 (N_3948,N_3672,N_3631);
xnor U3949 (N_3949,N_3765,N_3648);
or U3950 (N_3950,N_3665,N_3680);
and U3951 (N_3951,N_3645,N_3634);
nand U3952 (N_3952,N_3767,N_3703);
or U3953 (N_3953,N_3656,N_3658);
xor U3954 (N_3954,N_3608,N_3659);
nor U3955 (N_3955,N_3734,N_3643);
and U3956 (N_3956,N_3759,N_3788);
xor U3957 (N_3957,N_3778,N_3787);
and U3958 (N_3958,N_3654,N_3690);
nor U3959 (N_3959,N_3747,N_3668);
nand U3960 (N_3960,N_3774,N_3652);
xor U3961 (N_3961,N_3700,N_3709);
nor U3962 (N_3962,N_3743,N_3741);
or U3963 (N_3963,N_3665,N_3781);
nor U3964 (N_3964,N_3747,N_3695);
or U3965 (N_3965,N_3758,N_3706);
xnor U3966 (N_3966,N_3686,N_3792);
xor U3967 (N_3967,N_3767,N_3670);
or U3968 (N_3968,N_3613,N_3771);
and U3969 (N_3969,N_3662,N_3724);
nor U3970 (N_3970,N_3722,N_3708);
and U3971 (N_3971,N_3712,N_3646);
and U3972 (N_3972,N_3737,N_3662);
nor U3973 (N_3973,N_3600,N_3731);
nor U3974 (N_3974,N_3717,N_3616);
nor U3975 (N_3975,N_3744,N_3606);
and U3976 (N_3976,N_3674,N_3685);
or U3977 (N_3977,N_3656,N_3756);
xnor U3978 (N_3978,N_3695,N_3764);
nand U3979 (N_3979,N_3613,N_3733);
nand U3980 (N_3980,N_3677,N_3658);
or U3981 (N_3981,N_3665,N_3651);
nand U3982 (N_3982,N_3698,N_3674);
nor U3983 (N_3983,N_3764,N_3720);
xor U3984 (N_3984,N_3600,N_3728);
nor U3985 (N_3985,N_3679,N_3774);
or U3986 (N_3986,N_3648,N_3776);
xnor U3987 (N_3987,N_3673,N_3750);
or U3988 (N_3988,N_3746,N_3765);
nand U3989 (N_3989,N_3779,N_3672);
xnor U3990 (N_3990,N_3723,N_3642);
nor U3991 (N_3991,N_3604,N_3763);
xor U3992 (N_3992,N_3660,N_3767);
nand U3993 (N_3993,N_3600,N_3663);
xnor U3994 (N_3994,N_3730,N_3676);
nand U3995 (N_3995,N_3772,N_3796);
or U3996 (N_3996,N_3729,N_3681);
or U3997 (N_3997,N_3688,N_3662);
and U3998 (N_3998,N_3695,N_3703);
and U3999 (N_3999,N_3789,N_3651);
nand U4000 (N_4000,N_3879,N_3868);
nand U4001 (N_4001,N_3820,N_3874);
nor U4002 (N_4002,N_3881,N_3830);
nand U4003 (N_4003,N_3899,N_3989);
nand U4004 (N_4004,N_3951,N_3974);
or U4005 (N_4005,N_3913,N_3884);
and U4006 (N_4006,N_3885,N_3863);
and U4007 (N_4007,N_3990,N_3897);
or U4008 (N_4008,N_3815,N_3996);
nand U4009 (N_4009,N_3889,N_3936);
nand U4010 (N_4010,N_3825,N_3845);
nor U4011 (N_4011,N_3995,N_3966);
nor U4012 (N_4012,N_3887,N_3929);
xnor U4013 (N_4013,N_3924,N_3812);
nor U4014 (N_4014,N_3838,N_3828);
or U4015 (N_4015,N_3970,N_3920);
nor U4016 (N_4016,N_3803,N_3930);
nand U4017 (N_4017,N_3864,N_3928);
xnor U4018 (N_4018,N_3903,N_3985);
or U4019 (N_4019,N_3886,N_3827);
nand U4020 (N_4020,N_3988,N_3941);
xor U4021 (N_4021,N_3923,N_3817);
nor U4022 (N_4022,N_3823,N_3905);
xor U4023 (N_4023,N_3961,N_3898);
nand U4024 (N_4024,N_3832,N_3987);
xnor U4025 (N_4025,N_3869,N_3986);
nand U4026 (N_4026,N_3939,N_3944);
nand U4027 (N_4027,N_3818,N_3833);
or U4028 (N_4028,N_3846,N_3844);
xnor U4029 (N_4029,N_3811,N_3946);
or U4030 (N_4030,N_3906,N_3964);
nor U4031 (N_4031,N_3855,N_3993);
nand U4032 (N_4032,N_3947,N_3856);
and U4033 (N_4033,N_3819,N_3822);
nand U4034 (N_4034,N_3933,N_3813);
and U4035 (N_4035,N_3859,N_3872);
xnor U4036 (N_4036,N_3962,N_3850);
nor U4037 (N_4037,N_3840,N_3942);
nand U4038 (N_4038,N_3849,N_3922);
xor U4039 (N_4039,N_3911,N_3980);
and U4040 (N_4040,N_3901,N_3925);
or U4041 (N_4041,N_3918,N_3963);
or U4042 (N_4042,N_3867,N_3978);
nor U4043 (N_4043,N_3971,N_3842);
xnor U4044 (N_4044,N_3982,N_3919);
and U4045 (N_4045,N_3955,N_3871);
xnor U4046 (N_4046,N_3998,N_3976);
and U4047 (N_4047,N_3839,N_3853);
and U4048 (N_4048,N_3894,N_3824);
xnor U4049 (N_4049,N_3940,N_3854);
nor U4050 (N_4050,N_3882,N_3893);
or U4051 (N_4051,N_3956,N_3831);
xor U4052 (N_4052,N_3862,N_3847);
and U4053 (N_4053,N_3809,N_3959);
nor U4054 (N_4054,N_3965,N_3858);
nor U4055 (N_4055,N_3915,N_3851);
and U4056 (N_4056,N_3801,N_3878);
xor U4057 (N_4057,N_3900,N_3914);
and U4058 (N_4058,N_3890,N_3904);
or U4059 (N_4059,N_3958,N_3837);
nand U4060 (N_4060,N_3852,N_3891);
xnor U4061 (N_4061,N_3960,N_3836);
or U4062 (N_4062,N_3910,N_3861);
and U4063 (N_4063,N_3848,N_3877);
xnor U4064 (N_4064,N_3957,N_3808);
nor U4065 (N_4065,N_3934,N_3949);
nand U4066 (N_4066,N_3917,N_3938);
nand U4067 (N_4067,N_3950,N_3883);
nor U4068 (N_4068,N_3948,N_3991);
nand U4069 (N_4069,N_3943,N_3841);
nand U4070 (N_4070,N_3912,N_3892);
nor U4071 (N_4071,N_3829,N_3997);
nor U4072 (N_4072,N_3865,N_3834);
nor U4073 (N_4073,N_3866,N_3807);
nand U4074 (N_4074,N_3895,N_3805);
and U4075 (N_4075,N_3870,N_3975);
or U4076 (N_4076,N_3994,N_3814);
nand U4077 (N_4077,N_3896,N_3880);
or U4078 (N_4078,N_3927,N_3908);
nand U4079 (N_4079,N_3935,N_3875);
and U4080 (N_4080,N_3902,N_3857);
or U4081 (N_4081,N_3967,N_3953);
nor U4082 (N_4082,N_3873,N_3876);
and U4083 (N_4083,N_3952,N_3954);
and U4084 (N_4084,N_3802,N_3816);
and U4085 (N_4085,N_3810,N_3888);
nand U4086 (N_4086,N_3907,N_3968);
nand U4087 (N_4087,N_3826,N_3973);
or U4088 (N_4088,N_3992,N_3969);
and U4089 (N_4089,N_3983,N_3937);
and U4090 (N_4090,N_3800,N_3979);
nor U4091 (N_4091,N_3921,N_3945);
nand U4092 (N_4092,N_3821,N_3806);
nand U4093 (N_4093,N_3981,N_3835);
nand U4094 (N_4094,N_3999,N_3916);
xor U4095 (N_4095,N_3860,N_3972);
xnor U4096 (N_4096,N_3804,N_3909);
xnor U4097 (N_4097,N_3931,N_3926);
nand U4098 (N_4098,N_3984,N_3932);
xor U4099 (N_4099,N_3843,N_3977);
or U4100 (N_4100,N_3891,N_3984);
nor U4101 (N_4101,N_3986,N_3867);
nor U4102 (N_4102,N_3918,N_3827);
and U4103 (N_4103,N_3984,N_3841);
nor U4104 (N_4104,N_3921,N_3924);
nor U4105 (N_4105,N_3978,N_3807);
nand U4106 (N_4106,N_3826,N_3807);
xnor U4107 (N_4107,N_3862,N_3884);
nand U4108 (N_4108,N_3894,N_3911);
and U4109 (N_4109,N_3840,N_3991);
or U4110 (N_4110,N_3973,N_3904);
nand U4111 (N_4111,N_3991,N_3940);
nand U4112 (N_4112,N_3960,N_3994);
or U4113 (N_4113,N_3962,N_3807);
or U4114 (N_4114,N_3985,N_3975);
xnor U4115 (N_4115,N_3930,N_3839);
or U4116 (N_4116,N_3984,N_3994);
or U4117 (N_4117,N_3994,N_3975);
or U4118 (N_4118,N_3971,N_3856);
nand U4119 (N_4119,N_3999,N_3998);
or U4120 (N_4120,N_3915,N_3968);
nor U4121 (N_4121,N_3877,N_3870);
nand U4122 (N_4122,N_3980,N_3851);
nor U4123 (N_4123,N_3929,N_3907);
xnor U4124 (N_4124,N_3817,N_3879);
nor U4125 (N_4125,N_3910,N_3998);
and U4126 (N_4126,N_3919,N_3978);
nor U4127 (N_4127,N_3836,N_3904);
nor U4128 (N_4128,N_3985,N_3851);
or U4129 (N_4129,N_3849,N_3827);
and U4130 (N_4130,N_3805,N_3973);
and U4131 (N_4131,N_3985,N_3917);
xor U4132 (N_4132,N_3963,N_3917);
nor U4133 (N_4133,N_3820,N_3818);
or U4134 (N_4134,N_3916,N_3950);
and U4135 (N_4135,N_3853,N_3983);
xnor U4136 (N_4136,N_3922,N_3861);
and U4137 (N_4137,N_3979,N_3963);
or U4138 (N_4138,N_3820,N_3862);
nand U4139 (N_4139,N_3887,N_3853);
xnor U4140 (N_4140,N_3973,N_3917);
nand U4141 (N_4141,N_3884,N_3974);
xor U4142 (N_4142,N_3831,N_3855);
and U4143 (N_4143,N_3800,N_3886);
nand U4144 (N_4144,N_3961,N_3860);
or U4145 (N_4145,N_3977,N_3955);
and U4146 (N_4146,N_3886,N_3916);
xnor U4147 (N_4147,N_3833,N_3912);
and U4148 (N_4148,N_3894,N_3990);
nand U4149 (N_4149,N_3983,N_3965);
or U4150 (N_4150,N_3922,N_3988);
and U4151 (N_4151,N_3888,N_3921);
xor U4152 (N_4152,N_3952,N_3812);
nand U4153 (N_4153,N_3980,N_3967);
nand U4154 (N_4154,N_3896,N_3878);
and U4155 (N_4155,N_3997,N_3927);
or U4156 (N_4156,N_3842,N_3972);
nand U4157 (N_4157,N_3960,N_3815);
or U4158 (N_4158,N_3936,N_3833);
nand U4159 (N_4159,N_3901,N_3952);
nor U4160 (N_4160,N_3831,N_3840);
nand U4161 (N_4161,N_3966,N_3979);
xor U4162 (N_4162,N_3821,N_3932);
nand U4163 (N_4163,N_3829,N_3862);
nand U4164 (N_4164,N_3837,N_3939);
or U4165 (N_4165,N_3969,N_3929);
or U4166 (N_4166,N_3853,N_3981);
xor U4167 (N_4167,N_3818,N_3848);
xor U4168 (N_4168,N_3918,N_3969);
and U4169 (N_4169,N_3844,N_3906);
or U4170 (N_4170,N_3964,N_3989);
nor U4171 (N_4171,N_3818,N_3876);
and U4172 (N_4172,N_3938,N_3863);
and U4173 (N_4173,N_3943,N_3894);
nor U4174 (N_4174,N_3857,N_3989);
nand U4175 (N_4175,N_3883,N_3971);
xor U4176 (N_4176,N_3921,N_3942);
or U4177 (N_4177,N_3964,N_3806);
or U4178 (N_4178,N_3977,N_3963);
or U4179 (N_4179,N_3858,N_3857);
nand U4180 (N_4180,N_3976,N_3921);
nor U4181 (N_4181,N_3975,N_3890);
xor U4182 (N_4182,N_3938,N_3840);
or U4183 (N_4183,N_3866,N_3917);
or U4184 (N_4184,N_3846,N_3971);
or U4185 (N_4185,N_3899,N_3960);
nand U4186 (N_4186,N_3808,N_3993);
nor U4187 (N_4187,N_3957,N_3965);
xor U4188 (N_4188,N_3971,N_3892);
or U4189 (N_4189,N_3995,N_3933);
and U4190 (N_4190,N_3863,N_3837);
or U4191 (N_4191,N_3806,N_3824);
nor U4192 (N_4192,N_3908,N_3978);
nand U4193 (N_4193,N_3800,N_3844);
or U4194 (N_4194,N_3849,N_3980);
nor U4195 (N_4195,N_3940,N_3892);
and U4196 (N_4196,N_3953,N_3946);
nor U4197 (N_4197,N_3944,N_3812);
nand U4198 (N_4198,N_3907,N_3909);
nand U4199 (N_4199,N_3899,N_3907);
nor U4200 (N_4200,N_4125,N_4038);
nor U4201 (N_4201,N_4165,N_4056);
xnor U4202 (N_4202,N_4115,N_4029);
and U4203 (N_4203,N_4048,N_4066);
and U4204 (N_4204,N_4105,N_4121);
nand U4205 (N_4205,N_4124,N_4016);
or U4206 (N_4206,N_4156,N_4158);
nand U4207 (N_4207,N_4193,N_4055);
or U4208 (N_4208,N_4042,N_4039);
or U4209 (N_4209,N_4112,N_4089);
nand U4210 (N_4210,N_4059,N_4192);
or U4211 (N_4211,N_4131,N_4075);
nand U4212 (N_4212,N_4147,N_4187);
nand U4213 (N_4213,N_4134,N_4129);
and U4214 (N_4214,N_4043,N_4087);
or U4215 (N_4215,N_4139,N_4122);
nand U4216 (N_4216,N_4035,N_4199);
and U4217 (N_4217,N_4138,N_4024);
and U4218 (N_4218,N_4116,N_4068);
nand U4219 (N_4219,N_4054,N_4155);
or U4220 (N_4220,N_4197,N_4164);
xnor U4221 (N_4221,N_4081,N_4007);
and U4222 (N_4222,N_4119,N_4022);
or U4223 (N_4223,N_4108,N_4065);
nor U4224 (N_4224,N_4076,N_4078);
nand U4225 (N_4225,N_4195,N_4154);
and U4226 (N_4226,N_4003,N_4041);
nor U4227 (N_4227,N_4140,N_4030);
xnor U4228 (N_4228,N_4173,N_4194);
xnor U4229 (N_4229,N_4073,N_4118);
and U4230 (N_4230,N_4153,N_4188);
nor U4231 (N_4231,N_4049,N_4053);
nor U4232 (N_4232,N_4162,N_4143);
xnor U4233 (N_4233,N_4052,N_4036);
nor U4234 (N_4234,N_4080,N_4025);
and U4235 (N_4235,N_4114,N_4109);
nand U4236 (N_4236,N_4079,N_4050);
nand U4237 (N_4237,N_4060,N_4085);
nand U4238 (N_4238,N_4058,N_4002);
and U4239 (N_4239,N_4077,N_4033);
nand U4240 (N_4240,N_4104,N_4067);
and U4241 (N_4241,N_4127,N_4142);
xor U4242 (N_4242,N_4031,N_4026);
and U4243 (N_4243,N_4006,N_4062);
and U4244 (N_4244,N_4001,N_4189);
and U4245 (N_4245,N_4009,N_4100);
nand U4246 (N_4246,N_4094,N_4175);
nor U4247 (N_4247,N_4004,N_4013);
or U4248 (N_4248,N_4017,N_4064);
xor U4249 (N_4249,N_4027,N_4099);
nand U4250 (N_4250,N_4091,N_4040);
and U4251 (N_4251,N_4137,N_4092);
nand U4252 (N_4252,N_4190,N_4180);
xnor U4253 (N_4253,N_4069,N_4120);
xnor U4254 (N_4254,N_4141,N_4185);
or U4255 (N_4255,N_4135,N_4015);
nand U4256 (N_4256,N_4051,N_4186);
nand U4257 (N_4257,N_4084,N_4191);
nand U4258 (N_4258,N_4070,N_4000);
and U4259 (N_4259,N_4161,N_4019);
nand U4260 (N_4260,N_4157,N_4133);
or U4261 (N_4261,N_4095,N_4021);
nand U4262 (N_4262,N_4166,N_4014);
nand U4263 (N_4263,N_4107,N_4088);
or U4264 (N_4264,N_4151,N_4072);
and U4265 (N_4265,N_4083,N_4093);
and U4266 (N_4266,N_4012,N_4096);
and U4267 (N_4267,N_4179,N_4123);
nor U4268 (N_4268,N_4082,N_4028);
and U4269 (N_4269,N_4150,N_4103);
nor U4270 (N_4270,N_4171,N_4005);
nor U4271 (N_4271,N_4020,N_4182);
or U4272 (N_4272,N_4198,N_4011);
or U4273 (N_4273,N_4110,N_4044);
nand U4274 (N_4274,N_4117,N_4098);
nor U4275 (N_4275,N_4167,N_4046);
and U4276 (N_4276,N_4149,N_4163);
nor U4277 (N_4277,N_4111,N_4061);
and U4278 (N_4278,N_4071,N_4063);
nor U4279 (N_4279,N_4113,N_4160);
nor U4280 (N_4280,N_4183,N_4130);
nor U4281 (N_4281,N_4132,N_4174);
nand U4282 (N_4282,N_4159,N_4037);
xnor U4283 (N_4283,N_4106,N_4010);
nand U4284 (N_4284,N_4032,N_4148);
nor U4285 (N_4285,N_4136,N_4101);
or U4286 (N_4286,N_4047,N_4181);
xor U4287 (N_4287,N_4128,N_4184);
or U4288 (N_4288,N_4086,N_4102);
nor U4289 (N_4289,N_4196,N_4176);
nand U4290 (N_4290,N_4034,N_4057);
nand U4291 (N_4291,N_4008,N_4169);
or U4292 (N_4292,N_4177,N_4018);
or U4293 (N_4293,N_4097,N_4170);
and U4294 (N_4294,N_4152,N_4172);
or U4295 (N_4295,N_4126,N_4146);
nor U4296 (N_4296,N_4045,N_4074);
or U4297 (N_4297,N_4178,N_4168);
nand U4298 (N_4298,N_4144,N_4023);
and U4299 (N_4299,N_4145,N_4090);
or U4300 (N_4300,N_4141,N_4050);
and U4301 (N_4301,N_4053,N_4056);
or U4302 (N_4302,N_4135,N_4192);
and U4303 (N_4303,N_4048,N_4005);
xor U4304 (N_4304,N_4123,N_4033);
and U4305 (N_4305,N_4086,N_4014);
and U4306 (N_4306,N_4052,N_4001);
or U4307 (N_4307,N_4061,N_4137);
nor U4308 (N_4308,N_4172,N_4137);
nand U4309 (N_4309,N_4131,N_4176);
xnor U4310 (N_4310,N_4137,N_4174);
nand U4311 (N_4311,N_4090,N_4078);
and U4312 (N_4312,N_4066,N_4173);
xnor U4313 (N_4313,N_4027,N_4134);
and U4314 (N_4314,N_4109,N_4083);
nor U4315 (N_4315,N_4029,N_4106);
and U4316 (N_4316,N_4023,N_4047);
and U4317 (N_4317,N_4190,N_4073);
xnor U4318 (N_4318,N_4095,N_4146);
or U4319 (N_4319,N_4163,N_4087);
or U4320 (N_4320,N_4177,N_4049);
or U4321 (N_4321,N_4031,N_4027);
nand U4322 (N_4322,N_4092,N_4169);
or U4323 (N_4323,N_4106,N_4072);
nor U4324 (N_4324,N_4182,N_4017);
and U4325 (N_4325,N_4109,N_4104);
nor U4326 (N_4326,N_4065,N_4002);
and U4327 (N_4327,N_4194,N_4086);
and U4328 (N_4328,N_4030,N_4065);
nor U4329 (N_4329,N_4174,N_4038);
nand U4330 (N_4330,N_4038,N_4168);
nor U4331 (N_4331,N_4113,N_4125);
nor U4332 (N_4332,N_4144,N_4021);
or U4333 (N_4333,N_4119,N_4163);
and U4334 (N_4334,N_4140,N_4120);
nand U4335 (N_4335,N_4152,N_4087);
nand U4336 (N_4336,N_4006,N_4044);
nor U4337 (N_4337,N_4061,N_4038);
nor U4338 (N_4338,N_4179,N_4063);
xor U4339 (N_4339,N_4072,N_4165);
or U4340 (N_4340,N_4093,N_4127);
nand U4341 (N_4341,N_4040,N_4154);
nand U4342 (N_4342,N_4164,N_4096);
nand U4343 (N_4343,N_4001,N_4005);
nand U4344 (N_4344,N_4178,N_4130);
and U4345 (N_4345,N_4017,N_4151);
or U4346 (N_4346,N_4118,N_4151);
or U4347 (N_4347,N_4081,N_4115);
and U4348 (N_4348,N_4057,N_4193);
and U4349 (N_4349,N_4093,N_4034);
and U4350 (N_4350,N_4026,N_4033);
nor U4351 (N_4351,N_4171,N_4023);
nand U4352 (N_4352,N_4156,N_4088);
or U4353 (N_4353,N_4175,N_4153);
xor U4354 (N_4354,N_4066,N_4006);
nor U4355 (N_4355,N_4126,N_4156);
nand U4356 (N_4356,N_4092,N_4093);
and U4357 (N_4357,N_4150,N_4117);
xnor U4358 (N_4358,N_4079,N_4195);
or U4359 (N_4359,N_4035,N_4021);
and U4360 (N_4360,N_4176,N_4097);
or U4361 (N_4361,N_4128,N_4173);
or U4362 (N_4362,N_4173,N_4181);
nor U4363 (N_4363,N_4170,N_4193);
or U4364 (N_4364,N_4087,N_4011);
nor U4365 (N_4365,N_4107,N_4037);
nor U4366 (N_4366,N_4170,N_4184);
xor U4367 (N_4367,N_4180,N_4066);
nor U4368 (N_4368,N_4095,N_4072);
nand U4369 (N_4369,N_4090,N_4198);
nand U4370 (N_4370,N_4077,N_4088);
and U4371 (N_4371,N_4192,N_4007);
nand U4372 (N_4372,N_4032,N_4077);
nand U4373 (N_4373,N_4055,N_4010);
xor U4374 (N_4374,N_4118,N_4040);
nand U4375 (N_4375,N_4007,N_4182);
or U4376 (N_4376,N_4197,N_4093);
nor U4377 (N_4377,N_4048,N_4127);
and U4378 (N_4378,N_4073,N_4043);
or U4379 (N_4379,N_4177,N_4077);
nor U4380 (N_4380,N_4054,N_4136);
and U4381 (N_4381,N_4041,N_4168);
nor U4382 (N_4382,N_4182,N_4036);
nor U4383 (N_4383,N_4143,N_4187);
nor U4384 (N_4384,N_4058,N_4019);
xor U4385 (N_4385,N_4137,N_4133);
or U4386 (N_4386,N_4097,N_4096);
nand U4387 (N_4387,N_4117,N_4162);
or U4388 (N_4388,N_4141,N_4064);
and U4389 (N_4389,N_4172,N_4066);
nor U4390 (N_4390,N_4049,N_4059);
nand U4391 (N_4391,N_4165,N_4097);
and U4392 (N_4392,N_4163,N_4190);
nor U4393 (N_4393,N_4105,N_4077);
and U4394 (N_4394,N_4073,N_4180);
xnor U4395 (N_4395,N_4009,N_4062);
or U4396 (N_4396,N_4152,N_4187);
nand U4397 (N_4397,N_4164,N_4145);
xnor U4398 (N_4398,N_4024,N_4050);
or U4399 (N_4399,N_4092,N_4051);
or U4400 (N_4400,N_4334,N_4295);
nand U4401 (N_4401,N_4373,N_4283);
or U4402 (N_4402,N_4263,N_4298);
xnor U4403 (N_4403,N_4299,N_4228);
or U4404 (N_4404,N_4211,N_4313);
and U4405 (N_4405,N_4342,N_4218);
or U4406 (N_4406,N_4396,N_4365);
and U4407 (N_4407,N_4372,N_4268);
xor U4408 (N_4408,N_4371,N_4238);
nand U4409 (N_4409,N_4336,N_4387);
and U4410 (N_4410,N_4237,N_4343);
or U4411 (N_4411,N_4226,N_4254);
xor U4412 (N_4412,N_4265,N_4269);
nand U4413 (N_4413,N_4273,N_4395);
xnor U4414 (N_4414,N_4245,N_4366);
or U4415 (N_4415,N_4370,N_4275);
nand U4416 (N_4416,N_4256,N_4291);
xor U4417 (N_4417,N_4217,N_4337);
and U4418 (N_4418,N_4352,N_4332);
nor U4419 (N_4419,N_4346,N_4288);
or U4420 (N_4420,N_4322,N_4388);
nor U4421 (N_4421,N_4392,N_4203);
nor U4422 (N_4422,N_4207,N_4351);
and U4423 (N_4423,N_4390,N_4360);
nor U4424 (N_4424,N_4213,N_4230);
nand U4425 (N_4425,N_4356,N_4227);
nand U4426 (N_4426,N_4319,N_4277);
xor U4427 (N_4427,N_4232,N_4355);
xor U4428 (N_4428,N_4308,N_4339);
or U4429 (N_4429,N_4381,N_4310);
nor U4430 (N_4430,N_4267,N_4209);
nand U4431 (N_4431,N_4311,N_4240);
xnor U4432 (N_4432,N_4353,N_4302);
nand U4433 (N_4433,N_4234,N_4278);
nor U4434 (N_4434,N_4225,N_4201);
or U4435 (N_4435,N_4297,N_4309);
nor U4436 (N_4436,N_4363,N_4222);
and U4437 (N_4437,N_4255,N_4398);
xnor U4438 (N_4438,N_4214,N_4205);
xnor U4439 (N_4439,N_4202,N_4324);
or U4440 (N_4440,N_4321,N_4210);
and U4441 (N_4441,N_4250,N_4357);
nand U4442 (N_4442,N_4304,N_4271);
or U4443 (N_4443,N_4220,N_4243);
nor U4444 (N_4444,N_4258,N_4329);
and U4445 (N_4445,N_4391,N_4362);
xnor U4446 (N_4446,N_4219,N_4385);
or U4447 (N_4447,N_4380,N_4231);
nand U4448 (N_4448,N_4374,N_4368);
and U4449 (N_4449,N_4249,N_4248);
xnor U4450 (N_4450,N_4233,N_4253);
and U4451 (N_4451,N_4316,N_4252);
or U4452 (N_4452,N_4286,N_4384);
xnor U4453 (N_4453,N_4241,N_4208);
nand U4454 (N_4454,N_4364,N_4204);
nand U4455 (N_4455,N_4383,N_4206);
nand U4456 (N_4456,N_4312,N_4200);
and U4457 (N_4457,N_4314,N_4378);
and U4458 (N_4458,N_4320,N_4260);
nor U4459 (N_4459,N_4264,N_4292);
nand U4460 (N_4460,N_4326,N_4335);
and U4461 (N_4461,N_4303,N_4257);
or U4462 (N_4462,N_4327,N_4389);
and U4463 (N_4463,N_4282,N_4284);
xnor U4464 (N_4464,N_4377,N_4330);
nand U4465 (N_4465,N_4262,N_4293);
or U4466 (N_4466,N_4239,N_4358);
nor U4467 (N_4467,N_4386,N_4305);
and U4468 (N_4468,N_4247,N_4382);
or U4469 (N_4469,N_4235,N_4266);
or U4470 (N_4470,N_4317,N_4347);
xor U4471 (N_4471,N_4333,N_4307);
or U4472 (N_4472,N_4359,N_4375);
and U4473 (N_4473,N_4300,N_4242);
nor U4474 (N_4474,N_4224,N_4394);
or U4475 (N_4475,N_4367,N_4340);
or U4476 (N_4476,N_4341,N_4285);
nand U4477 (N_4477,N_4306,N_4251);
and U4478 (N_4478,N_4246,N_4296);
nor U4479 (N_4479,N_4279,N_4348);
and U4480 (N_4480,N_4274,N_4325);
xor U4481 (N_4481,N_4354,N_4290);
nand U4482 (N_4482,N_4236,N_4215);
nand U4483 (N_4483,N_4276,N_4244);
nand U4484 (N_4484,N_4223,N_4399);
and U4485 (N_4485,N_4272,N_4259);
or U4486 (N_4486,N_4361,N_4328);
or U4487 (N_4487,N_4315,N_4229);
or U4488 (N_4488,N_4280,N_4318);
or U4489 (N_4489,N_4261,N_4281);
or U4490 (N_4490,N_4287,N_4289);
xor U4491 (N_4491,N_4338,N_4345);
nand U4492 (N_4492,N_4369,N_4212);
or U4493 (N_4493,N_4393,N_4216);
xnor U4494 (N_4494,N_4221,N_4301);
nor U4495 (N_4495,N_4323,N_4294);
and U4496 (N_4496,N_4376,N_4349);
xor U4497 (N_4497,N_4379,N_4331);
and U4498 (N_4498,N_4397,N_4350);
xor U4499 (N_4499,N_4270,N_4344);
and U4500 (N_4500,N_4289,N_4328);
nor U4501 (N_4501,N_4399,N_4335);
and U4502 (N_4502,N_4200,N_4268);
nand U4503 (N_4503,N_4313,N_4200);
and U4504 (N_4504,N_4363,N_4373);
or U4505 (N_4505,N_4379,N_4304);
and U4506 (N_4506,N_4303,N_4228);
nor U4507 (N_4507,N_4223,N_4355);
or U4508 (N_4508,N_4283,N_4260);
xor U4509 (N_4509,N_4341,N_4300);
nor U4510 (N_4510,N_4216,N_4215);
and U4511 (N_4511,N_4227,N_4354);
and U4512 (N_4512,N_4338,N_4207);
nor U4513 (N_4513,N_4374,N_4284);
xor U4514 (N_4514,N_4239,N_4234);
and U4515 (N_4515,N_4212,N_4315);
xor U4516 (N_4516,N_4243,N_4272);
or U4517 (N_4517,N_4322,N_4283);
nor U4518 (N_4518,N_4359,N_4298);
and U4519 (N_4519,N_4391,N_4209);
or U4520 (N_4520,N_4206,N_4311);
or U4521 (N_4521,N_4299,N_4333);
xor U4522 (N_4522,N_4219,N_4248);
and U4523 (N_4523,N_4232,N_4394);
nor U4524 (N_4524,N_4220,N_4370);
or U4525 (N_4525,N_4384,N_4354);
and U4526 (N_4526,N_4235,N_4317);
nand U4527 (N_4527,N_4384,N_4328);
nand U4528 (N_4528,N_4342,N_4301);
nor U4529 (N_4529,N_4224,N_4211);
nand U4530 (N_4530,N_4343,N_4278);
and U4531 (N_4531,N_4222,N_4285);
nand U4532 (N_4532,N_4350,N_4263);
nor U4533 (N_4533,N_4308,N_4335);
nand U4534 (N_4534,N_4279,N_4219);
nand U4535 (N_4535,N_4207,N_4309);
and U4536 (N_4536,N_4308,N_4218);
and U4537 (N_4537,N_4396,N_4276);
or U4538 (N_4538,N_4353,N_4387);
nand U4539 (N_4539,N_4253,N_4366);
and U4540 (N_4540,N_4276,N_4332);
xor U4541 (N_4541,N_4282,N_4321);
nand U4542 (N_4542,N_4374,N_4388);
nor U4543 (N_4543,N_4239,N_4219);
nand U4544 (N_4544,N_4370,N_4351);
or U4545 (N_4545,N_4352,N_4310);
or U4546 (N_4546,N_4307,N_4253);
nor U4547 (N_4547,N_4338,N_4313);
xnor U4548 (N_4548,N_4237,N_4362);
and U4549 (N_4549,N_4228,N_4346);
or U4550 (N_4550,N_4213,N_4375);
or U4551 (N_4551,N_4309,N_4334);
nand U4552 (N_4552,N_4384,N_4386);
nand U4553 (N_4553,N_4296,N_4281);
or U4554 (N_4554,N_4209,N_4359);
or U4555 (N_4555,N_4396,N_4362);
nand U4556 (N_4556,N_4240,N_4317);
nor U4557 (N_4557,N_4214,N_4287);
nor U4558 (N_4558,N_4272,N_4360);
nor U4559 (N_4559,N_4286,N_4283);
nor U4560 (N_4560,N_4200,N_4355);
nand U4561 (N_4561,N_4333,N_4260);
xnor U4562 (N_4562,N_4362,N_4226);
or U4563 (N_4563,N_4245,N_4242);
nor U4564 (N_4564,N_4208,N_4270);
or U4565 (N_4565,N_4372,N_4339);
or U4566 (N_4566,N_4377,N_4323);
or U4567 (N_4567,N_4284,N_4219);
nand U4568 (N_4568,N_4292,N_4374);
or U4569 (N_4569,N_4272,N_4382);
or U4570 (N_4570,N_4245,N_4224);
or U4571 (N_4571,N_4313,N_4216);
and U4572 (N_4572,N_4277,N_4286);
xor U4573 (N_4573,N_4327,N_4215);
and U4574 (N_4574,N_4339,N_4351);
nor U4575 (N_4575,N_4259,N_4314);
nand U4576 (N_4576,N_4366,N_4306);
or U4577 (N_4577,N_4306,N_4315);
xor U4578 (N_4578,N_4269,N_4239);
or U4579 (N_4579,N_4298,N_4318);
and U4580 (N_4580,N_4384,N_4391);
nand U4581 (N_4581,N_4335,N_4312);
nand U4582 (N_4582,N_4372,N_4246);
nand U4583 (N_4583,N_4347,N_4383);
xnor U4584 (N_4584,N_4353,N_4206);
xnor U4585 (N_4585,N_4203,N_4299);
and U4586 (N_4586,N_4214,N_4225);
or U4587 (N_4587,N_4218,N_4265);
or U4588 (N_4588,N_4337,N_4224);
and U4589 (N_4589,N_4260,N_4369);
or U4590 (N_4590,N_4351,N_4225);
and U4591 (N_4591,N_4334,N_4395);
and U4592 (N_4592,N_4329,N_4381);
nand U4593 (N_4593,N_4315,N_4249);
nand U4594 (N_4594,N_4394,N_4273);
nor U4595 (N_4595,N_4249,N_4245);
or U4596 (N_4596,N_4288,N_4321);
xnor U4597 (N_4597,N_4250,N_4271);
nor U4598 (N_4598,N_4275,N_4271);
and U4599 (N_4599,N_4340,N_4264);
nand U4600 (N_4600,N_4428,N_4549);
or U4601 (N_4601,N_4439,N_4499);
nor U4602 (N_4602,N_4436,N_4533);
nor U4603 (N_4603,N_4490,N_4548);
xor U4604 (N_4604,N_4554,N_4411);
or U4605 (N_4605,N_4495,N_4587);
nand U4606 (N_4606,N_4522,N_4567);
and U4607 (N_4607,N_4445,N_4486);
xor U4608 (N_4608,N_4593,N_4412);
xnor U4609 (N_4609,N_4588,N_4598);
nor U4610 (N_4610,N_4413,N_4480);
or U4611 (N_4611,N_4547,N_4418);
nand U4612 (N_4612,N_4492,N_4539);
or U4613 (N_4613,N_4468,N_4419);
xnor U4614 (N_4614,N_4556,N_4502);
nor U4615 (N_4615,N_4520,N_4550);
and U4616 (N_4616,N_4458,N_4431);
or U4617 (N_4617,N_4465,N_4576);
xnor U4618 (N_4618,N_4561,N_4526);
and U4619 (N_4619,N_4475,N_4474);
and U4620 (N_4620,N_4479,N_4463);
or U4621 (N_4621,N_4421,N_4464);
or U4622 (N_4622,N_4519,N_4569);
nand U4623 (N_4623,N_4449,N_4581);
and U4624 (N_4624,N_4437,N_4500);
nor U4625 (N_4625,N_4594,N_4555);
xnor U4626 (N_4626,N_4585,N_4531);
and U4627 (N_4627,N_4451,N_4571);
nand U4628 (N_4628,N_4400,N_4444);
nand U4629 (N_4629,N_4524,N_4510);
nand U4630 (N_4630,N_4563,N_4470);
nor U4631 (N_4631,N_4434,N_4435);
or U4632 (N_4632,N_4511,N_4586);
or U4633 (N_4633,N_4532,N_4572);
xnor U4634 (N_4634,N_4438,N_4402);
and U4635 (N_4635,N_4557,N_4409);
xor U4636 (N_4636,N_4579,N_4501);
nor U4637 (N_4637,N_4405,N_4570);
xnor U4638 (N_4638,N_4427,N_4592);
xor U4639 (N_4639,N_4469,N_4454);
or U4640 (N_4640,N_4575,N_4414);
nor U4641 (N_4641,N_4433,N_4577);
nand U4642 (N_4642,N_4583,N_4591);
nor U4643 (N_4643,N_4599,N_4462);
and U4644 (N_4644,N_4455,N_4546);
nand U4645 (N_4645,N_4597,N_4516);
nand U4646 (N_4646,N_4416,N_4565);
xor U4647 (N_4647,N_4447,N_4542);
xor U4648 (N_4648,N_4530,N_4552);
nand U4649 (N_4649,N_4426,N_4521);
nand U4650 (N_4650,N_4472,N_4494);
xnor U4651 (N_4651,N_4482,N_4568);
nor U4652 (N_4652,N_4443,N_4446);
nand U4653 (N_4653,N_4448,N_4430);
or U4654 (N_4654,N_4525,N_4545);
or U4655 (N_4655,N_4429,N_4518);
nor U4656 (N_4656,N_4489,N_4453);
and U4657 (N_4657,N_4540,N_4582);
nor U4658 (N_4658,N_4408,N_4477);
nor U4659 (N_4659,N_4459,N_4504);
nand U4660 (N_4660,N_4422,N_4578);
xnor U4661 (N_4661,N_4544,N_4415);
nor U4662 (N_4662,N_4528,N_4509);
or U4663 (N_4663,N_4589,N_4508);
xnor U4664 (N_4664,N_4467,N_4432);
and U4665 (N_4665,N_4574,N_4410);
xor U4666 (N_4666,N_4481,N_4512);
and U4667 (N_4667,N_4513,N_4441);
and U4668 (N_4668,N_4553,N_4514);
and U4669 (N_4669,N_4425,N_4590);
or U4670 (N_4670,N_4584,N_4535);
xnor U4671 (N_4671,N_4560,N_4515);
nor U4672 (N_4672,N_4476,N_4420);
xnor U4673 (N_4673,N_4493,N_4595);
or U4674 (N_4674,N_4404,N_4491);
nand U4675 (N_4675,N_4407,N_4505);
and U4676 (N_4676,N_4406,N_4506);
and U4677 (N_4677,N_4503,N_4478);
xor U4678 (N_4678,N_4564,N_4471);
nand U4679 (N_4679,N_4442,N_4517);
or U4680 (N_4680,N_4497,N_4538);
xor U4681 (N_4681,N_4541,N_4562);
nand U4682 (N_4682,N_4498,N_4483);
or U4683 (N_4683,N_4473,N_4537);
or U4684 (N_4684,N_4401,N_4485);
nand U4685 (N_4685,N_4551,N_4457);
or U4686 (N_4686,N_4461,N_4529);
and U4687 (N_4687,N_4456,N_4596);
and U4688 (N_4688,N_4534,N_4487);
or U4689 (N_4689,N_4573,N_4466);
nor U4690 (N_4690,N_4484,N_4580);
nor U4691 (N_4691,N_4566,N_4417);
or U4692 (N_4692,N_4450,N_4460);
and U4693 (N_4693,N_4488,N_4452);
xor U4694 (N_4694,N_4496,N_4403);
nand U4695 (N_4695,N_4423,N_4543);
nand U4696 (N_4696,N_4523,N_4424);
or U4697 (N_4697,N_4527,N_4440);
xnor U4698 (N_4698,N_4507,N_4536);
nand U4699 (N_4699,N_4559,N_4558);
xor U4700 (N_4700,N_4585,N_4402);
xor U4701 (N_4701,N_4466,N_4559);
xnor U4702 (N_4702,N_4510,N_4457);
nand U4703 (N_4703,N_4587,N_4429);
and U4704 (N_4704,N_4554,N_4490);
or U4705 (N_4705,N_4466,N_4404);
or U4706 (N_4706,N_4479,N_4582);
nor U4707 (N_4707,N_4407,N_4441);
nand U4708 (N_4708,N_4405,N_4545);
nand U4709 (N_4709,N_4520,N_4542);
xor U4710 (N_4710,N_4465,N_4531);
and U4711 (N_4711,N_4508,N_4421);
xnor U4712 (N_4712,N_4403,N_4489);
nor U4713 (N_4713,N_4479,N_4543);
and U4714 (N_4714,N_4475,N_4476);
or U4715 (N_4715,N_4445,N_4515);
nor U4716 (N_4716,N_4587,N_4453);
or U4717 (N_4717,N_4506,N_4599);
nand U4718 (N_4718,N_4462,N_4568);
and U4719 (N_4719,N_4490,N_4491);
or U4720 (N_4720,N_4452,N_4461);
nor U4721 (N_4721,N_4554,N_4593);
and U4722 (N_4722,N_4549,N_4526);
or U4723 (N_4723,N_4479,N_4573);
nor U4724 (N_4724,N_4576,N_4571);
and U4725 (N_4725,N_4426,N_4462);
xor U4726 (N_4726,N_4405,N_4546);
nor U4727 (N_4727,N_4408,N_4526);
and U4728 (N_4728,N_4450,N_4464);
xnor U4729 (N_4729,N_4462,N_4566);
or U4730 (N_4730,N_4410,N_4414);
xnor U4731 (N_4731,N_4568,N_4471);
xor U4732 (N_4732,N_4577,N_4497);
and U4733 (N_4733,N_4534,N_4462);
nand U4734 (N_4734,N_4449,N_4572);
nand U4735 (N_4735,N_4498,N_4464);
xor U4736 (N_4736,N_4582,N_4556);
and U4737 (N_4737,N_4407,N_4577);
xnor U4738 (N_4738,N_4532,N_4534);
or U4739 (N_4739,N_4489,N_4470);
or U4740 (N_4740,N_4467,N_4597);
nand U4741 (N_4741,N_4492,N_4589);
and U4742 (N_4742,N_4445,N_4481);
and U4743 (N_4743,N_4420,N_4579);
xnor U4744 (N_4744,N_4436,N_4474);
nor U4745 (N_4745,N_4557,N_4545);
nor U4746 (N_4746,N_4583,N_4490);
or U4747 (N_4747,N_4552,N_4443);
nor U4748 (N_4748,N_4597,N_4598);
nor U4749 (N_4749,N_4449,N_4514);
nor U4750 (N_4750,N_4570,N_4597);
or U4751 (N_4751,N_4582,N_4532);
or U4752 (N_4752,N_4419,N_4522);
xnor U4753 (N_4753,N_4442,N_4526);
nor U4754 (N_4754,N_4530,N_4500);
xor U4755 (N_4755,N_4566,N_4483);
xor U4756 (N_4756,N_4551,N_4532);
xnor U4757 (N_4757,N_4521,N_4491);
and U4758 (N_4758,N_4524,N_4578);
nor U4759 (N_4759,N_4520,N_4586);
nor U4760 (N_4760,N_4420,N_4442);
nand U4761 (N_4761,N_4436,N_4493);
or U4762 (N_4762,N_4430,N_4416);
and U4763 (N_4763,N_4564,N_4545);
xor U4764 (N_4764,N_4403,N_4539);
xnor U4765 (N_4765,N_4566,N_4484);
nor U4766 (N_4766,N_4440,N_4410);
or U4767 (N_4767,N_4421,N_4546);
or U4768 (N_4768,N_4556,N_4480);
and U4769 (N_4769,N_4595,N_4547);
xor U4770 (N_4770,N_4434,N_4532);
and U4771 (N_4771,N_4482,N_4477);
nor U4772 (N_4772,N_4588,N_4550);
nand U4773 (N_4773,N_4421,N_4409);
nor U4774 (N_4774,N_4522,N_4424);
nor U4775 (N_4775,N_4445,N_4439);
or U4776 (N_4776,N_4502,N_4523);
nand U4777 (N_4777,N_4533,N_4591);
and U4778 (N_4778,N_4559,N_4496);
or U4779 (N_4779,N_4524,N_4550);
nor U4780 (N_4780,N_4549,N_4518);
xor U4781 (N_4781,N_4505,N_4530);
xnor U4782 (N_4782,N_4494,N_4581);
nand U4783 (N_4783,N_4513,N_4477);
nand U4784 (N_4784,N_4476,N_4536);
xor U4785 (N_4785,N_4523,N_4412);
or U4786 (N_4786,N_4450,N_4588);
and U4787 (N_4787,N_4580,N_4532);
nor U4788 (N_4788,N_4452,N_4411);
nor U4789 (N_4789,N_4599,N_4513);
nor U4790 (N_4790,N_4509,N_4576);
nor U4791 (N_4791,N_4573,N_4408);
xor U4792 (N_4792,N_4455,N_4451);
nand U4793 (N_4793,N_4580,N_4488);
xnor U4794 (N_4794,N_4501,N_4435);
xor U4795 (N_4795,N_4400,N_4506);
nor U4796 (N_4796,N_4499,N_4560);
and U4797 (N_4797,N_4422,N_4513);
nor U4798 (N_4798,N_4507,N_4477);
nor U4799 (N_4799,N_4521,N_4524);
nand U4800 (N_4800,N_4751,N_4772);
or U4801 (N_4801,N_4671,N_4764);
or U4802 (N_4802,N_4778,N_4741);
nor U4803 (N_4803,N_4626,N_4674);
and U4804 (N_4804,N_4783,N_4684);
nor U4805 (N_4805,N_4766,N_4683);
or U4806 (N_4806,N_4750,N_4738);
xnor U4807 (N_4807,N_4619,N_4655);
or U4808 (N_4808,N_4730,N_4668);
xnor U4809 (N_4809,N_4678,N_4698);
or U4810 (N_4810,N_4727,N_4679);
nand U4811 (N_4811,N_4696,N_4664);
nor U4812 (N_4812,N_4606,N_4615);
xnor U4813 (N_4813,N_4616,N_4692);
nand U4814 (N_4814,N_4700,N_4737);
xnor U4815 (N_4815,N_4601,N_4748);
nand U4816 (N_4816,N_4602,N_4680);
nand U4817 (N_4817,N_4688,N_4682);
xnor U4818 (N_4818,N_4621,N_4780);
nor U4819 (N_4819,N_4786,N_4745);
and U4820 (N_4820,N_4650,N_4790);
or U4821 (N_4821,N_4732,N_4627);
nand U4822 (N_4822,N_4793,N_4765);
xnor U4823 (N_4823,N_4726,N_4755);
xor U4824 (N_4824,N_4670,N_4695);
nand U4825 (N_4825,N_4631,N_4705);
nor U4826 (N_4826,N_4760,N_4753);
nor U4827 (N_4827,N_4667,N_4762);
nand U4828 (N_4828,N_4771,N_4623);
nand U4829 (N_4829,N_4644,N_4769);
nand U4830 (N_4830,N_4697,N_4653);
and U4831 (N_4831,N_4743,N_4673);
xnor U4832 (N_4832,N_4747,N_4716);
nand U4833 (N_4833,N_4740,N_4687);
and U4834 (N_4834,N_4691,N_4656);
xor U4835 (N_4835,N_4624,N_4686);
nand U4836 (N_4836,N_4757,N_4767);
nand U4837 (N_4837,N_4622,N_4669);
and U4838 (N_4838,N_4699,N_4675);
xnor U4839 (N_4839,N_4643,N_4611);
xor U4840 (N_4840,N_4648,N_4792);
xor U4841 (N_4841,N_4702,N_4666);
or U4842 (N_4842,N_4709,N_4756);
and U4843 (N_4843,N_4718,N_4629);
xor U4844 (N_4844,N_4662,N_4710);
and U4845 (N_4845,N_4725,N_4749);
or U4846 (N_4846,N_4768,N_4693);
or U4847 (N_4847,N_4609,N_4652);
xor U4848 (N_4848,N_4647,N_4707);
nand U4849 (N_4849,N_4719,N_4633);
xor U4850 (N_4850,N_4681,N_4798);
and U4851 (N_4851,N_4605,N_4796);
nand U4852 (N_4852,N_4638,N_4713);
nor U4853 (N_4853,N_4723,N_4781);
nand U4854 (N_4854,N_4636,N_4720);
xnor U4855 (N_4855,N_4690,N_4775);
or U4856 (N_4856,N_4618,N_4677);
and U4857 (N_4857,N_4722,N_4714);
and U4858 (N_4858,N_4608,N_4657);
nor U4859 (N_4859,N_4788,N_4641);
or U4860 (N_4860,N_4761,N_4637);
and U4861 (N_4861,N_4773,N_4782);
xnor U4862 (N_4862,N_4779,N_4704);
xnor U4863 (N_4863,N_4676,N_4607);
xnor U4864 (N_4864,N_4685,N_4752);
nand U4865 (N_4865,N_4634,N_4735);
or U4866 (N_4866,N_4632,N_4784);
nand U4867 (N_4867,N_4712,N_4724);
nand U4868 (N_4868,N_4642,N_4658);
and U4869 (N_4869,N_4785,N_4787);
nand U4870 (N_4870,N_4654,N_4663);
or U4871 (N_4871,N_4731,N_4661);
or U4872 (N_4872,N_4739,N_4717);
nor U4873 (N_4873,N_4614,N_4703);
nor U4874 (N_4874,N_4728,N_4721);
or U4875 (N_4875,N_4746,N_4799);
or U4876 (N_4876,N_4776,N_4635);
nand U4877 (N_4877,N_4742,N_4649);
and U4878 (N_4878,N_4612,N_4600);
xor U4879 (N_4879,N_4603,N_4645);
nor U4880 (N_4880,N_4770,N_4660);
or U4881 (N_4881,N_4689,N_4789);
and U4882 (N_4882,N_4754,N_4758);
and U4883 (N_4883,N_4706,N_4744);
or U4884 (N_4884,N_4639,N_4795);
and U4885 (N_4885,N_4617,N_4763);
or U4886 (N_4886,N_4777,N_4794);
xor U4887 (N_4887,N_4797,N_4672);
or U4888 (N_4888,N_4651,N_4774);
xnor U4889 (N_4889,N_4610,N_4701);
nor U4890 (N_4890,N_4630,N_4736);
nand U4891 (N_4891,N_4708,N_4659);
nand U4892 (N_4892,N_4694,N_4665);
nand U4893 (N_4893,N_4734,N_4613);
nand U4894 (N_4894,N_4733,N_4759);
or U4895 (N_4895,N_4625,N_4640);
nand U4896 (N_4896,N_4791,N_4729);
nand U4897 (N_4897,N_4711,N_4628);
xnor U4898 (N_4898,N_4715,N_4620);
or U4899 (N_4899,N_4604,N_4646);
or U4900 (N_4900,N_4749,N_4727);
or U4901 (N_4901,N_4612,N_4637);
nand U4902 (N_4902,N_4780,N_4601);
and U4903 (N_4903,N_4729,N_4670);
nand U4904 (N_4904,N_4678,N_4716);
and U4905 (N_4905,N_4786,N_4702);
or U4906 (N_4906,N_4625,N_4609);
nor U4907 (N_4907,N_4778,N_4739);
and U4908 (N_4908,N_4658,N_4647);
xor U4909 (N_4909,N_4606,N_4694);
nor U4910 (N_4910,N_4783,N_4695);
nor U4911 (N_4911,N_4626,N_4607);
nand U4912 (N_4912,N_4663,N_4622);
or U4913 (N_4913,N_4756,N_4748);
xor U4914 (N_4914,N_4642,N_4620);
or U4915 (N_4915,N_4789,N_4613);
and U4916 (N_4916,N_4607,N_4638);
xnor U4917 (N_4917,N_4661,N_4771);
nand U4918 (N_4918,N_4660,N_4687);
nor U4919 (N_4919,N_4700,N_4793);
nand U4920 (N_4920,N_4715,N_4651);
nand U4921 (N_4921,N_4702,N_4685);
and U4922 (N_4922,N_4625,N_4661);
and U4923 (N_4923,N_4722,N_4639);
or U4924 (N_4924,N_4744,N_4713);
or U4925 (N_4925,N_4752,N_4603);
nand U4926 (N_4926,N_4615,N_4688);
and U4927 (N_4927,N_4758,N_4624);
and U4928 (N_4928,N_4795,N_4645);
and U4929 (N_4929,N_4645,N_4654);
nor U4930 (N_4930,N_4740,N_4680);
nand U4931 (N_4931,N_4681,N_4704);
or U4932 (N_4932,N_4796,N_4693);
nor U4933 (N_4933,N_4737,N_4617);
or U4934 (N_4934,N_4772,N_4659);
or U4935 (N_4935,N_4633,N_4750);
or U4936 (N_4936,N_4739,N_4738);
nor U4937 (N_4937,N_4773,N_4647);
or U4938 (N_4938,N_4738,N_4778);
and U4939 (N_4939,N_4608,N_4669);
xnor U4940 (N_4940,N_4688,N_4774);
nand U4941 (N_4941,N_4712,N_4780);
xor U4942 (N_4942,N_4704,N_4705);
nor U4943 (N_4943,N_4653,N_4675);
xor U4944 (N_4944,N_4673,N_4612);
or U4945 (N_4945,N_4605,N_4787);
or U4946 (N_4946,N_4761,N_4712);
xnor U4947 (N_4947,N_4741,N_4752);
nor U4948 (N_4948,N_4604,N_4734);
or U4949 (N_4949,N_4651,N_4661);
and U4950 (N_4950,N_4700,N_4763);
or U4951 (N_4951,N_4671,N_4771);
and U4952 (N_4952,N_4772,N_4729);
nor U4953 (N_4953,N_4686,N_4627);
or U4954 (N_4954,N_4749,N_4759);
nand U4955 (N_4955,N_4746,N_4680);
nand U4956 (N_4956,N_4707,N_4724);
and U4957 (N_4957,N_4758,N_4750);
nor U4958 (N_4958,N_4615,N_4757);
xor U4959 (N_4959,N_4731,N_4774);
nand U4960 (N_4960,N_4610,N_4723);
nor U4961 (N_4961,N_4636,N_4716);
xnor U4962 (N_4962,N_4671,N_4746);
and U4963 (N_4963,N_4628,N_4716);
or U4964 (N_4964,N_4626,N_4786);
or U4965 (N_4965,N_4701,N_4674);
and U4966 (N_4966,N_4612,N_4770);
or U4967 (N_4967,N_4648,N_4799);
xor U4968 (N_4968,N_4734,N_4609);
xor U4969 (N_4969,N_4763,N_4645);
nand U4970 (N_4970,N_4764,N_4769);
nor U4971 (N_4971,N_4631,N_4679);
nand U4972 (N_4972,N_4787,N_4724);
and U4973 (N_4973,N_4758,N_4611);
xnor U4974 (N_4974,N_4704,N_4686);
xnor U4975 (N_4975,N_4710,N_4652);
xor U4976 (N_4976,N_4773,N_4665);
or U4977 (N_4977,N_4782,N_4609);
nand U4978 (N_4978,N_4711,N_4656);
or U4979 (N_4979,N_4738,N_4704);
and U4980 (N_4980,N_4754,N_4722);
xnor U4981 (N_4981,N_4693,N_4645);
xor U4982 (N_4982,N_4798,N_4635);
and U4983 (N_4983,N_4747,N_4761);
and U4984 (N_4984,N_4757,N_4754);
xnor U4985 (N_4985,N_4700,N_4732);
or U4986 (N_4986,N_4789,N_4686);
or U4987 (N_4987,N_4743,N_4611);
or U4988 (N_4988,N_4764,N_4606);
xor U4989 (N_4989,N_4649,N_4723);
nand U4990 (N_4990,N_4757,N_4678);
and U4991 (N_4991,N_4672,N_4772);
or U4992 (N_4992,N_4664,N_4617);
nand U4993 (N_4993,N_4644,N_4639);
or U4994 (N_4994,N_4796,N_4610);
and U4995 (N_4995,N_4683,N_4652);
or U4996 (N_4996,N_4747,N_4718);
nand U4997 (N_4997,N_4706,N_4758);
xor U4998 (N_4998,N_4616,N_4790);
nand U4999 (N_4999,N_4707,N_4651);
nand U5000 (N_5000,N_4897,N_4926);
xnor U5001 (N_5001,N_4850,N_4953);
and U5002 (N_5002,N_4949,N_4877);
nor U5003 (N_5003,N_4981,N_4823);
nand U5004 (N_5004,N_4844,N_4820);
and U5005 (N_5005,N_4995,N_4907);
and U5006 (N_5006,N_4848,N_4912);
and U5007 (N_5007,N_4982,N_4828);
or U5008 (N_5008,N_4904,N_4928);
nand U5009 (N_5009,N_4855,N_4806);
nor U5010 (N_5010,N_4961,N_4807);
xor U5011 (N_5011,N_4871,N_4888);
nor U5012 (N_5012,N_4868,N_4999);
and U5013 (N_5013,N_4860,N_4833);
or U5014 (N_5014,N_4822,N_4954);
and U5015 (N_5015,N_4834,N_4900);
and U5016 (N_5016,N_4908,N_4966);
nor U5017 (N_5017,N_4846,N_4958);
xnor U5018 (N_5018,N_4946,N_4903);
and U5019 (N_5019,N_4803,N_4826);
and U5020 (N_5020,N_4997,N_4976);
xor U5021 (N_5021,N_4998,N_4801);
nand U5022 (N_5022,N_4889,N_4873);
xor U5023 (N_5023,N_4964,N_4840);
or U5024 (N_5024,N_4913,N_4817);
nand U5025 (N_5025,N_4970,N_4906);
or U5026 (N_5026,N_4872,N_4879);
nand U5027 (N_5027,N_4957,N_4863);
nand U5028 (N_5028,N_4940,N_4925);
nand U5029 (N_5029,N_4808,N_4853);
nor U5030 (N_5030,N_4890,N_4869);
and U5031 (N_5031,N_4992,N_4810);
nor U5032 (N_5032,N_4951,N_4914);
or U5033 (N_5033,N_4852,N_4837);
nand U5034 (N_5034,N_4933,N_4994);
xor U5035 (N_5035,N_4993,N_4874);
nand U5036 (N_5036,N_4878,N_4839);
nor U5037 (N_5037,N_4934,N_4991);
nand U5038 (N_5038,N_4922,N_4980);
xor U5039 (N_5039,N_4930,N_4857);
nor U5040 (N_5040,N_4851,N_4841);
or U5041 (N_5041,N_4870,N_4990);
nor U5042 (N_5042,N_4819,N_4829);
nand U5043 (N_5043,N_4898,N_4832);
or U5044 (N_5044,N_4883,N_4895);
nor U5045 (N_5045,N_4974,N_4963);
or U5046 (N_5046,N_4996,N_4911);
nand U5047 (N_5047,N_4915,N_4866);
nor U5048 (N_5048,N_4917,N_4942);
or U5049 (N_5049,N_4856,N_4847);
and U5050 (N_5050,N_4927,N_4918);
nand U5051 (N_5051,N_4864,N_4821);
nand U5052 (N_5052,N_4919,N_4842);
nand U5053 (N_5053,N_4902,N_4838);
nor U5054 (N_5054,N_4984,N_4884);
nand U5055 (N_5055,N_4941,N_4955);
and U5056 (N_5056,N_4921,N_4891);
xor U5057 (N_5057,N_4950,N_4867);
nor U5058 (N_5058,N_4809,N_4825);
and U5059 (N_5059,N_4965,N_4929);
and U5060 (N_5060,N_4845,N_4830);
xor U5061 (N_5061,N_4945,N_4814);
or U5062 (N_5062,N_4875,N_4988);
nor U5063 (N_5063,N_4952,N_4862);
nand U5064 (N_5064,N_4849,N_4923);
nand U5065 (N_5065,N_4967,N_4983);
nor U5066 (N_5066,N_4824,N_4947);
and U5067 (N_5067,N_4944,N_4865);
and U5068 (N_5068,N_4811,N_4979);
xor U5069 (N_5069,N_4881,N_4827);
xnor U5070 (N_5070,N_4885,N_4939);
nand U5071 (N_5071,N_4835,N_4893);
nand U5072 (N_5072,N_4812,N_4948);
nand U5073 (N_5073,N_4876,N_4943);
nor U5074 (N_5074,N_4887,N_4920);
nor U5075 (N_5075,N_4989,N_4859);
xor U5076 (N_5076,N_4937,N_4858);
nand U5077 (N_5077,N_4836,N_4892);
or U5078 (N_5078,N_4899,N_4972);
nand U5079 (N_5079,N_4886,N_4971);
xnor U5080 (N_5080,N_4935,N_4931);
and U5081 (N_5081,N_4985,N_4924);
nor U5082 (N_5082,N_4978,N_4938);
or U5083 (N_5083,N_4910,N_4973);
and U5084 (N_5084,N_4861,N_4816);
nand U5085 (N_5085,N_4901,N_4896);
nand U5086 (N_5086,N_4815,N_4804);
xnor U5087 (N_5087,N_4932,N_4818);
nor U5088 (N_5088,N_4987,N_4813);
nor U5089 (N_5089,N_4975,N_4854);
or U5090 (N_5090,N_4960,N_4894);
nand U5091 (N_5091,N_4805,N_4802);
nand U5092 (N_5092,N_4959,N_4800);
nor U5093 (N_5093,N_4977,N_4962);
nor U5094 (N_5094,N_4909,N_4968);
xnor U5095 (N_5095,N_4986,N_4936);
and U5096 (N_5096,N_4969,N_4905);
or U5097 (N_5097,N_4956,N_4831);
xnor U5098 (N_5098,N_4880,N_4882);
and U5099 (N_5099,N_4843,N_4916);
or U5100 (N_5100,N_4829,N_4891);
nand U5101 (N_5101,N_4893,N_4898);
nand U5102 (N_5102,N_4801,N_4833);
nand U5103 (N_5103,N_4879,N_4889);
xnor U5104 (N_5104,N_4971,N_4873);
nor U5105 (N_5105,N_4897,N_4888);
nand U5106 (N_5106,N_4863,N_4939);
xor U5107 (N_5107,N_4910,N_4945);
or U5108 (N_5108,N_4874,N_4972);
nand U5109 (N_5109,N_4998,N_4893);
and U5110 (N_5110,N_4846,N_4909);
nor U5111 (N_5111,N_4942,N_4915);
nand U5112 (N_5112,N_4935,N_4827);
and U5113 (N_5113,N_4882,N_4894);
xor U5114 (N_5114,N_4844,N_4931);
and U5115 (N_5115,N_4875,N_4877);
and U5116 (N_5116,N_4900,N_4830);
xor U5117 (N_5117,N_4843,N_4922);
nor U5118 (N_5118,N_4813,N_4933);
nand U5119 (N_5119,N_4896,N_4931);
xor U5120 (N_5120,N_4938,N_4801);
xor U5121 (N_5121,N_4856,N_4850);
nor U5122 (N_5122,N_4885,N_4855);
nor U5123 (N_5123,N_4851,N_4862);
xor U5124 (N_5124,N_4845,N_4891);
xor U5125 (N_5125,N_4880,N_4905);
xor U5126 (N_5126,N_4977,N_4876);
xor U5127 (N_5127,N_4900,N_4891);
or U5128 (N_5128,N_4838,N_4863);
and U5129 (N_5129,N_4937,N_4939);
nor U5130 (N_5130,N_4892,N_4857);
xor U5131 (N_5131,N_4821,N_4884);
or U5132 (N_5132,N_4998,N_4982);
xor U5133 (N_5133,N_4802,N_4831);
xnor U5134 (N_5134,N_4804,N_4913);
xor U5135 (N_5135,N_4910,N_4954);
xor U5136 (N_5136,N_4925,N_4929);
xnor U5137 (N_5137,N_4801,N_4840);
nor U5138 (N_5138,N_4898,N_4981);
xor U5139 (N_5139,N_4989,N_4840);
nor U5140 (N_5140,N_4936,N_4912);
nor U5141 (N_5141,N_4830,N_4967);
or U5142 (N_5142,N_4927,N_4878);
and U5143 (N_5143,N_4811,N_4855);
or U5144 (N_5144,N_4870,N_4835);
nor U5145 (N_5145,N_4809,N_4977);
and U5146 (N_5146,N_4923,N_4940);
and U5147 (N_5147,N_4995,N_4892);
xnor U5148 (N_5148,N_4959,N_4848);
and U5149 (N_5149,N_4853,N_4913);
and U5150 (N_5150,N_4988,N_4843);
nor U5151 (N_5151,N_4946,N_4987);
or U5152 (N_5152,N_4948,N_4817);
and U5153 (N_5153,N_4897,N_4933);
nor U5154 (N_5154,N_4873,N_4978);
nand U5155 (N_5155,N_4928,N_4967);
xnor U5156 (N_5156,N_4898,N_4855);
and U5157 (N_5157,N_4800,N_4821);
nand U5158 (N_5158,N_4930,N_4917);
or U5159 (N_5159,N_4926,N_4893);
and U5160 (N_5160,N_4806,N_4972);
nand U5161 (N_5161,N_4844,N_4838);
or U5162 (N_5162,N_4881,N_4992);
and U5163 (N_5163,N_4854,N_4889);
and U5164 (N_5164,N_4968,N_4883);
nor U5165 (N_5165,N_4933,N_4978);
and U5166 (N_5166,N_4857,N_4997);
and U5167 (N_5167,N_4872,N_4854);
xnor U5168 (N_5168,N_4939,N_4878);
or U5169 (N_5169,N_4975,N_4823);
nand U5170 (N_5170,N_4968,N_4849);
nor U5171 (N_5171,N_4902,N_4800);
nand U5172 (N_5172,N_4966,N_4918);
xnor U5173 (N_5173,N_4845,N_4928);
xor U5174 (N_5174,N_4821,N_4897);
xor U5175 (N_5175,N_4815,N_4952);
or U5176 (N_5176,N_4834,N_4962);
and U5177 (N_5177,N_4931,N_4955);
nor U5178 (N_5178,N_4959,N_4852);
or U5179 (N_5179,N_4927,N_4888);
xor U5180 (N_5180,N_4905,N_4869);
nor U5181 (N_5181,N_4920,N_4947);
xnor U5182 (N_5182,N_4834,N_4931);
nor U5183 (N_5183,N_4947,N_4907);
and U5184 (N_5184,N_4873,N_4814);
xor U5185 (N_5185,N_4800,N_4872);
nand U5186 (N_5186,N_4853,N_4830);
nor U5187 (N_5187,N_4960,N_4956);
or U5188 (N_5188,N_4976,N_4959);
nor U5189 (N_5189,N_4869,N_4863);
and U5190 (N_5190,N_4864,N_4940);
and U5191 (N_5191,N_4802,N_4888);
or U5192 (N_5192,N_4818,N_4908);
xnor U5193 (N_5193,N_4985,N_4954);
and U5194 (N_5194,N_4944,N_4802);
or U5195 (N_5195,N_4994,N_4803);
nor U5196 (N_5196,N_4818,N_4886);
nor U5197 (N_5197,N_4955,N_4972);
nand U5198 (N_5198,N_4904,N_4877);
xnor U5199 (N_5199,N_4822,N_4854);
nand U5200 (N_5200,N_5152,N_5059);
or U5201 (N_5201,N_5010,N_5003);
xor U5202 (N_5202,N_5092,N_5142);
nor U5203 (N_5203,N_5013,N_5191);
xor U5204 (N_5204,N_5053,N_5115);
xor U5205 (N_5205,N_5033,N_5052);
nand U5206 (N_5206,N_5162,N_5019);
nand U5207 (N_5207,N_5025,N_5129);
and U5208 (N_5208,N_5176,N_5001);
and U5209 (N_5209,N_5096,N_5021);
nor U5210 (N_5210,N_5029,N_5193);
and U5211 (N_5211,N_5011,N_5143);
or U5212 (N_5212,N_5064,N_5043);
nand U5213 (N_5213,N_5095,N_5174);
nor U5214 (N_5214,N_5119,N_5007);
and U5215 (N_5215,N_5130,N_5135);
nand U5216 (N_5216,N_5114,N_5134);
nand U5217 (N_5217,N_5110,N_5044);
or U5218 (N_5218,N_5036,N_5113);
nand U5219 (N_5219,N_5136,N_5057);
or U5220 (N_5220,N_5189,N_5076);
nand U5221 (N_5221,N_5118,N_5006);
nand U5222 (N_5222,N_5054,N_5102);
nor U5223 (N_5223,N_5023,N_5050);
nor U5224 (N_5224,N_5172,N_5042);
or U5225 (N_5225,N_5038,N_5144);
nand U5226 (N_5226,N_5128,N_5037);
nand U5227 (N_5227,N_5131,N_5196);
and U5228 (N_5228,N_5195,N_5146);
nand U5229 (N_5229,N_5024,N_5156);
or U5230 (N_5230,N_5084,N_5069);
and U5231 (N_5231,N_5198,N_5139);
xnor U5232 (N_5232,N_5161,N_5032);
and U5233 (N_5233,N_5098,N_5170);
or U5234 (N_5234,N_5034,N_5192);
nand U5235 (N_5235,N_5080,N_5116);
nand U5236 (N_5236,N_5109,N_5111);
xor U5237 (N_5237,N_5167,N_5039);
xnor U5238 (N_5238,N_5027,N_5009);
and U5239 (N_5239,N_5062,N_5085);
or U5240 (N_5240,N_5046,N_5180);
and U5241 (N_5241,N_5017,N_5126);
and U5242 (N_5242,N_5079,N_5061);
and U5243 (N_5243,N_5040,N_5133);
xor U5244 (N_5244,N_5071,N_5022);
xor U5245 (N_5245,N_5179,N_5107);
or U5246 (N_5246,N_5028,N_5187);
and U5247 (N_5247,N_5141,N_5091);
nor U5248 (N_5248,N_5089,N_5164);
and U5249 (N_5249,N_5158,N_5138);
or U5250 (N_5250,N_5173,N_5030);
and U5251 (N_5251,N_5168,N_5145);
xnor U5252 (N_5252,N_5063,N_5016);
xnor U5253 (N_5253,N_5086,N_5125);
nand U5254 (N_5254,N_5122,N_5008);
nor U5255 (N_5255,N_5137,N_5002);
and U5256 (N_5256,N_5070,N_5171);
nor U5257 (N_5257,N_5188,N_5049);
nor U5258 (N_5258,N_5075,N_5081);
nand U5259 (N_5259,N_5154,N_5190);
xor U5260 (N_5260,N_5047,N_5093);
xor U5261 (N_5261,N_5060,N_5103);
or U5262 (N_5262,N_5150,N_5148);
nand U5263 (N_5263,N_5056,N_5014);
xnor U5264 (N_5264,N_5005,N_5072);
xor U5265 (N_5265,N_5157,N_5067);
nor U5266 (N_5266,N_5088,N_5087);
nor U5267 (N_5267,N_5048,N_5163);
xor U5268 (N_5268,N_5140,N_5101);
and U5269 (N_5269,N_5112,N_5151);
nor U5270 (N_5270,N_5020,N_5132);
xor U5271 (N_5271,N_5117,N_5159);
or U5272 (N_5272,N_5160,N_5199);
and U5273 (N_5273,N_5106,N_5155);
nand U5274 (N_5274,N_5082,N_5104);
and U5275 (N_5275,N_5066,N_5015);
and U5276 (N_5276,N_5012,N_5031);
nor U5277 (N_5277,N_5123,N_5058);
or U5278 (N_5278,N_5068,N_5073);
xor U5279 (N_5279,N_5120,N_5149);
and U5280 (N_5280,N_5184,N_5166);
nor U5281 (N_5281,N_5083,N_5026);
and U5282 (N_5282,N_5051,N_5035);
or U5283 (N_5283,N_5105,N_5165);
nand U5284 (N_5284,N_5153,N_5124);
and U5285 (N_5285,N_5147,N_5018);
or U5286 (N_5286,N_5181,N_5183);
nand U5287 (N_5287,N_5077,N_5108);
xor U5288 (N_5288,N_5041,N_5074);
nor U5289 (N_5289,N_5000,N_5097);
or U5290 (N_5290,N_5094,N_5169);
or U5291 (N_5291,N_5186,N_5178);
xnor U5292 (N_5292,N_5055,N_5197);
nand U5293 (N_5293,N_5127,N_5100);
and U5294 (N_5294,N_5175,N_5121);
nand U5295 (N_5295,N_5090,N_5185);
or U5296 (N_5296,N_5065,N_5194);
or U5297 (N_5297,N_5078,N_5182);
and U5298 (N_5298,N_5045,N_5177);
nand U5299 (N_5299,N_5099,N_5004);
nor U5300 (N_5300,N_5085,N_5111);
or U5301 (N_5301,N_5181,N_5003);
and U5302 (N_5302,N_5074,N_5159);
or U5303 (N_5303,N_5102,N_5129);
and U5304 (N_5304,N_5177,N_5103);
nand U5305 (N_5305,N_5092,N_5019);
nor U5306 (N_5306,N_5194,N_5115);
or U5307 (N_5307,N_5016,N_5185);
nand U5308 (N_5308,N_5182,N_5028);
nor U5309 (N_5309,N_5033,N_5118);
or U5310 (N_5310,N_5046,N_5192);
or U5311 (N_5311,N_5110,N_5013);
or U5312 (N_5312,N_5169,N_5084);
nor U5313 (N_5313,N_5012,N_5121);
or U5314 (N_5314,N_5101,N_5103);
xor U5315 (N_5315,N_5131,N_5063);
xnor U5316 (N_5316,N_5082,N_5154);
nor U5317 (N_5317,N_5044,N_5168);
or U5318 (N_5318,N_5108,N_5016);
nor U5319 (N_5319,N_5082,N_5064);
nand U5320 (N_5320,N_5193,N_5103);
and U5321 (N_5321,N_5008,N_5145);
and U5322 (N_5322,N_5069,N_5180);
xor U5323 (N_5323,N_5179,N_5097);
xnor U5324 (N_5324,N_5145,N_5084);
nor U5325 (N_5325,N_5011,N_5140);
or U5326 (N_5326,N_5034,N_5112);
and U5327 (N_5327,N_5079,N_5174);
and U5328 (N_5328,N_5077,N_5184);
nand U5329 (N_5329,N_5162,N_5088);
nand U5330 (N_5330,N_5153,N_5052);
nand U5331 (N_5331,N_5077,N_5042);
and U5332 (N_5332,N_5170,N_5102);
xnor U5333 (N_5333,N_5178,N_5029);
nor U5334 (N_5334,N_5149,N_5190);
nor U5335 (N_5335,N_5030,N_5056);
and U5336 (N_5336,N_5107,N_5162);
and U5337 (N_5337,N_5059,N_5052);
nor U5338 (N_5338,N_5073,N_5191);
nand U5339 (N_5339,N_5068,N_5016);
and U5340 (N_5340,N_5005,N_5040);
nor U5341 (N_5341,N_5096,N_5007);
xnor U5342 (N_5342,N_5174,N_5063);
and U5343 (N_5343,N_5139,N_5161);
and U5344 (N_5344,N_5051,N_5000);
xor U5345 (N_5345,N_5056,N_5063);
nand U5346 (N_5346,N_5148,N_5114);
nor U5347 (N_5347,N_5058,N_5065);
nand U5348 (N_5348,N_5168,N_5107);
nand U5349 (N_5349,N_5058,N_5170);
nor U5350 (N_5350,N_5161,N_5173);
xnor U5351 (N_5351,N_5097,N_5130);
xnor U5352 (N_5352,N_5096,N_5162);
and U5353 (N_5353,N_5194,N_5143);
nand U5354 (N_5354,N_5153,N_5149);
xor U5355 (N_5355,N_5142,N_5048);
nor U5356 (N_5356,N_5050,N_5068);
xor U5357 (N_5357,N_5158,N_5161);
xor U5358 (N_5358,N_5060,N_5154);
nand U5359 (N_5359,N_5137,N_5168);
and U5360 (N_5360,N_5039,N_5058);
or U5361 (N_5361,N_5063,N_5147);
or U5362 (N_5362,N_5167,N_5135);
and U5363 (N_5363,N_5096,N_5146);
xor U5364 (N_5364,N_5149,N_5176);
nand U5365 (N_5365,N_5129,N_5091);
xor U5366 (N_5366,N_5092,N_5031);
nand U5367 (N_5367,N_5030,N_5152);
xnor U5368 (N_5368,N_5150,N_5028);
or U5369 (N_5369,N_5067,N_5164);
nor U5370 (N_5370,N_5199,N_5171);
xnor U5371 (N_5371,N_5055,N_5090);
and U5372 (N_5372,N_5003,N_5076);
nor U5373 (N_5373,N_5145,N_5133);
or U5374 (N_5374,N_5065,N_5092);
xnor U5375 (N_5375,N_5153,N_5056);
nor U5376 (N_5376,N_5127,N_5012);
nor U5377 (N_5377,N_5027,N_5196);
nand U5378 (N_5378,N_5016,N_5156);
xor U5379 (N_5379,N_5176,N_5093);
xor U5380 (N_5380,N_5173,N_5059);
xnor U5381 (N_5381,N_5175,N_5178);
nor U5382 (N_5382,N_5194,N_5042);
or U5383 (N_5383,N_5046,N_5093);
nor U5384 (N_5384,N_5127,N_5168);
nor U5385 (N_5385,N_5131,N_5090);
nand U5386 (N_5386,N_5168,N_5094);
nand U5387 (N_5387,N_5147,N_5172);
or U5388 (N_5388,N_5038,N_5190);
and U5389 (N_5389,N_5156,N_5176);
nor U5390 (N_5390,N_5122,N_5050);
or U5391 (N_5391,N_5148,N_5046);
xor U5392 (N_5392,N_5068,N_5034);
nand U5393 (N_5393,N_5155,N_5095);
xor U5394 (N_5394,N_5108,N_5107);
or U5395 (N_5395,N_5130,N_5010);
nand U5396 (N_5396,N_5037,N_5160);
and U5397 (N_5397,N_5140,N_5175);
xor U5398 (N_5398,N_5070,N_5013);
nand U5399 (N_5399,N_5033,N_5120);
nor U5400 (N_5400,N_5354,N_5259);
nor U5401 (N_5401,N_5328,N_5262);
nor U5402 (N_5402,N_5324,N_5268);
xnor U5403 (N_5403,N_5247,N_5229);
nand U5404 (N_5404,N_5209,N_5206);
xnor U5405 (N_5405,N_5253,N_5356);
xnor U5406 (N_5406,N_5320,N_5234);
xor U5407 (N_5407,N_5362,N_5383);
or U5408 (N_5408,N_5303,N_5367);
nand U5409 (N_5409,N_5244,N_5302);
or U5410 (N_5410,N_5369,N_5271);
xor U5411 (N_5411,N_5387,N_5331);
xor U5412 (N_5412,N_5260,N_5222);
or U5413 (N_5413,N_5238,N_5360);
nand U5414 (N_5414,N_5230,N_5342);
xnor U5415 (N_5415,N_5295,N_5350);
or U5416 (N_5416,N_5364,N_5378);
and U5417 (N_5417,N_5339,N_5393);
or U5418 (N_5418,N_5207,N_5336);
nor U5419 (N_5419,N_5212,N_5266);
and U5420 (N_5420,N_5258,N_5214);
and U5421 (N_5421,N_5241,N_5312);
nor U5422 (N_5422,N_5300,N_5274);
or U5423 (N_5423,N_5231,N_5255);
nor U5424 (N_5424,N_5273,N_5397);
or U5425 (N_5425,N_5297,N_5308);
xor U5426 (N_5426,N_5293,N_5334);
xor U5427 (N_5427,N_5216,N_5371);
and U5428 (N_5428,N_5257,N_5326);
xnor U5429 (N_5429,N_5278,N_5385);
nor U5430 (N_5430,N_5279,N_5355);
nor U5431 (N_5431,N_5332,N_5347);
nand U5432 (N_5432,N_5346,N_5372);
nor U5433 (N_5433,N_5392,N_5205);
nand U5434 (N_5434,N_5237,N_5319);
or U5435 (N_5435,N_5269,N_5281);
xnor U5436 (N_5436,N_5323,N_5298);
and U5437 (N_5437,N_5314,N_5213);
or U5438 (N_5438,N_5275,N_5235);
and U5439 (N_5439,N_5317,N_5220);
and U5440 (N_5440,N_5313,N_5218);
xnor U5441 (N_5441,N_5363,N_5288);
nand U5442 (N_5442,N_5282,N_5223);
nand U5443 (N_5443,N_5370,N_5379);
or U5444 (N_5444,N_5345,N_5301);
nand U5445 (N_5445,N_5309,N_5228);
and U5446 (N_5446,N_5219,N_5264);
nor U5447 (N_5447,N_5325,N_5361);
nand U5448 (N_5448,N_5398,N_5399);
and U5449 (N_5449,N_5263,N_5359);
and U5450 (N_5450,N_5291,N_5307);
nand U5451 (N_5451,N_5208,N_5340);
xnor U5452 (N_5452,N_5210,N_5265);
xnor U5453 (N_5453,N_5284,N_5276);
xnor U5454 (N_5454,N_5344,N_5376);
nand U5455 (N_5455,N_5221,N_5246);
and U5456 (N_5456,N_5270,N_5261);
xnor U5457 (N_5457,N_5305,N_5202);
and U5458 (N_5458,N_5321,N_5335);
or U5459 (N_5459,N_5333,N_5351);
or U5460 (N_5460,N_5327,N_5232);
and U5461 (N_5461,N_5290,N_5352);
nand U5462 (N_5462,N_5343,N_5225);
nor U5463 (N_5463,N_5217,N_5233);
nor U5464 (N_5464,N_5294,N_5292);
and U5465 (N_5465,N_5373,N_5380);
or U5466 (N_5466,N_5330,N_5285);
and U5467 (N_5467,N_5318,N_5338);
xnor U5468 (N_5468,N_5315,N_5287);
xor U5469 (N_5469,N_5395,N_5267);
xor U5470 (N_5470,N_5322,N_5201);
or U5471 (N_5471,N_5224,N_5341);
and U5472 (N_5472,N_5375,N_5296);
nor U5473 (N_5473,N_5366,N_5388);
xnor U5474 (N_5474,N_5365,N_5240);
nand U5475 (N_5475,N_5353,N_5368);
and U5476 (N_5476,N_5283,N_5329);
or U5477 (N_5477,N_5250,N_5348);
nand U5478 (N_5478,N_5204,N_5299);
nand U5479 (N_5479,N_5272,N_5386);
and U5480 (N_5480,N_5389,N_5349);
nor U5481 (N_5481,N_5239,N_5256);
xor U5482 (N_5482,N_5396,N_5357);
nor U5483 (N_5483,N_5243,N_5203);
nand U5484 (N_5484,N_5252,N_5358);
nand U5485 (N_5485,N_5245,N_5311);
nand U5486 (N_5486,N_5211,N_5242);
nand U5487 (N_5487,N_5236,N_5254);
xnor U5488 (N_5488,N_5391,N_5374);
or U5489 (N_5489,N_5215,N_5251);
and U5490 (N_5490,N_5226,N_5227);
and U5491 (N_5491,N_5304,N_5249);
and U5492 (N_5492,N_5316,N_5384);
nor U5493 (N_5493,N_5382,N_5390);
or U5494 (N_5494,N_5377,N_5200);
nor U5495 (N_5495,N_5306,N_5310);
and U5496 (N_5496,N_5394,N_5248);
xor U5497 (N_5497,N_5337,N_5277);
nand U5498 (N_5498,N_5286,N_5280);
and U5499 (N_5499,N_5381,N_5289);
nand U5500 (N_5500,N_5285,N_5370);
and U5501 (N_5501,N_5332,N_5377);
or U5502 (N_5502,N_5292,N_5375);
and U5503 (N_5503,N_5378,N_5214);
xor U5504 (N_5504,N_5253,N_5298);
xnor U5505 (N_5505,N_5250,N_5342);
nand U5506 (N_5506,N_5374,N_5208);
or U5507 (N_5507,N_5220,N_5392);
nor U5508 (N_5508,N_5371,N_5240);
nand U5509 (N_5509,N_5258,N_5390);
or U5510 (N_5510,N_5339,N_5310);
and U5511 (N_5511,N_5390,N_5393);
nand U5512 (N_5512,N_5377,N_5387);
xnor U5513 (N_5513,N_5387,N_5218);
xor U5514 (N_5514,N_5327,N_5233);
or U5515 (N_5515,N_5228,N_5268);
nand U5516 (N_5516,N_5290,N_5204);
xnor U5517 (N_5517,N_5302,N_5231);
nor U5518 (N_5518,N_5358,N_5372);
and U5519 (N_5519,N_5304,N_5332);
or U5520 (N_5520,N_5354,N_5328);
xor U5521 (N_5521,N_5357,N_5223);
nand U5522 (N_5522,N_5248,N_5290);
and U5523 (N_5523,N_5301,N_5209);
xnor U5524 (N_5524,N_5321,N_5309);
nand U5525 (N_5525,N_5376,N_5322);
xor U5526 (N_5526,N_5342,N_5351);
nand U5527 (N_5527,N_5365,N_5310);
and U5528 (N_5528,N_5296,N_5367);
nand U5529 (N_5529,N_5212,N_5295);
nand U5530 (N_5530,N_5317,N_5330);
and U5531 (N_5531,N_5317,N_5324);
xnor U5532 (N_5532,N_5250,N_5253);
and U5533 (N_5533,N_5248,N_5316);
nor U5534 (N_5534,N_5362,N_5263);
xnor U5535 (N_5535,N_5287,N_5274);
and U5536 (N_5536,N_5224,N_5232);
xor U5537 (N_5537,N_5200,N_5348);
xnor U5538 (N_5538,N_5380,N_5206);
or U5539 (N_5539,N_5243,N_5397);
nand U5540 (N_5540,N_5320,N_5374);
or U5541 (N_5541,N_5367,N_5231);
or U5542 (N_5542,N_5296,N_5299);
or U5543 (N_5543,N_5268,N_5238);
and U5544 (N_5544,N_5249,N_5356);
nor U5545 (N_5545,N_5271,N_5337);
and U5546 (N_5546,N_5303,N_5217);
nor U5547 (N_5547,N_5224,N_5393);
nand U5548 (N_5548,N_5202,N_5303);
and U5549 (N_5549,N_5225,N_5299);
or U5550 (N_5550,N_5390,N_5319);
or U5551 (N_5551,N_5202,N_5380);
xnor U5552 (N_5552,N_5266,N_5366);
xor U5553 (N_5553,N_5340,N_5330);
xnor U5554 (N_5554,N_5233,N_5377);
xnor U5555 (N_5555,N_5257,N_5284);
nor U5556 (N_5556,N_5308,N_5396);
nand U5557 (N_5557,N_5249,N_5258);
or U5558 (N_5558,N_5291,N_5399);
and U5559 (N_5559,N_5324,N_5280);
xor U5560 (N_5560,N_5254,N_5367);
or U5561 (N_5561,N_5285,N_5286);
or U5562 (N_5562,N_5291,N_5336);
or U5563 (N_5563,N_5204,N_5262);
nor U5564 (N_5564,N_5339,N_5372);
or U5565 (N_5565,N_5232,N_5277);
nand U5566 (N_5566,N_5295,N_5346);
xor U5567 (N_5567,N_5226,N_5288);
nand U5568 (N_5568,N_5244,N_5358);
or U5569 (N_5569,N_5210,N_5232);
and U5570 (N_5570,N_5377,N_5345);
and U5571 (N_5571,N_5305,N_5352);
and U5572 (N_5572,N_5211,N_5295);
or U5573 (N_5573,N_5282,N_5239);
nor U5574 (N_5574,N_5317,N_5290);
xor U5575 (N_5575,N_5280,N_5255);
or U5576 (N_5576,N_5308,N_5238);
or U5577 (N_5577,N_5292,N_5394);
xor U5578 (N_5578,N_5246,N_5358);
nand U5579 (N_5579,N_5263,N_5351);
nand U5580 (N_5580,N_5252,N_5297);
xor U5581 (N_5581,N_5396,N_5265);
or U5582 (N_5582,N_5265,N_5280);
and U5583 (N_5583,N_5328,N_5338);
and U5584 (N_5584,N_5381,N_5301);
nor U5585 (N_5585,N_5254,N_5241);
xnor U5586 (N_5586,N_5326,N_5268);
and U5587 (N_5587,N_5323,N_5219);
xor U5588 (N_5588,N_5216,N_5261);
and U5589 (N_5589,N_5337,N_5335);
and U5590 (N_5590,N_5333,N_5384);
nand U5591 (N_5591,N_5251,N_5344);
nand U5592 (N_5592,N_5332,N_5249);
and U5593 (N_5593,N_5295,N_5332);
nand U5594 (N_5594,N_5347,N_5227);
or U5595 (N_5595,N_5229,N_5281);
nand U5596 (N_5596,N_5259,N_5384);
nor U5597 (N_5597,N_5305,N_5259);
nor U5598 (N_5598,N_5302,N_5292);
and U5599 (N_5599,N_5302,N_5298);
nand U5600 (N_5600,N_5598,N_5494);
or U5601 (N_5601,N_5566,N_5540);
and U5602 (N_5602,N_5544,N_5419);
and U5603 (N_5603,N_5523,N_5575);
nand U5604 (N_5604,N_5577,N_5509);
nor U5605 (N_5605,N_5556,N_5487);
nor U5606 (N_5606,N_5549,N_5465);
and U5607 (N_5607,N_5499,N_5470);
nand U5608 (N_5608,N_5587,N_5539);
xnor U5609 (N_5609,N_5408,N_5532);
xor U5610 (N_5610,N_5551,N_5489);
nand U5611 (N_5611,N_5564,N_5478);
nor U5612 (N_5612,N_5527,N_5582);
nor U5613 (N_5613,N_5520,N_5426);
and U5614 (N_5614,N_5525,N_5596);
nand U5615 (N_5615,N_5430,N_5568);
xnor U5616 (N_5616,N_5561,N_5448);
or U5617 (N_5617,N_5594,N_5407);
nor U5618 (N_5618,N_5546,N_5530);
nor U5619 (N_5619,N_5559,N_5591);
and U5620 (N_5620,N_5410,N_5438);
nor U5621 (N_5621,N_5421,N_5437);
or U5622 (N_5622,N_5483,N_5583);
and U5623 (N_5623,N_5581,N_5447);
and U5624 (N_5624,N_5496,N_5480);
and U5625 (N_5625,N_5428,N_5454);
nand U5626 (N_5626,N_5513,N_5506);
nor U5627 (N_5627,N_5567,N_5429);
or U5628 (N_5628,N_5536,N_5570);
or U5629 (N_5629,N_5555,N_5535);
nor U5630 (N_5630,N_5490,N_5473);
or U5631 (N_5631,N_5491,N_5467);
nor U5632 (N_5632,N_5456,N_5445);
xnor U5633 (N_5633,N_5413,N_5440);
xor U5634 (N_5634,N_5433,N_5443);
or U5635 (N_5635,N_5545,N_5446);
and U5636 (N_5636,N_5451,N_5526);
nand U5637 (N_5637,N_5484,N_5592);
and U5638 (N_5638,N_5458,N_5521);
and U5639 (N_5639,N_5431,N_5522);
nor U5640 (N_5640,N_5441,N_5524);
and U5641 (N_5641,N_5424,N_5574);
nand U5642 (N_5642,N_5404,N_5599);
or U5643 (N_5643,N_5512,N_5497);
or U5644 (N_5644,N_5455,N_5550);
xnor U5645 (N_5645,N_5541,N_5505);
nor U5646 (N_5646,N_5519,N_5427);
xor U5647 (N_5647,N_5481,N_5571);
nor U5648 (N_5648,N_5400,N_5469);
and U5649 (N_5649,N_5548,N_5460);
xor U5650 (N_5650,N_5444,N_5537);
and U5651 (N_5651,N_5529,N_5588);
nor U5652 (N_5652,N_5502,N_5517);
nor U5653 (N_5653,N_5500,N_5562);
or U5654 (N_5654,N_5403,N_5442);
nor U5655 (N_5655,N_5584,N_5472);
and U5656 (N_5656,N_5547,N_5563);
xnor U5657 (N_5657,N_5528,N_5569);
xnor U5658 (N_5658,N_5414,N_5420);
and U5659 (N_5659,N_5415,N_5501);
xnor U5660 (N_5660,N_5492,N_5516);
xor U5661 (N_5661,N_5507,N_5508);
or U5662 (N_5662,N_5538,N_5466);
xor U5663 (N_5663,N_5578,N_5423);
and U5664 (N_5664,N_5597,N_5461);
nor U5665 (N_5665,N_5504,N_5471);
xnor U5666 (N_5666,N_5495,N_5557);
nor U5667 (N_5667,N_5553,N_5560);
and U5668 (N_5668,N_5402,N_5439);
xor U5669 (N_5669,N_5543,N_5464);
xor U5670 (N_5670,N_5565,N_5449);
xor U5671 (N_5671,N_5452,N_5580);
and U5672 (N_5672,N_5450,N_5576);
and U5673 (N_5673,N_5476,N_5422);
nand U5674 (N_5674,N_5418,N_5409);
or U5675 (N_5675,N_5595,N_5585);
or U5676 (N_5676,N_5579,N_5416);
and U5677 (N_5677,N_5411,N_5453);
or U5678 (N_5678,N_5590,N_5531);
xor U5679 (N_5679,N_5417,N_5493);
nand U5680 (N_5680,N_5462,N_5482);
and U5681 (N_5681,N_5533,N_5510);
nor U5682 (N_5682,N_5435,N_5503);
and U5683 (N_5683,N_5586,N_5401);
xor U5684 (N_5684,N_5436,N_5552);
xnor U5685 (N_5685,N_5474,N_5488);
and U5686 (N_5686,N_5477,N_5554);
and U5687 (N_5687,N_5498,N_5558);
xor U5688 (N_5688,N_5486,N_5405);
and U5689 (N_5689,N_5542,N_5479);
xor U5690 (N_5690,N_5511,N_5572);
nor U5691 (N_5691,N_5534,N_5412);
and U5692 (N_5692,N_5432,N_5434);
nor U5693 (N_5693,N_5425,N_5463);
or U5694 (N_5694,N_5475,N_5457);
or U5695 (N_5695,N_5515,N_5573);
xnor U5696 (N_5696,N_5406,N_5593);
nand U5697 (N_5697,N_5468,N_5589);
xnor U5698 (N_5698,N_5518,N_5485);
xor U5699 (N_5699,N_5514,N_5459);
xnor U5700 (N_5700,N_5519,N_5494);
or U5701 (N_5701,N_5437,N_5560);
nor U5702 (N_5702,N_5515,N_5552);
or U5703 (N_5703,N_5539,N_5496);
nand U5704 (N_5704,N_5589,N_5457);
and U5705 (N_5705,N_5420,N_5488);
nand U5706 (N_5706,N_5413,N_5510);
or U5707 (N_5707,N_5576,N_5520);
nand U5708 (N_5708,N_5484,N_5486);
nand U5709 (N_5709,N_5539,N_5557);
and U5710 (N_5710,N_5573,N_5465);
xor U5711 (N_5711,N_5401,N_5416);
and U5712 (N_5712,N_5550,N_5557);
nor U5713 (N_5713,N_5551,N_5414);
and U5714 (N_5714,N_5594,N_5572);
nor U5715 (N_5715,N_5471,N_5554);
nor U5716 (N_5716,N_5408,N_5486);
and U5717 (N_5717,N_5410,N_5579);
and U5718 (N_5718,N_5489,N_5511);
nand U5719 (N_5719,N_5535,N_5482);
or U5720 (N_5720,N_5453,N_5554);
or U5721 (N_5721,N_5510,N_5485);
and U5722 (N_5722,N_5562,N_5452);
nor U5723 (N_5723,N_5448,N_5400);
nor U5724 (N_5724,N_5521,N_5477);
and U5725 (N_5725,N_5591,N_5588);
or U5726 (N_5726,N_5485,N_5486);
nor U5727 (N_5727,N_5470,N_5429);
xnor U5728 (N_5728,N_5414,N_5544);
or U5729 (N_5729,N_5595,N_5589);
nand U5730 (N_5730,N_5433,N_5473);
xor U5731 (N_5731,N_5595,N_5411);
xnor U5732 (N_5732,N_5480,N_5459);
and U5733 (N_5733,N_5506,N_5561);
or U5734 (N_5734,N_5433,N_5476);
or U5735 (N_5735,N_5527,N_5412);
xor U5736 (N_5736,N_5594,N_5423);
nand U5737 (N_5737,N_5495,N_5501);
or U5738 (N_5738,N_5528,N_5543);
or U5739 (N_5739,N_5562,N_5410);
xnor U5740 (N_5740,N_5482,N_5478);
xor U5741 (N_5741,N_5454,N_5471);
or U5742 (N_5742,N_5513,N_5458);
nand U5743 (N_5743,N_5507,N_5478);
xnor U5744 (N_5744,N_5548,N_5551);
or U5745 (N_5745,N_5560,N_5520);
and U5746 (N_5746,N_5424,N_5413);
nand U5747 (N_5747,N_5453,N_5501);
xnor U5748 (N_5748,N_5522,N_5523);
nand U5749 (N_5749,N_5453,N_5406);
nor U5750 (N_5750,N_5578,N_5440);
nor U5751 (N_5751,N_5424,N_5564);
nand U5752 (N_5752,N_5575,N_5508);
nor U5753 (N_5753,N_5455,N_5526);
xor U5754 (N_5754,N_5549,N_5472);
or U5755 (N_5755,N_5542,N_5455);
nor U5756 (N_5756,N_5451,N_5464);
and U5757 (N_5757,N_5479,N_5568);
and U5758 (N_5758,N_5437,N_5549);
xor U5759 (N_5759,N_5583,N_5530);
and U5760 (N_5760,N_5599,N_5493);
nand U5761 (N_5761,N_5409,N_5536);
and U5762 (N_5762,N_5552,N_5409);
xor U5763 (N_5763,N_5594,N_5555);
or U5764 (N_5764,N_5496,N_5578);
xnor U5765 (N_5765,N_5432,N_5487);
xnor U5766 (N_5766,N_5520,N_5590);
xor U5767 (N_5767,N_5580,N_5512);
or U5768 (N_5768,N_5594,N_5523);
xor U5769 (N_5769,N_5502,N_5506);
nand U5770 (N_5770,N_5496,N_5415);
xnor U5771 (N_5771,N_5477,N_5479);
nor U5772 (N_5772,N_5468,N_5410);
nand U5773 (N_5773,N_5500,N_5425);
xnor U5774 (N_5774,N_5494,N_5545);
nand U5775 (N_5775,N_5493,N_5509);
xor U5776 (N_5776,N_5561,N_5412);
and U5777 (N_5777,N_5466,N_5582);
nand U5778 (N_5778,N_5412,N_5422);
nand U5779 (N_5779,N_5575,N_5490);
or U5780 (N_5780,N_5448,N_5583);
xor U5781 (N_5781,N_5568,N_5521);
nor U5782 (N_5782,N_5566,N_5411);
nand U5783 (N_5783,N_5567,N_5540);
xnor U5784 (N_5784,N_5479,N_5464);
nor U5785 (N_5785,N_5457,N_5430);
nor U5786 (N_5786,N_5577,N_5442);
nor U5787 (N_5787,N_5477,N_5400);
and U5788 (N_5788,N_5454,N_5591);
or U5789 (N_5789,N_5466,N_5425);
nor U5790 (N_5790,N_5565,N_5560);
xnor U5791 (N_5791,N_5550,N_5564);
nor U5792 (N_5792,N_5416,N_5558);
and U5793 (N_5793,N_5506,N_5540);
nand U5794 (N_5794,N_5504,N_5415);
and U5795 (N_5795,N_5454,N_5481);
nand U5796 (N_5796,N_5432,N_5476);
nand U5797 (N_5797,N_5564,N_5403);
or U5798 (N_5798,N_5567,N_5568);
and U5799 (N_5799,N_5416,N_5580);
and U5800 (N_5800,N_5664,N_5682);
nor U5801 (N_5801,N_5652,N_5734);
or U5802 (N_5802,N_5780,N_5769);
and U5803 (N_5803,N_5707,N_5666);
and U5804 (N_5804,N_5612,N_5726);
nor U5805 (N_5805,N_5658,N_5686);
and U5806 (N_5806,N_5699,N_5669);
nor U5807 (N_5807,N_5733,N_5616);
and U5808 (N_5808,N_5798,N_5791);
nand U5809 (N_5809,N_5792,N_5725);
nor U5810 (N_5810,N_5774,N_5721);
xor U5811 (N_5811,N_5739,N_5723);
and U5812 (N_5812,N_5700,N_5709);
xnor U5813 (N_5813,N_5622,N_5683);
or U5814 (N_5814,N_5604,N_5633);
nand U5815 (N_5815,N_5790,N_5749);
or U5816 (N_5816,N_5777,N_5737);
xor U5817 (N_5817,N_5651,N_5753);
nor U5818 (N_5818,N_5718,N_5674);
nand U5819 (N_5819,N_5762,N_5659);
and U5820 (N_5820,N_5637,N_5771);
xor U5821 (N_5821,N_5759,N_5765);
nor U5822 (N_5822,N_5776,N_5758);
nor U5823 (N_5823,N_5678,N_5742);
nand U5824 (N_5824,N_5744,N_5665);
xor U5825 (N_5825,N_5614,N_5728);
and U5826 (N_5826,N_5796,N_5746);
or U5827 (N_5827,N_5773,N_5720);
or U5828 (N_5828,N_5706,N_5629);
and U5829 (N_5829,N_5602,N_5752);
and U5830 (N_5830,N_5626,N_5673);
or U5831 (N_5831,N_5679,N_5606);
xor U5832 (N_5832,N_5617,N_5600);
nor U5833 (N_5833,N_5741,N_5763);
nor U5834 (N_5834,N_5656,N_5645);
and U5835 (N_5835,N_5623,N_5687);
nand U5836 (N_5836,N_5670,N_5730);
xor U5837 (N_5837,N_5704,N_5624);
nand U5838 (N_5838,N_5722,N_5619);
or U5839 (N_5839,N_5740,N_5710);
xnor U5840 (N_5840,N_5605,N_5689);
xor U5841 (N_5841,N_5738,N_5748);
xor U5842 (N_5842,N_5768,N_5641);
or U5843 (N_5843,N_5672,N_5607);
nor U5844 (N_5844,N_5766,N_5787);
and U5845 (N_5845,N_5717,N_5654);
nand U5846 (N_5846,N_5799,N_5794);
nor U5847 (N_5847,N_5632,N_5712);
nand U5848 (N_5848,N_5745,N_5705);
or U5849 (N_5849,N_5714,N_5761);
xnor U5850 (N_5850,N_5713,N_5764);
and U5851 (N_5851,N_5630,N_5646);
and U5852 (N_5852,N_5751,N_5608);
nor U5853 (N_5853,N_5736,N_5634);
or U5854 (N_5854,N_5743,N_5628);
nor U5855 (N_5855,N_5681,N_5786);
xor U5856 (N_5856,N_5729,N_5701);
nand U5857 (N_5857,N_5639,N_5647);
nand U5858 (N_5858,N_5660,N_5711);
nor U5859 (N_5859,N_5603,N_5697);
nor U5860 (N_5860,N_5649,N_5620);
and U5861 (N_5861,N_5784,N_5653);
or U5862 (N_5862,N_5644,N_5662);
and U5863 (N_5863,N_5650,N_5657);
and U5864 (N_5864,N_5694,N_5750);
and U5865 (N_5865,N_5611,N_5783);
and U5866 (N_5866,N_5675,N_5690);
or U5867 (N_5867,N_5732,N_5724);
xor U5868 (N_5868,N_5655,N_5760);
nor U5869 (N_5869,N_5781,N_5716);
nor U5870 (N_5870,N_5668,N_5719);
and U5871 (N_5871,N_5770,N_5772);
nor U5872 (N_5872,N_5695,N_5703);
nor U5873 (N_5873,N_5667,N_5609);
xnor U5874 (N_5874,N_5642,N_5775);
nor U5875 (N_5875,N_5663,N_5688);
nor U5876 (N_5876,N_5708,N_5685);
and U5877 (N_5877,N_5613,N_5793);
xnor U5878 (N_5878,N_5767,N_5715);
xor U5879 (N_5879,N_5747,N_5782);
nor U5880 (N_5880,N_5635,N_5671);
nor U5881 (N_5881,N_5757,N_5684);
or U5882 (N_5882,N_5756,N_5702);
nand U5883 (N_5883,N_5610,N_5601);
or U5884 (N_5884,N_5789,N_5621);
xor U5885 (N_5885,N_5627,N_5680);
and U5886 (N_5886,N_5696,N_5640);
nand U5887 (N_5887,N_5691,N_5615);
or U5888 (N_5888,N_5638,N_5693);
nand U5889 (N_5889,N_5636,N_5797);
and U5890 (N_5890,N_5661,N_5779);
nor U5891 (N_5891,N_5648,N_5698);
or U5892 (N_5892,N_5755,N_5788);
nor U5893 (N_5893,N_5618,N_5785);
and U5894 (N_5894,N_5727,N_5631);
or U5895 (N_5895,N_5731,N_5692);
and U5896 (N_5896,N_5677,N_5754);
nor U5897 (N_5897,N_5778,N_5795);
nor U5898 (N_5898,N_5735,N_5643);
or U5899 (N_5899,N_5625,N_5676);
nand U5900 (N_5900,N_5667,N_5726);
or U5901 (N_5901,N_5614,N_5700);
and U5902 (N_5902,N_5649,N_5740);
and U5903 (N_5903,N_5622,N_5735);
nand U5904 (N_5904,N_5625,N_5636);
nand U5905 (N_5905,N_5630,N_5707);
xor U5906 (N_5906,N_5775,N_5641);
and U5907 (N_5907,N_5702,N_5644);
nand U5908 (N_5908,N_5778,N_5738);
or U5909 (N_5909,N_5697,N_5731);
and U5910 (N_5910,N_5794,N_5706);
or U5911 (N_5911,N_5665,N_5775);
xor U5912 (N_5912,N_5690,N_5624);
xnor U5913 (N_5913,N_5734,N_5643);
nor U5914 (N_5914,N_5705,N_5663);
nor U5915 (N_5915,N_5638,N_5743);
xnor U5916 (N_5916,N_5644,N_5700);
xor U5917 (N_5917,N_5602,N_5708);
or U5918 (N_5918,N_5602,N_5716);
nor U5919 (N_5919,N_5673,N_5700);
nand U5920 (N_5920,N_5725,N_5608);
nor U5921 (N_5921,N_5741,N_5757);
xnor U5922 (N_5922,N_5695,N_5694);
and U5923 (N_5923,N_5656,N_5724);
xor U5924 (N_5924,N_5639,N_5789);
nor U5925 (N_5925,N_5719,N_5722);
or U5926 (N_5926,N_5753,N_5744);
nor U5927 (N_5927,N_5697,N_5797);
and U5928 (N_5928,N_5795,N_5771);
nor U5929 (N_5929,N_5672,N_5798);
and U5930 (N_5930,N_5691,N_5760);
nor U5931 (N_5931,N_5789,N_5628);
or U5932 (N_5932,N_5695,N_5680);
nor U5933 (N_5933,N_5756,N_5610);
nand U5934 (N_5934,N_5741,N_5655);
and U5935 (N_5935,N_5631,N_5666);
and U5936 (N_5936,N_5663,N_5617);
or U5937 (N_5937,N_5733,N_5653);
nor U5938 (N_5938,N_5727,N_5757);
nand U5939 (N_5939,N_5773,N_5647);
or U5940 (N_5940,N_5600,N_5687);
nand U5941 (N_5941,N_5664,N_5795);
and U5942 (N_5942,N_5797,N_5773);
xor U5943 (N_5943,N_5794,N_5672);
and U5944 (N_5944,N_5660,N_5624);
and U5945 (N_5945,N_5713,N_5719);
nand U5946 (N_5946,N_5696,N_5780);
nand U5947 (N_5947,N_5671,N_5723);
nor U5948 (N_5948,N_5739,N_5772);
xnor U5949 (N_5949,N_5666,N_5778);
or U5950 (N_5950,N_5797,N_5736);
or U5951 (N_5951,N_5699,N_5779);
and U5952 (N_5952,N_5704,N_5758);
nand U5953 (N_5953,N_5701,N_5662);
nand U5954 (N_5954,N_5635,N_5737);
nand U5955 (N_5955,N_5784,N_5625);
and U5956 (N_5956,N_5708,N_5614);
nand U5957 (N_5957,N_5691,N_5786);
nor U5958 (N_5958,N_5713,N_5706);
xnor U5959 (N_5959,N_5726,N_5678);
nor U5960 (N_5960,N_5770,N_5617);
or U5961 (N_5961,N_5695,N_5686);
nand U5962 (N_5962,N_5630,N_5745);
or U5963 (N_5963,N_5685,N_5725);
nor U5964 (N_5964,N_5764,N_5657);
nor U5965 (N_5965,N_5673,N_5682);
and U5966 (N_5966,N_5722,N_5793);
or U5967 (N_5967,N_5783,N_5766);
nand U5968 (N_5968,N_5623,N_5600);
nand U5969 (N_5969,N_5633,N_5667);
nor U5970 (N_5970,N_5766,N_5750);
xor U5971 (N_5971,N_5680,N_5754);
or U5972 (N_5972,N_5635,N_5759);
or U5973 (N_5973,N_5751,N_5673);
nor U5974 (N_5974,N_5603,N_5600);
xor U5975 (N_5975,N_5638,N_5683);
nand U5976 (N_5976,N_5641,N_5761);
xnor U5977 (N_5977,N_5643,N_5674);
nand U5978 (N_5978,N_5779,N_5745);
or U5979 (N_5979,N_5646,N_5762);
nand U5980 (N_5980,N_5771,N_5782);
and U5981 (N_5981,N_5691,N_5747);
or U5982 (N_5982,N_5635,N_5763);
or U5983 (N_5983,N_5627,N_5687);
nand U5984 (N_5984,N_5769,N_5799);
or U5985 (N_5985,N_5611,N_5718);
or U5986 (N_5986,N_5781,N_5603);
nand U5987 (N_5987,N_5682,N_5709);
nor U5988 (N_5988,N_5649,N_5683);
nor U5989 (N_5989,N_5691,N_5677);
nand U5990 (N_5990,N_5636,N_5724);
nor U5991 (N_5991,N_5705,N_5762);
or U5992 (N_5992,N_5771,N_5752);
nand U5993 (N_5993,N_5795,N_5701);
nor U5994 (N_5994,N_5760,N_5667);
nor U5995 (N_5995,N_5750,N_5665);
nand U5996 (N_5996,N_5787,N_5627);
xnor U5997 (N_5997,N_5700,N_5772);
xor U5998 (N_5998,N_5736,N_5779);
nor U5999 (N_5999,N_5711,N_5728);
nor U6000 (N_6000,N_5842,N_5919);
and U6001 (N_6001,N_5858,N_5966);
nor U6002 (N_6002,N_5940,N_5934);
and U6003 (N_6003,N_5949,N_5849);
nor U6004 (N_6004,N_5972,N_5862);
xor U6005 (N_6005,N_5837,N_5938);
or U6006 (N_6006,N_5999,N_5816);
nand U6007 (N_6007,N_5846,N_5922);
nand U6008 (N_6008,N_5803,N_5825);
nand U6009 (N_6009,N_5833,N_5848);
or U6010 (N_6010,N_5933,N_5948);
nor U6011 (N_6011,N_5841,N_5988);
nand U6012 (N_6012,N_5958,N_5869);
and U6013 (N_6013,N_5900,N_5992);
nand U6014 (N_6014,N_5895,N_5804);
nor U6015 (N_6015,N_5979,N_5888);
xor U6016 (N_6016,N_5935,N_5964);
xor U6017 (N_6017,N_5822,N_5814);
and U6018 (N_6018,N_5856,N_5960);
and U6019 (N_6019,N_5823,N_5834);
nand U6020 (N_6020,N_5835,N_5830);
xnor U6021 (N_6021,N_5892,N_5886);
and U6022 (N_6022,N_5929,N_5985);
nor U6023 (N_6023,N_5957,N_5893);
nor U6024 (N_6024,N_5954,N_5991);
xnor U6025 (N_6025,N_5855,N_5916);
or U6026 (N_6026,N_5950,N_5800);
nand U6027 (N_6027,N_5959,N_5826);
or U6028 (N_6028,N_5824,N_5990);
xnor U6029 (N_6029,N_5889,N_5928);
nand U6030 (N_6030,N_5965,N_5801);
xor U6031 (N_6031,N_5831,N_5983);
nor U6032 (N_6032,N_5993,N_5820);
and U6033 (N_6033,N_5945,N_5807);
xor U6034 (N_6034,N_5978,N_5953);
nand U6035 (N_6035,N_5998,N_5894);
xor U6036 (N_6036,N_5989,N_5976);
nand U6037 (N_6037,N_5844,N_5917);
nor U6038 (N_6038,N_5829,N_5875);
nor U6039 (N_6039,N_5936,N_5802);
nor U6040 (N_6040,N_5840,N_5812);
nand U6041 (N_6041,N_5836,N_5977);
xor U6042 (N_6042,N_5881,N_5912);
nand U6043 (N_6043,N_5963,N_5969);
xnor U6044 (N_6044,N_5995,N_5974);
xnor U6045 (N_6045,N_5821,N_5808);
nand U6046 (N_6046,N_5868,N_5874);
and U6047 (N_6047,N_5890,N_5818);
xor U6048 (N_6048,N_5891,N_5904);
or U6049 (N_6049,N_5984,N_5975);
or U6050 (N_6050,N_5867,N_5902);
nand U6051 (N_6051,N_5806,N_5864);
and U6052 (N_6052,N_5878,N_5882);
and U6053 (N_6053,N_5817,N_5968);
nand U6054 (N_6054,N_5914,N_5896);
xor U6055 (N_6055,N_5986,N_5947);
nand U6056 (N_6056,N_5910,N_5982);
or U6057 (N_6057,N_5997,N_5839);
nand U6058 (N_6058,N_5926,N_5897);
and U6059 (N_6059,N_5908,N_5939);
and U6060 (N_6060,N_5981,N_5930);
and U6061 (N_6061,N_5887,N_5827);
and U6062 (N_6062,N_5944,N_5937);
nor U6063 (N_6063,N_5907,N_5845);
and U6064 (N_6064,N_5877,N_5927);
nand U6065 (N_6065,N_5838,N_5854);
or U6066 (N_6066,N_5946,N_5857);
nand U6067 (N_6067,N_5859,N_5961);
and U6068 (N_6068,N_5870,N_5925);
or U6069 (N_6069,N_5913,N_5880);
nand U6070 (N_6070,N_5819,N_5847);
xnor U6071 (N_6071,N_5885,N_5962);
or U6072 (N_6072,N_5941,N_5918);
and U6073 (N_6073,N_5852,N_5850);
or U6074 (N_6074,N_5865,N_5805);
and U6075 (N_6075,N_5876,N_5921);
nand U6076 (N_6076,N_5899,N_5905);
xor U6077 (N_6077,N_5923,N_5872);
or U6078 (N_6078,N_5873,N_5863);
xnor U6079 (N_6079,N_5903,N_5915);
and U6080 (N_6080,N_5898,N_5956);
or U6081 (N_6081,N_5860,N_5955);
nand U6082 (N_6082,N_5906,N_5951);
nand U6083 (N_6083,N_5815,N_5970);
or U6084 (N_6084,N_5920,N_5909);
nand U6085 (N_6085,N_5843,N_5943);
xor U6086 (N_6086,N_5996,N_5967);
and U6087 (N_6087,N_5942,N_5987);
nor U6088 (N_6088,N_5809,N_5811);
xor U6089 (N_6089,N_5813,N_5883);
nor U6090 (N_6090,N_5911,N_5871);
or U6091 (N_6091,N_5994,N_5932);
xnor U6092 (N_6092,N_5952,N_5879);
nand U6093 (N_6093,N_5971,N_5924);
nor U6094 (N_6094,N_5810,N_5901);
xnor U6095 (N_6095,N_5866,N_5973);
and U6096 (N_6096,N_5861,N_5884);
or U6097 (N_6097,N_5828,N_5980);
or U6098 (N_6098,N_5931,N_5853);
nor U6099 (N_6099,N_5832,N_5851);
and U6100 (N_6100,N_5942,N_5924);
xor U6101 (N_6101,N_5969,N_5812);
or U6102 (N_6102,N_5833,N_5980);
xor U6103 (N_6103,N_5851,N_5805);
xnor U6104 (N_6104,N_5806,N_5909);
and U6105 (N_6105,N_5927,N_5875);
and U6106 (N_6106,N_5818,N_5943);
and U6107 (N_6107,N_5952,N_5899);
or U6108 (N_6108,N_5930,N_5931);
and U6109 (N_6109,N_5968,N_5865);
xor U6110 (N_6110,N_5869,N_5851);
and U6111 (N_6111,N_5930,N_5824);
or U6112 (N_6112,N_5939,N_5896);
and U6113 (N_6113,N_5802,N_5814);
nor U6114 (N_6114,N_5875,N_5937);
nand U6115 (N_6115,N_5807,N_5995);
and U6116 (N_6116,N_5940,N_5888);
xor U6117 (N_6117,N_5887,N_5830);
xnor U6118 (N_6118,N_5942,N_5925);
xor U6119 (N_6119,N_5810,N_5941);
nor U6120 (N_6120,N_5850,N_5802);
nand U6121 (N_6121,N_5940,N_5821);
xnor U6122 (N_6122,N_5838,N_5885);
nor U6123 (N_6123,N_5854,N_5951);
nand U6124 (N_6124,N_5991,N_5992);
nor U6125 (N_6125,N_5922,N_5930);
nor U6126 (N_6126,N_5876,N_5810);
nor U6127 (N_6127,N_5879,N_5987);
or U6128 (N_6128,N_5899,N_5975);
nor U6129 (N_6129,N_5996,N_5810);
and U6130 (N_6130,N_5811,N_5954);
nand U6131 (N_6131,N_5894,N_5831);
or U6132 (N_6132,N_5819,N_5869);
nor U6133 (N_6133,N_5980,N_5979);
xnor U6134 (N_6134,N_5839,N_5988);
xor U6135 (N_6135,N_5933,N_5902);
and U6136 (N_6136,N_5873,N_5909);
nor U6137 (N_6137,N_5979,N_5977);
nand U6138 (N_6138,N_5821,N_5951);
or U6139 (N_6139,N_5871,N_5800);
xor U6140 (N_6140,N_5919,N_5924);
and U6141 (N_6141,N_5842,N_5947);
and U6142 (N_6142,N_5852,N_5821);
and U6143 (N_6143,N_5881,N_5846);
nand U6144 (N_6144,N_5985,N_5948);
and U6145 (N_6145,N_5801,N_5871);
or U6146 (N_6146,N_5837,N_5883);
nand U6147 (N_6147,N_5918,N_5858);
or U6148 (N_6148,N_5834,N_5964);
and U6149 (N_6149,N_5873,N_5858);
nand U6150 (N_6150,N_5898,N_5868);
nand U6151 (N_6151,N_5970,N_5906);
nor U6152 (N_6152,N_5810,N_5838);
nand U6153 (N_6153,N_5989,N_5862);
and U6154 (N_6154,N_5994,N_5922);
nor U6155 (N_6155,N_5972,N_5930);
nand U6156 (N_6156,N_5802,N_5867);
nor U6157 (N_6157,N_5857,N_5994);
nor U6158 (N_6158,N_5828,N_5863);
xor U6159 (N_6159,N_5873,N_5929);
or U6160 (N_6160,N_5963,N_5955);
nor U6161 (N_6161,N_5876,N_5959);
nand U6162 (N_6162,N_5952,N_5837);
or U6163 (N_6163,N_5995,N_5851);
or U6164 (N_6164,N_5965,N_5936);
nand U6165 (N_6165,N_5812,N_5982);
and U6166 (N_6166,N_5883,N_5976);
nand U6167 (N_6167,N_5831,N_5804);
or U6168 (N_6168,N_5890,N_5991);
or U6169 (N_6169,N_5887,N_5915);
nand U6170 (N_6170,N_5960,N_5902);
nor U6171 (N_6171,N_5902,N_5840);
xnor U6172 (N_6172,N_5955,N_5945);
nand U6173 (N_6173,N_5899,N_5902);
nor U6174 (N_6174,N_5931,N_5857);
xor U6175 (N_6175,N_5985,N_5811);
xor U6176 (N_6176,N_5883,N_5833);
nor U6177 (N_6177,N_5877,N_5806);
xor U6178 (N_6178,N_5946,N_5923);
nand U6179 (N_6179,N_5842,N_5971);
xor U6180 (N_6180,N_5991,N_5834);
nand U6181 (N_6181,N_5836,N_5930);
and U6182 (N_6182,N_5850,N_5812);
or U6183 (N_6183,N_5917,N_5835);
nor U6184 (N_6184,N_5990,N_5875);
or U6185 (N_6185,N_5829,N_5899);
or U6186 (N_6186,N_5894,N_5917);
nor U6187 (N_6187,N_5960,N_5853);
xor U6188 (N_6188,N_5829,N_5912);
nor U6189 (N_6189,N_5877,N_5836);
nand U6190 (N_6190,N_5924,N_5805);
xnor U6191 (N_6191,N_5955,N_5831);
xor U6192 (N_6192,N_5957,N_5830);
xor U6193 (N_6193,N_5979,N_5852);
xor U6194 (N_6194,N_5993,N_5865);
xnor U6195 (N_6195,N_5960,N_5835);
xnor U6196 (N_6196,N_5816,N_5957);
and U6197 (N_6197,N_5948,N_5958);
and U6198 (N_6198,N_5878,N_5991);
nor U6199 (N_6199,N_5995,N_5909);
and U6200 (N_6200,N_6174,N_6096);
and U6201 (N_6201,N_6143,N_6038);
nand U6202 (N_6202,N_6193,N_6065);
nor U6203 (N_6203,N_6135,N_6125);
nor U6204 (N_6204,N_6127,N_6072);
and U6205 (N_6205,N_6134,N_6025);
nand U6206 (N_6206,N_6045,N_6027);
or U6207 (N_6207,N_6163,N_6067);
nor U6208 (N_6208,N_6006,N_6020);
nor U6209 (N_6209,N_6001,N_6106);
and U6210 (N_6210,N_6121,N_6021);
or U6211 (N_6211,N_6153,N_6084);
xor U6212 (N_6212,N_6179,N_6026);
nand U6213 (N_6213,N_6181,N_6109);
or U6214 (N_6214,N_6172,N_6114);
nand U6215 (N_6215,N_6090,N_6036);
or U6216 (N_6216,N_6095,N_6047);
or U6217 (N_6217,N_6183,N_6008);
nand U6218 (N_6218,N_6080,N_6178);
or U6219 (N_6219,N_6137,N_6188);
nor U6220 (N_6220,N_6175,N_6159);
nor U6221 (N_6221,N_6037,N_6171);
and U6222 (N_6222,N_6165,N_6151);
nor U6223 (N_6223,N_6166,N_6197);
or U6224 (N_6224,N_6056,N_6030);
nor U6225 (N_6225,N_6075,N_6046);
nor U6226 (N_6226,N_6051,N_6004);
or U6227 (N_6227,N_6053,N_6060);
xor U6228 (N_6228,N_6156,N_6071);
nor U6229 (N_6229,N_6005,N_6083);
nand U6230 (N_6230,N_6070,N_6044);
xnor U6231 (N_6231,N_6140,N_6184);
xnor U6232 (N_6232,N_6032,N_6187);
xnor U6233 (N_6233,N_6118,N_6009);
nand U6234 (N_6234,N_6170,N_6113);
xnor U6235 (N_6235,N_6155,N_6150);
nand U6236 (N_6236,N_6099,N_6043);
nand U6237 (N_6237,N_6057,N_6198);
and U6238 (N_6238,N_6079,N_6119);
nor U6239 (N_6239,N_6182,N_6161);
xnor U6240 (N_6240,N_6112,N_6018);
nand U6241 (N_6241,N_6066,N_6139);
nor U6242 (N_6242,N_6128,N_6138);
xnor U6243 (N_6243,N_6039,N_6033);
xnor U6244 (N_6244,N_6035,N_6194);
xnor U6245 (N_6245,N_6063,N_6152);
xor U6246 (N_6246,N_6015,N_6048);
or U6247 (N_6247,N_6164,N_6074);
nor U6248 (N_6248,N_6031,N_6000);
and U6249 (N_6249,N_6133,N_6011);
nor U6250 (N_6250,N_6028,N_6185);
xor U6251 (N_6251,N_6107,N_6129);
xnor U6252 (N_6252,N_6052,N_6126);
or U6253 (N_6253,N_6042,N_6040);
xnor U6254 (N_6254,N_6029,N_6061);
or U6255 (N_6255,N_6136,N_6131);
nor U6256 (N_6256,N_6007,N_6154);
nor U6257 (N_6257,N_6017,N_6002);
nor U6258 (N_6258,N_6176,N_6013);
and U6259 (N_6259,N_6093,N_6191);
xnor U6260 (N_6260,N_6082,N_6014);
or U6261 (N_6261,N_6022,N_6196);
xnor U6262 (N_6262,N_6049,N_6024);
nand U6263 (N_6263,N_6087,N_6086);
nor U6264 (N_6264,N_6142,N_6160);
nor U6265 (N_6265,N_6089,N_6103);
nor U6266 (N_6266,N_6173,N_6162);
nand U6267 (N_6267,N_6100,N_6190);
xor U6268 (N_6268,N_6120,N_6122);
nor U6269 (N_6269,N_6157,N_6019);
and U6270 (N_6270,N_6034,N_6144);
and U6271 (N_6271,N_6199,N_6168);
or U6272 (N_6272,N_6062,N_6050);
nand U6273 (N_6273,N_6105,N_6077);
or U6274 (N_6274,N_6069,N_6055);
nand U6275 (N_6275,N_6016,N_6078);
and U6276 (N_6276,N_6130,N_6104);
and U6277 (N_6277,N_6085,N_6023);
and U6278 (N_6278,N_6041,N_6148);
nor U6279 (N_6279,N_6192,N_6094);
and U6280 (N_6280,N_6149,N_6064);
or U6281 (N_6281,N_6110,N_6097);
and U6282 (N_6282,N_6068,N_6124);
or U6283 (N_6283,N_6058,N_6054);
nor U6284 (N_6284,N_6088,N_6177);
nand U6285 (N_6285,N_6167,N_6146);
xnor U6286 (N_6286,N_6092,N_6081);
xor U6287 (N_6287,N_6117,N_6108);
xor U6288 (N_6288,N_6158,N_6180);
or U6289 (N_6289,N_6101,N_6141);
xor U6290 (N_6290,N_6116,N_6169);
nor U6291 (N_6291,N_6102,N_6145);
nor U6292 (N_6292,N_6147,N_6123);
xnor U6293 (N_6293,N_6059,N_6115);
or U6294 (N_6294,N_6076,N_6111);
xor U6295 (N_6295,N_6132,N_6186);
or U6296 (N_6296,N_6012,N_6091);
xnor U6297 (N_6297,N_6010,N_6003);
or U6298 (N_6298,N_6098,N_6195);
and U6299 (N_6299,N_6073,N_6189);
nand U6300 (N_6300,N_6131,N_6125);
and U6301 (N_6301,N_6091,N_6070);
and U6302 (N_6302,N_6081,N_6037);
xnor U6303 (N_6303,N_6104,N_6183);
xor U6304 (N_6304,N_6194,N_6083);
nand U6305 (N_6305,N_6173,N_6177);
or U6306 (N_6306,N_6033,N_6026);
nand U6307 (N_6307,N_6030,N_6017);
nand U6308 (N_6308,N_6116,N_6162);
or U6309 (N_6309,N_6143,N_6186);
nand U6310 (N_6310,N_6174,N_6159);
and U6311 (N_6311,N_6197,N_6009);
nor U6312 (N_6312,N_6141,N_6058);
xor U6313 (N_6313,N_6021,N_6195);
nor U6314 (N_6314,N_6173,N_6113);
xor U6315 (N_6315,N_6028,N_6076);
nor U6316 (N_6316,N_6147,N_6006);
xnor U6317 (N_6317,N_6005,N_6139);
or U6318 (N_6318,N_6164,N_6033);
or U6319 (N_6319,N_6189,N_6116);
xor U6320 (N_6320,N_6184,N_6034);
nand U6321 (N_6321,N_6192,N_6096);
nand U6322 (N_6322,N_6108,N_6114);
nor U6323 (N_6323,N_6108,N_6035);
nor U6324 (N_6324,N_6190,N_6135);
or U6325 (N_6325,N_6038,N_6083);
nand U6326 (N_6326,N_6066,N_6061);
nor U6327 (N_6327,N_6067,N_6049);
nand U6328 (N_6328,N_6137,N_6038);
or U6329 (N_6329,N_6089,N_6142);
and U6330 (N_6330,N_6143,N_6068);
nand U6331 (N_6331,N_6019,N_6058);
nand U6332 (N_6332,N_6025,N_6010);
xor U6333 (N_6333,N_6073,N_6066);
nand U6334 (N_6334,N_6083,N_6185);
xor U6335 (N_6335,N_6083,N_6091);
nor U6336 (N_6336,N_6108,N_6115);
nor U6337 (N_6337,N_6122,N_6117);
xnor U6338 (N_6338,N_6123,N_6048);
or U6339 (N_6339,N_6018,N_6081);
nand U6340 (N_6340,N_6022,N_6045);
and U6341 (N_6341,N_6084,N_6118);
nand U6342 (N_6342,N_6129,N_6152);
or U6343 (N_6343,N_6091,N_6082);
nand U6344 (N_6344,N_6194,N_6172);
or U6345 (N_6345,N_6036,N_6180);
xnor U6346 (N_6346,N_6178,N_6060);
xor U6347 (N_6347,N_6019,N_6163);
or U6348 (N_6348,N_6108,N_6052);
xor U6349 (N_6349,N_6036,N_6033);
or U6350 (N_6350,N_6120,N_6112);
and U6351 (N_6351,N_6131,N_6121);
nand U6352 (N_6352,N_6050,N_6098);
or U6353 (N_6353,N_6076,N_6167);
nor U6354 (N_6354,N_6119,N_6173);
and U6355 (N_6355,N_6004,N_6118);
xor U6356 (N_6356,N_6055,N_6039);
or U6357 (N_6357,N_6092,N_6084);
or U6358 (N_6358,N_6116,N_6049);
nand U6359 (N_6359,N_6015,N_6088);
or U6360 (N_6360,N_6118,N_6032);
or U6361 (N_6361,N_6024,N_6074);
nor U6362 (N_6362,N_6031,N_6170);
nor U6363 (N_6363,N_6036,N_6028);
nand U6364 (N_6364,N_6163,N_6168);
and U6365 (N_6365,N_6058,N_6084);
or U6366 (N_6366,N_6156,N_6045);
and U6367 (N_6367,N_6045,N_6021);
nand U6368 (N_6368,N_6115,N_6161);
nand U6369 (N_6369,N_6036,N_6056);
nand U6370 (N_6370,N_6028,N_6166);
xor U6371 (N_6371,N_6199,N_6083);
and U6372 (N_6372,N_6015,N_6130);
nor U6373 (N_6373,N_6106,N_6151);
nor U6374 (N_6374,N_6128,N_6168);
or U6375 (N_6375,N_6176,N_6112);
and U6376 (N_6376,N_6067,N_6150);
or U6377 (N_6377,N_6073,N_6053);
or U6378 (N_6378,N_6133,N_6042);
or U6379 (N_6379,N_6070,N_6004);
nand U6380 (N_6380,N_6072,N_6182);
nor U6381 (N_6381,N_6013,N_6050);
xnor U6382 (N_6382,N_6099,N_6018);
and U6383 (N_6383,N_6115,N_6020);
and U6384 (N_6384,N_6183,N_6128);
nor U6385 (N_6385,N_6038,N_6035);
nor U6386 (N_6386,N_6076,N_6164);
nand U6387 (N_6387,N_6048,N_6068);
or U6388 (N_6388,N_6088,N_6146);
or U6389 (N_6389,N_6058,N_6032);
or U6390 (N_6390,N_6188,N_6152);
and U6391 (N_6391,N_6077,N_6151);
nand U6392 (N_6392,N_6012,N_6110);
xor U6393 (N_6393,N_6146,N_6001);
nand U6394 (N_6394,N_6135,N_6155);
and U6395 (N_6395,N_6179,N_6137);
xnor U6396 (N_6396,N_6190,N_6169);
xnor U6397 (N_6397,N_6051,N_6176);
xor U6398 (N_6398,N_6184,N_6033);
or U6399 (N_6399,N_6177,N_6174);
and U6400 (N_6400,N_6207,N_6341);
nor U6401 (N_6401,N_6285,N_6383);
xnor U6402 (N_6402,N_6370,N_6240);
and U6403 (N_6403,N_6342,N_6313);
nor U6404 (N_6404,N_6312,N_6261);
xnor U6405 (N_6405,N_6388,N_6321);
nor U6406 (N_6406,N_6288,N_6319);
nand U6407 (N_6407,N_6354,N_6286);
nor U6408 (N_6408,N_6304,N_6332);
nand U6409 (N_6409,N_6396,N_6365);
nand U6410 (N_6410,N_6291,N_6367);
or U6411 (N_6411,N_6298,N_6376);
and U6412 (N_6412,N_6346,N_6248);
nand U6413 (N_6413,N_6275,N_6267);
nand U6414 (N_6414,N_6391,N_6315);
nand U6415 (N_6415,N_6379,N_6329);
nor U6416 (N_6416,N_6307,N_6395);
and U6417 (N_6417,N_6302,N_6347);
xor U6418 (N_6418,N_6293,N_6399);
and U6419 (N_6419,N_6340,N_6363);
or U6420 (N_6420,N_6299,N_6361);
nor U6421 (N_6421,N_6280,N_6355);
xnor U6422 (N_6422,N_6227,N_6328);
nand U6423 (N_6423,N_6330,N_6234);
and U6424 (N_6424,N_6331,N_6335);
and U6425 (N_6425,N_6366,N_6200);
and U6426 (N_6426,N_6238,N_6325);
xnor U6427 (N_6427,N_6343,N_6274);
nor U6428 (N_6428,N_6359,N_6231);
or U6429 (N_6429,N_6219,N_6271);
nor U6430 (N_6430,N_6289,N_6351);
nor U6431 (N_6431,N_6323,N_6392);
nand U6432 (N_6432,N_6226,N_6237);
nor U6433 (N_6433,N_6345,N_6389);
and U6434 (N_6434,N_6322,N_6386);
and U6435 (N_6435,N_6202,N_6301);
and U6436 (N_6436,N_6320,N_6239);
or U6437 (N_6437,N_6260,N_6310);
nor U6438 (N_6438,N_6225,N_6296);
or U6439 (N_6439,N_6308,N_6277);
or U6440 (N_6440,N_6352,N_6244);
and U6441 (N_6441,N_6327,N_6257);
nor U6442 (N_6442,N_6263,N_6201);
or U6443 (N_6443,N_6210,N_6373);
and U6444 (N_6444,N_6394,N_6372);
and U6445 (N_6445,N_6282,N_6243);
xnor U6446 (N_6446,N_6242,N_6316);
and U6447 (N_6447,N_6295,N_6269);
nand U6448 (N_6448,N_6259,N_6362);
nor U6449 (N_6449,N_6393,N_6306);
or U6450 (N_6450,N_6254,N_6297);
nor U6451 (N_6451,N_6222,N_6357);
nor U6452 (N_6452,N_6378,N_6369);
or U6453 (N_6453,N_6235,N_6223);
and U6454 (N_6454,N_6314,N_6266);
or U6455 (N_6455,N_6337,N_6236);
nand U6456 (N_6456,N_6245,N_6318);
or U6457 (N_6457,N_6317,N_6281);
and U6458 (N_6458,N_6270,N_6348);
or U6459 (N_6459,N_6387,N_6212);
nor U6460 (N_6460,N_6249,N_6265);
nand U6461 (N_6461,N_6213,N_6206);
nand U6462 (N_6462,N_6283,N_6349);
nor U6463 (N_6463,N_6217,N_6334);
nor U6464 (N_6464,N_6204,N_6233);
nor U6465 (N_6465,N_6374,N_6276);
xnor U6466 (N_6466,N_6264,N_6255);
and U6467 (N_6467,N_6303,N_6380);
nand U6468 (N_6468,N_6384,N_6272);
nor U6469 (N_6469,N_6398,N_6252);
xor U6470 (N_6470,N_6287,N_6230);
or U6471 (N_6471,N_6382,N_6333);
nand U6472 (N_6472,N_6368,N_6358);
nor U6473 (N_6473,N_6221,N_6326);
nand U6474 (N_6474,N_6256,N_6253);
and U6475 (N_6475,N_6350,N_6228);
xor U6476 (N_6476,N_6284,N_6375);
or U6477 (N_6477,N_6353,N_6209);
xnor U6478 (N_6478,N_6324,N_6279);
nand U6479 (N_6479,N_6339,N_6205);
and U6480 (N_6480,N_6220,N_6224);
xor U6481 (N_6481,N_6229,N_6397);
xnor U6482 (N_6482,N_6273,N_6338);
nand U6483 (N_6483,N_6294,N_6377);
nor U6484 (N_6484,N_6215,N_6216);
and U6485 (N_6485,N_6390,N_6246);
and U6486 (N_6486,N_6311,N_6344);
nand U6487 (N_6487,N_6211,N_6262);
nor U6488 (N_6488,N_6364,N_6300);
and U6489 (N_6489,N_6241,N_6305);
nor U6490 (N_6490,N_6203,N_6214);
and U6491 (N_6491,N_6232,N_6336);
xor U6492 (N_6492,N_6268,N_6371);
xnor U6493 (N_6493,N_6290,N_6356);
or U6494 (N_6494,N_6278,N_6292);
xor U6495 (N_6495,N_6251,N_6309);
xor U6496 (N_6496,N_6385,N_6258);
or U6497 (N_6497,N_6360,N_6250);
or U6498 (N_6498,N_6208,N_6247);
and U6499 (N_6499,N_6218,N_6381);
nand U6500 (N_6500,N_6251,N_6295);
xnor U6501 (N_6501,N_6240,N_6230);
nand U6502 (N_6502,N_6291,N_6256);
nor U6503 (N_6503,N_6212,N_6203);
and U6504 (N_6504,N_6341,N_6393);
and U6505 (N_6505,N_6354,N_6324);
and U6506 (N_6506,N_6204,N_6223);
xor U6507 (N_6507,N_6314,N_6262);
and U6508 (N_6508,N_6306,N_6297);
nand U6509 (N_6509,N_6267,N_6265);
nor U6510 (N_6510,N_6356,N_6203);
and U6511 (N_6511,N_6229,N_6360);
and U6512 (N_6512,N_6282,N_6335);
or U6513 (N_6513,N_6239,N_6389);
or U6514 (N_6514,N_6224,N_6334);
nand U6515 (N_6515,N_6292,N_6398);
nor U6516 (N_6516,N_6356,N_6347);
and U6517 (N_6517,N_6326,N_6238);
xor U6518 (N_6518,N_6243,N_6337);
and U6519 (N_6519,N_6205,N_6287);
or U6520 (N_6520,N_6263,N_6258);
xor U6521 (N_6521,N_6262,N_6321);
nand U6522 (N_6522,N_6289,N_6366);
or U6523 (N_6523,N_6270,N_6274);
nand U6524 (N_6524,N_6252,N_6217);
nand U6525 (N_6525,N_6396,N_6271);
nand U6526 (N_6526,N_6238,N_6319);
xnor U6527 (N_6527,N_6323,N_6373);
nor U6528 (N_6528,N_6367,N_6389);
nand U6529 (N_6529,N_6291,N_6331);
or U6530 (N_6530,N_6209,N_6260);
nor U6531 (N_6531,N_6201,N_6297);
and U6532 (N_6532,N_6380,N_6385);
nor U6533 (N_6533,N_6218,N_6345);
and U6534 (N_6534,N_6349,N_6336);
xnor U6535 (N_6535,N_6373,N_6221);
or U6536 (N_6536,N_6304,N_6352);
and U6537 (N_6537,N_6279,N_6317);
or U6538 (N_6538,N_6342,N_6347);
nor U6539 (N_6539,N_6231,N_6288);
nor U6540 (N_6540,N_6316,N_6284);
xnor U6541 (N_6541,N_6374,N_6205);
nor U6542 (N_6542,N_6386,N_6261);
xor U6543 (N_6543,N_6314,N_6272);
nor U6544 (N_6544,N_6292,N_6228);
nor U6545 (N_6545,N_6298,N_6290);
or U6546 (N_6546,N_6259,N_6384);
xnor U6547 (N_6547,N_6356,N_6298);
nand U6548 (N_6548,N_6313,N_6353);
nand U6549 (N_6549,N_6313,N_6330);
nor U6550 (N_6550,N_6226,N_6240);
and U6551 (N_6551,N_6215,N_6276);
xor U6552 (N_6552,N_6303,N_6295);
nor U6553 (N_6553,N_6364,N_6207);
or U6554 (N_6554,N_6339,N_6331);
or U6555 (N_6555,N_6210,N_6310);
xor U6556 (N_6556,N_6249,N_6202);
nor U6557 (N_6557,N_6241,N_6213);
or U6558 (N_6558,N_6207,N_6208);
or U6559 (N_6559,N_6302,N_6256);
or U6560 (N_6560,N_6240,N_6305);
nor U6561 (N_6561,N_6379,N_6284);
nand U6562 (N_6562,N_6327,N_6331);
or U6563 (N_6563,N_6232,N_6295);
or U6564 (N_6564,N_6200,N_6313);
and U6565 (N_6565,N_6397,N_6284);
or U6566 (N_6566,N_6384,N_6200);
or U6567 (N_6567,N_6338,N_6208);
nand U6568 (N_6568,N_6318,N_6398);
nand U6569 (N_6569,N_6308,N_6314);
and U6570 (N_6570,N_6311,N_6381);
and U6571 (N_6571,N_6223,N_6394);
nand U6572 (N_6572,N_6252,N_6230);
or U6573 (N_6573,N_6284,N_6355);
nor U6574 (N_6574,N_6381,N_6226);
and U6575 (N_6575,N_6340,N_6318);
nor U6576 (N_6576,N_6346,N_6387);
nor U6577 (N_6577,N_6245,N_6368);
and U6578 (N_6578,N_6340,N_6372);
and U6579 (N_6579,N_6294,N_6359);
nand U6580 (N_6580,N_6237,N_6212);
or U6581 (N_6581,N_6382,N_6244);
nor U6582 (N_6582,N_6332,N_6218);
xor U6583 (N_6583,N_6296,N_6216);
or U6584 (N_6584,N_6257,N_6359);
xnor U6585 (N_6585,N_6274,N_6301);
xnor U6586 (N_6586,N_6250,N_6396);
xnor U6587 (N_6587,N_6288,N_6334);
or U6588 (N_6588,N_6375,N_6257);
nand U6589 (N_6589,N_6276,N_6350);
nand U6590 (N_6590,N_6209,N_6225);
and U6591 (N_6591,N_6267,N_6309);
or U6592 (N_6592,N_6288,N_6209);
xor U6593 (N_6593,N_6209,N_6299);
and U6594 (N_6594,N_6297,N_6312);
nor U6595 (N_6595,N_6285,N_6330);
nand U6596 (N_6596,N_6337,N_6308);
or U6597 (N_6597,N_6258,N_6379);
and U6598 (N_6598,N_6365,N_6296);
and U6599 (N_6599,N_6336,N_6324);
and U6600 (N_6600,N_6556,N_6564);
xnor U6601 (N_6601,N_6565,N_6569);
xnor U6602 (N_6602,N_6487,N_6401);
xnor U6603 (N_6603,N_6438,N_6473);
nand U6604 (N_6604,N_6446,N_6496);
nor U6605 (N_6605,N_6493,N_6557);
and U6606 (N_6606,N_6509,N_6434);
nor U6607 (N_6607,N_6422,N_6583);
nor U6608 (N_6608,N_6550,N_6460);
xor U6609 (N_6609,N_6436,N_6406);
nand U6610 (N_6610,N_6539,N_6545);
and U6611 (N_6611,N_6408,N_6510);
nor U6612 (N_6612,N_6497,N_6423);
xor U6613 (N_6613,N_6536,N_6570);
xor U6614 (N_6614,N_6575,N_6532);
nor U6615 (N_6615,N_6471,N_6571);
nor U6616 (N_6616,N_6531,N_6538);
nand U6617 (N_6617,N_6498,N_6561);
and U6618 (N_6618,N_6594,N_6522);
xor U6619 (N_6619,N_6519,N_6502);
or U6620 (N_6620,N_6407,N_6439);
nor U6621 (N_6621,N_6530,N_6523);
xnor U6622 (N_6622,N_6574,N_6511);
and U6623 (N_6623,N_6578,N_6587);
or U6624 (N_6624,N_6433,N_6428);
xnor U6625 (N_6625,N_6430,N_6489);
nand U6626 (N_6626,N_6466,N_6485);
nor U6627 (N_6627,N_6567,N_6520);
nor U6628 (N_6628,N_6592,N_6475);
nand U6629 (N_6629,N_6589,N_6596);
xor U6630 (N_6630,N_6400,N_6590);
nand U6631 (N_6631,N_6529,N_6560);
xnor U6632 (N_6632,N_6413,N_6443);
nand U6633 (N_6633,N_6504,N_6426);
nor U6634 (N_6634,N_6593,N_6465);
xnor U6635 (N_6635,N_6459,N_6470);
nor U6636 (N_6636,N_6537,N_6432);
nand U6637 (N_6637,N_6444,N_6427);
xor U6638 (N_6638,N_6449,N_6452);
and U6639 (N_6639,N_6479,N_6552);
nand U6640 (N_6640,N_6492,N_6563);
xor U6641 (N_6641,N_6483,N_6597);
xor U6642 (N_6642,N_6464,N_6462);
nor U6643 (N_6643,N_6468,N_6453);
nand U6644 (N_6644,N_6541,N_6416);
nor U6645 (N_6645,N_6461,N_6458);
nor U6646 (N_6646,N_6418,N_6580);
and U6647 (N_6647,N_6481,N_6548);
nand U6648 (N_6648,N_6478,N_6573);
and U6649 (N_6649,N_6533,N_6424);
nor U6650 (N_6650,N_6405,N_6599);
and U6651 (N_6651,N_6513,N_6429);
nand U6652 (N_6652,N_6451,N_6534);
nand U6653 (N_6653,N_6546,N_6448);
nand U6654 (N_6654,N_6568,N_6577);
and U6655 (N_6655,N_6581,N_6445);
nand U6656 (N_6656,N_6467,N_6490);
nand U6657 (N_6657,N_6456,N_6566);
and U6658 (N_6658,N_6501,N_6525);
nand U6659 (N_6659,N_6527,N_6404);
nor U6660 (N_6660,N_6572,N_6480);
xor U6661 (N_6661,N_6421,N_6457);
and U6662 (N_6662,N_6559,N_6474);
xnor U6663 (N_6663,N_6584,N_6484);
nand U6664 (N_6664,N_6402,N_6516);
xor U6665 (N_6665,N_6505,N_6554);
nor U6666 (N_6666,N_6410,N_6476);
nor U6667 (N_6667,N_6591,N_6431);
or U6668 (N_6668,N_6549,N_6415);
nand U6669 (N_6669,N_6488,N_6555);
nor U6670 (N_6670,N_6435,N_6500);
or U6671 (N_6671,N_6437,N_6469);
and U6672 (N_6672,N_6544,N_6472);
or U6673 (N_6673,N_6455,N_6450);
and U6674 (N_6674,N_6526,N_6414);
and U6675 (N_6675,N_6576,N_6551);
or U6676 (N_6676,N_6442,N_6585);
xor U6677 (N_6677,N_6409,N_6558);
nor U6678 (N_6678,N_6412,N_6582);
xnor U6679 (N_6679,N_6507,N_6540);
and U6680 (N_6680,N_6528,N_6482);
nor U6681 (N_6681,N_6562,N_6420);
nand U6682 (N_6682,N_6588,N_6447);
xor U6683 (N_6683,N_6515,N_6411);
and U6684 (N_6684,N_6543,N_6579);
xor U6685 (N_6685,N_6495,N_6512);
or U6686 (N_6686,N_6506,N_6518);
xor U6687 (N_6687,N_6524,N_6598);
and U6688 (N_6688,N_6517,N_6441);
nor U6689 (N_6689,N_6494,N_6477);
xnor U6690 (N_6690,N_6542,N_6499);
or U6691 (N_6691,N_6503,N_6547);
and U6692 (N_6692,N_6486,N_6491);
nand U6693 (N_6693,N_6403,N_6595);
nor U6694 (N_6694,N_6508,N_6514);
or U6695 (N_6695,N_6425,N_6535);
and U6696 (N_6696,N_6553,N_6586);
nor U6697 (N_6697,N_6419,N_6463);
nor U6698 (N_6698,N_6521,N_6440);
or U6699 (N_6699,N_6454,N_6417);
or U6700 (N_6700,N_6598,N_6487);
nand U6701 (N_6701,N_6422,N_6410);
xnor U6702 (N_6702,N_6438,N_6572);
nand U6703 (N_6703,N_6458,N_6498);
and U6704 (N_6704,N_6450,N_6548);
nor U6705 (N_6705,N_6471,N_6516);
and U6706 (N_6706,N_6456,N_6401);
or U6707 (N_6707,N_6550,N_6490);
or U6708 (N_6708,N_6579,N_6544);
nor U6709 (N_6709,N_6566,N_6427);
nor U6710 (N_6710,N_6501,N_6493);
nor U6711 (N_6711,N_6562,N_6468);
xor U6712 (N_6712,N_6507,N_6452);
xor U6713 (N_6713,N_6521,N_6444);
nand U6714 (N_6714,N_6577,N_6549);
and U6715 (N_6715,N_6597,N_6519);
nand U6716 (N_6716,N_6577,N_6404);
nand U6717 (N_6717,N_6454,N_6573);
or U6718 (N_6718,N_6580,N_6431);
nor U6719 (N_6719,N_6593,N_6552);
xnor U6720 (N_6720,N_6582,N_6470);
and U6721 (N_6721,N_6449,N_6523);
and U6722 (N_6722,N_6545,N_6416);
and U6723 (N_6723,N_6429,N_6552);
and U6724 (N_6724,N_6523,N_6428);
nor U6725 (N_6725,N_6588,N_6506);
xnor U6726 (N_6726,N_6479,N_6489);
and U6727 (N_6727,N_6439,N_6539);
nor U6728 (N_6728,N_6586,N_6467);
nor U6729 (N_6729,N_6453,N_6488);
and U6730 (N_6730,N_6509,N_6598);
or U6731 (N_6731,N_6463,N_6579);
or U6732 (N_6732,N_6447,N_6415);
nor U6733 (N_6733,N_6507,N_6462);
and U6734 (N_6734,N_6430,N_6461);
nor U6735 (N_6735,N_6494,N_6404);
nor U6736 (N_6736,N_6520,N_6537);
or U6737 (N_6737,N_6574,N_6411);
xor U6738 (N_6738,N_6580,N_6591);
and U6739 (N_6739,N_6524,N_6406);
or U6740 (N_6740,N_6535,N_6424);
or U6741 (N_6741,N_6578,N_6584);
and U6742 (N_6742,N_6451,N_6456);
nand U6743 (N_6743,N_6499,N_6435);
nand U6744 (N_6744,N_6405,N_6588);
or U6745 (N_6745,N_6557,N_6506);
nor U6746 (N_6746,N_6528,N_6479);
and U6747 (N_6747,N_6546,N_6501);
and U6748 (N_6748,N_6432,N_6435);
or U6749 (N_6749,N_6455,N_6540);
xnor U6750 (N_6750,N_6473,N_6550);
nand U6751 (N_6751,N_6440,N_6451);
xnor U6752 (N_6752,N_6531,N_6583);
nand U6753 (N_6753,N_6524,N_6480);
or U6754 (N_6754,N_6481,N_6499);
nand U6755 (N_6755,N_6488,N_6464);
nor U6756 (N_6756,N_6453,N_6590);
xnor U6757 (N_6757,N_6548,N_6492);
xor U6758 (N_6758,N_6492,N_6431);
xnor U6759 (N_6759,N_6404,N_6405);
or U6760 (N_6760,N_6507,N_6420);
nand U6761 (N_6761,N_6574,N_6460);
and U6762 (N_6762,N_6400,N_6553);
nor U6763 (N_6763,N_6449,N_6496);
nand U6764 (N_6764,N_6520,N_6577);
and U6765 (N_6765,N_6470,N_6597);
xor U6766 (N_6766,N_6517,N_6458);
and U6767 (N_6767,N_6402,N_6469);
nand U6768 (N_6768,N_6406,N_6433);
nand U6769 (N_6769,N_6410,N_6432);
nor U6770 (N_6770,N_6570,N_6411);
and U6771 (N_6771,N_6553,N_6560);
xor U6772 (N_6772,N_6560,N_6444);
nand U6773 (N_6773,N_6419,N_6552);
nand U6774 (N_6774,N_6462,N_6495);
and U6775 (N_6775,N_6449,N_6573);
xor U6776 (N_6776,N_6591,N_6469);
nand U6777 (N_6777,N_6417,N_6446);
xor U6778 (N_6778,N_6585,N_6548);
and U6779 (N_6779,N_6463,N_6470);
and U6780 (N_6780,N_6545,N_6419);
nand U6781 (N_6781,N_6531,N_6404);
nor U6782 (N_6782,N_6573,N_6419);
and U6783 (N_6783,N_6456,N_6534);
or U6784 (N_6784,N_6557,N_6483);
or U6785 (N_6785,N_6446,N_6419);
and U6786 (N_6786,N_6417,N_6559);
nor U6787 (N_6787,N_6550,N_6486);
nor U6788 (N_6788,N_6529,N_6400);
nand U6789 (N_6789,N_6417,N_6514);
or U6790 (N_6790,N_6461,N_6515);
or U6791 (N_6791,N_6598,N_6547);
or U6792 (N_6792,N_6503,N_6538);
nand U6793 (N_6793,N_6533,N_6416);
xor U6794 (N_6794,N_6467,N_6492);
and U6795 (N_6795,N_6560,N_6504);
and U6796 (N_6796,N_6450,N_6558);
or U6797 (N_6797,N_6494,N_6585);
nand U6798 (N_6798,N_6427,N_6440);
nand U6799 (N_6799,N_6513,N_6599);
and U6800 (N_6800,N_6662,N_6693);
or U6801 (N_6801,N_6698,N_6629);
nor U6802 (N_6802,N_6737,N_6679);
nor U6803 (N_6803,N_6744,N_6617);
and U6804 (N_6804,N_6779,N_6695);
nand U6805 (N_6805,N_6752,N_6783);
nand U6806 (N_6806,N_6720,N_6606);
nor U6807 (N_6807,N_6631,N_6602);
and U6808 (N_6808,N_6769,N_6672);
or U6809 (N_6809,N_6622,N_6642);
or U6810 (N_6810,N_6691,N_6674);
nor U6811 (N_6811,N_6635,N_6730);
xor U6812 (N_6812,N_6636,N_6670);
nand U6813 (N_6813,N_6768,N_6664);
xor U6814 (N_6814,N_6657,N_6767);
nor U6815 (N_6815,N_6648,N_6639);
nand U6816 (N_6816,N_6682,N_6790);
nor U6817 (N_6817,N_6608,N_6623);
xor U6818 (N_6818,N_6668,N_6794);
or U6819 (N_6819,N_6604,N_6641);
and U6820 (N_6820,N_6796,N_6758);
or U6821 (N_6821,N_6683,N_6746);
or U6822 (N_6822,N_6703,N_6605);
or U6823 (N_6823,N_6678,N_6745);
nor U6824 (N_6824,N_6741,N_6694);
nand U6825 (N_6825,N_6675,N_6760);
nor U6826 (N_6826,N_6729,N_6613);
and U6827 (N_6827,N_6786,N_6616);
nand U6828 (N_6828,N_6643,N_6785);
or U6829 (N_6829,N_6721,N_6724);
nor U6830 (N_6830,N_6640,N_6633);
or U6831 (N_6831,N_6625,N_6632);
and U6832 (N_6832,N_6634,N_6663);
and U6833 (N_6833,N_6763,N_6773);
nand U6834 (N_6834,N_6772,N_6621);
nand U6835 (N_6835,N_6777,N_6726);
and U6836 (N_6836,N_6660,N_6601);
nor U6837 (N_6837,N_6793,N_6699);
and U6838 (N_6838,N_6686,N_6781);
or U6839 (N_6839,N_6650,N_6787);
or U6840 (N_6840,N_6620,N_6771);
or U6841 (N_6841,N_6754,N_6669);
and U6842 (N_6842,N_6762,N_6731);
nand U6843 (N_6843,N_6784,N_6713);
xor U6844 (N_6844,N_6655,N_6659);
nor U6845 (N_6845,N_6749,N_6658);
nor U6846 (N_6846,N_6736,N_6709);
nand U6847 (N_6847,N_6614,N_6701);
xnor U6848 (N_6848,N_6696,N_6755);
and U6849 (N_6849,N_6732,N_6638);
and U6850 (N_6850,N_6750,N_6677);
nand U6851 (N_6851,N_6795,N_6710);
xor U6852 (N_6852,N_6766,N_6645);
xor U6853 (N_6853,N_6765,N_6733);
nand U6854 (N_6854,N_6611,N_6619);
or U6855 (N_6855,N_6774,N_6742);
nand U6856 (N_6856,N_6782,N_6692);
xnor U6857 (N_6857,N_6609,N_6735);
nor U6858 (N_6858,N_6707,N_6652);
nand U6859 (N_6859,N_6646,N_6757);
or U6860 (N_6860,N_6676,N_6798);
and U6861 (N_6861,N_6705,N_6761);
or U6862 (N_6862,N_6725,N_6667);
or U6863 (N_6863,N_6708,N_6797);
and U6864 (N_6864,N_6715,N_6788);
and U6865 (N_6865,N_6789,N_6759);
nor U6866 (N_6866,N_6689,N_6690);
or U6867 (N_6867,N_6647,N_6756);
xor U6868 (N_6868,N_6716,N_6780);
and U6869 (N_6869,N_6747,N_6680);
and U6870 (N_6870,N_6706,N_6791);
and U6871 (N_6871,N_6775,N_6753);
xor U6872 (N_6872,N_6704,N_6656);
nand U6873 (N_6873,N_6697,N_6700);
and U6874 (N_6874,N_6711,N_6684);
and U6875 (N_6875,N_6734,N_6624);
or U6876 (N_6876,N_6612,N_6628);
and U6877 (N_6877,N_6740,N_6666);
nand U6878 (N_6878,N_6653,N_6630);
or U6879 (N_6879,N_6681,N_6649);
or U6880 (N_6880,N_6714,N_6615);
nand U6881 (N_6881,N_6685,N_6727);
and U6882 (N_6882,N_6626,N_6723);
nand U6883 (N_6883,N_6776,N_6687);
or U6884 (N_6884,N_6751,N_6702);
or U6885 (N_6885,N_6610,N_6792);
nor U6886 (N_6886,N_6718,N_6618);
and U6887 (N_6887,N_6661,N_6603);
xor U6888 (N_6888,N_6607,N_6717);
or U6889 (N_6889,N_6637,N_6770);
nand U6890 (N_6890,N_6665,N_6748);
or U6891 (N_6891,N_6739,N_6743);
and U6892 (N_6892,N_6671,N_6600);
and U6893 (N_6893,N_6627,N_6712);
nor U6894 (N_6894,N_6799,N_6688);
or U6895 (N_6895,N_6673,N_6654);
or U6896 (N_6896,N_6778,N_6719);
nand U6897 (N_6897,N_6728,N_6644);
nand U6898 (N_6898,N_6764,N_6738);
or U6899 (N_6899,N_6651,N_6722);
xor U6900 (N_6900,N_6710,N_6717);
xnor U6901 (N_6901,N_6794,N_6786);
or U6902 (N_6902,N_6732,N_6778);
and U6903 (N_6903,N_6637,N_6701);
nand U6904 (N_6904,N_6645,N_6768);
nor U6905 (N_6905,N_6680,N_6686);
or U6906 (N_6906,N_6725,N_6702);
or U6907 (N_6907,N_6686,N_6760);
nor U6908 (N_6908,N_6611,N_6777);
or U6909 (N_6909,N_6729,N_6601);
nor U6910 (N_6910,N_6772,N_6697);
nor U6911 (N_6911,N_6733,N_6770);
nand U6912 (N_6912,N_6762,N_6674);
or U6913 (N_6913,N_6640,N_6770);
nand U6914 (N_6914,N_6703,N_6739);
and U6915 (N_6915,N_6683,N_6688);
xnor U6916 (N_6916,N_6768,N_6652);
xor U6917 (N_6917,N_6788,N_6689);
nand U6918 (N_6918,N_6735,N_6651);
xnor U6919 (N_6919,N_6751,N_6612);
or U6920 (N_6920,N_6630,N_6766);
or U6921 (N_6921,N_6767,N_6614);
nand U6922 (N_6922,N_6754,N_6685);
xor U6923 (N_6923,N_6706,N_6701);
xnor U6924 (N_6924,N_6746,N_6713);
and U6925 (N_6925,N_6713,N_6718);
nor U6926 (N_6926,N_6764,N_6640);
or U6927 (N_6927,N_6621,N_6614);
xor U6928 (N_6928,N_6794,N_6628);
xnor U6929 (N_6929,N_6610,N_6674);
xnor U6930 (N_6930,N_6795,N_6786);
xor U6931 (N_6931,N_6768,N_6779);
and U6932 (N_6932,N_6632,N_6652);
or U6933 (N_6933,N_6761,N_6734);
or U6934 (N_6934,N_6787,N_6741);
xnor U6935 (N_6935,N_6690,N_6755);
or U6936 (N_6936,N_6686,N_6667);
nor U6937 (N_6937,N_6607,N_6702);
nor U6938 (N_6938,N_6664,N_6769);
and U6939 (N_6939,N_6797,N_6763);
nor U6940 (N_6940,N_6695,N_6764);
and U6941 (N_6941,N_6651,N_6738);
nand U6942 (N_6942,N_6643,N_6743);
xor U6943 (N_6943,N_6700,N_6667);
or U6944 (N_6944,N_6606,N_6748);
xor U6945 (N_6945,N_6692,N_6735);
and U6946 (N_6946,N_6637,N_6725);
nand U6947 (N_6947,N_6754,N_6613);
nor U6948 (N_6948,N_6765,N_6652);
and U6949 (N_6949,N_6747,N_6635);
xnor U6950 (N_6950,N_6725,N_6708);
or U6951 (N_6951,N_6672,N_6747);
nor U6952 (N_6952,N_6603,N_6706);
nand U6953 (N_6953,N_6752,N_6788);
nor U6954 (N_6954,N_6601,N_6790);
and U6955 (N_6955,N_6717,N_6656);
or U6956 (N_6956,N_6647,N_6686);
xor U6957 (N_6957,N_6700,N_6685);
nand U6958 (N_6958,N_6623,N_6761);
or U6959 (N_6959,N_6661,N_6618);
or U6960 (N_6960,N_6669,N_6684);
and U6961 (N_6961,N_6730,N_6673);
or U6962 (N_6962,N_6798,N_6799);
xnor U6963 (N_6963,N_6756,N_6733);
or U6964 (N_6964,N_6773,N_6609);
xor U6965 (N_6965,N_6796,N_6651);
nand U6966 (N_6966,N_6782,N_6601);
nor U6967 (N_6967,N_6765,N_6759);
and U6968 (N_6968,N_6646,N_6792);
and U6969 (N_6969,N_6649,N_6615);
nand U6970 (N_6970,N_6778,N_6785);
and U6971 (N_6971,N_6784,N_6743);
or U6972 (N_6972,N_6624,N_6600);
nor U6973 (N_6973,N_6647,N_6645);
or U6974 (N_6974,N_6784,N_6765);
xor U6975 (N_6975,N_6606,N_6688);
nor U6976 (N_6976,N_6765,N_6783);
or U6977 (N_6977,N_6796,N_6739);
xnor U6978 (N_6978,N_6717,N_6612);
xor U6979 (N_6979,N_6729,N_6713);
nand U6980 (N_6980,N_6706,N_6637);
xor U6981 (N_6981,N_6741,N_6625);
xor U6982 (N_6982,N_6656,N_6620);
or U6983 (N_6983,N_6775,N_6787);
and U6984 (N_6984,N_6672,N_6606);
nor U6985 (N_6985,N_6735,N_6642);
or U6986 (N_6986,N_6661,N_6740);
or U6987 (N_6987,N_6699,N_6788);
nand U6988 (N_6988,N_6670,N_6766);
and U6989 (N_6989,N_6752,N_6751);
nor U6990 (N_6990,N_6636,N_6757);
xor U6991 (N_6991,N_6605,N_6663);
nor U6992 (N_6992,N_6799,N_6706);
nor U6993 (N_6993,N_6685,N_6757);
or U6994 (N_6994,N_6769,N_6647);
xnor U6995 (N_6995,N_6675,N_6679);
or U6996 (N_6996,N_6646,N_6750);
and U6997 (N_6997,N_6692,N_6673);
or U6998 (N_6998,N_6715,N_6796);
or U6999 (N_6999,N_6661,N_6602);
and U7000 (N_7000,N_6916,N_6901);
and U7001 (N_7001,N_6909,N_6872);
nor U7002 (N_7002,N_6883,N_6974);
xor U7003 (N_7003,N_6999,N_6933);
nor U7004 (N_7004,N_6813,N_6960);
nand U7005 (N_7005,N_6935,N_6804);
or U7006 (N_7006,N_6862,N_6851);
and U7007 (N_7007,N_6989,N_6975);
nor U7008 (N_7008,N_6983,N_6915);
nand U7009 (N_7009,N_6811,N_6866);
xor U7010 (N_7010,N_6986,N_6905);
or U7011 (N_7011,N_6832,N_6856);
and U7012 (N_7012,N_6839,N_6895);
nand U7013 (N_7013,N_6814,N_6877);
xnor U7014 (N_7014,N_6863,N_6853);
xnor U7015 (N_7015,N_6812,N_6858);
xor U7016 (N_7016,N_6950,N_6988);
or U7017 (N_7017,N_6807,N_6821);
and U7018 (N_7018,N_6990,N_6910);
nor U7019 (N_7019,N_6860,N_6857);
or U7020 (N_7020,N_6947,N_6932);
and U7021 (N_7021,N_6865,N_6875);
nand U7022 (N_7022,N_6835,N_6845);
and U7023 (N_7023,N_6802,N_6847);
xnor U7024 (N_7024,N_6876,N_6881);
or U7025 (N_7025,N_6819,N_6955);
nand U7026 (N_7026,N_6920,N_6861);
or U7027 (N_7027,N_6911,N_6997);
or U7028 (N_7028,N_6852,N_6973);
nand U7029 (N_7029,N_6886,N_6976);
nor U7030 (N_7030,N_6979,N_6918);
and U7031 (N_7031,N_6800,N_6937);
and U7032 (N_7032,N_6904,N_6823);
nor U7033 (N_7033,N_6956,N_6885);
nand U7034 (N_7034,N_6834,N_6964);
and U7035 (N_7035,N_6954,N_6816);
or U7036 (N_7036,N_6923,N_6928);
or U7037 (N_7037,N_6844,N_6870);
xnor U7038 (N_7038,N_6815,N_6913);
or U7039 (N_7039,N_6878,N_6934);
xnor U7040 (N_7040,N_6842,N_6958);
and U7041 (N_7041,N_6831,N_6890);
nor U7042 (N_7042,N_6926,N_6891);
nor U7043 (N_7043,N_6946,N_6828);
and U7044 (N_7044,N_6981,N_6882);
xor U7045 (N_7045,N_6836,N_6971);
nand U7046 (N_7046,N_6874,N_6889);
xor U7047 (N_7047,N_6985,N_6826);
xor U7048 (N_7048,N_6849,N_6887);
nand U7049 (N_7049,N_6867,N_6818);
nand U7050 (N_7050,N_6941,N_6898);
xor U7051 (N_7051,N_6879,N_6957);
nor U7052 (N_7052,N_6966,N_6902);
nand U7053 (N_7053,N_6830,N_6808);
nand U7054 (N_7054,N_6833,N_6817);
nor U7055 (N_7055,N_6963,N_6942);
nand U7056 (N_7056,N_6892,N_6893);
nand U7057 (N_7057,N_6925,N_6930);
xor U7058 (N_7058,N_6924,N_6864);
or U7059 (N_7059,N_6995,N_6912);
nor U7060 (N_7060,N_6919,N_6907);
and U7061 (N_7061,N_6899,N_6801);
nor U7062 (N_7062,N_6953,N_6998);
nand U7063 (N_7063,N_6982,N_6900);
xnor U7064 (N_7064,N_6810,N_6848);
xnor U7065 (N_7065,N_6914,N_6938);
xor U7066 (N_7066,N_6970,N_6896);
nand U7067 (N_7067,N_6951,N_6838);
nor U7068 (N_7068,N_6837,N_6880);
and U7069 (N_7069,N_6903,N_6945);
xnor U7070 (N_7070,N_6850,N_6917);
and U7071 (N_7071,N_6884,N_6843);
nor U7072 (N_7072,N_6962,N_6869);
xor U7073 (N_7073,N_6978,N_6922);
and U7074 (N_7074,N_6977,N_6868);
nor U7075 (N_7075,N_6972,N_6803);
nor U7076 (N_7076,N_6987,N_6906);
nand U7077 (N_7077,N_6936,N_6859);
or U7078 (N_7078,N_6927,N_6829);
nand U7079 (N_7079,N_6940,N_6806);
xnor U7080 (N_7080,N_6980,N_6943);
xor U7081 (N_7081,N_6888,N_6840);
nor U7082 (N_7082,N_6984,N_6894);
nand U7083 (N_7083,N_6827,N_6992);
or U7084 (N_7084,N_6961,N_6965);
nor U7085 (N_7085,N_6939,N_6841);
or U7086 (N_7086,N_6871,N_6929);
and U7087 (N_7087,N_6908,N_6921);
and U7088 (N_7088,N_6873,N_6854);
and U7089 (N_7089,N_6820,N_6809);
nor U7090 (N_7090,N_6967,N_6952);
nand U7091 (N_7091,N_6968,N_6825);
xor U7092 (N_7092,N_6993,N_6824);
or U7093 (N_7093,N_6959,N_6948);
xnor U7094 (N_7094,N_6846,N_6991);
nor U7095 (N_7095,N_6897,N_6931);
and U7096 (N_7096,N_6994,N_6944);
nor U7097 (N_7097,N_6855,N_6996);
nor U7098 (N_7098,N_6822,N_6969);
xor U7099 (N_7099,N_6805,N_6949);
nand U7100 (N_7100,N_6806,N_6932);
xor U7101 (N_7101,N_6853,N_6981);
and U7102 (N_7102,N_6805,N_6864);
xor U7103 (N_7103,N_6877,N_6950);
nor U7104 (N_7104,N_6856,N_6999);
nor U7105 (N_7105,N_6885,N_6960);
nor U7106 (N_7106,N_6845,N_6850);
nor U7107 (N_7107,N_6924,N_6973);
nand U7108 (N_7108,N_6963,N_6882);
and U7109 (N_7109,N_6918,N_6819);
nor U7110 (N_7110,N_6847,N_6850);
and U7111 (N_7111,N_6876,N_6960);
xnor U7112 (N_7112,N_6956,N_6921);
nand U7113 (N_7113,N_6871,N_6879);
nor U7114 (N_7114,N_6831,N_6847);
nor U7115 (N_7115,N_6870,N_6857);
or U7116 (N_7116,N_6984,N_6873);
nor U7117 (N_7117,N_6886,N_6823);
or U7118 (N_7118,N_6839,N_6921);
nor U7119 (N_7119,N_6932,N_6830);
or U7120 (N_7120,N_6931,N_6924);
nor U7121 (N_7121,N_6948,N_6803);
nand U7122 (N_7122,N_6995,N_6891);
or U7123 (N_7123,N_6896,N_6820);
nor U7124 (N_7124,N_6985,N_6900);
nand U7125 (N_7125,N_6903,N_6834);
xor U7126 (N_7126,N_6891,N_6943);
nor U7127 (N_7127,N_6882,N_6909);
and U7128 (N_7128,N_6858,N_6852);
nand U7129 (N_7129,N_6924,N_6813);
and U7130 (N_7130,N_6947,N_6847);
xnor U7131 (N_7131,N_6854,N_6859);
nor U7132 (N_7132,N_6903,N_6865);
nand U7133 (N_7133,N_6807,N_6862);
nor U7134 (N_7134,N_6847,N_6982);
and U7135 (N_7135,N_6942,N_6824);
and U7136 (N_7136,N_6878,N_6921);
nand U7137 (N_7137,N_6969,N_6892);
and U7138 (N_7138,N_6809,N_6825);
and U7139 (N_7139,N_6985,N_6849);
or U7140 (N_7140,N_6913,N_6915);
xor U7141 (N_7141,N_6923,N_6868);
nand U7142 (N_7142,N_6887,N_6916);
and U7143 (N_7143,N_6863,N_6960);
xor U7144 (N_7144,N_6927,N_6973);
nor U7145 (N_7145,N_6959,N_6818);
xnor U7146 (N_7146,N_6883,N_6889);
nor U7147 (N_7147,N_6854,N_6984);
xnor U7148 (N_7148,N_6848,N_6815);
and U7149 (N_7149,N_6997,N_6900);
nand U7150 (N_7150,N_6935,N_6819);
xnor U7151 (N_7151,N_6886,N_6935);
nand U7152 (N_7152,N_6812,N_6938);
xnor U7153 (N_7153,N_6940,N_6818);
xnor U7154 (N_7154,N_6963,N_6828);
and U7155 (N_7155,N_6885,N_6949);
nor U7156 (N_7156,N_6843,N_6941);
nand U7157 (N_7157,N_6938,N_6879);
nand U7158 (N_7158,N_6867,N_6946);
xor U7159 (N_7159,N_6924,N_6868);
and U7160 (N_7160,N_6968,N_6846);
nor U7161 (N_7161,N_6960,N_6842);
or U7162 (N_7162,N_6842,N_6937);
or U7163 (N_7163,N_6803,N_6844);
nand U7164 (N_7164,N_6981,N_6908);
nand U7165 (N_7165,N_6878,N_6822);
nand U7166 (N_7166,N_6815,N_6973);
nor U7167 (N_7167,N_6959,N_6968);
and U7168 (N_7168,N_6971,N_6991);
and U7169 (N_7169,N_6819,N_6922);
nor U7170 (N_7170,N_6821,N_6917);
and U7171 (N_7171,N_6827,N_6846);
and U7172 (N_7172,N_6857,N_6983);
or U7173 (N_7173,N_6806,N_6918);
xor U7174 (N_7174,N_6823,N_6986);
nor U7175 (N_7175,N_6921,N_6806);
nand U7176 (N_7176,N_6955,N_6813);
nand U7177 (N_7177,N_6937,N_6810);
nor U7178 (N_7178,N_6944,N_6980);
or U7179 (N_7179,N_6958,N_6880);
xnor U7180 (N_7180,N_6959,N_6978);
or U7181 (N_7181,N_6970,N_6995);
xnor U7182 (N_7182,N_6902,N_6925);
xnor U7183 (N_7183,N_6853,N_6857);
nand U7184 (N_7184,N_6871,N_6824);
or U7185 (N_7185,N_6954,N_6886);
or U7186 (N_7186,N_6908,N_6955);
xor U7187 (N_7187,N_6961,N_6880);
nor U7188 (N_7188,N_6886,N_6974);
nand U7189 (N_7189,N_6848,N_6872);
and U7190 (N_7190,N_6829,N_6989);
nor U7191 (N_7191,N_6938,N_6827);
xnor U7192 (N_7192,N_6802,N_6843);
xor U7193 (N_7193,N_6835,N_6923);
nor U7194 (N_7194,N_6972,N_6816);
nand U7195 (N_7195,N_6983,N_6938);
and U7196 (N_7196,N_6879,N_6949);
or U7197 (N_7197,N_6906,N_6814);
nor U7198 (N_7198,N_6812,N_6866);
xor U7199 (N_7199,N_6942,N_6925);
nor U7200 (N_7200,N_7113,N_7144);
nand U7201 (N_7201,N_7066,N_7123);
nor U7202 (N_7202,N_7057,N_7079);
xnor U7203 (N_7203,N_7019,N_7087);
nor U7204 (N_7204,N_7086,N_7196);
nand U7205 (N_7205,N_7088,N_7151);
and U7206 (N_7206,N_7036,N_7055);
nor U7207 (N_7207,N_7083,N_7153);
xor U7208 (N_7208,N_7075,N_7002);
nor U7209 (N_7209,N_7160,N_7116);
xnor U7210 (N_7210,N_7010,N_7016);
nor U7211 (N_7211,N_7171,N_7195);
or U7212 (N_7212,N_7070,N_7076);
or U7213 (N_7213,N_7004,N_7053);
nand U7214 (N_7214,N_7112,N_7141);
nor U7215 (N_7215,N_7154,N_7110);
nor U7216 (N_7216,N_7176,N_7121);
or U7217 (N_7217,N_7047,N_7185);
nand U7218 (N_7218,N_7078,N_7025);
nor U7219 (N_7219,N_7006,N_7148);
or U7220 (N_7220,N_7106,N_7027);
nand U7221 (N_7221,N_7089,N_7009);
and U7222 (N_7222,N_7026,N_7126);
nand U7223 (N_7223,N_7068,N_7011);
nor U7224 (N_7224,N_7105,N_7133);
xor U7225 (N_7225,N_7090,N_7150);
nand U7226 (N_7226,N_7164,N_7092);
nand U7227 (N_7227,N_7035,N_7031);
xnor U7228 (N_7228,N_7188,N_7040);
nor U7229 (N_7229,N_7174,N_7041);
and U7230 (N_7230,N_7137,N_7140);
or U7231 (N_7231,N_7043,N_7061);
nand U7232 (N_7232,N_7170,N_7048);
xor U7233 (N_7233,N_7108,N_7054);
nor U7234 (N_7234,N_7177,N_7189);
and U7235 (N_7235,N_7056,N_7022);
nor U7236 (N_7236,N_7038,N_7082);
nand U7237 (N_7237,N_7186,N_7073);
and U7238 (N_7238,N_7149,N_7097);
nand U7239 (N_7239,N_7034,N_7190);
nand U7240 (N_7240,N_7030,N_7168);
nand U7241 (N_7241,N_7096,N_7180);
or U7242 (N_7242,N_7098,N_7199);
xor U7243 (N_7243,N_7187,N_7143);
or U7244 (N_7244,N_7039,N_7102);
nor U7245 (N_7245,N_7119,N_7109);
or U7246 (N_7246,N_7095,N_7050);
or U7247 (N_7247,N_7049,N_7181);
xor U7248 (N_7248,N_7007,N_7044);
nor U7249 (N_7249,N_7194,N_7064);
and U7250 (N_7250,N_7145,N_7099);
nand U7251 (N_7251,N_7156,N_7067);
xnor U7252 (N_7252,N_7069,N_7000);
nand U7253 (N_7253,N_7028,N_7003);
or U7254 (N_7254,N_7134,N_7081);
and U7255 (N_7255,N_7147,N_7001);
xnor U7256 (N_7256,N_7167,N_7124);
nand U7257 (N_7257,N_7072,N_7018);
or U7258 (N_7258,N_7198,N_7114);
nand U7259 (N_7259,N_7062,N_7193);
nor U7260 (N_7260,N_7012,N_7046);
and U7261 (N_7261,N_7103,N_7132);
nand U7262 (N_7262,N_7118,N_7084);
or U7263 (N_7263,N_7152,N_7192);
and U7264 (N_7264,N_7080,N_7015);
or U7265 (N_7265,N_7191,N_7104);
and U7266 (N_7266,N_7128,N_7122);
and U7267 (N_7267,N_7091,N_7197);
nand U7268 (N_7268,N_7052,N_7100);
and U7269 (N_7269,N_7142,N_7173);
nor U7270 (N_7270,N_7131,N_7013);
xor U7271 (N_7271,N_7032,N_7125);
and U7272 (N_7272,N_7017,N_7085);
and U7273 (N_7273,N_7014,N_7165);
nor U7274 (N_7274,N_7120,N_7161);
xor U7275 (N_7275,N_7020,N_7063);
xor U7276 (N_7276,N_7139,N_7101);
or U7277 (N_7277,N_7138,N_7042);
xnor U7278 (N_7278,N_7058,N_7024);
or U7279 (N_7279,N_7158,N_7071);
nand U7280 (N_7280,N_7021,N_7051);
xor U7281 (N_7281,N_7175,N_7077);
xor U7282 (N_7282,N_7115,N_7146);
and U7283 (N_7283,N_7136,N_7179);
or U7284 (N_7284,N_7172,N_7178);
or U7285 (N_7285,N_7163,N_7059);
and U7286 (N_7286,N_7093,N_7111);
and U7287 (N_7287,N_7065,N_7135);
nand U7288 (N_7288,N_7094,N_7169);
and U7289 (N_7289,N_7033,N_7130);
and U7290 (N_7290,N_7074,N_7183);
and U7291 (N_7291,N_7005,N_7159);
nand U7292 (N_7292,N_7129,N_7107);
nor U7293 (N_7293,N_7157,N_7184);
nor U7294 (N_7294,N_7029,N_7060);
and U7295 (N_7295,N_7117,N_7008);
and U7296 (N_7296,N_7162,N_7182);
nor U7297 (N_7297,N_7037,N_7127);
nor U7298 (N_7298,N_7045,N_7023);
nand U7299 (N_7299,N_7155,N_7166);
or U7300 (N_7300,N_7058,N_7133);
xnor U7301 (N_7301,N_7130,N_7058);
nand U7302 (N_7302,N_7068,N_7115);
or U7303 (N_7303,N_7178,N_7129);
and U7304 (N_7304,N_7163,N_7047);
nand U7305 (N_7305,N_7070,N_7155);
nor U7306 (N_7306,N_7184,N_7094);
or U7307 (N_7307,N_7044,N_7033);
nand U7308 (N_7308,N_7098,N_7017);
xnor U7309 (N_7309,N_7098,N_7087);
nor U7310 (N_7310,N_7145,N_7136);
or U7311 (N_7311,N_7138,N_7161);
nor U7312 (N_7312,N_7027,N_7085);
or U7313 (N_7313,N_7099,N_7184);
and U7314 (N_7314,N_7180,N_7159);
nor U7315 (N_7315,N_7037,N_7082);
nand U7316 (N_7316,N_7116,N_7054);
xor U7317 (N_7317,N_7140,N_7089);
xor U7318 (N_7318,N_7101,N_7146);
and U7319 (N_7319,N_7180,N_7093);
xor U7320 (N_7320,N_7088,N_7118);
nor U7321 (N_7321,N_7063,N_7117);
nor U7322 (N_7322,N_7091,N_7110);
nand U7323 (N_7323,N_7034,N_7009);
or U7324 (N_7324,N_7053,N_7037);
or U7325 (N_7325,N_7135,N_7130);
xor U7326 (N_7326,N_7169,N_7123);
nor U7327 (N_7327,N_7151,N_7034);
nand U7328 (N_7328,N_7185,N_7089);
or U7329 (N_7329,N_7174,N_7104);
and U7330 (N_7330,N_7075,N_7092);
xnor U7331 (N_7331,N_7109,N_7020);
nand U7332 (N_7332,N_7147,N_7095);
nor U7333 (N_7333,N_7105,N_7169);
and U7334 (N_7334,N_7056,N_7114);
xnor U7335 (N_7335,N_7066,N_7190);
and U7336 (N_7336,N_7096,N_7017);
xor U7337 (N_7337,N_7007,N_7074);
xnor U7338 (N_7338,N_7080,N_7010);
and U7339 (N_7339,N_7085,N_7177);
nand U7340 (N_7340,N_7158,N_7033);
nor U7341 (N_7341,N_7001,N_7196);
xor U7342 (N_7342,N_7176,N_7059);
or U7343 (N_7343,N_7105,N_7026);
nor U7344 (N_7344,N_7044,N_7194);
and U7345 (N_7345,N_7188,N_7035);
and U7346 (N_7346,N_7034,N_7006);
nor U7347 (N_7347,N_7033,N_7159);
or U7348 (N_7348,N_7018,N_7109);
nand U7349 (N_7349,N_7071,N_7103);
and U7350 (N_7350,N_7131,N_7161);
xnor U7351 (N_7351,N_7083,N_7197);
or U7352 (N_7352,N_7044,N_7001);
xnor U7353 (N_7353,N_7113,N_7137);
or U7354 (N_7354,N_7136,N_7113);
and U7355 (N_7355,N_7085,N_7002);
xnor U7356 (N_7356,N_7102,N_7025);
nand U7357 (N_7357,N_7159,N_7041);
nand U7358 (N_7358,N_7122,N_7077);
nor U7359 (N_7359,N_7199,N_7177);
or U7360 (N_7360,N_7014,N_7116);
xnor U7361 (N_7361,N_7072,N_7188);
nor U7362 (N_7362,N_7086,N_7081);
and U7363 (N_7363,N_7106,N_7119);
and U7364 (N_7364,N_7119,N_7125);
or U7365 (N_7365,N_7084,N_7112);
or U7366 (N_7366,N_7019,N_7117);
or U7367 (N_7367,N_7198,N_7059);
xor U7368 (N_7368,N_7021,N_7158);
nand U7369 (N_7369,N_7040,N_7081);
and U7370 (N_7370,N_7126,N_7069);
or U7371 (N_7371,N_7128,N_7162);
and U7372 (N_7372,N_7091,N_7086);
and U7373 (N_7373,N_7085,N_7061);
and U7374 (N_7374,N_7036,N_7054);
nor U7375 (N_7375,N_7017,N_7117);
and U7376 (N_7376,N_7181,N_7179);
or U7377 (N_7377,N_7038,N_7078);
xor U7378 (N_7378,N_7153,N_7042);
and U7379 (N_7379,N_7040,N_7065);
xor U7380 (N_7380,N_7146,N_7033);
xor U7381 (N_7381,N_7116,N_7085);
nor U7382 (N_7382,N_7067,N_7024);
xor U7383 (N_7383,N_7173,N_7073);
and U7384 (N_7384,N_7092,N_7107);
xnor U7385 (N_7385,N_7026,N_7084);
or U7386 (N_7386,N_7120,N_7192);
xor U7387 (N_7387,N_7198,N_7166);
or U7388 (N_7388,N_7102,N_7120);
xnor U7389 (N_7389,N_7095,N_7167);
or U7390 (N_7390,N_7005,N_7106);
and U7391 (N_7391,N_7179,N_7082);
or U7392 (N_7392,N_7044,N_7131);
or U7393 (N_7393,N_7159,N_7134);
or U7394 (N_7394,N_7034,N_7018);
xor U7395 (N_7395,N_7043,N_7052);
nand U7396 (N_7396,N_7188,N_7076);
and U7397 (N_7397,N_7108,N_7087);
nor U7398 (N_7398,N_7191,N_7081);
nor U7399 (N_7399,N_7120,N_7113);
or U7400 (N_7400,N_7312,N_7325);
and U7401 (N_7401,N_7288,N_7267);
or U7402 (N_7402,N_7358,N_7215);
nor U7403 (N_7403,N_7253,N_7249);
xnor U7404 (N_7404,N_7350,N_7289);
nand U7405 (N_7405,N_7373,N_7268);
nand U7406 (N_7406,N_7303,N_7355);
xor U7407 (N_7407,N_7379,N_7371);
or U7408 (N_7408,N_7338,N_7359);
nand U7409 (N_7409,N_7220,N_7310);
nand U7410 (N_7410,N_7211,N_7240);
or U7411 (N_7411,N_7243,N_7244);
nand U7412 (N_7412,N_7327,N_7386);
xor U7413 (N_7413,N_7368,N_7213);
nand U7414 (N_7414,N_7382,N_7278);
nor U7415 (N_7415,N_7313,N_7326);
and U7416 (N_7416,N_7230,N_7236);
xor U7417 (N_7417,N_7218,N_7214);
and U7418 (N_7418,N_7205,N_7206);
or U7419 (N_7419,N_7239,N_7300);
and U7420 (N_7420,N_7224,N_7258);
nor U7421 (N_7421,N_7250,N_7307);
nand U7422 (N_7422,N_7262,N_7271);
and U7423 (N_7423,N_7329,N_7290);
or U7424 (N_7424,N_7385,N_7391);
or U7425 (N_7425,N_7248,N_7361);
xnor U7426 (N_7426,N_7301,N_7212);
xnor U7427 (N_7427,N_7324,N_7294);
or U7428 (N_7428,N_7337,N_7265);
and U7429 (N_7429,N_7252,N_7319);
nand U7430 (N_7430,N_7384,N_7261);
nor U7431 (N_7431,N_7357,N_7340);
xnor U7432 (N_7432,N_7226,N_7237);
nand U7433 (N_7433,N_7365,N_7304);
nor U7434 (N_7434,N_7296,N_7395);
nor U7435 (N_7435,N_7347,N_7269);
or U7436 (N_7436,N_7394,N_7397);
xnor U7437 (N_7437,N_7229,N_7351);
xnor U7438 (N_7438,N_7275,N_7398);
and U7439 (N_7439,N_7280,N_7388);
nand U7440 (N_7440,N_7341,N_7393);
and U7441 (N_7441,N_7318,N_7260);
and U7442 (N_7442,N_7376,N_7202);
or U7443 (N_7443,N_7223,N_7374);
or U7444 (N_7444,N_7335,N_7323);
and U7445 (N_7445,N_7298,N_7241);
nand U7446 (N_7446,N_7367,N_7346);
or U7447 (N_7447,N_7336,N_7334);
nand U7448 (N_7448,N_7315,N_7345);
and U7449 (N_7449,N_7293,N_7272);
or U7450 (N_7450,N_7210,N_7291);
nand U7451 (N_7451,N_7227,N_7277);
and U7452 (N_7452,N_7228,N_7221);
nor U7453 (N_7453,N_7364,N_7207);
nor U7454 (N_7454,N_7235,N_7270);
xor U7455 (N_7455,N_7344,N_7375);
nand U7456 (N_7456,N_7320,N_7363);
xnor U7457 (N_7457,N_7348,N_7273);
xor U7458 (N_7458,N_7309,N_7245);
nor U7459 (N_7459,N_7282,N_7263);
or U7460 (N_7460,N_7330,N_7321);
nand U7461 (N_7461,N_7225,N_7266);
or U7462 (N_7462,N_7259,N_7208);
or U7463 (N_7463,N_7200,N_7231);
and U7464 (N_7464,N_7264,N_7378);
and U7465 (N_7465,N_7286,N_7292);
and U7466 (N_7466,N_7285,N_7284);
and U7467 (N_7467,N_7295,N_7281);
and U7468 (N_7468,N_7396,N_7287);
nand U7469 (N_7469,N_7369,N_7390);
nor U7470 (N_7470,N_7246,N_7308);
or U7471 (N_7471,N_7311,N_7362);
or U7472 (N_7472,N_7366,N_7322);
or U7473 (N_7473,N_7203,N_7209);
nand U7474 (N_7474,N_7370,N_7217);
and U7475 (N_7475,N_7314,N_7305);
and U7476 (N_7476,N_7380,N_7238);
xnor U7477 (N_7477,N_7387,N_7354);
nand U7478 (N_7478,N_7381,N_7222);
nor U7479 (N_7479,N_7232,N_7276);
and U7480 (N_7480,N_7201,N_7356);
xnor U7481 (N_7481,N_7219,N_7343);
nand U7482 (N_7482,N_7274,N_7306);
nand U7483 (N_7483,N_7251,N_7216);
xor U7484 (N_7484,N_7377,N_7360);
xor U7485 (N_7485,N_7302,N_7256);
or U7486 (N_7486,N_7297,N_7372);
or U7487 (N_7487,N_7316,N_7255);
or U7488 (N_7488,N_7339,N_7389);
nor U7489 (N_7489,N_7392,N_7254);
nand U7490 (N_7490,N_7352,N_7333);
and U7491 (N_7491,N_7328,N_7247);
or U7492 (N_7492,N_7332,N_7257);
xnor U7493 (N_7493,N_7383,N_7204);
nor U7494 (N_7494,N_7353,N_7242);
or U7495 (N_7495,N_7279,N_7283);
nor U7496 (N_7496,N_7342,N_7317);
nor U7497 (N_7497,N_7299,N_7234);
nor U7498 (N_7498,N_7349,N_7331);
nand U7499 (N_7499,N_7399,N_7233);
xor U7500 (N_7500,N_7355,N_7315);
nor U7501 (N_7501,N_7275,N_7211);
nor U7502 (N_7502,N_7303,N_7360);
nor U7503 (N_7503,N_7222,N_7348);
xor U7504 (N_7504,N_7392,N_7357);
and U7505 (N_7505,N_7218,N_7252);
xor U7506 (N_7506,N_7248,N_7231);
and U7507 (N_7507,N_7230,N_7381);
nand U7508 (N_7508,N_7305,N_7361);
or U7509 (N_7509,N_7349,N_7355);
or U7510 (N_7510,N_7202,N_7233);
nand U7511 (N_7511,N_7284,N_7321);
nand U7512 (N_7512,N_7388,N_7374);
nor U7513 (N_7513,N_7398,N_7259);
nand U7514 (N_7514,N_7330,N_7277);
and U7515 (N_7515,N_7229,N_7250);
or U7516 (N_7516,N_7345,N_7357);
or U7517 (N_7517,N_7282,N_7215);
and U7518 (N_7518,N_7283,N_7281);
and U7519 (N_7519,N_7376,N_7360);
nor U7520 (N_7520,N_7214,N_7337);
nor U7521 (N_7521,N_7210,N_7382);
or U7522 (N_7522,N_7203,N_7384);
or U7523 (N_7523,N_7287,N_7384);
nand U7524 (N_7524,N_7326,N_7239);
xor U7525 (N_7525,N_7257,N_7328);
xor U7526 (N_7526,N_7298,N_7231);
nand U7527 (N_7527,N_7224,N_7337);
or U7528 (N_7528,N_7371,N_7334);
or U7529 (N_7529,N_7391,N_7375);
nor U7530 (N_7530,N_7254,N_7227);
and U7531 (N_7531,N_7311,N_7383);
nor U7532 (N_7532,N_7375,N_7323);
or U7533 (N_7533,N_7254,N_7395);
nand U7534 (N_7534,N_7260,N_7379);
nand U7535 (N_7535,N_7358,N_7300);
nand U7536 (N_7536,N_7316,N_7243);
nor U7537 (N_7537,N_7246,N_7293);
and U7538 (N_7538,N_7274,N_7397);
nand U7539 (N_7539,N_7343,N_7204);
or U7540 (N_7540,N_7293,N_7318);
nor U7541 (N_7541,N_7212,N_7302);
nor U7542 (N_7542,N_7363,N_7239);
xnor U7543 (N_7543,N_7207,N_7375);
or U7544 (N_7544,N_7208,N_7234);
and U7545 (N_7545,N_7292,N_7325);
nor U7546 (N_7546,N_7332,N_7380);
xor U7547 (N_7547,N_7337,N_7234);
or U7548 (N_7548,N_7296,N_7349);
and U7549 (N_7549,N_7247,N_7258);
nor U7550 (N_7550,N_7232,N_7328);
nor U7551 (N_7551,N_7351,N_7384);
xor U7552 (N_7552,N_7365,N_7211);
nand U7553 (N_7553,N_7333,N_7311);
xnor U7554 (N_7554,N_7254,N_7316);
nand U7555 (N_7555,N_7255,N_7232);
nand U7556 (N_7556,N_7330,N_7204);
or U7557 (N_7557,N_7322,N_7203);
and U7558 (N_7558,N_7234,N_7388);
and U7559 (N_7559,N_7377,N_7214);
or U7560 (N_7560,N_7327,N_7218);
xor U7561 (N_7561,N_7258,N_7338);
and U7562 (N_7562,N_7219,N_7392);
nor U7563 (N_7563,N_7297,N_7205);
nor U7564 (N_7564,N_7239,N_7351);
nor U7565 (N_7565,N_7298,N_7257);
or U7566 (N_7566,N_7326,N_7207);
and U7567 (N_7567,N_7301,N_7388);
or U7568 (N_7568,N_7396,N_7288);
nor U7569 (N_7569,N_7286,N_7265);
nor U7570 (N_7570,N_7227,N_7366);
or U7571 (N_7571,N_7337,N_7346);
or U7572 (N_7572,N_7244,N_7364);
or U7573 (N_7573,N_7350,N_7216);
xnor U7574 (N_7574,N_7226,N_7356);
nor U7575 (N_7575,N_7330,N_7237);
and U7576 (N_7576,N_7359,N_7337);
nand U7577 (N_7577,N_7372,N_7235);
nand U7578 (N_7578,N_7254,N_7269);
or U7579 (N_7579,N_7212,N_7268);
and U7580 (N_7580,N_7353,N_7320);
or U7581 (N_7581,N_7372,N_7234);
or U7582 (N_7582,N_7286,N_7362);
or U7583 (N_7583,N_7205,N_7317);
xor U7584 (N_7584,N_7233,N_7355);
xor U7585 (N_7585,N_7205,N_7340);
nand U7586 (N_7586,N_7358,N_7272);
or U7587 (N_7587,N_7382,N_7315);
and U7588 (N_7588,N_7245,N_7381);
or U7589 (N_7589,N_7295,N_7296);
and U7590 (N_7590,N_7233,N_7383);
nor U7591 (N_7591,N_7391,N_7297);
or U7592 (N_7592,N_7277,N_7338);
nor U7593 (N_7593,N_7232,N_7370);
nand U7594 (N_7594,N_7393,N_7276);
or U7595 (N_7595,N_7286,N_7282);
or U7596 (N_7596,N_7218,N_7392);
and U7597 (N_7597,N_7244,N_7217);
nand U7598 (N_7598,N_7240,N_7216);
nand U7599 (N_7599,N_7321,N_7242);
and U7600 (N_7600,N_7565,N_7543);
or U7601 (N_7601,N_7503,N_7568);
nand U7602 (N_7602,N_7445,N_7471);
nor U7603 (N_7603,N_7490,N_7414);
or U7604 (N_7604,N_7438,N_7401);
nor U7605 (N_7605,N_7572,N_7519);
xor U7606 (N_7606,N_7421,N_7402);
nor U7607 (N_7607,N_7561,N_7514);
and U7608 (N_7608,N_7433,N_7475);
nand U7609 (N_7609,N_7518,N_7560);
or U7610 (N_7610,N_7586,N_7407);
or U7611 (N_7611,N_7509,N_7582);
nand U7612 (N_7612,N_7530,N_7547);
or U7613 (N_7613,N_7521,N_7567);
or U7614 (N_7614,N_7527,N_7511);
or U7615 (N_7615,N_7469,N_7546);
or U7616 (N_7616,N_7544,N_7574);
nand U7617 (N_7617,N_7489,N_7566);
and U7618 (N_7618,N_7406,N_7472);
or U7619 (N_7619,N_7466,N_7411);
nor U7620 (N_7620,N_7464,N_7431);
nand U7621 (N_7621,N_7555,N_7426);
and U7622 (N_7622,N_7444,N_7470);
nand U7623 (N_7623,N_7473,N_7592);
xor U7624 (N_7624,N_7501,N_7559);
nand U7625 (N_7625,N_7597,N_7595);
and U7626 (N_7626,N_7493,N_7537);
nor U7627 (N_7627,N_7474,N_7434);
nor U7628 (N_7628,N_7562,N_7556);
or U7629 (N_7629,N_7428,N_7494);
and U7630 (N_7630,N_7545,N_7548);
xnor U7631 (N_7631,N_7517,N_7409);
nand U7632 (N_7632,N_7456,N_7539);
nand U7633 (N_7633,N_7558,N_7476);
xnor U7634 (N_7634,N_7570,N_7596);
and U7635 (N_7635,N_7432,N_7583);
nand U7636 (N_7636,N_7510,N_7495);
or U7637 (N_7637,N_7533,N_7478);
xor U7638 (N_7638,N_7576,N_7578);
nor U7639 (N_7639,N_7553,N_7451);
nor U7640 (N_7640,N_7523,N_7429);
nand U7641 (N_7641,N_7599,N_7507);
nor U7642 (N_7642,N_7492,N_7458);
or U7643 (N_7643,N_7526,N_7424);
nor U7644 (N_7644,N_7551,N_7508);
nand U7645 (N_7645,N_7557,N_7400);
nand U7646 (N_7646,N_7487,N_7404);
nor U7647 (N_7647,N_7482,N_7455);
nand U7648 (N_7648,N_7590,N_7485);
nand U7649 (N_7649,N_7587,N_7410);
nand U7650 (N_7650,N_7446,N_7422);
or U7651 (N_7651,N_7536,N_7497);
xor U7652 (N_7652,N_7593,N_7412);
xnor U7653 (N_7653,N_7486,N_7573);
and U7654 (N_7654,N_7598,N_7580);
nor U7655 (N_7655,N_7591,N_7427);
nor U7656 (N_7656,N_7425,N_7405);
and U7657 (N_7657,N_7534,N_7529);
or U7658 (N_7658,N_7538,N_7443);
or U7659 (N_7659,N_7447,N_7450);
or U7660 (N_7660,N_7468,N_7516);
and U7661 (N_7661,N_7499,N_7408);
xnor U7662 (N_7662,N_7564,N_7463);
nand U7663 (N_7663,N_7436,N_7528);
nor U7664 (N_7664,N_7435,N_7535);
or U7665 (N_7665,N_7418,N_7480);
nand U7666 (N_7666,N_7577,N_7419);
nor U7667 (N_7667,N_7457,N_7415);
and U7668 (N_7668,N_7512,N_7417);
nand U7669 (N_7669,N_7403,N_7479);
nor U7670 (N_7670,N_7484,N_7515);
and U7671 (N_7671,N_7588,N_7505);
xnor U7672 (N_7672,N_7461,N_7552);
or U7673 (N_7673,N_7542,N_7522);
nand U7674 (N_7674,N_7440,N_7467);
or U7675 (N_7675,N_7524,N_7430);
and U7676 (N_7676,N_7532,N_7437);
xnor U7677 (N_7677,N_7420,N_7498);
nand U7678 (N_7678,N_7477,N_7453);
xnor U7679 (N_7679,N_7525,N_7442);
nand U7680 (N_7680,N_7481,N_7449);
and U7681 (N_7681,N_7502,N_7488);
and U7682 (N_7682,N_7520,N_7589);
xor U7683 (N_7683,N_7571,N_7454);
nand U7684 (N_7684,N_7439,N_7500);
xor U7685 (N_7685,N_7554,N_7504);
and U7686 (N_7686,N_7594,N_7579);
or U7687 (N_7687,N_7483,N_7462);
xor U7688 (N_7688,N_7441,N_7491);
nor U7689 (N_7689,N_7452,N_7585);
xor U7690 (N_7690,N_7448,N_7513);
and U7691 (N_7691,N_7575,N_7569);
and U7692 (N_7692,N_7540,N_7584);
and U7693 (N_7693,N_7416,N_7496);
nand U7694 (N_7694,N_7459,N_7563);
nor U7695 (N_7695,N_7581,N_7549);
nand U7696 (N_7696,N_7531,N_7506);
or U7697 (N_7697,N_7460,N_7413);
nor U7698 (N_7698,N_7550,N_7423);
nor U7699 (N_7699,N_7541,N_7465);
and U7700 (N_7700,N_7567,N_7565);
nor U7701 (N_7701,N_7412,N_7455);
nor U7702 (N_7702,N_7577,N_7598);
nand U7703 (N_7703,N_7509,N_7480);
xor U7704 (N_7704,N_7412,N_7405);
xor U7705 (N_7705,N_7578,N_7448);
xnor U7706 (N_7706,N_7569,N_7539);
and U7707 (N_7707,N_7471,N_7483);
or U7708 (N_7708,N_7579,N_7421);
nand U7709 (N_7709,N_7424,N_7563);
or U7710 (N_7710,N_7424,N_7559);
nor U7711 (N_7711,N_7407,N_7543);
or U7712 (N_7712,N_7531,N_7466);
nand U7713 (N_7713,N_7593,N_7462);
xor U7714 (N_7714,N_7434,N_7471);
xnor U7715 (N_7715,N_7440,N_7557);
nor U7716 (N_7716,N_7511,N_7468);
nor U7717 (N_7717,N_7407,N_7587);
and U7718 (N_7718,N_7417,N_7490);
nor U7719 (N_7719,N_7431,N_7580);
nor U7720 (N_7720,N_7493,N_7406);
xor U7721 (N_7721,N_7438,N_7553);
nor U7722 (N_7722,N_7403,N_7416);
xor U7723 (N_7723,N_7448,N_7496);
or U7724 (N_7724,N_7545,N_7416);
nand U7725 (N_7725,N_7537,N_7566);
nand U7726 (N_7726,N_7440,N_7478);
xnor U7727 (N_7727,N_7468,N_7447);
xnor U7728 (N_7728,N_7598,N_7424);
xnor U7729 (N_7729,N_7548,N_7542);
and U7730 (N_7730,N_7490,N_7585);
nor U7731 (N_7731,N_7455,N_7543);
nor U7732 (N_7732,N_7501,N_7591);
nand U7733 (N_7733,N_7510,N_7599);
xnor U7734 (N_7734,N_7468,N_7400);
or U7735 (N_7735,N_7542,N_7563);
nor U7736 (N_7736,N_7479,N_7579);
xor U7737 (N_7737,N_7452,N_7460);
xnor U7738 (N_7738,N_7442,N_7584);
and U7739 (N_7739,N_7462,N_7422);
or U7740 (N_7740,N_7588,N_7442);
xnor U7741 (N_7741,N_7485,N_7497);
nor U7742 (N_7742,N_7550,N_7554);
or U7743 (N_7743,N_7528,N_7424);
xnor U7744 (N_7744,N_7429,N_7536);
nand U7745 (N_7745,N_7402,N_7532);
and U7746 (N_7746,N_7589,N_7585);
xnor U7747 (N_7747,N_7570,N_7537);
nand U7748 (N_7748,N_7523,N_7572);
or U7749 (N_7749,N_7551,N_7412);
or U7750 (N_7750,N_7400,N_7566);
xnor U7751 (N_7751,N_7511,N_7584);
or U7752 (N_7752,N_7567,N_7490);
nand U7753 (N_7753,N_7463,N_7518);
nor U7754 (N_7754,N_7575,N_7418);
nor U7755 (N_7755,N_7565,N_7505);
xor U7756 (N_7756,N_7541,N_7559);
nor U7757 (N_7757,N_7561,N_7473);
nand U7758 (N_7758,N_7444,N_7598);
nand U7759 (N_7759,N_7497,N_7592);
xnor U7760 (N_7760,N_7465,N_7429);
or U7761 (N_7761,N_7510,N_7555);
or U7762 (N_7762,N_7557,N_7423);
and U7763 (N_7763,N_7409,N_7585);
xnor U7764 (N_7764,N_7572,N_7476);
xnor U7765 (N_7765,N_7596,N_7473);
and U7766 (N_7766,N_7442,N_7530);
xnor U7767 (N_7767,N_7436,N_7566);
nor U7768 (N_7768,N_7532,N_7525);
xnor U7769 (N_7769,N_7578,N_7493);
nor U7770 (N_7770,N_7500,N_7554);
and U7771 (N_7771,N_7588,N_7591);
nand U7772 (N_7772,N_7472,N_7485);
xnor U7773 (N_7773,N_7508,N_7586);
xor U7774 (N_7774,N_7430,N_7465);
and U7775 (N_7775,N_7503,N_7453);
nand U7776 (N_7776,N_7415,N_7587);
xor U7777 (N_7777,N_7469,N_7447);
nand U7778 (N_7778,N_7549,N_7588);
or U7779 (N_7779,N_7576,N_7426);
and U7780 (N_7780,N_7523,N_7500);
and U7781 (N_7781,N_7543,N_7484);
and U7782 (N_7782,N_7576,N_7470);
or U7783 (N_7783,N_7405,N_7522);
nor U7784 (N_7784,N_7506,N_7461);
xnor U7785 (N_7785,N_7442,N_7593);
xnor U7786 (N_7786,N_7539,N_7574);
nor U7787 (N_7787,N_7472,N_7568);
or U7788 (N_7788,N_7522,N_7424);
nor U7789 (N_7789,N_7444,N_7440);
and U7790 (N_7790,N_7534,N_7550);
and U7791 (N_7791,N_7438,N_7555);
and U7792 (N_7792,N_7596,N_7572);
and U7793 (N_7793,N_7410,N_7427);
nand U7794 (N_7794,N_7408,N_7486);
xor U7795 (N_7795,N_7457,N_7456);
xor U7796 (N_7796,N_7537,N_7432);
and U7797 (N_7797,N_7481,N_7422);
nand U7798 (N_7798,N_7514,N_7519);
nand U7799 (N_7799,N_7545,N_7550);
nor U7800 (N_7800,N_7714,N_7651);
or U7801 (N_7801,N_7681,N_7792);
and U7802 (N_7802,N_7771,N_7673);
xor U7803 (N_7803,N_7656,N_7689);
nand U7804 (N_7804,N_7757,N_7767);
and U7805 (N_7805,N_7600,N_7669);
xnor U7806 (N_7806,N_7632,N_7791);
and U7807 (N_7807,N_7675,N_7758);
or U7808 (N_7808,N_7618,N_7684);
xor U7809 (N_7809,N_7652,N_7690);
and U7810 (N_7810,N_7727,N_7664);
or U7811 (N_7811,N_7647,N_7609);
and U7812 (N_7812,N_7703,N_7614);
nor U7813 (N_7813,N_7639,N_7697);
nand U7814 (N_7814,N_7627,N_7672);
nor U7815 (N_7815,N_7794,N_7665);
nor U7816 (N_7816,N_7744,N_7724);
and U7817 (N_7817,N_7606,N_7650);
or U7818 (N_7818,N_7713,N_7751);
and U7819 (N_7819,N_7787,N_7776);
nor U7820 (N_7820,N_7737,N_7763);
or U7821 (N_7821,N_7701,N_7643);
nor U7822 (N_7822,N_7641,N_7754);
or U7823 (N_7823,N_7633,N_7790);
xnor U7824 (N_7824,N_7685,N_7608);
or U7825 (N_7825,N_7691,N_7765);
nor U7826 (N_7826,N_7774,N_7613);
nor U7827 (N_7827,N_7789,N_7726);
and U7828 (N_7828,N_7710,N_7780);
xor U7829 (N_7829,N_7721,N_7680);
xor U7830 (N_7830,N_7785,N_7707);
or U7831 (N_7831,N_7629,N_7702);
nand U7832 (N_7832,N_7745,N_7706);
and U7833 (N_7833,N_7730,N_7646);
and U7834 (N_7834,N_7693,N_7786);
and U7835 (N_7835,N_7612,N_7781);
nor U7836 (N_7836,N_7782,N_7621);
nand U7837 (N_7837,N_7750,N_7637);
xor U7838 (N_7838,N_7741,N_7759);
nor U7839 (N_7839,N_7679,N_7766);
xor U7840 (N_7840,N_7625,N_7762);
or U7841 (N_7841,N_7734,N_7749);
and U7842 (N_7842,N_7626,N_7764);
xnor U7843 (N_7843,N_7715,N_7699);
xnor U7844 (N_7844,N_7668,N_7700);
nand U7845 (N_7845,N_7663,N_7716);
nor U7846 (N_7846,N_7686,N_7772);
nor U7847 (N_7847,N_7622,N_7746);
nand U7848 (N_7848,N_7666,N_7718);
nand U7849 (N_7849,N_7687,N_7773);
nand U7850 (N_7850,N_7640,N_7692);
xnor U7851 (N_7851,N_7796,N_7628);
and U7852 (N_7852,N_7683,N_7729);
or U7853 (N_7853,N_7719,N_7738);
nor U7854 (N_7854,N_7682,N_7660);
or U7855 (N_7855,N_7797,N_7658);
nand U7856 (N_7856,N_7717,N_7617);
and U7857 (N_7857,N_7634,N_7615);
nor U7858 (N_7858,N_7695,N_7778);
nand U7859 (N_7859,N_7694,N_7638);
and U7860 (N_7860,N_7708,N_7648);
nor U7861 (N_7861,N_7616,N_7756);
xor U7862 (N_7862,N_7644,N_7631);
nand U7863 (N_7863,N_7661,N_7655);
nand U7864 (N_7864,N_7667,N_7720);
xor U7865 (N_7865,N_7688,N_7732);
and U7866 (N_7866,N_7671,N_7676);
nor U7867 (N_7867,N_7799,N_7740);
xnor U7868 (N_7868,N_7783,N_7705);
xor U7869 (N_7869,N_7624,N_7739);
and U7870 (N_7870,N_7748,N_7788);
nand U7871 (N_7871,N_7736,N_7678);
nor U7872 (N_7872,N_7798,N_7743);
or U7873 (N_7873,N_7620,N_7610);
nor U7874 (N_7874,N_7649,N_7601);
nand U7875 (N_7875,N_7795,N_7752);
and U7876 (N_7876,N_7696,N_7604);
xnor U7877 (N_7877,N_7731,N_7722);
and U7878 (N_7878,N_7635,N_7755);
xnor U7879 (N_7879,N_7760,N_7770);
xnor U7880 (N_7880,N_7769,N_7623);
nand U7881 (N_7881,N_7728,N_7659);
and U7882 (N_7882,N_7742,N_7636);
nor U7883 (N_7883,N_7654,N_7602);
and U7884 (N_7884,N_7725,N_7777);
nor U7885 (N_7885,N_7747,N_7630);
nor U7886 (N_7886,N_7619,N_7733);
nand U7887 (N_7887,N_7662,N_7677);
nor U7888 (N_7888,N_7698,N_7761);
nor U7889 (N_7889,N_7779,N_7603);
xnor U7890 (N_7890,N_7607,N_7670);
and U7891 (N_7891,N_7642,N_7645);
and U7892 (N_7892,N_7712,N_7753);
nand U7893 (N_7893,N_7723,N_7784);
nand U7894 (N_7894,N_7768,N_7711);
nand U7895 (N_7895,N_7704,N_7709);
nand U7896 (N_7896,N_7611,N_7605);
nand U7897 (N_7897,N_7653,N_7674);
nor U7898 (N_7898,N_7793,N_7775);
nand U7899 (N_7899,N_7657,N_7735);
and U7900 (N_7900,N_7724,N_7648);
nand U7901 (N_7901,N_7675,N_7679);
xnor U7902 (N_7902,N_7793,N_7641);
or U7903 (N_7903,N_7765,N_7711);
nor U7904 (N_7904,N_7674,N_7666);
or U7905 (N_7905,N_7767,N_7614);
nor U7906 (N_7906,N_7630,N_7727);
xor U7907 (N_7907,N_7618,N_7613);
or U7908 (N_7908,N_7697,N_7782);
and U7909 (N_7909,N_7773,N_7748);
or U7910 (N_7910,N_7737,N_7627);
and U7911 (N_7911,N_7744,N_7795);
xor U7912 (N_7912,N_7614,N_7661);
nand U7913 (N_7913,N_7637,N_7662);
nor U7914 (N_7914,N_7692,N_7777);
nand U7915 (N_7915,N_7661,N_7710);
nor U7916 (N_7916,N_7757,N_7739);
and U7917 (N_7917,N_7784,N_7694);
xnor U7918 (N_7918,N_7739,N_7756);
nand U7919 (N_7919,N_7730,N_7720);
nor U7920 (N_7920,N_7666,N_7618);
nand U7921 (N_7921,N_7773,N_7685);
nor U7922 (N_7922,N_7612,N_7696);
or U7923 (N_7923,N_7726,N_7621);
xor U7924 (N_7924,N_7789,N_7754);
and U7925 (N_7925,N_7677,N_7756);
and U7926 (N_7926,N_7796,N_7733);
and U7927 (N_7927,N_7697,N_7709);
or U7928 (N_7928,N_7744,N_7746);
or U7929 (N_7929,N_7684,N_7718);
and U7930 (N_7930,N_7772,N_7784);
nand U7931 (N_7931,N_7614,N_7686);
nor U7932 (N_7932,N_7682,N_7772);
and U7933 (N_7933,N_7695,N_7682);
nand U7934 (N_7934,N_7678,N_7695);
or U7935 (N_7935,N_7644,N_7611);
or U7936 (N_7936,N_7715,N_7771);
and U7937 (N_7937,N_7674,N_7768);
nand U7938 (N_7938,N_7706,N_7720);
and U7939 (N_7939,N_7795,N_7725);
and U7940 (N_7940,N_7745,N_7724);
xor U7941 (N_7941,N_7752,N_7703);
or U7942 (N_7942,N_7642,N_7652);
and U7943 (N_7943,N_7761,N_7616);
or U7944 (N_7944,N_7654,N_7652);
nor U7945 (N_7945,N_7646,N_7615);
nor U7946 (N_7946,N_7603,N_7609);
nor U7947 (N_7947,N_7719,N_7688);
nand U7948 (N_7948,N_7612,N_7690);
or U7949 (N_7949,N_7753,N_7716);
nor U7950 (N_7950,N_7784,N_7779);
and U7951 (N_7951,N_7777,N_7690);
nor U7952 (N_7952,N_7621,N_7640);
xnor U7953 (N_7953,N_7643,N_7655);
and U7954 (N_7954,N_7744,N_7678);
nor U7955 (N_7955,N_7683,N_7779);
and U7956 (N_7956,N_7752,N_7770);
nand U7957 (N_7957,N_7621,N_7607);
nor U7958 (N_7958,N_7728,N_7673);
nor U7959 (N_7959,N_7659,N_7677);
xnor U7960 (N_7960,N_7718,N_7733);
nand U7961 (N_7961,N_7792,N_7738);
nand U7962 (N_7962,N_7681,N_7604);
and U7963 (N_7963,N_7641,N_7785);
and U7964 (N_7964,N_7661,N_7765);
nand U7965 (N_7965,N_7635,N_7681);
xnor U7966 (N_7966,N_7683,N_7731);
nor U7967 (N_7967,N_7690,N_7643);
and U7968 (N_7968,N_7756,N_7663);
nand U7969 (N_7969,N_7774,N_7667);
and U7970 (N_7970,N_7699,N_7665);
xor U7971 (N_7971,N_7676,N_7769);
nand U7972 (N_7972,N_7672,N_7616);
xor U7973 (N_7973,N_7642,N_7786);
nand U7974 (N_7974,N_7604,N_7726);
nor U7975 (N_7975,N_7797,N_7739);
or U7976 (N_7976,N_7722,N_7716);
or U7977 (N_7977,N_7733,N_7779);
nor U7978 (N_7978,N_7765,N_7780);
or U7979 (N_7979,N_7685,N_7795);
nand U7980 (N_7980,N_7666,N_7743);
nor U7981 (N_7981,N_7627,N_7717);
xnor U7982 (N_7982,N_7697,N_7746);
xnor U7983 (N_7983,N_7619,N_7729);
and U7984 (N_7984,N_7795,N_7630);
and U7985 (N_7985,N_7689,N_7643);
nand U7986 (N_7986,N_7689,N_7684);
xor U7987 (N_7987,N_7710,N_7615);
or U7988 (N_7988,N_7699,N_7628);
and U7989 (N_7989,N_7758,N_7655);
nand U7990 (N_7990,N_7634,N_7730);
nor U7991 (N_7991,N_7648,N_7626);
nor U7992 (N_7992,N_7610,N_7632);
nor U7993 (N_7993,N_7624,N_7646);
and U7994 (N_7994,N_7652,N_7792);
xnor U7995 (N_7995,N_7636,N_7710);
or U7996 (N_7996,N_7714,N_7672);
or U7997 (N_7997,N_7694,N_7752);
nor U7998 (N_7998,N_7796,N_7760);
and U7999 (N_7999,N_7666,N_7687);
or U8000 (N_8000,N_7936,N_7914);
xnor U8001 (N_8001,N_7805,N_7855);
and U8002 (N_8002,N_7909,N_7815);
nand U8003 (N_8003,N_7854,N_7835);
xor U8004 (N_8004,N_7957,N_7942);
nand U8005 (N_8005,N_7965,N_7924);
xor U8006 (N_8006,N_7919,N_7865);
nor U8007 (N_8007,N_7853,N_7923);
or U8008 (N_8008,N_7991,N_7838);
nand U8009 (N_8009,N_7849,N_7820);
xnor U8010 (N_8010,N_7932,N_7943);
nor U8011 (N_8011,N_7883,N_7902);
nand U8012 (N_8012,N_7968,N_7867);
nand U8013 (N_8013,N_7900,N_7920);
xor U8014 (N_8014,N_7964,N_7947);
or U8015 (N_8015,N_7903,N_7904);
or U8016 (N_8016,N_7847,N_7983);
and U8017 (N_8017,N_7810,N_7801);
or U8018 (N_8018,N_7871,N_7921);
and U8019 (N_8019,N_7831,N_7858);
nor U8020 (N_8020,N_7963,N_7825);
nand U8021 (N_8021,N_7892,N_7861);
nor U8022 (N_8022,N_7982,N_7966);
or U8023 (N_8023,N_7811,N_7999);
xnor U8024 (N_8024,N_7972,N_7954);
and U8025 (N_8025,N_7944,N_7852);
xor U8026 (N_8026,N_7864,N_7851);
xor U8027 (N_8027,N_7818,N_7837);
nand U8028 (N_8028,N_7971,N_7830);
or U8029 (N_8029,N_7819,N_7875);
and U8030 (N_8030,N_7806,N_7908);
nand U8031 (N_8031,N_7891,N_7812);
and U8032 (N_8032,N_7824,N_7984);
nand U8033 (N_8033,N_7844,N_7856);
nand U8034 (N_8034,N_7846,N_7868);
nand U8035 (N_8035,N_7906,N_7990);
nand U8036 (N_8036,N_7840,N_7836);
nand U8037 (N_8037,N_7960,N_7809);
xnor U8038 (N_8038,N_7981,N_7933);
nand U8039 (N_8039,N_7834,N_7860);
or U8040 (N_8040,N_7962,N_7956);
and U8041 (N_8041,N_7877,N_7827);
and U8042 (N_8042,N_7918,N_7881);
xor U8043 (N_8043,N_7833,N_7959);
xor U8044 (N_8044,N_7803,N_7970);
nor U8045 (N_8045,N_7872,N_7882);
nor U8046 (N_8046,N_7922,N_7988);
nand U8047 (N_8047,N_7961,N_7949);
and U8048 (N_8048,N_7886,N_7866);
nor U8049 (N_8049,N_7980,N_7925);
nor U8050 (N_8050,N_7814,N_7989);
nor U8051 (N_8051,N_7994,N_7895);
nor U8052 (N_8052,N_7884,N_7841);
xnor U8053 (N_8053,N_7978,N_7829);
nor U8054 (N_8054,N_7817,N_7905);
nor U8055 (N_8055,N_7993,N_7889);
nand U8056 (N_8056,N_7870,N_7941);
xor U8057 (N_8057,N_7823,N_7985);
or U8058 (N_8058,N_7930,N_7907);
xor U8059 (N_8059,N_7850,N_7939);
or U8060 (N_8060,N_7979,N_7808);
or U8061 (N_8061,N_7948,N_7816);
xor U8062 (N_8062,N_7926,N_7931);
xor U8063 (N_8063,N_7952,N_7896);
and U8064 (N_8064,N_7927,N_7928);
and U8065 (N_8065,N_7813,N_7910);
or U8066 (N_8066,N_7987,N_7826);
and U8067 (N_8067,N_7888,N_7951);
nor U8068 (N_8068,N_7832,N_7958);
nand U8069 (N_8069,N_7975,N_7974);
or U8070 (N_8070,N_7953,N_7899);
or U8071 (N_8071,N_7992,N_7822);
nor U8072 (N_8072,N_7885,N_7879);
xnor U8073 (N_8073,N_7901,N_7940);
or U8074 (N_8074,N_7839,N_7898);
nand U8075 (N_8075,N_7912,N_7845);
and U8076 (N_8076,N_7874,N_7955);
xor U8077 (N_8077,N_7828,N_7913);
xor U8078 (N_8078,N_7973,N_7998);
xnor U8079 (N_8079,N_7807,N_7915);
or U8080 (N_8080,N_7911,N_7946);
nand U8081 (N_8081,N_7976,N_7929);
nor U8082 (N_8082,N_7862,N_7917);
or U8083 (N_8083,N_7937,N_7880);
xor U8084 (N_8084,N_7945,N_7997);
and U8085 (N_8085,N_7863,N_7800);
and U8086 (N_8086,N_7857,N_7938);
xnor U8087 (N_8087,N_7996,N_7950);
or U8088 (N_8088,N_7977,N_7842);
or U8089 (N_8089,N_7859,N_7995);
nor U8090 (N_8090,N_7893,N_7876);
xor U8091 (N_8091,N_7869,N_7848);
and U8092 (N_8092,N_7890,N_7821);
nor U8093 (N_8093,N_7887,N_7967);
nor U8094 (N_8094,N_7894,N_7986);
or U8095 (N_8095,N_7897,N_7969);
xnor U8096 (N_8096,N_7916,N_7804);
nand U8097 (N_8097,N_7843,N_7802);
nand U8098 (N_8098,N_7873,N_7935);
xnor U8099 (N_8099,N_7878,N_7934);
nand U8100 (N_8100,N_7904,N_7997);
nor U8101 (N_8101,N_7814,N_7832);
and U8102 (N_8102,N_7939,N_7998);
nand U8103 (N_8103,N_7812,N_7925);
nor U8104 (N_8104,N_7940,N_7978);
or U8105 (N_8105,N_7839,N_7974);
xor U8106 (N_8106,N_7863,N_7841);
nor U8107 (N_8107,N_7956,N_7957);
and U8108 (N_8108,N_7841,N_7836);
or U8109 (N_8109,N_7848,N_7986);
nor U8110 (N_8110,N_7872,N_7900);
nor U8111 (N_8111,N_7940,N_7914);
and U8112 (N_8112,N_7929,N_7868);
nand U8113 (N_8113,N_7815,N_7896);
xnor U8114 (N_8114,N_7842,N_7867);
xnor U8115 (N_8115,N_7992,N_7859);
nand U8116 (N_8116,N_7862,N_7827);
xnor U8117 (N_8117,N_7925,N_7873);
nand U8118 (N_8118,N_7922,N_7886);
nand U8119 (N_8119,N_7893,N_7826);
nand U8120 (N_8120,N_7883,N_7984);
nand U8121 (N_8121,N_7964,N_7874);
or U8122 (N_8122,N_7966,N_7913);
nor U8123 (N_8123,N_7895,N_7808);
or U8124 (N_8124,N_7903,N_7965);
xnor U8125 (N_8125,N_7926,N_7846);
xnor U8126 (N_8126,N_7901,N_7855);
nand U8127 (N_8127,N_7848,N_7812);
nand U8128 (N_8128,N_7872,N_7865);
or U8129 (N_8129,N_7890,N_7916);
xnor U8130 (N_8130,N_7930,N_7874);
nor U8131 (N_8131,N_7994,N_7876);
nand U8132 (N_8132,N_7892,N_7846);
xor U8133 (N_8133,N_7917,N_7999);
and U8134 (N_8134,N_7837,N_7839);
nor U8135 (N_8135,N_7879,N_7899);
xnor U8136 (N_8136,N_7803,N_7831);
xor U8137 (N_8137,N_7866,N_7977);
nand U8138 (N_8138,N_7945,N_7857);
nand U8139 (N_8139,N_7871,N_7878);
and U8140 (N_8140,N_7968,N_7906);
and U8141 (N_8141,N_7801,N_7914);
and U8142 (N_8142,N_7904,N_7901);
or U8143 (N_8143,N_7800,N_7820);
xor U8144 (N_8144,N_7921,N_7919);
xor U8145 (N_8145,N_7916,N_7802);
nor U8146 (N_8146,N_7997,N_7814);
or U8147 (N_8147,N_7890,N_7989);
nor U8148 (N_8148,N_7840,N_7967);
or U8149 (N_8149,N_7834,N_7911);
and U8150 (N_8150,N_7827,N_7834);
xor U8151 (N_8151,N_7858,N_7852);
or U8152 (N_8152,N_7909,N_7866);
or U8153 (N_8153,N_7945,N_7993);
nand U8154 (N_8154,N_7997,N_7834);
or U8155 (N_8155,N_7828,N_7838);
nand U8156 (N_8156,N_7965,N_7917);
nor U8157 (N_8157,N_7825,N_7988);
or U8158 (N_8158,N_7866,N_7851);
and U8159 (N_8159,N_7985,N_7863);
or U8160 (N_8160,N_7957,N_7961);
nand U8161 (N_8161,N_7982,N_7981);
xor U8162 (N_8162,N_7883,N_7859);
nor U8163 (N_8163,N_7999,N_7957);
xnor U8164 (N_8164,N_7858,N_7838);
xor U8165 (N_8165,N_7812,N_7939);
nor U8166 (N_8166,N_7872,N_7911);
and U8167 (N_8167,N_7908,N_7966);
xnor U8168 (N_8168,N_7996,N_7932);
xnor U8169 (N_8169,N_7855,N_7998);
and U8170 (N_8170,N_7901,N_7824);
nand U8171 (N_8171,N_7911,N_7805);
xnor U8172 (N_8172,N_7866,N_7925);
nor U8173 (N_8173,N_7895,N_7851);
xor U8174 (N_8174,N_7878,N_7900);
or U8175 (N_8175,N_7935,N_7870);
nor U8176 (N_8176,N_7854,N_7955);
or U8177 (N_8177,N_7875,N_7835);
nand U8178 (N_8178,N_7845,N_7989);
and U8179 (N_8179,N_7870,N_7896);
nor U8180 (N_8180,N_7939,N_7938);
nor U8181 (N_8181,N_7930,N_7942);
nand U8182 (N_8182,N_7898,N_7880);
nand U8183 (N_8183,N_7906,N_7833);
or U8184 (N_8184,N_7921,N_7934);
xor U8185 (N_8185,N_7973,N_7962);
and U8186 (N_8186,N_7841,N_7885);
or U8187 (N_8187,N_7811,N_7993);
xor U8188 (N_8188,N_7987,N_7950);
and U8189 (N_8189,N_7866,N_7979);
or U8190 (N_8190,N_7853,N_7970);
xnor U8191 (N_8191,N_7802,N_7969);
or U8192 (N_8192,N_7972,N_7889);
nand U8193 (N_8193,N_7852,N_7966);
nand U8194 (N_8194,N_7876,N_7827);
and U8195 (N_8195,N_7884,N_7991);
and U8196 (N_8196,N_7915,N_7857);
and U8197 (N_8197,N_7922,N_7953);
or U8198 (N_8198,N_7979,N_7904);
or U8199 (N_8199,N_7861,N_7849);
xnor U8200 (N_8200,N_8173,N_8029);
xnor U8201 (N_8201,N_8060,N_8034);
nand U8202 (N_8202,N_8136,N_8083);
nor U8203 (N_8203,N_8115,N_8021);
xnor U8204 (N_8204,N_8050,N_8061);
and U8205 (N_8205,N_8056,N_8195);
nor U8206 (N_8206,N_8129,N_8080);
xor U8207 (N_8207,N_8069,N_8166);
nand U8208 (N_8208,N_8110,N_8030);
nand U8209 (N_8209,N_8108,N_8118);
or U8210 (N_8210,N_8087,N_8172);
and U8211 (N_8211,N_8179,N_8145);
nand U8212 (N_8212,N_8123,N_8001);
xnor U8213 (N_8213,N_8192,N_8152);
nor U8214 (N_8214,N_8103,N_8187);
nor U8215 (N_8215,N_8081,N_8065);
nor U8216 (N_8216,N_8183,N_8093);
xnor U8217 (N_8217,N_8137,N_8160);
and U8218 (N_8218,N_8007,N_8058);
xnor U8219 (N_8219,N_8059,N_8119);
nand U8220 (N_8220,N_8150,N_8185);
and U8221 (N_8221,N_8017,N_8113);
or U8222 (N_8222,N_8067,N_8116);
nor U8223 (N_8223,N_8042,N_8146);
xnor U8224 (N_8224,N_8157,N_8178);
nand U8225 (N_8225,N_8043,N_8097);
xnor U8226 (N_8226,N_8182,N_8151);
nand U8227 (N_8227,N_8165,N_8154);
nor U8228 (N_8228,N_8031,N_8163);
nand U8229 (N_8229,N_8088,N_8077);
nand U8230 (N_8230,N_8133,N_8010);
and U8231 (N_8231,N_8106,N_8144);
xnor U8232 (N_8232,N_8057,N_8134);
and U8233 (N_8233,N_8068,N_8082);
or U8234 (N_8234,N_8120,N_8096);
nand U8235 (N_8235,N_8126,N_8090);
xor U8236 (N_8236,N_8111,N_8175);
or U8237 (N_8237,N_8070,N_8194);
or U8238 (N_8238,N_8078,N_8180);
nand U8239 (N_8239,N_8009,N_8184);
and U8240 (N_8240,N_8188,N_8064);
nor U8241 (N_8241,N_8045,N_8041);
and U8242 (N_8242,N_8162,N_8117);
and U8243 (N_8243,N_8100,N_8135);
or U8244 (N_8244,N_8053,N_8038);
nor U8245 (N_8245,N_8156,N_8148);
nor U8246 (N_8246,N_8142,N_8084);
nor U8247 (N_8247,N_8073,N_8141);
xnor U8248 (N_8248,N_8048,N_8107);
nand U8249 (N_8249,N_8066,N_8189);
or U8250 (N_8250,N_8130,N_8072);
or U8251 (N_8251,N_8006,N_8159);
xnor U8252 (N_8252,N_8023,N_8000);
nor U8253 (N_8253,N_8051,N_8170);
nand U8254 (N_8254,N_8075,N_8005);
nand U8255 (N_8255,N_8062,N_8104);
nor U8256 (N_8256,N_8013,N_8197);
nand U8257 (N_8257,N_8138,N_8158);
and U8258 (N_8258,N_8124,N_8025);
or U8259 (N_8259,N_8019,N_8109);
or U8260 (N_8260,N_8004,N_8012);
xnor U8261 (N_8261,N_8168,N_8063);
xor U8262 (N_8262,N_8121,N_8085);
nand U8263 (N_8263,N_8127,N_8054);
nor U8264 (N_8264,N_8149,N_8139);
nor U8265 (N_8265,N_8055,N_8174);
and U8266 (N_8266,N_8052,N_8186);
xnor U8267 (N_8267,N_8022,N_8177);
or U8268 (N_8268,N_8181,N_8015);
nor U8269 (N_8269,N_8176,N_8089);
and U8270 (N_8270,N_8128,N_8105);
or U8271 (N_8271,N_8016,N_8102);
nand U8272 (N_8272,N_8114,N_8079);
nor U8273 (N_8273,N_8026,N_8171);
nand U8274 (N_8274,N_8037,N_8169);
or U8275 (N_8275,N_8143,N_8167);
or U8276 (N_8276,N_8147,N_8035);
or U8277 (N_8277,N_8036,N_8091);
or U8278 (N_8278,N_8086,N_8011);
nor U8279 (N_8279,N_8018,N_8024);
nor U8280 (N_8280,N_8027,N_8020);
or U8281 (N_8281,N_8122,N_8199);
or U8282 (N_8282,N_8155,N_8071);
and U8283 (N_8283,N_8098,N_8161);
nor U8284 (N_8284,N_8196,N_8125);
nor U8285 (N_8285,N_8140,N_8076);
xnor U8286 (N_8286,N_8074,N_8132);
and U8287 (N_8287,N_8014,N_8095);
nand U8288 (N_8288,N_8101,N_8112);
and U8289 (N_8289,N_8099,N_8008);
nand U8290 (N_8290,N_8049,N_8040);
or U8291 (N_8291,N_8044,N_8193);
xnor U8292 (N_8292,N_8032,N_8033);
and U8293 (N_8293,N_8164,N_8047);
nor U8294 (N_8294,N_8131,N_8153);
xnor U8295 (N_8295,N_8003,N_8198);
nor U8296 (N_8296,N_8092,N_8094);
nand U8297 (N_8297,N_8191,N_8190);
or U8298 (N_8298,N_8039,N_8002);
xor U8299 (N_8299,N_8028,N_8046);
and U8300 (N_8300,N_8022,N_8009);
or U8301 (N_8301,N_8161,N_8189);
nor U8302 (N_8302,N_8142,N_8114);
xnor U8303 (N_8303,N_8173,N_8188);
and U8304 (N_8304,N_8026,N_8194);
xor U8305 (N_8305,N_8133,N_8186);
and U8306 (N_8306,N_8050,N_8046);
xnor U8307 (N_8307,N_8192,N_8118);
nor U8308 (N_8308,N_8071,N_8003);
nand U8309 (N_8309,N_8052,N_8040);
nor U8310 (N_8310,N_8199,N_8019);
nand U8311 (N_8311,N_8070,N_8025);
nand U8312 (N_8312,N_8052,N_8097);
nand U8313 (N_8313,N_8101,N_8013);
xor U8314 (N_8314,N_8073,N_8055);
or U8315 (N_8315,N_8032,N_8066);
and U8316 (N_8316,N_8016,N_8198);
and U8317 (N_8317,N_8050,N_8004);
nor U8318 (N_8318,N_8191,N_8061);
xor U8319 (N_8319,N_8187,N_8162);
nand U8320 (N_8320,N_8167,N_8042);
or U8321 (N_8321,N_8145,N_8028);
or U8322 (N_8322,N_8161,N_8107);
or U8323 (N_8323,N_8107,N_8149);
and U8324 (N_8324,N_8114,N_8078);
or U8325 (N_8325,N_8091,N_8167);
nand U8326 (N_8326,N_8077,N_8010);
and U8327 (N_8327,N_8078,N_8152);
nor U8328 (N_8328,N_8182,N_8028);
and U8329 (N_8329,N_8186,N_8044);
nor U8330 (N_8330,N_8112,N_8158);
and U8331 (N_8331,N_8119,N_8189);
nand U8332 (N_8332,N_8053,N_8018);
nand U8333 (N_8333,N_8000,N_8127);
or U8334 (N_8334,N_8138,N_8051);
xor U8335 (N_8335,N_8171,N_8142);
or U8336 (N_8336,N_8175,N_8104);
and U8337 (N_8337,N_8129,N_8058);
or U8338 (N_8338,N_8103,N_8174);
or U8339 (N_8339,N_8055,N_8037);
nand U8340 (N_8340,N_8064,N_8161);
xor U8341 (N_8341,N_8119,N_8023);
or U8342 (N_8342,N_8052,N_8162);
and U8343 (N_8343,N_8164,N_8023);
nor U8344 (N_8344,N_8110,N_8166);
nand U8345 (N_8345,N_8145,N_8095);
nor U8346 (N_8346,N_8057,N_8152);
nor U8347 (N_8347,N_8142,N_8105);
and U8348 (N_8348,N_8060,N_8130);
xnor U8349 (N_8349,N_8082,N_8027);
nand U8350 (N_8350,N_8044,N_8074);
or U8351 (N_8351,N_8124,N_8094);
xor U8352 (N_8352,N_8186,N_8132);
or U8353 (N_8353,N_8035,N_8190);
xor U8354 (N_8354,N_8137,N_8109);
nor U8355 (N_8355,N_8142,N_8194);
or U8356 (N_8356,N_8178,N_8066);
or U8357 (N_8357,N_8071,N_8056);
or U8358 (N_8358,N_8026,N_8122);
nand U8359 (N_8359,N_8047,N_8050);
xnor U8360 (N_8360,N_8024,N_8062);
xnor U8361 (N_8361,N_8066,N_8185);
or U8362 (N_8362,N_8191,N_8044);
or U8363 (N_8363,N_8034,N_8008);
and U8364 (N_8364,N_8131,N_8013);
xor U8365 (N_8365,N_8088,N_8198);
xnor U8366 (N_8366,N_8194,N_8054);
nand U8367 (N_8367,N_8143,N_8173);
xor U8368 (N_8368,N_8112,N_8094);
xnor U8369 (N_8369,N_8118,N_8107);
or U8370 (N_8370,N_8132,N_8150);
nor U8371 (N_8371,N_8073,N_8037);
or U8372 (N_8372,N_8053,N_8139);
and U8373 (N_8373,N_8088,N_8156);
xnor U8374 (N_8374,N_8154,N_8125);
and U8375 (N_8375,N_8107,N_8124);
and U8376 (N_8376,N_8132,N_8002);
nand U8377 (N_8377,N_8151,N_8112);
nor U8378 (N_8378,N_8116,N_8096);
nor U8379 (N_8379,N_8137,N_8077);
nor U8380 (N_8380,N_8096,N_8046);
and U8381 (N_8381,N_8067,N_8180);
xnor U8382 (N_8382,N_8080,N_8191);
xor U8383 (N_8383,N_8062,N_8177);
xnor U8384 (N_8384,N_8146,N_8019);
nor U8385 (N_8385,N_8001,N_8081);
xnor U8386 (N_8386,N_8153,N_8107);
xor U8387 (N_8387,N_8131,N_8162);
nand U8388 (N_8388,N_8189,N_8129);
xor U8389 (N_8389,N_8106,N_8038);
xor U8390 (N_8390,N_8171,N_8061);
and U8391 (N_8391,N_8111,N_8126);
xnor U8392 (N_8392,N_8058,N_8015);
xnor U8393 (N_8393,N_8047,N_8180);
xnor U8394 (N_8394,N_8022,N_8111);
nor U8395 (N_8395,N_8019,N_8041);
and U8396 (N_8396,N_8154,N_8041);
nor U8397 (N_8397,N_8094,N_8130);
xnor U8398 (N_8398,N_8012,N_8187);
or U8399 (N_8399,N_8089,N_8019);
and U8400 (N_8400,N_8330,N_8356);
nand U8401 (N_8401,N_8345,N_8386);
nand U8402 (N_8402,N_8397,N_8375);
or U8403 (N_8403,N_8202,N_8266);
or U8404 (N_8404,N_8370,N_8372);
nor U8405 (N_8405,N_8265,N_8312);
and U8406 (N_8406,N_8389,N_8220);
or U8407 (N_8407,N_8213,N_8247);
or U8408 (N_8408,N_8333,N_8344);
nor U8409 (N_8409,N_8218,N_8359);
and U8410 (N_8410,N_8297,N_8373);
or U8411 (N_8411,N_8355,N_8200);
nand U8412 (N_8412,N_8233,N_8270);
xnor U8413 (N_8413,N_8276,N_8310);
or U8414 (N_8414,N_8380,N_8206);
and U8415 (N_8415,N_8352,N_8399);
nor U8416 (N_8416,N_8201,N_8240);
xor U8417 (N_8417,N_8319,N_8304);
or U8418 (N_8418,N_8347,N_8298);
xor U8419 (N_8419,N_8314,N_8289);
and U8420 (N_8420,N_8362,N_8396);
xnor U8421 (N_8421,N_8290,N_8209);
nor U8422 (N_8422,N_8281,N_8221);
and U8423 (N_8423,N_8274,N_8231);
nor U8424 (N_8424,N_8350,N_8217);
xor U8425 (N_8425,N_8249,N_8394);
xor U8426 (N_8426,N_8339,N_8280);
and U8427 (N_8427,N_8351,N_8207);
nor U8428 (N_8428,N_8368,N_8239);
xor U8429 (N_8429,N_8353,N_8210);
or U8430 (N_8430,N_8323,N_8387);
nand U8431 (N_8431,N_8367,N_8252);
nor U8432 (N_8432,N_8328,N_8301);
xnor U8433 (N_8433,N_8235,N_8379);
nor U8434 (N_8434,N_8322,N_8300);
xor U8435 (N_8435,N_8237,N_8326);
xor U8436 (N_8436,N_8325,N_8234);
and U8437 (N_8437,N_8268,N_8261);
and U8438 (N_8438,N_8294,N_8243);
nand U8439 (N_8439,N_8321,N_8285);
nor U8440 (N_8440,N_8263,N_8226);
xor U8441 (N_8441,N_8264,N_8222);
xor U8442 (N_8442,N_8331,N_8324);
nand U8443 (N_8443,N_8296,N_8377);
nor U8444 (N_8444,N_8305,N_8346);
xnor U8445 (N_8445,N_8215,N_8267);
and U8446 (N_8446,N_8291,N_8395);
and U8447 (N_8447,N_8251,N_8336);
nand U8448 (N_8448,N_8241,N_8259);
nand U8449 (N_8449,N_8306,N_8364);
nand U8450 (N_8450,N_8230,N_8371);
nand U8451 (N_8451,N_8303,N_8316);
xor U8452 (N_8452,N_8273,N_8392);
nand U8453 (N_8453,N_8309,N_8388);
xnor U8454 (N_8454,N_8385,N_8258);
or U8455 (N_8455,N_8256,N_8382);
or U8456 (N_8456,N_8216,N_8320);
or U8457 (N_8457,N_8302,N_8378);
nor U8458 (N_8458,N_8229,N_8327);
nand U8459 (N_8459,N_8342,N_8269);
xor U8460 (N_8460,N_8376,N_8204);
nor U8461 (N_8461,N_8246,N_8255);
xnor U8462 (N_8462,N_8203,N_8363);
and U8463 (N_8463,N_8260,N_8253);
or U8464 (N_8464,N_8236,N_8393);
nor U8465 (N_8465,N_8348,N_8248);
nor U8466 (N_8466,N_8299,N_8313);
and U8467 (N_8467,N_8288,N_8357);
nor U8468 (N_8468,N_8374,N_8225);
or U8469 (N_8469,N_8343,N_8383);
nand U8470 (N_8470,N_8272,N_8334);
nor U8471 (N_8471,N_8337,N_8354);
nand U8472 (N_8472,N_8295,N_8232);
nor U8473 (N_8473,N_8315,N_8384);
or U8474 (N_8474,N_8242,N_8358);
and U8475 (N_8475,N_8398,N_8293);
xor U8476 (N_8476,N_8365,N_8341);
nand U8477 (N_8477,N_8271,N_8279);
nor U8478 (N_8478,N_8244,N_8257);
nand U8479 (N_8479,N_8292,N_8283);
and U8480 (N_8480,N_8286,N_8211);
and U8481 (N_8481,N_8282,N_8390);
nor U8482 (N_8482,N_8349,N_8318);
nor U8483 (N_8483,N_8278,N_8338);
xnor U8484 (N_8484,N_8238,N_8205);
and U8485 (N_8485,N_8332,N_8275);
and U8486 (N_8486,N_8311,N_8340);
nand U8487 (N_8487,N_8219,N_8245);
nor U8488 (N_8488,N_8381,N_8277);
or U8489 (N_8489,N_8227,N_8369);
nor U8490 (N_8490,N_8223,N_8214);
or U8491 (N_8491,N_8212,N_8317);
nor U8492 (N_8492,N_8366,N_8308);
nand U8493 (N_8493,N_8335,N_8361);
xnor U8494 (N_8494,N_8262,N_8284);
xnor U8495 (N_8495,N_8224,N_8307);
or U8496 (N_8496,N_8208,N_8250);
nand U8497 (N_8497,N_8391,N_8254);
nor U8498 (N_8498,N_8287,N_8329);
nand U8499 (N_8499,N_8360,N_8228);
or U8500 (N_8500,N_8253,N_8204);
nor U8501 (N_8501,N_8221,N_8252);
or U8502 (N_8502,N_8323,N_8282);
and U8503 (N_8503,N_8215,N_8368);
nand U8504 (N_8504,N_8333,N_8308);
and U8505 (N_8505,N_8227,N_8371);
nor U8506 (N_8506,N_8210,N_8366);
and U8507 (N_8507,N_8218,N_8352);
and U8508 (N_8508,N_8252,N_8394);
nor U8509 (N_8509,N_8306,N_8279);
xor U8510 (N_8510,N_8334,N_8269);
xor U8511 (N_8511,N_8391,N_8276);
nor U8512 (N_8512,N_8270,N_8325);
and U8513 (N_8513,N_8298,N_8348);
xor U8514 (N_8514,N_8202,N_8291);
xnor U8515 (N_8515,N_8312,N_8294);
or U8516 (N_8516,N_8395,N_8250);
nand U8517 (N_8517,N_8264,N_8356);
nand U8518 (N_8518,N_8280,N_8307);
nand U8519 (N_8519,N_8318,N_8328);
or U8520 (N_8520,N_8355,N_8241);
xnor U8521 (N_8521,N_8327,N_8267);
nand U8522 (N_8522,N_8381,N_8307);
nand U8523 (N_8523,N_8221,N_8228);
nand U8524 (N_8524,N_8224,N_8303);
nor U8525 (N_8525,N_8299,N_8230);
nor U8526 (N_8526,N_8308,N_8324);
xnor U8527 (N_8527,N_8310,N_8322);
or U8528 (N_8528,N_8329,N_8394);
or U8529 (N_8529,N_8273,N_8211);
nor U8530 (N_8530,N_8277,N_8291);
nand U8531 (N_8531,N_8329,N_8278);
nand U8532 (N_8532,N_8307,N_8232);
and U8533 (N_8533,N_8397,N_8204);
or U8534 (N_8534,N_8359,N_8394);
xnor U8535 (N_8535,N_8374,N_8369);
xnor U8536 (N_8536,N_8221,N_8292);
and U8537 (N_8537,N_8308,N_8375);
or U8538 (N_8538,N_8394,N_8374);
xor U8539 (N_8539,N_8346,N_8254);
and U8540 (N_8540,N_8381,N_8317);
nor U8541 (N_8541,N_8200,N_8398);
nor U8542 (N_8542,N_8346,N_8210);
and U8543 (N_8543,N_8349,N_8369);
nand U8544 (N_8544,N_8223,N_8203);
nand U8545 (N_8545,N_8361,N_8365);
xnor U8546 (N_8546,N_8335,N_8360);
xor U8547 (N_8547,N_8214,N_8308);
or U8548 (N_8548,N_8272,N_8389);
nor U8549 (N_8549,N_8308,N_8263);
nand U8550 (N_8550,N_8243,N_8273);
nand U8551 (N_8551,N_8206,N_8356);
or U8552 (N_8552,N_8280,N_8399);
nand U8553 (N_8553,N_8296,N_8209);
xor U8554 (N_8554,N_8308,N_8265);
or U8555 (N_8555,N_8395,N_8234);
xor U8556 (N_8556,N_8231,N_8354);
xnor U8557 (N_8557,N_8263,N_8220);
or U8558 (N_8558,N_8322,N_8258);
xor U8559 (N_8559,N_8380,N_8217);
xor U8560 (N_8560,N_8205,N_8258);
and U8561 (N_8561,N_8342,N_8238);
nor U8562 (N_8562,N_8202,N_8314);
xnor U8563 (N_8563,N_8305,N_8238);
xnor U8564 (N_8564,N_8270,N_8394);
xnor U8565 (N_8565,N_8207,N_8263);
xnor U8566 (N_8566,N_8284,N_8308);
xor U8567 (N_8567,N_8257,N_8311);
or U8568 (N_8568,N_8390,N_8223);
xor U8569 (N_8569,N_8310,N_8359);
nand U8570 (N_8570,N_8316,N_8318);
and U8571 (N_8571,N_8289,N_8395);
or U8572 (N_8572,N_8323,N_8286);
nand U8573 (N_8573,N_8318,N_8282);
xor U8574 (N_8574,N_8262,N_8396);
nor U8575 (N_8575,N_8382,N_8200);
nand U8576 (N_8576,N_8231,N_8223);
nor U8577 (N_8577,N_8352,N_8262);
and U8578 (N_8578,N_8240,N_8304);
and U8579 (N_8579,N_8358,N_8255);
or U8580 (N_8580,N_8316,N_8240);
nor U8581 (N_8581,N_8259,N_8218);
nor U8582 (N_8582,N_8398,N_8260);
or U8583 (N_8583,N_8242,N_8301);
and U8584 (N_8584,N_8399,N_8273);
nor U8585 (N_8585,N_8215,N_8296);
xor U8586 (N_8586,N_8317,N_8304);
nor U8587 (N_8587,N_8268,N_8283);
xnor U8588 (N_8588,N_8331,N_8378);
nand U8589 (N_8589,N_8289,N_8349);
nor U8590 (N_8590,N_8337,N_8280);
nor U8591 (N_8591,N_8364,N_8348);
xor U8592 (N_8592,N_8335,N_8318);
or U8593 (N_8593,N_8388,N_8300);
and U8594 (N_8594,N_8294,N_8382);
nor U8595 (N_8595,N_8363,N_8306);
xnor U8596 (N_8596,N_8216,N_8369);
or U8597 (N_8597,N_8345,N_8226);
xnor U8598 (N_8598,N_8391,N_8320);
or U8599 (N_8599,N_8378,N_8219);
or U8600 (N_8600,N_8589,N_8488);
nor U8601 (N_8601,N_8424,N_8422);
or U8602 (N_8602,N_8481,N_8474);
and U8603 (N_8603,N_8456,N_8453);
nand U8604 (N_8604,N_8597,N_8554);
or U8605 (N_8605,N_8490,N_8509);
nor U8606 (N_8606,N_8530,N_8418);
xor U8607 (N_8607,N_8493,N_8556);
and U8608 (N_8608,N_8403,N_8502);
and U8609 (N_8609,N_8516,N_8494);
nand U8610 (N_8610,N_8568,N_8455);
nor U8611 (N_8611,N_8436,N_8433);
xnor U8612 (N_8612,N_8435,N_8434);
nand U8613 (N_8613,N_8461,N_8573);
nand U8614 (N_8614,N_8599,N_8536);
xor U8615 (N_8615,N_8503,N_8552);
or U8616 (N_8616,N_8404,N_8457);
xor U8617 (N_8617,N_8441,N_8498);
or U8618 (N_8618,N_8505,N_8548);
nor U8619 (N_8619,N_8432,N_8480);
nor U8620 (N_8620,N_8588,N_8533);
nor U8621 (N_8621,N_8585,N_8529);
nand U8622 (N_8622,N_8586,N_8521);
xnor U8623 (N_8623,N_8473,N_8511);
xnor U8624 (N_8624,N_8469,N_8566);
xor U8625 (N_8625,N_8517,N_8584);
and U8626 (N_8626,N_8581,N_8537);
or U8627 (N_8627,N_8567,N_8497);
and U8628 (N_8628,N_8528,N_8541);
xnor U8629 (N_8629,N_8564,N_8510);
nand U8630 (N_8630,N_8519,N_8466);
xor U8631 (N_8631,N_8592,N_8414);
or U8632 (N_8632,N_8487,N_8460);
nand U8633 (N_8633,N_8405,N_8587);
nor U8634 (N_8634,N_8580,N_8440);
nor U8635 (N_8635,N_8472,N_8544);
nand U8636 (N_8636,N_8458,N_8508);
or U8637 (N_8637,N_8525,N_8479);
nand U8638 (N_8638,N_8527,N_8468);
nand U8639 (N_8639,N_8565,N_8448);
nor U8640 (N_8640,N_8524,N_8450);
or U8641 (N_8641,N_8591,N_8596);
or U8642 (N_8642,N_8431,N_8410);
and U8643 (N_8643,N_8492,N_8495);
xnor U8644 (N_8644,N_8579,N_8491);
nand U8645 (N_8645,N_8484,N_8421);
xnor U8646 (N_8646,N_8412,N_8423);
and U8647 (N_8647,N_8439,N_8583);
and U8648 (N_8648,N_8478,N_8542);
or U8649 (N_8649,N_8416,N_8430);
or U8650 (N_8650,N_8415,N_8520);
xor U8651 (N_8651,N_8593,N_8595);
xnor U8652 (N_8652,N_8406,N_8476);
nand U8653 (N_8653,N_8578,N_8535);
or U8654 (N_8654,N_8522,N_8549);
and U8655 (N_8655,N_8428,N_8558);
nand U8656 (N_8656,N_8545,N_8411);
and U8657 (N_8657,N_8553,N_8470);
or U8658 (N_8658,N_8485,N_8506);
or U8659 (N_8659,N_8429,N_8482);
nor U8660 (N_8660,N_8594,N_8486);
nand U8661 (N_8661,N_8402,N_8452);
nor U8662 (N_8662,N_8409,N_8417);
xnor U8663 (N_8663,N_8445,N_8561);
or U8664 (N_8664,N_8513,N_8538);
xnor U8665 (N_8665,N_8504,N_8570);
and U8666 (N_8666,N_8475,N_8489);
nor U8667 (N_8667,N_8562,N_8575);
xor U8668 (N_8668,N_8534,N_8467);
and U8669 (N_8669,N_8557,N_8569);
nor U8670 (N_8670,N_8571,N_8420);
and U8671 (N_8671,N_8427,N_8576);
or U8672 (N_8672,N_8419,N_8463);
xnor U8673 (N_8673,N_8526,N_8514);
and U8674 (N_8674,N_8449,N_8437);
nand U8675 (N_8675,N_8512,N_8446);
and U8676 (N_8676,N_8413,N_8559);
nand U8677 (N_8677,N_8543,N_8507);
nand U8678 (N_8678,N_8400,N_8515);
nand U8679 (N_8679,N_8451,N_8539);
nor U8680 (N_8680,N_8532,N_8501);
xor U8681 (N_8681,N_8518,N_8551);
nand U8682 (N_8682,N_8598,N_8438);
and U8683 (N_8683,N_8577,N_8499);
nor U8684 (N_8684,N_8550,N_8540);
nand U8685 (N_8685,N_8471,N_8500);
xnor U8686 (N_8686,N_8425,N_8531);
nor U8687 (N_8687,N_8408,N_8401);
xor U8688 (N_8688,N_8582,N_8442);
xor U8689 (N_8689,N_8443,N_8523);
nor U8690 (N_8690,N_8459,N_8462);
and U8691 (N_8691,N_8444,N_8563);
nand U8692 (N_8692,N_8464,N_8574);
nand U8693 (N_8693,N_8465,N_8447);
nand U8694 (N_8694,N_8590,N_8547);
nor U8695 (N_8695,N_8483,N_8572);
or U8696 (N_8696,N_8426,N_8407);
nor U8697 (N_8697,N_8546,N_8496);
and U8698 (N_8698,N_8560,N_8454);
and U8699 (N_8699,N_8477,N_8555);
nand U8700 (N_8700,N_8512,N_8458);
nand U8701 (N_8701,N_8504,N_8563);
nor U8702 (N_8702,N_8496,N_8419);
or U8703 (N_8703,N_8501,N_8544);
or U8704 (N_8704,N_8581,N_8438);
and U8705 (N_8705,N_8458,N_8423);
nand U8706 (N_8706,N_8582,N_8488);
and U8707 (N_8707,N_8405,N_8531);
or U8708 (N_8708,N_8555,N_8498);
nor U8709 (N_8709,N_8405,N_8582);
and U8710 (N_8710,N_8446,N_8416);
xor U8711 (N_8711,N_8480,N_8415);
and U8712 (N_8712,N_8426,N_8531);
or U8713 (N_8713,N_8500,N_8416);
nand U8714 (N_8714,N_8440,N_8562);
xor U8715 (N_8715,N_8584,N_8547);
xor U8716 (N_8716,N_8519,N_8537);
xor U8717 (N_8717,N_8532,N_8567);
and U8718 (N_8718,N_8518,N_8474);
nand U8719 (N_8719,N_8575,N_8421);
and U8720 (N_8720,N_8419,N_8461);
nand U8721 (N_8721,N_8581,N_8559);
and U8722 (N_8722,N_8404,N_8506);
or U8723 (N_8723,N_8468,N_8559);
nor U8724 (N_8724,N_8510,N_8539);
and U8725 (N_8725,N_8548,N_8516);
and U8726 (N_8726,N_8488,N_8555);
or U8727 (N_8727,N_8456,N_8468);
xnor U8728 (N_8728,N_8505,N_8405);
nor U8729 (N_8729,N_8519,N_8576);
and U8730 (N_8730,N_8537,N_8450);
nand U8731 (N_8731,N_8507,N_8442);
xnor U8732 (N_8732,N_8525,N_8437);
xor U8733 (N_8733,N_8492,N_8599);
xor U8734 (N_8734,N_8532,N_8536);
nor U8735 (N_8735,N_8438,N_8491);
or U8736 (N_8736,N_8484,N_8585);
nand U8737 (N_8737,N_8474,N_8578);
nand U8738 (N_8738,N_8422,N_8563);
nor U8739 (N_8739,N_8536,N_8424);
xor U8740 (N_8740,N_8441,N_8518);
or U8741 (N_8741,N_8454,N_8497);
or U8742 (N_8742,N_8486,N_8453);
nor U8743 (N_8743,N_8436,N_8539);
xor U8744 (N_8744,N_8558,N_8484);
or U8745 (N_8745,N_8434,N_8594);
nand U8746 (N_8746,N_8560,N_8586);
xor U8747 (N_8747,N_8516,N_8474);
and U8748 (N_8748,N_8455,N_8490);
xnor U8749 (N_8749,N_8529,N_8527);
xnor U8750 (N_8750,N_8432,N_8565);
nand U8751 (N_8751,N_8413,N_8506);
and U8752 (N_8752,N_8545,N_8422);
and U8753 (N_8753,N_8514,N_8598);
or U8754 (N_8754,N_8576,N_8459);
or U8755 (N_8755,N_8527,N_8444);
or U8756 (N_8756,N_8486,N_8508);
nand U8757 (N_8757,N_8422,N_8576);
nor U8758 (N_8758,N_8402,N_8571);
xor U8759 (N_8759,N_8487,N_8493);
and U8760 (N_8760,N_8421,N_8449);
xnor U8761 (N_8761,N_8422,N_8526);
nor U8762 (N_8762,N_8584,N_8465);
nor U8763 (N_8763,N_8558,N_8413);
xor U8764 (N_8764,N_8430,N_8466);
xnor U8765 (N_8765,N_8502,N_8413);
and U8766 (N_8766,N_8406,N_8457);
and U8767 (N_8767,N_8470,N_8598);
and U8768 (N_8768,N_8575,N_8412);
nand U8769 (N_8769,N_8449,N_8573);
nor U8770 (N_8770,N_8471,N_8534);
nor U8771 (N_8771,N_8493,N_8477);
nor U8772 (N_8772,N_8447,N_8575);
nand U8773 (N_8773,N_8590,N_8422);
xnor U8774 (N_8774,N_8459,N_8518);
nor U8775 (N_8775,N_8455,N_8585);
and U8776 (N_8776,N_8570,N_8595);
nor U8777 (N_8777,N_8478,N_8434);
nand U8778 (N_8778,N_8498,N_8503);
xor U8779 (N_8779,N_8586,N_8561);
nand U8780 (N_8780,N_8510,N_8574);
xor U8781 (N_8781,N_8412,N_8571);
nand U8782 (N_8782,N_8422,N_8544);
or U8783 (N_8783,N_8415,N_8459);
and U8784 (N_8784,N_8513,N_8583);
nor U8785 (N_8785,N_8422,N_8597);
nand U8786 (N_8786,N_8482,N_8556);
nor U8787 (N_8787,N_8545,N_8520);
nor U8788 (N_8788,N_8510,N_8443);
nand U8789 (N_8789,N_8519,N_8445);
nand U8790 (N_8790,N_8489,N_8554);
or U8791 (N_8791,N_8473,N_8566);
xor U8792 (N_8792,N_8543,N_8497);
nand U8793 (N_8793,N_8564,N_8407);
nand U8794 (N_8794,N_8560,N_8543);
nand U8795 (N_8795,N_8483,N_8518);
nor U8796 (N_8796,N_8567,N_8463);
nor U8797 (N_8797,N_8483,N_8407);
and U8798 (N_8798,N_8554,N_8508);
xnor U8799 (N_8799,N_8514,N_8474);
and U8800 (N_8800,N_8780,N_8727);
nand U8801 (N_8801,N_8729,N_8734);
or U8802 (N_8802,N_8708,N_8761);
nand U8803 (N_8803,N_8781,N_8688);
xnor U8804 (N_8804,N_8742,N_8655);
or U8805 (N_8805,N_8726,N_8782);
nor U8806 (N_8806,N_8722,N_8715);
or U8807 (N_8807,N_8653,N_8717);
nand U8808 (N_8808,N_8654,N_8793);
or U8809 (N_8809,N_8606,N_8643);
and U8810 (N_8810,N_8667,N_8757);
and U8811 (N_8811,N_8670,N_8640);
or U8812 (N_8812,N_8783,N_8773);
and U8813 (N_8813,N_8601,N_8701);
nor U8814 (N_8814,N_8768,N_8625);
or U8815 (N_8815,N_8650,N_8692);
or U8816 (N_8816,N_8745,N_8634);
and U8817 (N_8817,N_8718,N_8686);
nor U8818 (N_8818,N_8671,N_8621);
and U8819 (N_8819,N_8681,N_8623);
or U8820 (N_8820,N_8635,N_8751);
or U8821 (N_8821,N_8787,N_8679);
nor U8822 (N_8822,N_8744,N_8663);
nor U8823 (N_8823,N_8728,N_8784);
xor U8824 (N_8824,N_8767,N_8713);
and U8825 (N_8825,N_8719,N_8774);
nand U8826 (N_8826,N_8697,N_8611);
or U8827 (N_8827,N_8772,N_8645);
and U8828 (N_8828,N_8624,N_8705);
or U8829 (N_8829,N_8736,N_8788);
nor U8830 (N_8830,N_8602,N_8740);
or U8831 (N_8831,N_8677,N_8732);
or U8832 (N_8832,N_8615,N_8730);
xor U8833 (N_8833,N_8676,N_8723);
xnor U8834 (N_8834,N_8661,N_8797);
nor U8835 (N_8835,N_8646,N_8741);
xor U8836 (N_8836,N_8669,N_8603);
nand U8837 (N_8837,N_8648,N_8796);
xor U8838 (N_8838,N_8785,N_8725);
and U8839 (N_8839,N_8629,N_8694);
and U8840 (N_8840,N_8765,N_8613);
or U8841 (N_8841,N_8651,N_8746);
nor U8842 (N_8842,N_8610,N_8660);
xor U8843 (N_8843,N_8620,N_8658);
nand U8844 (N_8844,N_8747,N_8657);
nand U8845 (N_8845,N_8752,N_8743);
or U8846 (N_8846,N_8710,N_8798);
nand U8847 (N_8847,N_8627,N_8724);
nand U8848 (N_8848,N_8763,N_8619);
nor U8849 (N_8849,N_8790,N_8644);
nor U8850 (N_8850,N_8605,N_8604);
nor U8851 (N_8851,N_8673,N_8614);
nor U8852 (N_8852,N_8711,N_8685);
nor U8853 (N_8853,N_8699,N_8665);
and U8854 (N_8854,N_8687,N_8700);
or U8855 (N_8855,N_8759,N_8631);
nor U8856 (N_8856,N_8664,N_8617);
nor U8857 (N_8857,N_8612,N_8749);
or U8858 (N_8858,N_8758,N_8652);
and U8859 (N_8859,N_8760,N_8666);
and U8860 (N_8860,N_8756,N_8690);
nor U8861 (N_8861,N_8632,N_8794);
or U8862 (N_8862,N_8786,N_8739);
xnor U8863 (N_8863,N_8695,N_8778);
nand U8864 (N_8864,N_8639,N_8600);
nor U8865 (N_8865,N_8795,N_8714);
or U8866 (N_8866,N_8642,N_8616);
and U8867 (N_8867,N_8703,N_8704);
and U8868 (N_8868,N_8608,N_8647);
nand U8869 (N_8869,N_8707,N_8769);
and U8870 (N_8870,N_8637,N_8737);
nor U8871 (N_8871,N_8755,N_8641);
and U8872 (N_8872,N_8748,N_8712);
or U8873 (N_8873,N_8656,N_8789);
nand U8874 (N_8874,N_8630,N_8733);
nand U8875 (N_8875,N_8674,N_8696);
nor U8876 (N_8876,N_8678,N_8702);
xnor U8877 (N_8877,N_8609,N_8799);
or U8878 (N_8878,N_8633,N_8716);
or U8879 (N_8879,N_8779,N_8775);
or U8880 (N_8880,N_8698,N_8766);
nor U8881 (N_8881,N_8738,N_8776);
or U8882 (N_8882,N_8662,N_8680);
and U8883 (N_8883,N_8706,N_8649);
and U8884 (N_8884,N_8618,N_8675);
xor U8885 (N_8885,N_8735,N_8659);
nand U8886 (N_8886,N_8684,N_8791);
xor U8887 (N_8887,N_8622,N_8709);
xnor U8888 (N_8888,N_8626,N_8682);
and U8889 (N_8889,N_8754,N_8731);
nand U8890 (N_8890,N_8628,N_8672);
or U8891 (N_8891,N_8636,N_8770);
or U8892 (N_8892,N_8777,N_8683);
and U8893 (N_8893,N_8668,N_8689);
xnor U8894 (N_8894,N_8750,N_8638);
nor U8895 (N_8895,N_8693,N_8762);
nand U8896 (N_8896,N_8720,N_8721);
nor U8897 (N_8897,N_8753,N_8771);
xor U8898 (N_8898,N_8792,N_8607);
or U8899 (N_8899,N_8691,N_8764);
and U8900 (N_8900,N_8608,N_8744);
nand U8901 (N_8901,N_8752,N_8606);
xnor U8902 (N_8902,N_8620,N_8662);
or U8903 (N_8903,N_8673,N_8748);
or U8904 (N_8904,N_8664,N_8724);
or U8905 (N_8905,N_8720,N_8645);
and U8906 (N_8906,N_8679,N_8695);
nand U8907 (N_8907,N_8792,N_8615);
xnor U8908 (N_8908,N_8626,N_8662);
and U8909 (N_8909,N_8679,N_8707);
nand U8910 (N_8910,N_8656,N_8738);
or U8911 (N_8911,N_8677,N_8767);
or U8912 (N_8912,N_8639,N_8644);
and U8913 (N_8913,N_8605,N_8710);
xor U8914 (N_8914,N_8667,N_8685);
or U8915 (N_8915,N_8762,N_8691);
or U8916 (N_8916,N_8617,N_8624);
xor U8917 (N_8917,N_8642,N_8615);
nor U8918 (N_8918,N_8792,N_8777);
or U8919 (N_8919,N_8691,N_8694);
nor U8920 (N_8920,N_8786,N_8751);
nor U8921 (N_8921,N_8778,N_8652);
and U8922 (N_8922,N_8645,N_8678);
or U8923 (N_8923,N_8611,N_8715);
nand U8924 (N_8924,N_8630,N_8729);
and U8925 (N_8925,N_8656,N_8609);
xor U8926 (N_8926,N_8613,N_8657);
xor U8927 (N_8927,N_8709,N_8684);
nand U8928 (N_8928,N_8788,N_8628);
nor U8929 (N_8929,N_8745,N_8622);
xor U8930 (N_8930,N_8701,N_8695);
nor U8931 (N_8931,N_8723,N_8664);
nand U8932 (N_8932,N_8623,N_8665);
nand U8933 (N_8933,N_8617,N_8666);
xnor U8934 (N_8934,N_8722,N_8763);
and U8935 (N_8935,N_8635,N_8602);
or U8936 (N_8936,N_8701,N_8731);
xnor U8937 (N_8937,N_8680,N_8605);
xor U8938 (N_8938,N_8624,N_8686);
nand U8939 (N_8939,N_8645,N_8665);
xor U8940 (N_8940,N_8603,N_8743);
nand U8941 (N_8941,N_8786,N_8744);
nor U8942 (N_8942,N_8636,N_8600);
nor U8943 (N_8943,N_8712,N_8681);
nor U8944 (N_8944,N_8704,N_8622);
nand U8945 (N_8945,N_8776,N_8793);
xor U8946 (N_8946,N_8619,N_8674);
and U8947 (N_8947,N_8653,N_8618);
nor U8948 (N_8948,N_8659,N_8765);
and U8949 (N_8949,N_8749,N_8609);
nand U8950 (N_8950,N_8640,N_8797);
xnor U8951 (N_8951,N_8659,N_8632);
nand U8952 (N_8952,N_8610,N_8678);
nand U8953 (N_8953,N_8642,N_8766);
and U8954 (N_8954,N_8779,N_8610);
nor U8955 (N_8955,N_8793,N_8725);
and U8956 (N_8956,N_8729,N_8764);
or U8957 (N_8957,N_8696,N_8791);
or U8958 (N_8958,N_8613,N_8772);
and U8959 (N_8959,N_8718,N_8700);
and U8960 (N_8960,N_8733,N_8793);
or U8961 (N_8961,N_8765,N_8654);
nand U8962 (N_8962,N_8744,N_8645);
nand U8963 (N_8963,N_8727,N_8656);
or U8964 (N_8964,N_8795,N_8712);
nor U8965 (N_8965,N_8726,N_8610);
xor U8966 (N_8966,N_8641,N_8637);
and U8967 (N_8967,N_8754,N_8777);
or U8968 (N_8968,N_8634,N_8747);
nand U8969 (N_8969,N_8612,N_8622);
xnor U8970 (N_8970,N_8619,N_8658);
nand U8971 (N_8971,N_8661,N_8728);
nand U8972 (N_8972,N_8625,N_8761);
nor U8973 (N_8973,N_8619,N_8634);
and U8974 (N_8974,N_8710,N_8683);
or U8975 (N_8975,N_8762,N_8779);
and U8976 (N_8976,N_8756,N_8749);
nor U8977 (N_8977,N_8796,N_8698);
nand U8978 (N_8978,N_8797,N_8639);
or U8979 (N_8979,N_8778,N_8605);
xnor U8980 (N_8980,N_8649,N_8643);
xor U8981 (N_8981,N_8663,N_8743);
and U8982 (N_8982,N_8649,N_8707);
nor U8983 (N_8983,N_8662,N_8642);
and U8984 (N_8984,N_8623,N_8725);
and U8985 (N_8985,N_8685,N_8680);
xnor U8986 (N_8986,N_8734,N_8703);
or U8987 (N_8987,N_8633,N_8775);
or U8988 (N_8988,N_8602,N_8616);
nand U8989 (N_8989,N_8752,N_8782);
or U8990 (N_8990,N_8771,N_8670);
nand U8991 (N_8991,N_8655,N_8603);
nand U8992 (N_8992,N_8717,N_8686);
nor U8993 (N_8993,N_8745,N_8685);
xnor U8994 (N_8994,N_8745,N_8763);
xnor U8995 (N_8995,N_8752,N_8672);
and U8996 (N_8996,N_8778,N_8715);
or U8997 (N_8997,N_8767,N_8603);
nand U8998 (N_8998,N_8781,N_8637);
and U8999 (N_8999,N_8788,N_8672);
or U9000 (N_9000,N_8842,N_8910);
nor U9001 (N_9001,N_8813,N_8846);
or U9002 (N_9002,N_8825,N_8974);
and U9003 (N_9003,N_8890,N_8864);
nor U9004 (N_9004,N_8936,N_8957);
xnor U9005 (N_9005,N_8970,N_8990);
nor U9006 (N_9006,N_8838,N_8851);
xnor U9007 (N_9007,N_8853,N_8837);
nor U9008 (N_9008,N_8942,N_8963);
or U9009 (N_9009,N_8832,N_8988);
nand U9010 (N_9010,N_8860,N_8894);
and U9011 (N_9011,N_8997,N_8918);
and U9012 (N_9012,N_8952,N_8850);
nand U9013 (N_9013,N_8919,N_8872);
and U9014 (N_9014,N_8969,N_8950);
and U9015 (N_9015,N_8935,N_8960);
and U9016 (N_9016,N_8930,N_8839);
nand U9017 (N_9017,N_8912,N_8947);
and U9018 (N_9018,N_8873,N_8958);
nand U9019 (N_9019,N_8941,N_8923);
nor U9020 (N_9020,N_8827,N_8931);
nand U9021 (N_9021,N_8906,N_8845);
and U9022 (N_9022,N_8975,N_8849);
or U9023 (N_9023,N_8878,N_8835);
or U9024 (N_9024,N_8895,N_8892);
and U9025 (N_9025,N_8857,N_8980);
nor U9026 (N_9026,N_8877,N_8945);
xor U9027 (N_9027,N_8962,N_8946);
or U9028 (N_9028,N_8982,N_8949);
xnor U9029 (N_9029,N_8961,N_8831);
and U9030 (N_9030,N_8843,N_8991);
xor U9031 (N_9031,N_8834,N_8989);
nand U9032 (N_9032,N_8927,N_8866);
or U9033 (N_9033,N_8995,N_8828);
nor U9034 (N_9034,N_8998,N_8848);
nor U9035 (N_9035,N_8926,N_8818);
nor U9036 (N_9036,N_8869,N_8889);
and U9037 (N_9037,N_8829,N_8993);
nor U9038 (N_9038,N_8992,N_8983);
nand U9039 (N_9039,N_8925,N_8984);
xnor U9040 (N_9040,N_8943,N_8868);
and U9041 (N_9041,N_8977,N_8884);
nor U9042 (N_9042,N_8922,N_8804);
xor U9043 (N_9043,N_8819,N_8886);
xor U9044 (N_9044,N_8938,N_8921);
nor U9045 (N_9045,N_8844,N_8814);
or U9046 (N_9046,N_8913,N_8914);
or U9047 (N_9047,N_8966,N_8898);
and U9048 (N_9048,N_8917,N_8978);
nand U9049 (N_9049,N_8859,N_8862);
or U9050 (N_9050,N_8953,N_8883);
nor U9051 (N_9051,N_8816,N_8880);
xor U9052 (N_9052,N_8973,N_8901);
nor U9053 (N_9053,N_8903,N_8882);
or U9054 (N_9054,N_8905,N_8968);
or U9055 (N_9055,N_8879,N_8854);
nor U9056 (N_9056,N_8800,N_8897);
and U9057 (N_9057,N_8817,N_8824);
nand U9058 (N_9058,N_8944,N_8871);
xor U9059 (N_9059,N_8933,N_8826);
and U9060 (N_9060,N_8948,N_8801);
xor U9061 (N_9061,N_8833,N_8858);
or U9062 (N_9062,N_8909,N_8803);
nand U9063 (N_9063,N_8876,N_8855);
nor U9064 (N_9064,N_8881,N_8810);
nand U9065 (N_9065,N_8928,N_8867);
and U9066 (N_9066,N_8976,N_8870);
xnor U9067 (N_9067,N_8924,N_8929);
or U9068 (N_9068,N_8811,N_8994);
and U9069 (N_9069,N_8999,N_8856);
nor U9070 (N_9070,N_8891,N_8956);
xor U9071 (N_9071,N_8986,N_8887);
nand U9072 (N_9072,N_8954,N_8916);
nor U9073 (N_9073,N_8874,N_8805);
xnor U9074 (N_9074,N_8996,N_8852);
and U9075 (N_9075,N_8939,N_8981);
nor U9076 (N_9076,N_8979,N_8821);
xor U9077 (N_9077,N_8822,N_8967);
nand U9078 (N_9078,N_8830,N_8841);
xnor U9079 (N_9079,N_8840,N_8865);
and U9080 (N_9080,N_8985,N_8900);
or U9081 (N_9081,N_8806,N_8802);
or U9082 (N_9082,N_8847,N_8965);
xor U9083 (N_9083,N_8920,N_8888);
xor U9084 (N_9084,N_8955,N_8885);
and U9085 (N_9085,N_8907,N_8987);
nand U9086 (N_9086,N_8932,N_8899);
xor U9087 (N_9087,N_8908,N_8836);
nand U9088 (N_9088,N_8896,N_8861);
or U9089 (N_9089,N_8915,N_8934);
or U9090 (N_9090,N_8911,N_8808);
or U9091 (N_9091,N_8812,N_8904);
or U9092 (N_9092,N_8959,N_8893);
nand U9093 (N_9093,N_8815,N_8940);
nand U9094 (N_9094,N_8820,N_8964);
nand U9095 (N_9095,N_8951,N_8902);
nor U9096 (N_9096,N_8809,N_8971);
nor U9097 (N_9097,N_8972,N_8863);
nor U9098 (N_9098,N_8937,N_8875);
nor U9099 (N_9099,N_8807,N_8823);
or U9100 (N_9100,N_8907,N_8943);
or U9101 (N_9101,N_8896,N_8841);
or U9102 (N_9102,N_8849,N_8968);
nor U9103 (N_9103,N_8806,N_8849);
nor U9104 (N_9104,N_8835,N_8886);
and U9105 (N_9105,N_8864,N_8807);
nor U9106 (N_9106,N_8818,N_8990);
nor U9107 (N_9107,N_8975,N_8957);
nor U9108 (N_9108,N_8944,N_8905);
or U9109 (N_9109,N_8829,N_8866);
and U9110 (N_9110,N_8981,N_8851);
nand U9111 (N_9111,N_8913,N_8948);
xnor U9112 (N_9112,N_8937,N_8866);
or U9113 (N_9113,N_8825,N_8868);
and U9114 (N_9114,N_8936,N_8857);
nand U9115 (N_9115,N_8909,N_8843);
and U9116 (N_9116,N_8980,N_8806);
and U9117 (N_9117,N_8804,N_8898);
and U9118 (N_9118,N_8927,N_8983);
or U9119 (N_9119,N_8966,N_8971);
nand U9120 (N_9120,N_8950,N_8811);
or U9121 (N_9121,N_8876,N_8853);
nor U9122 (N_9122,N_8981,N_8985);
and U9123 (N_9123,N_8901,N_8839);
nor U9124 (N_9124,N_8902,N_8831);
xor U9125 (N_9125,N_8814,N_8859);
or U9126 (N_9126,N_8937,N_8929);
nand U9127 (N_9127,N_8893,N_8896);
nand U9128 (N_9128,N_8800,N_8931);
nor U9129 (N_9129,N_8896,N_8856);
and U9130 (N_9130,N_8966,N_8890);
nand U9131 (N_9131,N_8809,N_8965);
nor U9132 (N_9132,N_8934,N_8942);
nor U9133 (N_9133,N_8886,N_8992);
and U9134 (N_9134,N_8908,N_8942);
and U9135 (N_9135,N_8906,N_8990);
nand U9136 (N_9136,N_8966,N_8817);
xor U9137 (N_9137,N_8864,N_8926);
xor U9138 (N_9138,N_8985,N_8840);
and U9139 (N_9139,N_8856,N_8821);
and U9140 (N_9140,N_8975,N_8978);
xor U9141 (N_9141,N_8833,N_8937);
and U9142 (N_9142,N_8916,N_8891);
nand U9143 (N_9143,N_8932,N_8910);
xnor U9144 (N_9144,N_8821,N_8963);
xnor U9145 (N_9145,N_8983,N_8809);
nand U9146 (N_9146,N_8943,N_8935);
and U9147 (N_9147,N_8872,N_8848);
nor U9148 (N_9148,N_8824,N_8829);
nand U9149 (N_9149,N_8881,N_8910);
xnor U9150 (N_9150,N_8843,N_8860);
and U9151 (N_9151,N_8916,N_8922);
and U9152 (N_9152,N_8835,N_8980);
or U9153 (N_9153,N_8985,N_8980);
or U9154 (N_9154,N_8856,N_8914);
and U9155 (N_9155,N_8855,N_8896);
and U9156 (N_9156,N_8955,N_8847);
xor U9157 (N_9157,N_8804,N_8914);
and U9158 (N_9158,N_8935,N_8998);
or U9159 (N_9159,N_8898,N_8850);
xor U9160 (N_9160,N_8975,N_8966);
or U9161 (N_9161,N_8842,N_8926);
or U9162 (N_9162,N_8988,N_8952);
and U9163 (N_9163,N_8810,N_8804);
nand U9164 (N_9164,N_8969,N_8961);
or U9165 (N_9165,N_8872,N_8947);
nor U9166 (N_9166,N_8857,N_8899);
nor U9167 (N_9167,N_8886,N_8865);
nor U9168 (N_9168,N_8970,N_8800);
xnor U9169 (N_9169,N_8810,N_8901);
and U9170 (N_9170,N_8903,N_8935);
nand U9171 (N_9171,N_8856,N_8992);
xor U9172 (N_9172,N_8884,N_8946);
nand U9173 (N_9173,N_8862,N_8895);
nor U9174 (N_9174,N_8995,N_8980);
nand U9175 (N_9175,N_8809,N_8939);
nand U9176 (N_9176,N_8822,N_8821);
and U9177 (N_9177,N_8933,N_8902);
and U9178 (N_9178,N_8809,N_8859);
or U9179 (N_9179,N_8920,N_8832);
xor U9180 (N_9180,N_8923,N_8840);
nand U9181 (N_9181,N_8982,N_8871);
and U9182 (N_9182,N_8873,N_8820);
nor U9183 (N_9183,N_8847,N_8964);
and U9184 (N_9184,N_8913,N_8934);
and U9185 (N_9185,N_8891,N_8973);
xnor U9186 (N_9186,N_8882,N_8992);
nor U9187 (N_9187,N_8896,N_8913);
and U9188 (N_9188,N_8986,N_8867);
and U9189 (N_9189,N_8881,N_8993);
nand U9190 (N_9190,N_8805,N_8895);
xor U9191 (N_9191,N_8859,N_8954);
or U9192 (N_9192,N_8849,N_8967);
xor U9193 (N_9193,N_8870,N_8871);
xor U9194 (N_9194,N_8845,N_8847);
and U9195 (N_9195,N_8815,N_8893);
nand U9196 (N_9196,N_8810,N_8820);
xor U9197 (N_9197,N_8893,N_8805);
or U9198 (N_9198,N_8921,N_8997);
nand U9199 (N_9199,N_8847,N_8823);
nor U9200 (N_9200,N_9044,N_9139);
or U9201 (N_9201,N_9121,N_9064);
xnor U9202 (N_9202,N_9067,N_9039);
nand U9203 (N_9203,N_9007,N_9034);
or U9204 (N_9204,N_9119,N_9052);
and U9205 (N_9205,N_9094,N_9015);
nand U9206 (N_9206,N_9079,N_9153);
xnor U9207 (N_9207,N_9161,N_9159);
and U9208 (N_9208,N_9131,N_9125);
nand U9209 (N_9209,N_9018,N_9118);
xor U9210 (N_9210,N_9177,N_9113);
nand U9211 (N_9211,N_9077,N_9008);
or U9212 (N_9212,N_9162,N_9041);
nand U9213 (N_9213,N_9195,N_9104);
nand U9214 (N_9214,N_9089,N_9100);
nor U9215 (N_9215,N_9108,N_9149);
and U9216 (N_9216,N_9133,N_9076);
or U9217 (N_9217,N_9009,N_9132);
and U9218 (N_9218,N_9087,N_9170);
nand U9219 (N_9219,N_9166,N_9112);
and U9220 (N_9220,N_9182,N_9151);
nor U9221 (N_9221,N_9168,N_9055);
xor U9222 (N_9222,N_9152,N_9114);
and U9223 (N_9223,N_9107,N_9126);
nor U9224 (N_9224,N_9096,N_9117);
nand U9225 (N_9225,N_9124,N_9024);
or U9226 (N_9226,N_9173,N_9140);
nand U9227 (N_9227,N_9156,N_9084);
xor U9228 (N_9228,N_9020,N_9190);
nand U9229 (N_9229,N_9122,N_9172);
or U9230 (N_9230,N_9105,N_9081);
nand U9231 (N_9231,N_9144,N_9061);
nor U9232 (N_9232,N_9127,N_9062);
and U9233 (N_9233,N_9187,N_9048);
nand U9234 (N_9234,N_9155,N_9176);
nor U9235 (N_9235,N_9196,N_9142);
or U9236 (N_9236,N_9082,N_9188);
nor U9237 (N_9237,N_9134,N_9160);
nand U9238 (N_9238,N_9088,N_9111);
nor U9239 (N_9239,N_9185,N_9000);
nand U9240 (N_9240,N_9057,N_9179);
and U9241 (N_9241,N_9045,N_9189);
and U9242 (N_9242,N_9085,N_9198);
and U9243 (N_9243,N_9005,N_9030);
xor U9244 (N_9244,N_9136,N_9080);
or U9245 (N_9245,N_9091,N_9137);
xor U9246 (N_9246,N_9028,N_9116);
xnor U9247 (N_9247,N_9042,N_9138);
nand U9248 (N_9248,N_9167,N_9106);
nand U9249 (N_9249,N_9099,N_9004);
xor U9250 (N_9250,N_9180,N_9003);
or U9251 (N_9251,N_9016,N_9092);
xor U9252 (N_9252,N_9135,N_9154);
or U9253 (N_9253,N_9035,N_9019);
and U9254 (N_9254,N_9191,N_9147);
nor U9255 (N_9255,N_9072,N_9075);
nand U9256 (N_9256,N_9199,N_9037);
or U9257 (N_9257,N_9120,N_9186);
xnor U9258 (N_9258,N_9184,N_9097);
and U9259 (N_9259,N_9036,N_9054);
and U9260 (N_9260,N_9164,N_9183);
and U9261 (N_9261,N_9059,N_9025);
and U9262 (N_9262,N_9049,N_9123);
nand U9263 (N_9263,N_9078,N_9073);
and U9264 (N_9264,N_9101,N_9023);
nand U9265 (N_9265,N_9090,N_9065);
xor U9266 (N_9266,N_9157,N_9102);
nor U9267 (N_9267,N_9141,N_9051);
and U9268 (N_9268,N_9074,N_9006);
and U9269 (N_9269,N_9109,N_9027);
xor U9270 (N_9270,N_9001,N_9014);
nor U9271 (N_9271,N_9022,N_9069);
nor U9272 (N_9272,N_9031,N_9150);
and U9273 (N_9273,N_9086,N_9129);
xnor U9274 (N_9274,N_9130,N_9098);
xor U9275 (N_9275,N_9046,N_9197);
nand U9276 (N_9276,N_9128,N_9012);
nor U9277 (N_9277,N_9192,N_9146);
xnor U9278 (N_9278,N_9169,N_9175);
and U9279 (N_9279,N_9010,N_9013);
nand U9280 (N_9280,N_9017,N_9071);
nand U9281 (N_9281,N_9068,N_9083);
xor U9282 (N_9282,N_9002,N_9056);
or U9283 (N_9283,N_9032,N_9115);
xnor U9284 (N_9284,N_9058,N_9011);
and U9285 (N_9285,N_9171,N_9066);
xnor U9286 (N_9286,N_9193,N_9174);
nor U9287 (N_9287,N_9143,N_9043);
or U9288 (N_9288,N_9095,N_9033);
nand U9289 (N_9289,N_9070,N_9040);
xnor U9290 (N_9290,N_9060,N_9178);
nor U9291 (N_9291,N_9158,N_9110);
xor U9292 (N_9292,N_9021,N_9063);
xnor U9293 (N_9293,N_9165,N_9038);
nor U9294 (N_9294,N_9050,N_9047);
xnor U9295 (N_9295,N_9103,N_9181);
nor U9296 (N_9296,N_9145,N_9026);
or U9297 (N_9297,N_9053,N_9163);
nor U9298 (N_9298,N_9194,N_9029);
and U9299 (N_9299,N_9148,N_9093);
nor U9300 (N_9300,N_9166,N_9007);
nand U9301 (N_9301,N_9030,N_9008);
nor U9302 (N_9302,N_9068,N_9161);
and U9303 (N_9303,N_9175,N_9168);
nand U9304 (N_9304,N_9181,N_9198);
xnor U9305 (N_9305,N_9125,N_9001);
xnor U9306 (N_9306,N_9161,N_9133);
or U9307 (N_9307,N_9138,N_9125);
nand U9308 (N_9308,N_9066,N_9108);
nand U9309 (N_9309,N_9141,N_9014);
nand U9310 (N_9310,N_9034,N_9073);
nand U9311 (N_9311,N_9015,N_9067);
nand U9312 (N_9312,N_9068,N_9037);
or U9313 (N_9313,N_9122,N_9113);
or U9314 (N_9314,N_9003,N_9073);
or U9315 (N_9315,N_9151,N_9152);
and U9316 (N_9316,N_9111,N_9142);
and U9317 (N_9317,N_9192,N_9141);
and U9318 (N_9318,N_9159,N_9187);
and U9319 (N_9319,N_9081,N_9093);
nor U9320 (N_9320,N_9194,N_9124);
or U9321 (N_9321,N_9140,N_9101);
and U9322 (N_9322,N_9191,N_9056);
nor U9323 (N_9323,N_9157,N_9131);
or U9324 (N_9324,N_9112,N_9034);
nand U9325 (N_9325,N_9107,N_9102);
and U9326 (N_9326,N_9185,N_9127);
nor U9327 (N_9327,N_9187,N_9178);
nand U9328 (N_9328,N_9002,N_9053);
xor U9329 (N_9329,N_9030,N_9161);
and U9330 (N_9330,N_9134,N_9162);
nand U9331 (N_9331,N_9186,N_9020);
nor U9332 (N_9332,N_9197,N_9067);
nand U9333 (N_9333,N_9024,N_9093);
or U9334 (N_9334,N_9032,N_9191);
or U9335 (N_9335,N_9091,N_9022);
or U9336 (N_9336,N_9052,N_9063);
nand U9337 (N_9337,N_9189,N_9033);
nor U9338 (N_9338,N_9135,N_9124);
nor U9339 (N_9339,N_9019,N_9054);
xor U9340 (N_9340,N_9092,N_9122);
or U9341 (N_9341,N_9160,N_9150);
nand U9342 (N_9342,N_9080,N_9071);
xnor U9343 (N_9343,N_9021,N_9024);
nor U9344 (N_9344,N_9151,N_9125);
or U9345 (N_9345,N_9120,N_9082);
xnor U9346 (N_9346,N_9059,N_9017);
nor U9347 (N_9347,N_9057,N_9199);
nor U9348 (N_9348,N_9035,N_9121);
nor U9349 (N_9349,N_9024,N_9188);
nor U9350 (N_9350,N_9104,N_9188);
xnor U9351 (N_9351,N_9077,N_9070);
nor U9352 (N_9352,N_9035,N_9054);
xor U9353 (N_9353,N_9005,N_9110);
nand U9354 (N_9354,N_9133,N_9084);
nand U9355 (N_9355,N_9049,N_9104);
xnor U9356 (N_9356,N_9199,N_9035);
and U9357 (N_9357,N_9113,N_9183);
or U9358 (N_9358,N_9121,N_9014);
xor U9359 (N_9359,N_9044,N_9127);
nor U9360 (N_9360,N_9003,N_9115);
xor U9361 (N_9361,N_9053,N_9081);
nand U9362 (N_9362,N_9047,N_9178);
or U9363 (N_9363,N_9002,N_9106);
or U9364 (N_9364,N_9114,N_9079);
nor U9365 (N_9365,N_9017,N_9193);
xnor U9366 (N_9366,N_9048,N_9063);
or U9367 (N_9367,N_9188,N_9071);
and U9368 (N_9368,N_9126,N_9186);
and U9369 (N_9369,N_9004,N_9137);
or U9370 (N_9370,N_9000,N_9079);
nor U9371 (N_9371,N_9049,N_9103);
or U9372 (N_9372,N_9001,N_9162);
nor U9373 (N_9373,N_9028,N_9177);
and U9374 (N_9374,N_9175,N_9115);
nor U9375 (N_9375,N_9141,N_9065);
or U9376 (N_9376,N_9082,N_9083);
and U9377 (N_9377,N_9091,N_9101);
or U9378 (N_9378,N_9001,N_9106);
xnor U9379 (N_9379,N_9172,N_9062);
or U9380 (N_9380,N_9191,N_9027);
and U9381 (N_9381,N_9102,N_9148);
nor U9382 (N_9382,N_9057,N_9189);
or U9383 (N_9383,N_9177,N_9148);
nor U9384 (N_9384,N_9163,N_9198);
nand U9385 (N_9385,N_9132,N_9139);
nand U9386 (N_9386,N_9105,N_9018);
nand U9387 (N_9387,N_9158,N_9026);
nor U9388 (N_9388,N_9050,N_9121);
nor U9389 (N_9389,N_9106,N_9081);
and U9390 (N_9390,N_9070,N_9060);
nor U9391 (N_9391,N_9091,N_9159);
nand U9392 (N_9392,N_9161,N_9083);
xor U9393 (N_9393,N_9120,N_9123);
xnor U9394 (N_9394,N_9183,N_9042);
xnor U9395 (N_9395,N_9106,N_9099);
nand U9396 (N_9396,N_9112,N_9095);
nand U9397 (N_9397,N_9116,N_9077);
nand U9398 (N_9398,N_9013,N_9015);
xnor U9399 (N_9399,N_9164,N_9028);
and U9400 (N_9400,N_9310,N_9215);
or U9401 (N_9401,N_9299,N_9226);
nor U9402 (N_9402,N_9268,N_9317);
nor U9403 (N_9403,N_9375,N_9331);
xnor U9404 (N_9404,N_9386,N_9260);
nor U9405 (N_9405,N_9265,N_9239);
nor U9406 (N_9406,N_9258,N_9291);
nand U9407 (N_9407,N_9303,N_9343);
nor U9408 (N_9408,N_9253,N_9286);
and U9409 (N_9409,N_9398,N_9349);
nor U9410 (N_9410,N_9217,N_9372);
xnor U9411 (N_9411,N_9245,N_9231);
nor U9412 (N_9412,N_9344,N_9249);
and U9413 (N_9413,N_9298,N_9233);
nand U9414 (N_9414,N_9353,N_9238);
or U9415 (N_9415,N_9305,N_9315);
nand U9416 (N_9416,N_9211,N_9352);
nand U9417 (N_9417,N_9208,N_9246);
xor U9418 (N_9418,N_9325,N_9380);
nor U9419 (N_9419,N_9210,N_9393);
xor U9420 (N_9420,N_9250,N_9314);
nor U9421 (N_9421,N_9385,N_9356);
or U9422 (N_9422,N_9369,N_9327);
and U9423 (N_9423,N_9259,N_9228);
nand U9424 (N_9424,N_9261,N_9201);
and U9425 (N_9425,N_9323,N_9360);
or U9426 (N_9426,N_9256,N_9373);
xor U9427 (N_9427,N_9363,N_9362);
nand U9428 (N_9428,N_9220,N_9374);
xor U9429 (N_9429,N_9326,N_9371);
nor U9430 (N_9430,N_9296,N_9392);
or U9431 (N_9431,N_9350,N_9288);
xnor U9432 (N_9432,N_9236,N_9244);
nor U9433 (N_9433,N_9294,N_9359);
and U9434 (N_9434,N_9219,N_9287);
nor U9435 (N_9435,N_9252,N_9394);
nor U9436 (N_9436,N_9355,N_9284);
and U9437 (N_9437,N_9365,N_9309);
or U9438 (N_9438,N_9387,N_9263);
nand U9439 (N_9439,N_9395,N_9379);
nand U9440 (N_9440,N_9312,N_9273);
nand U9441 (N_9441,N_9235,N_9329);
nor U9442 (N_9442,N_9311,N_9336);
nor U9443 (N_9443,N_9358,N_9318);
xor U9444 (N_9444,N_9262,N_9376);
or U9445 (N_9445,N_9242,N_9357);
nand U9446 (N_9446,N_9307,N_9274);
and U9447 (N_9447,N_9330,N_9378);
or U9448 (N_9448,N_9351,N_9308);
nor U9449 (N_9449,N_9266,N_9254);
nor U9450 (N_9450,N_9290,N_9206);
nand U9451 (N_9451,N_9205,N_9204);
and U9452 (N_9452,N_9324,N_9396);
or U9453 (N_9453,N_9342,N_9289);
or U9454 (N_9454,N_9335,N_9279);
xor U9455 (N_9455,N_9281,N_9280);
or U9456 (N_9456,N_9292,N_9370);
nand U9457 (N_9457,N_9399,N_9270);
and U9458 (N_9458,N_9214,N_9213);
nand U9459 (N_9459,N_9295,N_9221);
nand U9460 (N_9460,N_9302,N_9383);
nor U9461 (N_9461,N_9332,N_9237);
xnor U9462 (N_9462,N_9267,N_9255);
xor U9463 (N_9463,N_9277,N_9382);
or U9464 (N_9464,N_9320,N_9367);
nor U9465 (N_9465,N_9346,N_9234);
or U9466 (N_9466,N_9271,N_9269);
nor U9467 (N_9467,N_9203,N_9202);
nand U9468 (N_9468,N_9248,N_9240);
nor U9469 (N_9469,N_9209,N_9278);
nand U9470 (N_9470,N_9200,N_9364);
nand U9471 (N_9471,N_9377,N_9306);
xnor U9472 (N_9472,N_9264,N_9276);
and U9473 (N_9473,N_9300,N_9339);
nand U9474 (N_9474,N_9338,N_9225);
or U9475 (N_9475,N_9247,N_9272);
nand U9476 (N_9476,N_9229,N_9297);
or U9477 (N_9477,N_9354,N_9316);
nand U9478 (N_9478,N_9293,N_9334);
xnor U9479 (N_9479,N_9361,N_9384);
or U9480 (N_9480,N_9207,N_9251);
nor U9481 (N_9481,N_9345,N_9223);
and U9482 (N_9482,N_9322,N_9224);
nor U9483 (N_9483,N_9241,N_9366);
or U9484 (N_9484,N_9218,N_9341);
xor U9485 (N_9485,N_9243,N_9347);
and U9486 (N_9486,N_9222,N_9319);
nor U9487 (N_9487,N_9388,N_9313);
and U9488 (N_9488,N_9390,N_9232);
and U9489 (N_9489,N_9301,N_9348);
nor U9490 (N_9490,N_9391,N_9257);
xnor U9491 (N_9491,N_9368,N_9285);
nand U9492 (N_9492,N_9397,N_9230);
nand U9493 (N_9493,N_9283,N_9321);
nand U9494 (N_9494,N_9340,N_9337);
or U9495 (N_9495,N_9212,N_9282);
xnor U9496 (N_9496,N_9216,N_9227);
xnor U9497 (N_9497,N_9275,N_9333);
xor U9498 (N_9498,N_9381,N_9389);
nand U9499 (N_9499,N_9304,N_9328);
nand U9500 (N_9500,N_9262,N_9282);
or U9501 (N_9501,N_9367,N_9338);
and U9502 (N_9502,N_9390,N_9271);
nand U9503 (N_9503,N_9270,N_9284);
nor U9504 (N_9504,N_9382,N_9280);
and U9505 (N_9505,N_9214,N_9271);
xor U9506 (N_9506,N_9230,N_9270);
xor U9507 (N_9507,N_9237,N_9372);
nand U9508 (N_9508,N_9336,N_9348);
and U9509 (N_9509,N_9286,N_9292);
nand U9510 (N_9510,N_9342,N_9393);
or U9511 (N_9511,N_9284,N_9318);
or U9512 (N_9512,N_9321,N_9287);
or U9513 (N_9513,N_9361,N_9260);
and U9514 (N_9514,N_9223,N_9210);
nor U9515 (N_9515,N_9256,N_9325);
or U9516 (N_9516,N_9257,N_9237);
and U9517 (N_9517,N_9326,N_9316);
xor U9518 (N_9518,N_9367,N_9285);
nand U9519 (N_9519,N_9208,N_9325);
nand U9520 (N_9520,N_9332,N_9323);
xor U9521 (N_9521,N_9397,N_9209);
nand U9522 (N_9522,N_9203,N_9346);
xor U9523 (N_9523,N_9397,N_9239);
xnor U9524 (N_9524,N_9230,N_9399);
nand U9525 (N_9525,N_9270,N_9382);
and U9526 (N_9526,N_9276,N_9229);
nand U9527 (N_9527,N_9334,N_9391);
nand U9528 (N_9528,N_9215,N_9340);
or U9529 (N_9529,N_9296,N_9286);
nand U9530 (N_9530,N_9261,N_9217);
nand U9531 (N_9531,N_9331,N_9376);
nand U9532 (N_9532,N_9373,N_9240);
or U9533 (N_9533,N_9332,N_9325);
xnor U9534 (N_9534,N_9303,N_9322);
xnor U9535 (N_9535,N_9248,N_9327);
xnor U9536 (N_9536,N_9364,N_9310);
xor U9537 (N_9537,N_9347,N_9321);
nor U9538 (N_9538,N_9373,N_9227);
and U9539 (N_9539,N_9289,N_9201);
xnor U9540 (N_9540,N_9268,N_9271);
nand U9541 (N_9541,N_9271,N_9316);
and U9542 (N_9542,N_9338,N_9340);
and U9543 (N_9543,N_9373,N_9272);
xor U9544 (N_9544,N_9233,N_9289);
or U9545 (N_9545,N_9234,N_9331);
and U9546 (N_9546,N_9386,N_9394);
xnor U9547 (N_9547,N_9275,N_9392);
nor U9548 (N_9548,N_9229,N_9355);
and U9549 (N_9549,N_9289,N_9348);
nor U9550 (N_9550,N_9356,N_9351);
nor U9551 (N_9551,N_9320,N_9256);
and U9552 (N_9552,N_9303,N_9358);
or U9553 (N_9553,N_9313,N_9216);
xor U9554 (N_9554,N_9221,N_9323);
nor U9555 (N_9555,N_9264,N_9387);
nand U9556 (N_9556,N_9366,N_9330);
and U9557 (N_9557,N_9386,N_9326);
xor U9558 (N_9558,N_9315,N_9261);
nor U9559 (N_9559,N_9335,N_9342);
or U9560 (N_9560,N_9328,N_9279);
nor U9561 (N_9561,N_9243,N_9278);
or U9562 (N_9562,N_9299,N_9242);
nand U9563 (N_9563,N_9233,N_9256);
or U9564 (N_9564,N_9304,N_9367);
nor U9565 (N_9565,N_9395,N_9334);
nor U9566 (N_9566,N_9252,N_9297);
nand U9567 (N_9567,N_9316,N_9280);
nand U9568 (N_9568,N_9272,N_9269);
nand U9569 (N_9569,N_9246,N_9278);
or U9570 (N_9570,N_9298,N_9251);
nor U9571 (N_9571,N_9234,N_9397);
and U9572 (N_9572,N_9389,N_9221);
xor U9573 (N_9573,N_9329,N_9228);
nor U9574 (N_9574,N_9345,N_9255);
nor U9575 (N_9575,N_9273,N_9201);
or U9576 (N_9576,N_9266,N_9297);
nand U9577 (N_9577,N_9366,N_9285);
nor U9578 (N_9578,N_9292,N_9296);
or U9579 (N_9579,N_9271,N_9356);
and U9580 (N_9580,N_9217,N_9342);
or U9581 (N_9581,N_9385,N_9309);
and U9582 (N_9582,N_9204,N_9352);
xnor U9583 (N_9583,N_9354,N_9257);
and U9584 (N_9584,N_9313,N_9324);
nand U9585 (N_9585,N_9395,N_9290);
xnor U9586 (N_9586,N_9279,N_9341);
and U9587 (N_9587,N_9338,N_9351);
and U9588 (N_9588,N_9219,N_9220);
or U9589 (N_9589,N_9388,N_9392);
xnor U9590 (N_9590,N_9207,N_9213);
and U9591 (N_9591,N_9227,N_9364);
and U9592 (N_9592,N_9223,N_9384);
nor U9593 (N_9593,N_9248,N_9323);
nor U9594 (N_9594,N_9214,N_9332);
or U9595 (N_9595,N_9227,N_9384);
or U9596 (N_9596,N_9305,N_9222);
nand U9597 (N_9597,N_9297,N_9347);
or U9598 (N_9598,N_9364,N_9289);
nor U9599 (N_9599,N_9217,N_9237);
and U9600 (N_9600,N_9471,N_9552);
and U9601 (N_9601,N_9554,N_9546);
and U9602 (N_9602,N_9480,N_9509);
or U9603 (N_9603,N_9523,N_9524);
nand U9604 (N_9604,N_9521,N_9559);
nand U9605 (N_9605,N_9528,N_9578);
xnor U9606 (N_9606,N_9537,N_9597);
or U9607 (N_9607,N_9527,N_9446);
and U9608 (N_9608,N_9539,N_9491);
or U9609 (N_9609,N_9584,N_9500);
nand U9610 (N_9610,N_9447,N_9529);
nor U9611 (N_9611,N_9404,N_9416);
or U9612 (N_9612,N_9568,N_9443);
xnor U9613 (N_9613,N_9533,N_9587);
or U9614 (N_9614,N_9534,N_9430);
nand U9615 (N_9615,N_9427,N_9538);
xor U9616 (N_9616,N_9501,N_9588);
and U9617 (N_9617,N_9519,N_9576);
xnor U9618 (N_9618,N_9580,N_9425);
xor U9619 (N_9619,N_9531,N_9567);
and U9620 (N_9620,N_9417,N_9437);
xnor U9621 (N_9621,N_9517,N_9545);
xnor U9622 (N_9622,N_9406,N_9401);
nor U9623 (N_9623,N_9467,N_9595);
and U9624 (N_9624,N_9540,N_9449);
nor U9625 (N_9625,N_9423,N_9564);
and U9626 (N_9626,N_9455,N_9553);
xnor U9627 (N_9627,N_9503,N_9507);
and U9628 (N_9628,N_9478,N_9452);
nor U9629 (N_9629,N_9535,N_9543);
xor U9630 (N_9630,N_9571,N_9436);
nand U9631 (N_9631,N_9432,N_9558);
or U9632 (N_9632,N_9515,N_9496);
or U9633 (N_9633,N_9561,N_9458);
nor U9634 (N_9634,N_9569,N_9573);
xor U9635 (N_9635,N_9518,N_9591);
nor U9636 (N_9636,N_9488,N_9439);
or U9637 (N_9637,N_9441,N_9494);
and U9638 (N_9638,N_9555,N_9566);
nand U9639 (N_9639,N_9419,N_9596);
or U9640 (N_9640,N_9482,N_9589);
and U9641 (N_9641,N_9409,N_9477);
nand U9642 (N_9642,N_9570,N_9565);
nor U9643 (N_9643,N_9444,N_9408);
or U9644 (N_9644,N_9465,N_9481);
and U9645 (N_9645,N_9457,N_9572);
xnor U9646 (N_9646,N_9547,N_9505);
nor U9647 (N_9647,N_9487,N_9504);
or U9648 (N_9648,N_9495,N_9476);
nor U9649 (N_9649,N_9426,N_9562);
and U9650 (N_9650,N_9557,N_9499);
or U9651 (N_9651,N_9563,N_9442);
and U9652 (N_9652,N_9464,N_9440);
nand U9653 (N_9653,N_9418,N_9410);
or U9654 (N_9654,N_9431,N_9593);
nand U9655 (N_9655,N_9462,N_9474);
nand U9656 (N_9656,N_9450,N_9469);
nor U9657 (N_9657,N_9549,N_9590);
or U9658 (N_9658,N_9498,N_9516);
nor U9659 (N_9659,N_9403,N_9502);
nor U9660 (N_9660,N_9550,N_9424);
xnor U9661 (N_9661,N_9448,N_9400);
nand U9662 (N_9662,N_9506,N_9433);
nand U9663 (N_9663,N_9598,N_9434);
nand U9664 (N_9664,N_9575,N_9479);
xor U9665 (N_9665,N_9421,N_9411);
and U9666 (N_9666,N_9536,N_9560);
nand U9667 (N_9667,N_9599,N_9513);
or U9668 (N_9668,N_9508,N_9414);
nand U9669 (N_9669,N_9520,N_9454);
nand U9670 (N_9670,N_9473,N_9582);
and U9671 (N_9671,N_9493,N_9405);
nand U9672 (N_9672,N_9428,N_9420);
and U9673 (N_9673,N_9463,N_9407);
or U9674 (N_9674,N_9510,N_9461);
and U9675 (N_9675,N_9435,N_9592);
or U9676 (N_9676,N_9514,N_9451);
nor U9677 (N_9677,N_9551,N_9415);
nor U9678 (N_9678,N_9438,N_9453);
or U9679 (N_9679,N_9475,N_9460);
nor U9680 (N_9680,N_9459,N_9492);
xor U9681 (N_9681,N_9489,N_9429);
and U9682 (N_9682,N_9544,N_9472);
nor U9683 (N_9683,N_9556,N_9594);
nand U9684 (N_9684,N_9586,N_9490);
and U9685 (N_9685,N_9583,N_9530);
xor U9686 (N_9686,N_9577,N_9402);
and U9687 (N_9687,N_9522,N_9413);
nand U9688 (N_9688,N_9585,N_9466);
or U9689 (N_9689,N_9486,N_9581);
and U9690 (N_9690,N_9548,N_9542);
xor U9691 (N_9691,N_9470,N_9468);
nand U9692 (N_9692,N_9511,N_9412);
or U9693 (N_9693,N_9483,N_9532);
nor U9694 (N_9694,N_9512,N_9456);
xnor U9695 (N_9695,N_9579,N_9525);
nand U9696 (N_9696,N_9445,N_9497);
xnor U9697 (N_9697,N_9485,N_9422);
nand U9698 (N_9698,N_9574,N_9484);
xor U9699 (N_9699,N_9526,N_9541);
nor U9700 (N_9700,N_9501,N_9447);
and U9701 (N_9701,N_9560,N_9576);
nor U9702 (N_9702,N_9427,N_9559);
nand U9703 (N_9703,N_9582,N_9597);
nand U9704 (N_9704,N_9484,N_9481);
and U9705 (N_9705,N_9571,N_9599);
nor U9706 (N_9706,N_9596,N_9577);
xor U9707 (N_9707,N_9526,N_9497);
nor U9708 (N_9708,N_9564,N_9464);
or U9709 (N_9709,N_9428,N_9472);
nand U9710 (N_9710,N_9544,N_9535);
or U9711 (N_9711,N_9597,N_9420);
nand U9712 (N_9712,N_9505,N_9432);
nand U9713 (N_9713,N_9526,N_9594);
nor U9714 (N_9714,N_9580,N_9504);
and U9715 (N_9715,N_9424,N_9512);
nand U9716 (N_9716,N_9545,N_9570);
xor U9717 (N_9717,N_9527,N_9537);
xnor U9718 (N_9718,N_9494,N_9589);
and U9719 (N_9719,N_9526,N_9459);
or U9720 (N_9720,N_9508,N_9567);
nor U9721 (N_9721,N_9480,N_9428);
nor U9722 (N_9722,N_9564,N_9443);
nor U9723 (N_9723,N_9439,N_9502);
or U9724 (N_9724,N_9508,N_9595);
nor U9725 (N_9725,N_9413,N_9546);
xnor U9726 (N_9726,N_9406,N_9462);
nor U9727 (N_9727,N_9562,N_9450);
and U9728 (N_9728,N_9562,N_9478);
nor U9729 (N_9729,N_9487,N_9451);
nand U9730 (N_9730,N_9588,N_9589);
nor U9731 (N_9731,N_9577,N_9543);
and U9732 (N_9732,N_9453,N_9599);
or U9733 (N_9733,N_9540,N_9545);
nor U9734 (N_9734,N_9532,N_9434);
or U9735 (N_9735,N_9543,N_9454);
nand U9736 (N_9736,N_9420,N_9509);
nand U9737 (N_9737,N_9490,N_9454);
nand U9738 (N_9738,N_9549,N_9524);
nor U9739 (N_9739,N_9586,N_9465);
nor U9740 (N_9740,N_9556,N_9546);
or U9741 (N_9741,N_9486,N_9449);
and U9742 (N_9742,N_9418,N_9477);
and U9743 (N_9743,N_9581,N_9460);
xnor U9744 (N_9744,N_9407,N_9441);
or U9745 (N_9745,N_9415,N_9561);
xnor U9746 (N_9746,N_9538,N_9507);
and U9747 (N_9747,N_9475,N_9428);
nand U9748 (N_9748,N_9564,N_9433);
and U9749 (N_9749,N_9513,N_9454);
and U9750 (N_9750,N_9483,N_9432);
nand U9751 (N_9751,N_9402,N_9411);
xor U9752 (N_9752,N_9480,N_9510);
nand U9753 (N_9753,N_9528,N_9569);
nand U9754 (N_9754,N_9484,N_9467);
xor U9755 (N_9755,N_9517,N_9422);
or U9756 (N_9756,N_9485,N_9426);
or U9757 (N_9757,N_9457,N_9470);
or U9758 (N_9758,N_9592,N_9554);
nand U9759 (N_9759,N_9592,N_9452);
or U9760 (N_9760,N_9563,N_9586);
or U9761 (N_9761,N_9548,N_9579);
xnor U9762 (N_9762,N_9461,N_9580);
xnor U9763 (N_9763,N_9589,N_9509);
xnor U9764 (N_9764,N_9474,N_9451);
and U9765 (N_9765,N_9451,N_9507);
nor U9766 (N_9766,N_9552,N_9495);
xor U9767 (N_9767,N_9421,N_9452);
xnor U9768 (N_9768,N_9411,N_9581);
and U9769 (N_9769,N_9528,N_9476);
or U9770 (N_9770,N_9508,N_9421);
nor U9771 (N_9771,N_9536,N_9444);
nor U9772 (N_9772,N_9548,N_9504);
nor U9773 (N_9773,N_9592,N_9539);
nand U9774 (N_9774,N_9506,N_9420);
xnor U9775 (N_9775,N_9414,N_9481);
xnor U9776 (N_9776,N_9570,N_9497);
xor U9777 (N_9777,N_9447,N_9584);
nor U9778 (N_9778,N_9583,N_9536);
xor U9779 (N_9779,N_9472,N_9416);
or U9780 (N_9780,N_9571,N_9574);
or U9781 (N_9781,N_9489,N_9482);
and U9782 (N_9782,N_9501,N_9436);
and U9783 (N_9783,N_9509,N_9545);
nand U9784 (N_9784,N_9550,N_9502);
nand U9785 (N_9785,N_9467,N_9413);
or U9786 (N_9786,N_9575,N_9436);
nor U9787 (N_9787,N_9429,N_9515);
and U9788 (N_9788,N_9495,N_9402);
xor U9789 (N_9789,N_9495,N_9575);
nand U9790 (N_9790,N_9586,N_9413);
or U9791 (N_9791,N_9506,N_9479);
nor U9792 (N_9792,N_9570,N_9580);
nor U9793 (N_9793,N_9435,N_9569);
and U9794 (N_9794,N_9431,N_9507);
nor U9795 (N_9795,N_9470,N_9456);
and U9796 (N_9796,N_9531,N_9404);
nand U9797 (N_9797,N_9596,N_9439);
xnor U9798 (N_9798,N_9523,N_9597);
nand U9799 (N_9799,N_9504,N_9458);
nand U9800 (N_9800,N_9658,N_9674);
nor U9801 (N_9801,N_9734,N_9661);
and U9802 (N_9802,N_9640,N_9739);
xnor U9803 (N_9803,N_9796,N_9719);
xor U9804 (N_9804,N_9659,N_9604);
nor U9805 (N_9805,N_9682,N_9688);
xnor U9806 (N_9806,N_9632,N_9681);
xor U9807 (N_9807,N_9652,N_9744);
nor U9808 (N_9808,N_9678,N_9643);
xnor U9809 (N_9809,N_9720,N_9731);
and U9810 (N_9810,N_9639,N_9730);
xor U9811 (N_9811,N_9711,N_9685);
nand U9812 (N_9812,N_9627,N_9779);
nand U9813 (N_9813,N_9713,N_9783);
or U9814 (N_9814,N_9668,N_9715);
nand U9815 (N_9815,N_9707,N_9697);
nand U9816 (N_9816,N_9614,N_9723);
or U9817 (N_9817,N_9653,N_9757);
and U9818 (N_9818,N_9737,N_9655);
xnor U9819 (N_9819,N_9773,N_9645);
nor U9820 (N_9820,N_9728,N_9642);
or U9821 (N_9821,N_9666,N_9698);
or U9822 (N_9822,N_9798,N_9662);
or U9823 (N_9823,N_9751,N_9628);
and U9824 (N_9824,N_9791,N_9743);
nand U9825 (N_9825,N_9741,N_9786);
or U9826 (N_9826,N_9616,N_9733);
nor U9827 (N_9827,N_9745,N_9761);
nor U9828 (N_9828,N_9726,N_9683);
and U9829 (N_9829,N_9625,N_9793);
and U9830 (N_9830,N_9747,N_9615);
and U9831 (N_9831,N_9699,N_9738);
xor U9832 (N_9832,N_9759,N_9732);
and U9833 (N_9833,N_9649,N_9772);
nor U9834 (N_9834,N_9650,N_9603);
xnor U9835 (N_9835,N_9705,N_9670);
nor U9836 (N_9836,N_9644,N_9607);
and U9837 (N_9837,N_9690,N_9634);
and U9838 (N_9838,N_9752,N_9777);
and U9839 (N_9839,N_9609,N_9619);
or U9840 (N_9840,N_9789,N_9673);
and U9841 (N_9841,N_9784,N_9750);
and U9842 (N_9842,N_9657,N_9702);
or U9843 (N_9843,N_9780,N_9792);
xnor U9844 (N_9844,N_9675,N_9621);
xnor U9845 (N_9845,N_9693,N_9701);
xor U9846 (N_9846,N_9630,N_9680);
or U9847 (N_9847,N_9729,N_9765);
nor U9848 (N_9848,N_9749,N_9714);
xnor U9849 (N_9849,N_9770,N_9696);
or U9850 (N_9850,N_9691,N_9785);
xor U9851 (N_9851,N_9762,N_9646);
xnor U9852 (N_9852,N_9764,N_9663);
nand U9853 (N_9853,N_9727,N_9606);
xor U9854 (N_9854,N_9799,N_9664);
and U9855 (N_9855,N_9794,N_9736);
and U9856 (N_9856,N_9648,N_9710);
nor U9857 (N_9857,N_9651,N_9712);
nor U9858 (N_9858,N_9654,N_9671);
xor U9859 (N_9859,N_9618,N_9638);
and U9860 (N_9860,N_9740,N_9612);
or U9861 (N_9861,N_9629,N_9776);
and U9862 (N_9862,N_9753,N_9692);
nor U9863 (N_9863,N_9600,N_9660);
xor U9864 (N_9864,N_9790,N_9724);
and U9865 (N_9865,N_9775,N_9672);
nor U9866 (N_9866,N_9722,N_9620);
nor U9867 (N_9867,N_9611,N_9746);
nor U9868 (N_9868,N_9778,N_9686);
or U9869 (N_9869,N_9610,N_9706);
or U9870 (N_9870,N_9613,N_9624);
and U9871 (N_9871,N_9656,N_9669);
or U9872 (N_9872,N_9700,N_9771);
nor U9873 (N_9873,N_9665,N_9769);
nor U9874 (N_9874,N_9703,N_9637);
or U9875 (N_9875,N_9754,N_9647);
xor U9876 (N_9876,N_9718,N_9601);
nor U9877 (N_9877,N_9768,N_9763);
or U9878 (N_9878,N_9758,N_9795);
nor U9879 (N_9879,N_9756,N_9689);
or U9880 (N_9880,N_9709,N_9602);
xnor U9881 (N_9881,N_9748,N_9787);
nor U9882 (N_9882,N_9742,N_9635);
nor U9883 (N_9883,N_9716,N_9617);
nor U9884 (N_9884,N_9608,N_9684);
nand U9885 (N_9885,N_9695,N_9766);
nand U9886 (N_9886,N_9781,N_9623);
nor U9887 (N_9887,N_9767,N_9782);
or U9888 (N_9888,N_9631,N_9677);
and U9889 (N_9889,N_9626,N_9788);
or U9890 (N_9890,N_9725,N_9721);
xnor U9891 (N_9891,N_9605,N_9641);
and U9892 (N_9892,N_9708,N_9676);
xnor U9893 (N_9893,N_9636,N_9667);
and U9894 (N_9894,N_9755,N_9774);
xnor U9895 (N_9895,N_9687,N_9735);
and U9896 (N_9896,N_9694,N_9679);
and U9897 (N_9897,N_9633,N_9797);
nor U9898 (N_9898,N_9717,N_9704);
xor U9899 (N_9899,N_9622,N_9760);
and U9900 (N_9900,N_9658,N_9766);
and U9901 (N_9901,N_9634,N_9657);
or U9902 (N_9902,N_9667,N_9659);
and U9903 (N_9903,N_9633,N_9699);
nor U9904 (N_9904,N_9609,N_9737);
nor U9905 (N_9905,N_9787,N_9668);
xnor U9906 (N_9906,N_9644,N_9642);
and U9907 (N_9907,N_9776,N_9795);
nand U9908 (N_9908,N_9684,N_9775);
nor U9909 (N_9909,N_9611,N_9646);
nand U9910 (N_9910,N_9670,N_9799);
nor U9911 (N_9911,N_9662,N_9703);
or U9912 (N_9912,N_9687,N_9707);
nor U9913 (N_9913,N_9661,N_9682);
or U9914 (N_9914,N_9616,N_9663);
xnor U9915 (N_9915,N_9745,N_9636);
nand U9916 (N_9916,N_9798,N_9680);
nand U9917 (N_9917,N_9768,N_9660);
or U9918 (N_9918,N_9779,N_9761);
xnor U9919 (N_9919,N_9766,N_9735);
and U9920 (N_9920,N_9713,N_9738);
and U9921 (N_9921,N_9661,N_9735);
or U9922 (N_9922,N_9673,N_9651);
or U9923 (N_9923,N_9631,N_9787);
or U9924 (N_9924,N_9767,N_9766);
nor U9925 (N_9925,N_9760,N_9783);
and U9926 (N_9926,N_9715,N_9655);
nand U9927 (N_9927,N_9696,N_9759);
and U9928 (N_9928,N_9771,N_9767);
nand U9929 (N_9929,N_9732,N_9738);
xor U9930 (N_9930,N_9790,N_9715);
or U9931 (N_9931,N_9750,N_9635);
and U9932 (N_9932,N_9797,N_9732);
and U9933 (N_9933,N_9734,N_9639);
nor U9934 (N_9934,N_9667,N_9656);
nand U9935 (N_9935,N_9681,N_9728);
and U9936 (N_9936,N_9793,N_9683);
nand U9937 (N_9937,N_9676,N_9612);
or U9938 (N_9938,N_9648,N_9730);
nor U9939 (N_9939,N_9787,N_9700);
or U9940 (N_9940,N_9770,N_9750);
xnor U9941 (N_9941,N_9606,N_9739);
nor U9942 (N_9942,N_9707,N_9675);
and U9943 (N_9943,N_9678,N_9632);
nor U9944 (N_9944,N_9763,N_9790);
nand U9945 (N_9945,N_9726,N_9724);
and U9946 (N_9946,N_9760,N_9732);
or U9947 (N_9947,N_9669,N_9640);
xor U9948 (N_9948,N_9729,N_9746);
nand U9949 (N_9949,N_9761,N_9725);
xnor U9950 (N_9950,N_9712,N_9680);
and U9951 (N_9951,N_9751,N_9782);
or U9952 (N_9952,N_9605,N_9735);
and U9953 (N_9953,N_9773,N_9649);
nand U9954 (N_9954,N_9713,N_9714);
nor U9955 (N_9955,N_9738,N_9745);
nor U9956 (N_9956,N_9759,N_9788);
nor U9957 (N_9957,N_9619,N_9677);
nand U9958 (N_9958,N_9787,N_9656);
nor U9959 (N_9959,N_9643,N_9649);
nand U9960 (N_9960,N_9665,N_9678);
xnor U9961 (N_9961,N_9687,N_9732);
nor U9962 (N_9962,N_9731,N_9687);
nor U9963 (N_9963,N_9634,N_9647);
and U9964 (N_9964,N_9741,N_9658);
xor U9965 (N_9965,N_9645,N_9774);
xnor U9966 (N_9966,N_9669,N_9734);
xor U9967 (N_9967,N_9631,N_9607);
nand U9968 (N_9968,N_9714,N_9669);
nand U9969 (N_9969,N_9781,N_9733);
nor U9970 (N_9970,N_9613,N_9697);
xor U9971 (N_9971,N_9640,N_9737);
and U9972 (N_9972,N_9664,N_9669);
or U9973 (N_9973,N_9795,N_9735);
or U9974 (N_9974,N_9710,N_9733);
and U9975 (N_9975,N_9779,N_9604);
or U9976 (N_9976,N_9780,N_9630);
or U9977 (N_9977,N_9718,N_9614);
and U9978 (N_9978,N_9682,N_9600);
nand U9979 (N_9979,N_9760,N_9705);
xnor U9980 (N_9980,N_9606,N_9784);
or U9981 (N_9981,N_9638,N_9737);
nand U9982 (N_9982,N_9644,N_9757);
or U9983 (N_9983,N_9632,N_9649);
nor U9984 (N_9984,N_9741,N_9771);
or U9985 (N_9985,N_9748,N_9705);
nor U9986 (N_9986,N_9615,N_9667);
and U9987 (N_9987,N_9656,N_9684);
xnor U9988 (N_9988,N_9706,N_9750);
nand U9989 (N_9989,N_9615,N_9645);
nand U9990 (N_9990,N_9776,N_9757);
and U9991 (N_9991,N_9726,N_9645);
or U9992 (N_9992,N_9614,N_9619);
nand U9993 (N_9993,N_9623,N_9707);
nor U9994 (N_9994,N_9767,N_9778);
or U9995 (N_9995,N_9639,N_9621);
nand U9996 (N_9996,N_9767,N_9604);
nand U9997 (N_9997,N_9762,N_9784);
nand U9998 (N_9998,N_9737,N_9664);
nor U9999 (N_9999,N_9622,N_9660);
and UO_0 (O_0,N_9879,N_9857);
or UO_1 (O_1,N_9889,N_9835);
nand UO_2 (O_2,N_9850,N_9979);
nand UO_3 (O_3,N_9815,N_9853);
xnor UO_4 (O_4,N_9817,N_9859);
or UO_5 (O_5,N_9975,N_9892);
and UO_6 (O_6,N_9897,N_9810);
and UO_7 (O_7,N_9869,N_9944);
or UO_8 (O_8,N_9865,N_9968);
nand UO_9 (O_9,N_9824,N_9894);
nor UO_10 (O_10,N_9898,N_9915);
and UO_11 (O_11,N_9809,N_9996);
nand UO_12 (O_12,N_9871,N_9829);
and UO_13 (O_13,N_9937,N_9941);
nor UO_14 (O_14,N_9812,N_9973);
xnor UO_15 (O_15,N_9914,N_9805);
or UO_16 (O_16,N_9920,N_9934);
or UO_17 (O_17,N_9802,N_9856);
nand UO_18 (O_18,N_9807,N_9885);
xor UO_19 (O_19,N_9819,N_9945);
or UO_20 (O_20,N_9860,N_9884);
xnor UO_21 (O_21,N_9950,N_9982);
nor UO_22 (O_22,N_9958,N_9938);
xor UO_23 (O_23,N_9956,N_9965);
nand UO_24 (O_24,N_9844,N_9904);
nand UO_25 (O_25,N_9988,N_9926);
nor UO_26 (O_26,N_9836,N_9999);
nor UO_27 (O_27,N_9800,N_9907);
nor UO_28 (O_28,N_9964,N_9966);
and UO_29 (O_29,N_9822,N_9972);
or UO_30 (O_30,N_9881,N_9962);
nand UO_31 (O_31,N_9995,N_9909);
xor UO_32 (O_32,N_9905,N_9935);
nand UO_33 (O_33,N_9946,N_9883);
nand UO_34 (O_34,N_9895,N_9942);
nand UO_35 (O_35,N_9963,N_9910);
nand UO_36 (O_36,N_9870,N_9983);
nor UO_37 (O_37,N_9970,N_9936);
and UO_38 (O_38,N_9971,N_9900);
nand UO_39 (O_39,N_9980,N_9833);
nor UO_40 (O_40,N_9876,N_9823);
xnor UO_41 (O_41,N_9985,N_9967);
nor UO_42 (O_42,N_9811,N_9954);
or UO_43 (O_43,N_9991,N_9924);
and UO_44 (O_44,N_9801,N_9891);
and UO_45 (O_45,N_9955,N_9830);
nand UO_46 (O_46,N_9940,N_9843);
or UO_47 (O_47,N_9851,N_9989);
and UO_48 (O_48,N_9804,N_9858);
xnor UO_49 (O_49,N_9877,N_9957);
nand UO_50 (O_50,N_9960,N_9847);
xor UO_51 (O_51,N_9948,N_9931);
nor UO_52 (O_52,N_9976,N_9814);
or UO_53 (O_53,N_9855,N_9947);
nor UO_54 (O_54,N_9906,N_9925);
nand UO_55 (O_55,N_9826,N_9854);
xor UO_56 (O_56,N_9816,N_9923);
xnor UO_57 (O_57,N_9899,N_9828);
nand UO_58 (O_58,N_9808,N_9866);
nor UO_59 (O_59,N_9867,N_9997);
nor UO_60 (O_60,N_9803,N_9821);
xor UO_61 (O_61,N_9882,N_9825);
and UO_62 (O_62,N_9943,N_9813);
xor UO_63 (O_63,N_9919,N_9911);
and UO_64 (O_64,N_9951,N_9986);
or UO_65 (O_65,N_9834,N_9827);
nand UO_66 (O_66,N_9921,N_9922);
or UO_67 (O_67,N_9974,N_9952);
or UO_68 (O_68,N_9933,N_9852);
nor UO_69 (O_69,N_9978,N_9896);
and UO_70 (O_70,N_9929,N_9875);
and UO_71 (O_71,N_9837,N_9874);
and UO_72 (O_72,N_9878,N_9918);
nand UO_73 (O_73,N_9949,N_9903);
and UO_74 (O_74,N_9863,N_9873);
xor UO_75 (O_75,N_9932,N_9901);
nor UO_76 (O_76,N_9806,N_9908);
and UO_77 (O_77,N_9994,N_9845);
nor UO_78 (O_78,N_9953,N_9888);
nor UO_79 (O_79,N_9939,N_9886);
xor UO_80 (O_80,N_9820,N_9831);
xnor UO_81 (O_81,N_9981,N_9977);
or UO_82 (O_82,N_9998,N_9927);
nor UO_83 (O_83,N_9832,N_9839);
xor UO_84 (O_84,N_9849,N_9917);
nor UO_85 (O_85,N_9864,N_9928);
or UO_86 (O_86,N_9868,N_9916);
nand UO_87 (O_87,N_9838,N_9959);
or UO_88 (O_88,N_9887,N_9880);
nand UO_89 (O_89,N_9848,N_9993);
nor UO_90 (O_90,N_9912,N_9984);
and UO_91 (O_91,N_9842,N_9987);
and UO_92 (O_92,N_9893,N_9961);
nor UO_93 (O_93,N_9840,N_9913);
and UO_94 (O_94,N_9862,N_9846);
xnor UO_95 (O_95,N_9818,N_9969);
nor UO_96 (O_96,N_9930,N_9890);
xor UO_97 (O_97,N_9990,N_9872);
or UO_98 (O_98,N_9902,N_9861);
xnor UO_99 (O_99,N_9992,N_9841);
or UO_100 (O_100,N_9836,N_9950);
or UO_101 (O_101,N_9965,N_9916);
nor UO_102 (O_102,N_9953,N_9965);
and UO_103 (O_103,N_9909,N_9878);
xor UO_104 (O_104,N_9815,N_9954);
and UO_105 (O_105,N_9994,N_9882);
nand UO_106 (O_106,N_9800,N_9816);
or UO_107 (O_107,N_9910,N_9827);
or UO_108 (O_108,N_9850,N_9972);
xnor UO_109 (O_109,N_9842,N_9955);
nand UO_110 (O_110,N_9860,N_9944);
nand UO_111 (O_111,N_9953,N_9821);
or UO_112 (O_112,N_9938,N_9998);
xnor UO_113 (O_113,N_9956,N_9861);
and UO_114 (O_114,N_9971,N_9801);
xor UO_115 (O_115,N_9915,N_9899);
and UO_116 (O_116,N_9866,N_9811);
or UO_117 (O_117,N_9960,N_9874);
xor UO_118 (O_118,N_9893,N_9836);
or UO_119 (O_119,N_9815,N_9991);
nand UO_120 (O_120,N_9967,N_9975);
nor UO_121 (O_121,N_9925,N_9852);
xor UO_122 (O_122,N_9803,N_9858);
and UO_123 (O_123,N_9850,N_9983);
nor UO_124 (O_124,N_9824,N_9838);
or UO_125 (O_125,N_9937,N_9958);
nor UO_126 (O_126,N_9815,N_9985);
nand UO_127 (O_127,N_9926,N_9845);
nand UO_128 (O_128,N_9987,N_9818);
and UO_129 (O_129,N_9901,N_9960);
or UO_130 (O_130,N_9857,N_9848);
nand UO_131 (O_131,N_9956,N_9905);
and UO_132 (O_132,N_9916,N_9933);
or UO_133 (O_133,N_9971,N_9836);
nor UO_134 (O_134,N_9946,N_9827);
xnor UO_135 (O_135,N_9838,N_9835);
nor UO_136 (O_136,N_9969,N_9961);
xor UO_137 (O_137,N_9914,N_9816);
nand UO_138 (O_138,N_9868,N_9972);
xnor UO_139 (O_139,N_9965,N_9888);
xor UO_140 (O_140,N_9863,N_9973);
or UO_141 (O_141,N_9989,N_9947);
nand UO_142 (O_142,N_9815,N_9893);
and UO_143 (O_143,N_9815,N_9869);
or UO_144 (O_144,N_9922,N_9826);
and UO_145 (O_145,N_9921,N_9981);
xnor UO_146 (O_146,N_9875,N_9871);
xnor UO_147 (O_147,N_9967,N_9863);
nor UO_148 (O_148,N_9803,N_9871);
xor UO_149 (O_149,N_9889,N_9837);
xor UO_150 (O_150,N_9943,N_9883);
nor UO_151 (O_151,N_9955,N_9939);
or UO_152 (O_152,N_9897,N_9898);
or UO_153 (O_153,N_9807,N_9953);
and UO_154 (O_154,N_9994,N_9800);
nand UO_155 (O_155,N_9868,N_9886);
xor UO_156 (O_156,N_9810,N_9819);
xnor UO_157 (O_157,N_9800,N_9896);
and UO_158 (O_158,N_9966,N_9871);
nor UO_159 (O_159,N_9871,N_9986);
or UO_160 (O_160,N_9831,N_9967);
nand UO_161 (O_161,N_9822,N_9949);
nor UO_162 (O_162,N_9941,N_9863);
xnor UO_163 (O_163,N_9908,N_9873);
or UO_164 (O_164,N_9834,N_9803);
or UO_165 (O_165,N_9839,N_9874);
or UO_166 (O_166,N_9936,N_9960);
nand UO_167 (O_167,N_9968,N_9875);
and UO_168 (O_168,N_9826,N_9950);
nor UO_169 (O_169,N_9950,N_9926);
nor UO_170 (O_170,N_9841,N_9853);
nor UO_171 (O_171,N_9928,N_9865);
or UO_172 (O_172,N_9912,N_9801);
xnor UO_173 (O_173,N_9966,N_9960);
nor UO_174 (O_174,N_9896,N_9933);
xor UO_175 (O_175,N_9951,N_9868);
nor UO_176 (O_176,N_9975,N_9884);
nand UO_177 (O_177,N_9877,N_9968);
or UO_178 (O_178,N_9862,N_9991);
nand UO_179 (O_179,N_9917,N_9829);
nand UO_180 (O_180,N_9947,N_9821);
or UO_181 (O_181,N_9946,N_9910);
and UO_182 (O_182,N_9892,N_9891);
and UO_183 (O_183,N_9965,N_9968);
nand UO_184 (O_184,N_9948,N_9801);
and UO_185 (O_185,N_9940,N_9825);
xor UO_186 (O_186,N_9881,N_9928);
nor UO_187 (O_187,N_9859,N_9934);
and UO_188 (O_188,N_9839,N_9923);
and UO_189 (O_189,N_9837,N_9844);
and UO_190 (O_190,N_9899,N_9802);
and UO_191 (O_191,N_9959,N_9812);
nor UO_192 (O_192,N_9824,N_9866);
xor UO_193 (O_193,N_9872,N_9819);
nand UO_194 (O_194,N_9958,N_9869);
nand UO_195 (O_195,N_9977,N_9806);
nand UO_196 (O_196,N_9888,N_9864);
nor UO_197 (O_197,N_9913,N_9842);
nor UO_198 (O_198,N_9840,N_9936);
and UO_199 (O_199,N_9854,N_9985);
nand UO_200 (O_200,N_9814,N_9917);
xor UO_201 (O_201,N_9872,N_9943);
xor UO_202 (O_202,N_9976,N_9811);
nand UO_203 (O_203,N_9814,N_9937);
nor UO_204 (O_204,N_9917,N_9950);
nand UO_205 (O_205,N_9846,N_9929);
nor UO_206 (O_206,N_9825,N_9905);
or UO_207 (O_207,N_9924,N_9891);
xnor UO_208 (O_208,N_9803,N_9801);
and UO_209 (O_209,N_9908,N_9955);
nor UO_210 (O_210,N_9913,N_9947);
xor UO_211 (O_211,N_9919,N_9856);
xnor UO_212 (O_212,N_9923,N_9829);
or UO_213 (O_213,N_9840,N_9811);
and UO_214 (O_214,N_9833,N_9824);
xor UO_215 (O_215,N_9842,N_9964);
nor UO_216 (O_216,N_9883,N_9927);
nand UO_217 (O_217,N_9976,N_9816);
nand UO_218 (O_218,N_9984,N_9914);
or UO_219 (O_219,N_9885,N_9902);
xor UO_220 (O_220,N_9867,N_9818);
nor UO_221 (O_221,N_9814,N_9868);
and UO_222 (O_222,N_9911,N_9871);
and UO_223 (O_223,N_9940,N_9844);
nor UO_224 (O_224,N_9810,N_9998);
or UO_225 (O_225,N_9928,N_9812);
nand UO_226 (O_226,N_9974,N_9815);
and UO_227 (O_227,N_9978,N_9938);
nor UO_228 (O_228,N_9994,N_9970);
and UO_229 (O_229,N_9981,N_9885);
nand UO_230 (O_230,N_9855,N_9975);
nor UO_231 (O_231,N_9970,N_9904);
nand UO_232 (O_232,N_9929,N_9926);
nand UO_233 (O_233,N_9962,N_9987);
or UO_234 (O_234,N_9861,N_9975);
nor UO_235 (O_235,N_9901,N_9872);
and UO_236 (O_236,N_9987,N_9959);
and UO_237 (O_237,N_9981,N_9892);
xor UO_238 (O_238,N_9829,N_9889);
nand UO_239 (O_239,N_9845,N_9839);
nand UO_240 (O_240,N_9826,N_9949);
nor UO_241 (O_241,N_9807,N_9847);
or UO_242 (O_242,N_9914,N_9808);
nand UO_243 (O_243,N_9908,N_9931);
or UO_244 (O_244,N_9860,N_9845);
nand UO_245 (O_245,N_9906,N_9975);
xnor UO_246 (O_246,N_9803,N_9889);
nor UO_247 (O_247,N_9936,N_9813);
xor UO_248 (O_248,N_9922,N_9935);
or UO_249 (O_249,N_9919,N_9845);
or UO_250 (O_250,N_9946,N_9840);
or UO_251 (O_251,N_9843,N_9925);
and UO_252 (O_252,N_9996,N_9992);
nor UO_253 (O_253,N_9982,N_9900);
and UO_254 (O_254,N_9835,N_9987);
or UO_255 (O_255,N_9873,N_9987);
nor UO_256 (O_256,N_9831,N_9864);
and UO_257 (O_257,N_9875,N_9911);
or UO_258 (O_258,N_9876,N_9847);
nor UO_259 (O_259,N_9970,N_9851);
nand UO_260 (O_260,N_9850,N_9897);
nand UO_261 (O_261,N_9827,N_9932);
nand UO_262 (O_262,N_9920,N_9937);
nand UO_263 (O_263,N_9909,N_9970);
nor UO_264 (O_264,N_9977,N_9852);
nor UO_265 (O_265,N_9920,N_9940);
nand UO_266 (O_266,N_9900,N_9849);
nand UO_267 (O_267,N_9802,N_9906);
nor UO_268 (O_268,N_9962,N_9991);
nor UO_269 (O_269,N_9865,N_9989);
nand UO_270 (O_270,N_9963,N_9935);
nor UO_271 (O_271,N_9816,N_9951);
nand UO_272 (O_272,N_9958,N_9864);
nor UO_273 (O_273,N_9802,N_9888);
and UO_274 (O_274,N_9958,N_9934);
xnor UO_275 (O_275,N_9825,N_9845);
nand UO_276 (O_276,N_9869,N_9977);
or UO_277 (O_277,N_9893,N_9942);
and UO_278 (O_278,N_9845,N_9868);
nor UO_279 (O_279,N_9855,N_9934);
nand UO_280 (O_280,N_9944,N_9829);
or UO_281 (O_281,N_9871,N_9998);
xnor UO_282 (O_282,N_9906,N_9853);
nand UO_283 (O_283,N_9926,N_9833);
nor UO_284 (O_284,N_9883,N_9986);
or UO_285 (O_285,N_9874,N_9968);
nor UO_286 (O_286,N_9962,N_9956);
and UO_287 (O_287,N_9948,N_9932);
xnor UO_288 (O_288,N_9988,N_9872);
or UO_289 (O_289,N_9956,N_9822);
or UO_290 (O_290,N_9914,N_9965);
or UO_291 (O_291,N_9902,N_9981);
nor UO_292 (O_292,N_9884,N_9940);
xnor UO_293 (O_293,N_9994,N_9875);
nand UO_294 (O_294,N_9988,N_9826);
nor UO_295 (O_295,N_9990,N_9942);
or UO_296 (O_296,N_9831,N_9977);
xnor UO_297 (O_297,N_9952,N_9917);
and UO_298 (O_298,N_9991,N_9910);
xnor UO_299 (O_299,N_9829,N_9899);
or UO_300 (O_300,N_9930,N_9831);
nor UO_301 (O_301,N_9909,N_9829);
xnor UO_302 (O_302,N_9961,N_9807);
nor UO_303 (O_303,N_9876,N_9996);
or UO_304 (O_304,N_9978,N_9833);
nor UO_305 (O_305,N_9867,N_9849);
and UO_306 (O_306,N_9879,N_9846);
nor UO_307 (O_307,N_9848,N_9844);
nor UO_308 (O_308,N_9880,N_9830);
or UO_309 (O_309,N_9851,N_9975);
xnor UO_310 (O_310,N_9831,N_9950);
nor UO_311 (O_311,N_9866,N_9863);
and UO_312 (O_312,N_9945,N_9961);
nand UO_313 (O_313,N_9859,N_9899);
nand UO_314 (O_314,N_9837,N_9834);
xnor UO_315 (O_315,N_9906,N_9915);
nor UO_316 (O_316,N_9846,N_9802);
and UO_317 (O_317,N_9892,N_9908);
xor UO_318 (O_318,N_9821,N_9835);
nand UO_319 (O_319,N_9953,N_9963);
xnor UO_320 (O_320,N_9887,N_9822);
and UO_321 (O_321,N_9855,N_9964);
and UO_322 (O_322,N_9824,N_9860);
or UO_323 (O_323,N_9808,N_9903);
nor UO_324 (O_324,N_9856,N_9916);
and UO_325 (O_325,N_9818,N_9898);
nor UO_326 (O_326,N_9899,N_9911);
or UO_327 (O_327,N_9914,N_9970);
nor UO_328 (O_328,N_9986,N_9940);
and UO_329 (O_329,N_9928,N_9914);
nor UO_330 (O_330,N_9817,N_9906);
nand UO_331 (O_331,N_9866,N_9918);
nor UO_332 (O_332,N_9977,N_9894);
nor UO_333 (O_333,N_9844,N_9872);
and UO_334 (O_334,N_9805,N_9990);
nor UO_335 (O_335,N_9986,N_9947);
and UO_336 (O_336,N_9838,N_9854);
xnor UO_337 (O_337,N_9954,N_9802);
xnor UO_338 (O_338,N_9862,N_9894);
or UO_339 (O_339,N_9834,N_9962);
or UO_340 (O_340,N_9868,N_9809);
nor UO_341 (O_341,N_9909,N_9936);
and UO_342 (O_342,N_9855,N_9830);
and UO_343 (O_343,N_9856,N_9840);
nand UO_344 (O_344,N_9932,N_9829);
or UO_345 (O_345,N_9851,N_9811);
nor UO_346 (O_346,N_9944,N_9843);
nand UO_347 (O_347,N_9803,N_9951);
or UO_348 (O_348,N_9811,N_9824);
and UO_349 (O_349,N_9924,N_9818);
xnor UO_350 (O_350,N_9811,N_9898);
or UO_351 (O_351,N_9985,N_9919);
xnor UO_352 (O_352,N_9965,N_9943);
nor UO_353 (O_353,N_9957,N_9850);
xor UO_354 (O_354,N_9850,N_9821);
nor UO_355 (O_355,N_9900,N_9972);
and UO_356 (O_356,N_9882,N_9812);
xnor UO_357 (O_357,N_9941,N_9873);
or UO_358 (O_358,N_9933,N_9968);
nor UO_359 (O_359,N_9844,N_9891);
nand UO_360 (O_360,N_9877,N_9857);
nor UO_361 (O_361,N_9987,N_9863);
or UO_362 (O_362,N_9823,N_9981);
nand UO_363 (O_363,N_9921,N_9962);
and UO_364 (O_364,N_9927,N_9920);
xnor UO_365 (O_365,N_9982,N_9963);
xor UO_366 (O_366,N_9857,N_9852);
xor UO_367 (O_367,N_9917,N_9823);
or UO_368 (O_368,N_9996,N_9824);
and UO_369 (O_369,N_9812,N_9993);
or UO_370 (O_370,N_9919,N_9950);
nor UO_371 (O_371,N_9857,N_9907);
xor UO_372 (O_372,N_9922,N_9996);
and UO_373 (O_373,N_9895,N_9959);
or UO_374 (O_374,N_9932,N_9830);
nand UO_375 (O_375,N_9929,N_9936);
nand UO_376 (O_376,N_9824,N_9862);
nand UO_377 (O_377,N_9984,N_9870);
xor UO_378 (O_378,N_9838,N_9944);
nand UO_379 (O_379,N_9876,N_9932);
or UO_380 (O_380,N_9998,N_9906);
xor UO_381 (O_381,N_9841,N_9974);
and UO_382 (O_382,N_9860,N_9974);
nor UO_383 (O_383,N_9961,N_9845);
or UO_384 (O_384,N_9813,N_9938);
or UO_385 (O_385,N_9859,N_9976);
or UO_386 (O_386,N_9959,N_9851);
xor UO_387 (O_387,N_9840,N_9845);
nor UO_388 (O_388,N_9912,N_9919);
and UO_389 (O_389,N_9821,N_9889);
and UO_390 (O_390,N_9961,N_9931);
xnor UO_391 (O_391,N_9862,N_9930);
nand UO_392 (O_392,N_9849,N_9933);
or UO_393 (O_393,N_9941,N_9835);
nand UO_394 (O_394,N_9817,N_9982);
nor UO_395 (O_395,N_9929,N_9907);
and UO_396 (O_396,N_9835,N_9939);
and UO_397 (O_397,N_9844,N_9987);
and UO_398 (O_398,N_9983,N_9811);
xor UO_399 (O_399,N_9822,N_9930);
nor UO_400 (O_400,N_9822,N_9883);
nor UO_401 (O_401,N_9877,N_9841);
or UO_402 (O_402,N_9900,N_9901);
or UO_403 (O_403,N_9844,N_9878);
xor UO_404 (O_404,N_9869,N_9892);
or UO_405 (O_405,N_9809,N_9937);
nor UO_406 (O_406,N_9972,N_9851);
nand UO_407 (O_407,N_9905,N_9848);
and UO_408 (O_408,N_9871,N_9858);
nand UO_409 (O_409,N_9894,N_9965);
and UO_410 (O_410,N_9931,N_9806);
and UO_411 (O_411,N_9940,N_9956);
nand UO_412 (O_412,N_9979,N_9905);
or UO_413 (O_413,N_9834,N_9812);
nand UO_414 (O_414,N_9813,N_9984);
xor UO_415 (O_415,N_9828,N_9997);
nor UO_416 (O_416,N_9914,N_9958);
and UO_417 (O_417,N_9890,N_9975);
and UO_418 (O_418,N_9836,N_9809);
nor UO_419 (O_419,N_9857,N_9843);
nand UO_420 (O_420,N_9877,N_9896);
and UO_421 (O_421,N_9806,N_9866);
or UO_422 (O_422,N_9901,N_9863);
or UO_423 (O_423,N_9964,N_9997);
nand UO_424 (O_424,N_9808,N_9891);
nor UO_425 (O_425,N_9822,N_9810);
nand UO_426 (O_426,N_9873,N_9967);
nand UO_427 (O_427,N_9938,N_9997);
nand UO_428 (O_428,N_9878,N_9863);
and UO_429 (O_429,N_9939,N_9946);
xor UO_430 (O_430,N_9887,N_9895);
xnor UO_431 (O_431,N_9947,N_9978);
or UO_432 (O_432,N_9856,N_9920);
and UO_433 (O_433,N_9820,N_9932);
nand UO_434 (O_434,N_9936,N_9846);
nand UO_435 (O_435,N_9893,N_9892);
xnor UO_436 (O_436,N_9869,N_9834);
nand UO_437 (O_437,N_9800,N_9846);
nand UO_438 (O_438,N_9955,N_9993);
and UO_439 (O_439,N_9811,N_9947);
nand UO_440 (O_440,N_9976,N_9963);
or UO_441 (O_441,N_9939,N_9993);
xor UO_442 (O_442,N_9903,N_9857);
nand UO_443 (O_443,N_9901,N_9876);
and UO_444 (O_444,N_9809,N_9899);
nand UO_445 (O_445,N_9807,N_9808);
or UO_446 (O_446,N_9977,N_9942);
nand UO_447 (O_447,N_9993,N_9933);
and UO_448 (O_448,N_9944,N_9970);
nor UO_449 (O_449,N_9875,N_9973);
nor UO_450 (O_450,N_9802,N_9835);
xor UO_451 (O_451,N_9992,N_9825);
xor UO_452 (O_452,N_9916,N_9915);
xor UO_453 (O_453,N_9828,N_9884);
nor UO_454 (O_454,N_9891,N_9839);
or UO_455 (O_455,N_9813,N_9958);
and UO_456 (O_456,N_9918,N_9905);
xor UO_457 (O_457,N_9926,N_9881);
xnor UO_458 (O_458,N_9826,N_9905);
nand UO_459 (O_459,N_9905,N_9928);
and UO_460 (O_460,N_9897,N_9885);
nor UO_461 (O_461,N_9965,N_9932);
xor UO_462 (O_462,N_9974,N_9835);
or UO_463 (O_463,N_9807,N_9882);
nand UO_464 (O_464,N_9880,N_9907);
nand UO_465 (O_465,N_9876,N_9931);
or UO_466 (O_466,N_9827,N_9861);
nor UO_467 (O_467,N_9854,N_9970);
xor UO_468 (O_468,N_9989,N_9858);
and UO_469 (O_469,N_9916,N_9810);
xnor UO_470 (O_470,N_9831,N_9861);
xnor UO_471 (O_471,N_9939,N_9839);
or UO_472 (O_472,N_9902,N_9993);
xor UO_473 (O_473,N_9907,N_9892);
and UO_474 (O_474,N_9809,N_9993);
nand UO_475 (O_475,N_9843,N_9880);
xnor UO_476 (O_476,N_9906,N_9871);
or UO_477 (O_477,N_9817,N_9803);
or UO_478 (O_478,N_9999,N_9851);
or UO_479 (O_479,N_9952,N_9980);
and UO_480 (O_480,N_9943,N_9876);
nor UO_481 (O_481,N_9849,N_9996);
or UO_482 (O_482,N_9870,N_9907);
xnor UO_483 (O_483,N_9986,N_9900);
and UO_484 (O_484,N_9957,N_9946);
xor UO_485 (O_485,N_9936,N_9897);
or UO_486 (O_486,N_9846,N_9911);
xnor UO_487 (O_487,N_9833,N_9852);
nor UO_488 (O_488,N_9876,N_9862);
and UO_489 (O_489,N_9880,N_9862);
or UO_490 (O_490,N_9807,N_9816);
nor UO_491 (O_491,N_9800,N_9943);
or UO_492 (O_492,N_9870,N_9846);
nand UO_493 (O_493,N_9844,N_9958);
nor UO_494 (O_494,N_9953,N_9856);
nand UO_495 (O_495,N_9986,N_9966);
nand UO_496 (O_496,N_9910,N_9995);
nand UO_497 (O_497,N_9816,N_9866);
nor UO_498 (O_498,N_9815,N_9875);
or UO_499 (O_499,N_9930,N_9833);
or UO_500 (O_500,N_9875,N_9806);
or UO_501 (O_501,N_9841,N_9908);
and UO_502 (O_502,N_9934,N_9947);
and UO_503 (O_503,N_9904,N_9827);
or UO_504 (O_504,N_9873,N_9929);
nand UO_505 (O_505,N_9946,N_9829);
nor UO_506 (O_506,N_9865,N_9971);
nand UO_507 (O_507,N_9842,N_9888);
xor UO_508 (O_508,N_9816,N_9811);
nand UO_509 (O_509,N_9841,N_9813);
nor UO_510 (O_510,N_9988,N_9898);
and UO_511 (O_511,N_9972,N_9817);
nor UO_512 (O_512,N_9978,N_9858);
and UO_513 (O_513,N_9918,N_9885);
nor UO_514 (O_514,N_9952,N_9987);
xor UO_515 (O_515,N_9847,N_9901);
nand UO_516 (O_516,N_9985,N_9946);
and UO_517 (O_517,N_9831,N_9946);
or UO_518 (O_518,N_9861,N_9803);
xor UO_519 (O_519,N_9989,N_9828);
and UO_520 (O_520,N_9969,N_9970);
nand UO_521 (O_521,N_9907,N_9841);
nand UO_522 (O_522,N_9982,N_9831);
xor UO_523 (O_523,N_9907,N_9898);
or UO_524 (O_524,N_9886,N_9972);
nand UO_525 (O_525,N_9858,N_9856);
and UO_526 (O_526,N_9976,N_9959);
and UO_527 (O_527,N_9956,N_9989);
xor UO_528 (O_528,N_9952,N_9861);
xor UO_529 (O_529,N_9939,N_9856);
nand UO_530 (O_530,N_9881,N_9862);
nand UO_531 (O_531,N_9836,N_9927);
xnor UO_532 (O_532,N_9961,N_9947);
and UO_533 (O_533,N_9826,N_9953);
nor UO_534 (O_534,N_9919,N_9905);
or UO_535 (O_535,N_9923,N_9948);
or UO_536 (O_536,N_9978,N_9864);
nand UO_537 (O_537,N_9916,N_9904);
nand UO_538 (O_538,N_9848,N_9858);
nor UO_539 (O_539,N_9892,N_9831);
nor UO_540 (O_540,N_9855,N_9989);
nor UO_541 (O_541,N_9814,N_9961);
xor UO_542 (O_542,N_9883,N_9980);
nand UO_543 (O_543,N_9858,N_9863);
or UO_544 (O_544,N_9874,N_9875);
xor UO_545 (O_545,N_9875,N_9812);
nand UO_546 (O_546,N_9936,N_9986);
nor UO_547 (O_547,N_9924,N_9867);
nand UO_548 (O_548,N_9972,N_9879);
nor UO_549 (O_549,N_9887,N_9910);
or UO_550 (O_550,N_9860,N_9960);
nand UO_551 (O_551,N_9912,N_9913);
xor UO_552 (O_552,N_9901,N_9846);
xor UO_553 (O_553,N_9887,N_9818);
nor UO_554 (O_554,N_9962,N_9810);
nor UO_555 (O_555,N_9850,N_9872);
nor UO_556 (O_556,N_9826,N_9967);
xnor UO_557 (O_557,N_9841,N_9995);
xor UO_558 (O_558,N_9808,N_9872);
and UO_559 (O_559,N_9997,N_9915);
xor UO_560 (O_560,N_9876,N_9965);
nor UO_561 (O_561,N_9908,N_9867);
or UO_562 (O_562,N_9818,N_9870);
or UO_563 (O_563,N_9811,N_9975);
and UO_564 (O_564,N_9952,N_9944);
and UO_565 (O_565,N_9850,N_9964);
or UO_566 (O_566,N_9941,N_9933);
and UO_567 (O_567,N_9984,N_9882);
xor UO_568 (O_568,N_9910,N_9943);
and UO_569 (O_569,N_9848,N_9998);
xor UO_570 (O_570,N_9947,N_9854);
nor UO_571 (O_571,N_9929,N_9976);
nand UO_572 (O_572,N_9886,N_9857);
or UO_573 (O_573,N_9819,N_9903);
and UO_574 (O_574,N_9972,N_9865);
and UO_575 (O_575,N_9920,N_9852);
nand UO_576 (O_576,N_9866,N_9953);
nand UO_577 (O_577,N_9945,N_9920);
xor UO_578 (O_578,N_9800,N_9843);
xor UO_579 (O_579,N_9919,N_9862);
and UO_580 (O_580,N_9882,N_9815);
and UO_581 (O_581,N_9921,N_9940);
nor UO_582 (O_582,N_9903,N_9858);
nand UO_583 (O_583,N_9960,N_9988);
or UO_584 (O_584,N_9867,N_9931);
or UO_585 (O_585,N_9966,N_9934);
xnor UO_586 (O_586,N_9832,N_9942);
xnor UO_587 (O_587,N_9848,N_9840);
nor UO_588 (O_588,N_9826,N_9937);
and UO_589 (O_589,N_9843,N_9965);
xor UO_590 (O_590,N_9960,N_9989);
nand UO_591 (O_591,N_9981,N_9811);
xor UO_592 (O_592,N_9976,N_9893);
nand UO_593 (O_593,N_9803,N_9868);
or UO_594 (O_594,N_9843,N_9990);
and UO_595 (O_595,N_9991,N_9860);
nand UO_596 (O_596,N_9852,N_9817);
nand UO_597 (O_597,N_9967,N_9916);
and UO_598 (O_598,N_9993,N_9846);
xor UO_599 (O_599,N_9960,N_9930);
or UO_600 (O_600,N_9936,N_9979);
nand UO_601 (O_601,N_9918,N_9998);
or UO_602 (O_602,N_9818,N_9941);
nand UO_603 (O_603,N_9830,N_9867);
xor UO_604 (O_604,N_9841,N_9862);
and UO_605 (O_605,N_9920,N_9811);
or UO_606 (O_606,N_9859,N_9806);
nand UO_607 (O_607,N_9804,N_9950);
and UO_608 (O_608,N_9899,N_9874);
or UO_609 (O_609,N_9995,N_9908);
or UO_610 (O_610,N_9926,N_9863);
xnor UO_611 (O_611,N_9806,N_9920);
nand UO_612 (O_612,N_9861,N_9875);
and UO_613 (O_613,N_9824,N_9922);
xor UO_614 (O_614,N_9908,N_9839);
or UO_615 (O_615,N_9910,N_9972);
nor UO_616 (O_616,N_9988,N_9940);
and UO_617 (O_617,N_9874,N_9832);
nand UO_618 (O_618,N_9911,N_9802);
or UO_619 (O_619,N_9926,N_9928);
xor UO_620 (O_620,N_9927,N_9903);
nor UO_621 (O_621,N_9980,N_9818);
and UO_622 (O_622,N_9898,N_9837);
nor UO_623 (O_623,N_9853,N_9834);
xnor UO_624 (O_624,N_9843,N_9998);
or UO_625 (O_625,N_9890,N_9928);
xor UO_626 (O_626,N_9971,N_9933);
nor UO_627 (O_627,N_9992,N_9872);
and UO_628 (O_628,N_9894,N_9934);
nor UO_629 (O_629,N_9970,N_9830);
and UO_630 (O_630,N_9993,N_9888);
xnor UO_631 (O_631,N_9975,N_9887);
xnor UO_632 (O_632,N_9999,N_9868);
and UO_633 (O_633,N_9918,N_9845);
and UO_634 (O_634,N_9929,N_9843);
and UO_635 (O_635,N_9892,N_9937);
nor UO_636 (O_636,N_9871,N_9872);
and UO_637 (O_637,N_9847,N_9835);
xnor UO_638 (O_638,N_9933,N_9984);
xor UO_639 (O_639,N_9989,N_9819);
nor UO_640 (O_640,N_9891,N_9905);
and UO_641 (O_641,N_9993,N_9926);
or UO_642 (O_642,N_9859,N_9904);
nand UO_643 (O_643,N_9837,N_9977);
nand UO_644 (O_644,N_9893,N_9971);
and UO_645 (O_645,N_9920,N_9922);
nand UO_646 (O_646,N_9838,N_9833);
or UO_647 (O_647,N_9800,N_9992);
nand UO_648 (O_648,N_9957,N_9927);
or UO_649 (O_649,N_9863,N_9922);
xnor UO_650 (O_650,N_9890,N_9885);
xor UO_651 (O_651,N_9944,N_9965);
nand UO_652 (O_652,N_9995,N_9856);
xor UO_653 (O_653,N_9805,N_9908);
and UO_654 (O_654,N_9843,N_9881);
nand UO_655 (O_655,N_9805,N_9850);
and UO_656 (O_656,N_9840,N_9975);
nor UO_657 (O_657,N_9982,N_9810);
xnor UO_658 (O_658,N_9968,N_9958);
xnor UO_659 (O_659,N_9927,N_9982);
or UO_660 (O_660,N_9928,N_9842);
or UO_661 (O_661,N_9818,N_9819);
or UO_662 (O_662,N_9909,N_9825);
nor UO_663 (O_663,N_9828,N_9960);
and UO_664 (O_664,N_9919,N_9810);
xnor UO_665 (O_665,N_9902,N_9960);
nand UO_666 (O_666,N_9903,N_9936);
xor UO_667 (O_667,N_9836,N_9904);
and UO_668 (O_668,N_9817,N_9836);
and UO_669 (O_669,N_9858,N_9958);
or UO_670 (O_670,N_9881,N_9886);
and UO_671 (O_671,N_9931,N_9951);
and UO_672 (O_672,N_9931,N_9877);
nor UO_673 (O_673,N_9941,N_9801);
or UO_674 (O_674,N_9983,N_9959);
nor UO_675 (O_675,N_9835,N_9828);
or UO_676 (O_676,N_9990,N_9820);
nand UO_677 (O_677,N_9804,N_9811);
nand UO_678 (O_678,N_9806,N_9878);
or UO_679 (O_679,N_9953,N_9935);
xor UO_680 (O_680,N_9808,N_9845);
and UO_681 (O_681,N_9862,N_9892);
nor UO_682 (O_682,N_9864,N_9972);
and UO_683 (O_683,N_9970,N_9814);
nand UO_684 (O_684,N_9832,N_9834);
and UO_685 (O_685,N_9837,N_9900);
or UO_686 (O_686,N_9985,N_9846);
nor UO_687 (O_687,N_9868,N_9900);
nand UO_688 (O_688,N_9956,N_9863);
nor UO_689 (O_689,N_9897,N_9961);
or UO_690 (O_690,N_9822,N_9950);
nor UO_691 (O_691,N_9920,N_9981);
or UO_692 (O_692,N_9909,N_9954);
xnor UO_693 (O_693,N_9842,N_9927);
xor UO_694 (O_694,N_9921,N_9877);
nor UO_695 (O_695,N_9819,N_9953);
xor UO_696 (O_696,N_9816,N_9863);
xor UO_697 (O_697,N_9863,N_9840);
nor UO_698 (O_698,N_9976,N_9800);
xnor UO_699 (O_699,N_9926,N_9861);
nor UO_700 (O_700,N_9822,N_9968);
and UO_701 (O_701,N_9960,N_9807);
nand UO_702 (O_702,N_9876,N_9875);
nand UO_703 (O_703,N_9916,N_9887);
and UO_704 (O_704,N_9861,N_9818);
nor UO_705 (O_705,N_9851,N_9940);
or UO_706 (O_706,N_9845,N_9822);
and UO_707 (O_707,N_9863,N_9892);
and UO_708 (O_708,N_9975,N_9844);
or UO_709 (O_709,N_9866,N_9978);
nand UO_710 (O_710,N_9827,N_9846);
or UO_711 (O_711,N_9881,N_9978);
xnor UO_712 (O_712,N_9970,N_9852);
and UO_713 (O_713,N_9937,N_9911);
xor UO_714 (O_714,N_9980,N_9857);
nand UO_715 (O_715,N_9824,N_9963);
nor UO_716 (O_716,N_9888,N_9916);
nor UO_717 (O_717,N_9926,N_9857);
nor UO_718 (O_718,N_9953,N_9956);
nand UO_719 (O_719,N_9842,N_9828);
nor UO_720 (O_720,N_9881,N_9870);
nor UO_721 (O_721,N_9906,N_9889);
nor UO_722 (O_722,N_9838,N_9902);
and UO_723 (O_723,N_9812,N_9807);
nor UO_724 (O_724,N_9837,N_9932);
xnor UO_725 (O_725,N_9884,N_9937);
nor UO_726 (O_726,N_9897,N_9976);
nor UO_727 (O_727,N_9995,N_9866);
nand UO_728 (O_728,N_9975,N_9866);
xor UO_729 (O_729,N_9828,N_9973);
or UO_730 (O_730,N_9899,N_9882);
xor UO_731 (O_731,N_9967,N_9973);
xor UO_732 (O_732,N_9844,N_9809);
nand UO_733 (O_733,N_9907,N_9918);
nand UO_734 (O_734,N_9847,N_9991);
nand UO_735 (O_735,N_9874,N_9806);
or UO_736 (O_736,N_9881,N_9942);
nor UO_737 (O_737,N_9956,N_9846);
nor UO_738 (O_738,N_9962,N_9928);
xnor UO_739 (O_739,N_9988,N_9808);
xnor UO_740 (O_740,N_9849,N_9882);
nor UO_741 (O_741,N_9847,N_9858);
xnor UO_742 (O_742,N_9987,N_9920);
nor UO_743 (O_743,N_9984,N_9932);
nand UO_744 (O_744,N_9992,N_9889);
and UO_745 (O_745,N_9847,N_9905);
nor UO_746 (O_746,N_9855,N_9974);
nor UO_747 (O_747,N_9873,N_9806);
nand UO_748 (O_748,N_9989,N_9908);
or UO_749 (O_749,N_9976,N_9887);
xnor UO_750 (O_750,N_9949,N_9901);
nor UO_751 (O_751,N_9828,N_9848);
or UO_752 (O_752,N_9931,N_9847);
and UO_753 (O_753,N_9869,N_9947);
nand UO_754 (O_754,N_9970,N_9813);
and UO_755 (O_755,N_9837,N_9922);
xor UO_756 (O_756,N_9969,N_9897);
and UO_757 (O_757,N_9955,N_9834);
nor UO_758 (O_758,N_9943,N_9994);
nor UO_759 (O_759,N_9859,N_9832);
nand UO_760 (O_760,N_9866,N_9946);
and UO_761 (O_761,N_9850,N_9961);
xor UO_762 (O_762,N_9992,N_9873);
xor UO_763 (O_763,N_9942,N_9842);
nor UO_764 (O_764,N_9834,N_9948);
and UO_765 (O_765,N_9858,N_9965);
or UO_766 (O_766,N_9894,N_9864);
or UO_767 (O_767,N_9808,N_9925);
or UO_768 (O_768,N_9925,N_9833);
nand UO_769 (O_769,N_9829,N_9872);
and UO_770 (O_770,N_9829,N_9888);
and UO_771 (O_771,N_9865,N_9878);
and UO_772 (O_772,N_9974,N_9883);
and UO_773 (O_773,N_9983,N_9996);
xnor UO_774 (O_774,N_9908,N_9869);
xnor UO_775 (O_775,N_9907,N_9976);
xor UO_776 (O_776,N_9823,N_9859);
and UO_777 (O_777,N_9902,N_9982);
or UO_778 (O_778,N_9875,N_9930);
nand UO_779 (O_779,N_9912,N_9986);
and UO_780 (O_780,N_9956,N_9992);
nor UO_781 (O_781,N_9804,N_9902);
xor UO_782 (O_782,N_9852,N_9844);
nand UO_783 (O_783,N_9896,N_9834);
or UO_784 (O_784,N_9801,N_9800);
or UO_785 (O_785,N_9934,N_9921);
nor UO_786 (O_786,N_9970,N_9897);
xor UO_787 (O_787,N_9812,N_9981);
and UO_788 (O_788,N_9836,N_9990);
nand UO_789 (O_789,N_9883,N_9820);
nand UO_790 (O_790,N_9932,N_9970);
nand UO_791 (O_791,N_9911,N_9881);
nand UO_792 (O_792,N_9984,N_9902);
nor UO_793 (O_793,N_9848,N_9884);
and UO_794 (O_794,N_9812,N_9879);
and UO_795 (O_795,N_9924,N_9957);
or UO_796 (O_796,N_9836,N_9820);
and UO_797 (O_797,N_9811,N_9859);
and UO_798 (O_798,N_9871,N_9835);
and UO_799 (O_799,N_9887,N_9954);
nor UO_800 (O_800,N_9801,N_9862);
nor UO_801 (O_801,N_9836,N_9936);
xor UO_802 (O_802,N_9970,N_9922);
nand UO_803 (O_803,N_9867,N_9813);
or UO_804 (O_804,N_9990,N_9875);
nor UO_805 (O_805,N_9983,N_9992);
and UO_806 (O_806,N_9934,N_9899);
or UO_807 (O_807,N_9927,N_9977);
and UO_808 (O_808,N_9914,N_9861);
or UO_809 (O_809,N_9921,N_9846);
and UO_810 (O_810,N_9992,N_9802);
or UO_811 (O_811,N_9919,N_9873);
and UO_812 (O_812,N_9940,N_9811);
nor UO_813 (O_813,N_9894,N_9962);
or UO_814 (O_814,N_9836,N_9918);
nor UO_815 (O_815,N_9832,N_9829);
nand UO_816 (O_816,N_9823,N_9944);
or UO_817 (O_817,N_9865,N_9891);
or UO_818 (O_818,N_9959,N_9820);
and UO_819 (O_819,N_9815,N_9850);
or UO_820 (O_820,N_9802,N_9925);
nor UO_821 (O_821,N_9921,N_9842);
or UO_822 (O_822,N_9885,N_9837);
or UO_823 (O_823,N_9992,N_9963);
nand UO_824 (O_824,N_9897,N_9941);
or UO_825 (O_825,N_9938,N_9854);
and UO_826 (O_826,N_9912,N_9827);
nor UO_827 (O_827,N_9945,N_9998);
or UO_828 (O_828,N_9982,N_9952);
nand UO_829 (O_829,N_9957,N_9829);
nor UO_830 (O_830,N_9822,N_9923);
xor UO_831 (O_831,N_9984,N_9947);
or UO_832 (O_832,N_9901,N_9991);
xor UO_833 (O_833,N_9950,N_9949);
nor UO_834 (O_834,N_9803,N_9978);
nand UO_835 (O_835,N_9843,N_9996);
nand UO_836 (O_836,N_9807,N_9906);
nor UO_837 (O_837,N_9868,N_9961);
nand UO_838 (O_838,N_9916,N_9919);
nor UO_839 (O_839,N_9920,N_9885);
and UO_840 (O_840,N_9951,N_9978);
nand UO_841 (O_841,N_9904,N_9865);
nand UO_842 (O_842,N_9924,N_9802);
nor UO_843 (O_843,N_9944,N_9954);
nor UO_844 (O_844,N_9970,N_9952);
xnor UO_845 (O_845,N_9813,N_9874);
and UO_846 (O_846,N_9822,N_9894);
xnor UO_847 (O_847,N_9809,N_9834);
nand UO_848 (O_848,N_9874,N_9939);
xor UO_849 (O_849,N_9829,N_9881);
xnor UO_850 (O_850,N_9807,N_9860);
nand UO_851 (O_851,N_9946,N_9876);
or UO_852 (O_852,N_9823,N_9950);
nand UO_853 (O_853,N_9858,N_9822);
nor UO_854 (O_854,N_9876,N_9857);
nand UO_855 (O_855,N_9817,N_9992);
xnor UO_856 (O_856,N_9857,N_9953);
nor UO_857 (O_857,N_9961,N_9817);
nor UO_858 (O_858,N_9915,N_9846);
and UO_859 (O_859,N_9916,N_9822);
or UO_860 (O_860,N_9809,N_9821);
nor UO_861 (O_861,N_9811,N_9930);
nand UO_862 (O_862,N_9846,N_9905);
xor UO_863 (O_863,N_9828,N_9810);
xnor UO_864 (O_864,N_9891,N_9850);
and UO_865 (O_865,N_9826,N_9850);
and UO_866 (O_866,N_9901,N_9810);
and UO_867 (O_867,N_9932,N_9818);
nand UO_868 (O_868,N_9833,N_9907);
and UO_869 (O_869,N_9891,N_9984);
xor UO_870 (O_870,N_9862,N_9970);
and UO_871 (O_871,N_9836,N_9807);
nand UO_872 (O_872,N_9974,N_9981);
nor UO_873 (O_873,N_9860,N_9871);
xnor UO_874 (O_874,N_9889,N_9932);
and UO_875 (O_875,N_9970,N_9947);
or UO_876 (O_876,N_9890,N_9963);
or UO_877 (O_877,N_9977,N_9851);
or UO_878 (O_878,N_9828,N_9886);
nor UO_879 (O_879,N_9871,N_9964);
xor UO_880 (O_880,N_9832,N_9909);
nand UO_881 (O_881,N_9994,N_9936);
or UO_882 (O_882,N_9882,N_9964);
nand UO_883 (O_883,N_9821,N_9921);
xnor UO_884 (O_884,N_9961,N_9912);
and UO_885 (O_885,N_9883,N_9918);
xnor UO_886 (O_886,N_9968,N_9889);
nor UO_887 (O_887,N_9812,N_9860);
nand UO_888 (O_888,N_9826,N_9845);
nand UO_889 (O_889,N_9968,N_9915);
xnor UO_890 (O_890,N_9910,N_9862);
and UO_891 (O_891,N_9992,N_9810);
nand UO_892 (O_892,N_9932,N_9874);
nand UO_893 (O_893,N_9970,N_9946);
xor UO_894 (O_894,N_9863,N_9995);
and UO_895 (O_895,N_9999,N_9973);
nor UO_896 (O_896,N_9814,N_9880);
and UO_897 (O_897,N_9995,N_9921);
xnor UO_898 (O_898,N_9951,N_9852);
nor UO_899 (O_899,N_9870,N_9814);
and UO_900 (O_900,N_9802,N_9951);
nor UO_901 (O_901,N_9868,N_9995);
nand UO_902 (O_902,N_9876,N_9806);
xor UO_903 (O_903,N_9882,N_9821);
and UO_904 (O_904,N_9873,N_9817);
or UO_905 (O_905,N_9989,N_9967);
nor UO_906 (O_906,N_9902,N_9990);
or UO_907 (O_907,N_9821,N_9898);
nor UO_908 (O_908,N_9876,N_9893);
nand UO_909 (O_909,N_9858,N_9929);
or UO_910 (O_910,N_9962,N_9945);
and UO_911 (O_911,N_9838,N_9965);
xnor UO_912 (O_912,N_9910,N_9816);
nand UO_913 (O_913,N_9865,N_9902);
nand UO_914 (O_914,N_9846,N_9821);
or UO_915 (O_915,N_9841,N_9868);
nand UO_916 (O_916,N_9939,N_9843);
xnor UO_917 (O_917,N_9966,N_9858);
or UO_918 (O_918,N_9938,N_9924);
nand UO_919 (O_919,N_9990,N_9934);
nand UO_920 (O_920,N_9923,N_9922);
nor UO_921 (O_921,N_9811,N_9906);
or UO_922 (O_922,N_9984,N_9893);
or UO_923 (O_923,N_9851,N_9949);
nand UO_924 (O_924,N_9992,N_9803);
and UO_925 (O_925,N_9971,N_9939);
and UO_926 (O_926,N_9993,N_9842);
nor UO_927 (O_927,N_9978,N_9940);
and UO_928 (O_928,N_9934,N_9830);
nand UO_929 (O_929,N_9802,N_9996);
nand UO_930 (O_930,N_9832,N_9856);
xor UO_931 (O_931,N_9895,N_9840);
xnor UO_932 (O_932,N_9867,N_9891);
or UO_933 (O_933,N_9872,N_9938);
nor UO_934 (O_934,N_9887,N_9960);
nand UO_935 (O_935,N_9965,N_9930);
xnor UO_936 (O_936,N_9820,N_9824);
and UO_937 (O_937,N_9876,N_9963);
and UO_938 (O_938,N_9946,N_9976);
or UO_939 (O_939,N_9886,N_9895);
nand UO_940 (O_940,N_9913,N_9960);
nor UO_941 (O_941,N_9829,N_9996);
and UO_942 (O_942,N_9935,N_9926);
nand UO_943 (O_943,N_9931,N_9815);
and UO_944 (O_944,N_9986,N_9803);
xnor UO_945 (O_945,N_9953,N_9982);
nor UO_946 (O_946,N_9833,N_9888);
xor UO_947 (O_947,N_9806,N_9877);
or UO_948 (O_948,N_9841,N_9893);
and UO_949 (O_949,N_9838,N_9810);
or UO_950 (O_950,N_9909,N_9989);
or UO_951 (O_951,N_9856,N_9889);
nand UO_952 (O_952,N_9906,N_9968);
or UO_953 (O_953,N_9810,N_9880);
xnor UO_954 (O_954,N_9891,N_9915);
nand UO_955 (O_955,N_9939,N_9847);
nand UO_956 (O_956,N_9874,N_9938);
or UO_957 (O_957,N_9825,N_9924);
and UO_958 (O_958,N_9984,N_9812);
xnor UO_959 (O_959,N_9849,N_9990);
xor UO_960 (O_960,N_9801,N_9817);
nand UO_961 (O_961,N_9824,N_9893);
nor UO_962 (O_962,N_9817,N_9823);
nand UO_963 (O_963,N_9936,N_9820);
xnor UO_964 (O_964,N_9898,N_9810);
or UO_965 (O_965,N_9971,N_9802);
and UO_966 (O_966,N_9980,N_9984);
nor UO_967 (O_967,N_9996,N_9993);
and UO_968 (O_968,N_9867,N_9902);
nor UO_969 (O_969,N_9938,N_9825);
and UO_970 (O_970,N_9844,N_9888);
xor UO_971 (O_971,N_9844,N_9982);
xnor UO_972 (O_972,N_9834,N_9846);
or UO_973 (O_973,N_9979,N_9895);
or UO_974 (O_974,N_9957,N_9802);
nor UO_975 (O_975,N_9953,N_9921);
nor UO_976 (O_976,N_9897,N_9902);
and UO_977 (O_977,N_9836,N_9869);
and UO_978 (O_978,N_9835,N_9856);
xnor UO_979 (O_979,N_9959,N_9901);
nor UO_980 (O_980,N_9825,N_9982);
and UO_981 (O_981,N_9870,N_9850);
nor UO_982 (O_982,N_9999,N_9853);
nand UO_983 (O_983,N_9958,N_9875);
xnor UO_984 (O_984,N_9941,N_9859);
xor UO_985 (O_985,N_9967,N_9823);
xor UO_986 (O_986,N_9915,N_9926);
nand UO_987 (O_987,N_9837,N_9969);
nand UO_988 (O_988,N_9919,N_9910);
xor UO_989 (O_989,N_9888,N_9848);
xnor UO_990 (O_990,N_9975,N_9954);
and UO_991 (O_991,N_9810,N_9952);
xnor UO_992 (O_992,N_9998,N_9820);
and UO_993 (O_993,N_9926,N_9977);
nand UO_994 (O_994,N_9826,N_9811);
xor UO_995 (O_995,N_9845,N_9894);
or UO_996 (O_996,N_9813,N_9807);
xnor UO_997 (O_997,N_9888,N_9934);
xnor UO_998 (O_998,N_9908,N_9963);
xnor UO_999 (O_999,N_9951,N_9835);
nand UO_1000 (O_1000,N_9821,N_9807);
nand UO_1001 (O_1001,N_9914,N_9837);
xor UO_1002 (O_1002,N_9980,N_9835);
or UO_1003 (O_1003,N_9931,N_9833);
and UO_1004 (O_1004,N_9971,N_9874);
nor UO_1005 (O_1005,N_9992,N_9910);
and UO_1006 (O_1006,N_9962,N_9819);
and UO_1007 (O_1007,N_9809,N_9924);
xnor UO_1008 (O_1008,N_9849,N_9801);
or UO_1009 (O_1009,N_9890,N_9956);
nor UO_1010 (O_1010,N_9822,N_9882);
and UO_1011 (O_1011,N_9815,N_9960);
or UO_1012 (O_1012,N_9940,N_9806);
xor UO_1013 (O_1013,N_9800,N_9956);
and UO_1014 (O_1014,N_9809,N_9833);
and UO_1015 (O_1015,N_9815,N_9809);
and UO_1016 (O_1016,N_9870,N_9922);
xor UO_1017 (O_1017,N_9955,N_9975);
or UO_1018 (O_1018,N_9996,N_9948);
nor UO_1019 (O_1019,N_9930,N_9839);
nor UO_1020 (O_1020,N_9868,N_9925);
or UO_1021 (O_1021,N_9894,N_9968);
or UO_1022 (O_1022,N_9911,N_9975);
nand UO_1023 (O_1023,N_9833,N_9999);
and UO_1024 (O_1024,N_9814,N_9816);
xnor UO_1025 (O_1025,N_9902,N_9986);
nand UO_1026 (O_1026,N_9934,N_9891);
nand UO_1027 (O_1027,N_9991,N_9914);
nand UO_1028 (O_1028,N_9934,N_9970);
nor UO_1029 (O_1029,N_9920,N_9848);
and UO_1030 (O_1030,N_9967,N_9802);
nand UO_1031 (O_1031,N_9803,N_9816);
or UO_1032 (O_1032,N_9818,N_9936);
nand UO_1033 (O_1033,N_9835,N_9830);
nor UO_1034 (O_1034,N_9936,N_9805);
nor UO_1035 (O_1035,N_9944,N_9873);
or UO_1036 (O_1036,N_9984,N_9879);
and UO_1037 (O_1037,N_9855,N_9988);
xor UO_1038 (O_1038,N_9851,N_9908);
and UO_1039 (O_1039,N_9883,N_9949);
and UO_1040 (O_1040,N_9803,N_9955);
nor UO_1041 (O_1041,N_9892,N_9927);
or UO_1042 (O_1042,N_9840,N_9921);
and UO_1043 (O_1043,N_9883,N_9987);
nor UO_1044 (O_1044,N_9809,N_9888);
nand UO_1045 (O_1045,N_9801,N_9961);
nand UO_1046 (O_1046,N_9943,N_9901);
xnor UO_1047 (O_1047,N_9923,N_9889);
and UO_1048 (O_1048,N_9814,N_9807);
and UO_1049 (O_1049,N_9826,N_9976);
or UO_1050 (O_1050,N_9852,N_9937);
or UO_1051 (O_1051,N_9945,N_9828);
nor UO_1052 (O_1052,N_9960,N_9970);
and UO_1053 (O_1053,N_9872,N_9903);
and UO_1054 (O_1054,N_9917,N_9800);
nor UO_1055 (O_1055,N_9834,N_9927);
nand UO_1056 (O_1056,N_9867,N_9825);
or UO_1057 (O_1057,N_9820,N_9832);
nor UO_1058 (O_1058,N_9992,N_9976);
nand UO_1059 (O_1059,N_9931,N_9842);
or UO_1060 (O_1060,N_9950,N_9946);
xnor UO_1061 (O_1061,N_9860,N_9942);
and UO_1062 (O_1062,N_9886,N_9992);
or UO_1063 (O_1063,N_9941,N_9842);
xnor UO_1064 (O_1064,N_9881,N_9801);
or UO_1065 (O_1065,N_9904,N_9803);
nor UO_1066 (O_1066,N_9972,N_9948);
nor UO_1067 (O_1067,N_9972,N_9831);
xnor UO_1068 (O_1068,N_9983,N_9869);
and UO_1069 (O_1069,N_9853,N_9913);
nand UO_1070 (O_1070,N_9912,N_9943);
or UO_1071 (O_1071,N_9871,N_9913);
nor UO_1072 (O_1072,N_9800,N_9818);
or UO_1073 (O_1073,N_9899,N_9879);
and UO_1074 (O_1074,N_9840,N_9992);
nor UO_1075 (O_1075,N_9825,N_9839);
and UO_1076 (O_1076,N_9800,N_9933);
nor UO_1077 (O_1077,N_9870,N_9837);
xnor UO_1078 (O_1078,N_9816,N_9911);
nor UO_1079 (O_1079,N_9987,N_9894);
or UO_1080 (O_1080,N_9859,N_9920);
xor UO_1081 (O_1081,N_9838,N_9816);
nor UO_1082 (O_1082,N_9849,N_9951);
and UO_1083 (O_1083,N_9899,N_9801);
and UO_1084 (O_1084,N_9988,N_9999);
or UO_1085 (O_1085,N_9877,N_9952);
and UO_1086 (O_1086,N_9810,N_9879);
xor UO_1087 (O_1087,N_9826,N_9941);
nand UO_1088 (O_1088,N_9973,N_9835);
and UO_1089 (O_1089,N_9907,N_9926);
nor UO_1090 (O_1090,N_9988,N_9966);
and UO_1091 (O_1091,N_9808,N_9955);
xnor UO_1092 (O_1092,N_9859,N_9916);
nor UO_1093 (O_1093,N_9923,N_9900);
nand UO_1094 (O_1094,N_9994,N_9865);
xor UO_1095 (O_1095,N_9862,N_9999);
nor UO_1096 (O_1096,N_9823,N_9851);
nor UO_1097 (O_1097,N_9821,N_9948);
and UO_1098 (O_1098,N_9975,N_9934);
xnor UO_1099 (O_1099,N_9960,N_9839);
and UO_1100 (O_1100,N_9925,N_9893);
nor UO_1101 (O_1101,N_9832,N_9900);
nor UO_1102 (O_1102,N_9965,N_9907);
xnor UO_1103 (O_1103,N_9951,N_9867);
nor UO_1104 (O_1104,N_9875,N_9932);
and UO_1105 (O_1105,N_9997,N_9936);
nor UO_1106 (O_1106,N_9856,N_9932);
or UO_1107 (O_1107,N_9910,N_9980);
nor UO_1108 (O_1108,N_9816,N_9899);
nor UO_1109 (O_1109,N_9866,N_9948);
nand UO_1110 (O_1110,N_9973,N_9971);
nor UO_1111 (O_1111,N_9923,N_9914);
nor UO_1112 (O_1112,N_9912,N_9832);
or UO_1113 (O_1113,N_9916,N_9940);
nor UO_1114 (O_1114,N_9804,N_9992);
and UO_1115 (O_1115,N_9865,N_9981);
xnor UO_1116 (O_1116,N_9950,N_9945);
nand UO_1117 (O_1117,N_9857,N_9917);
or UO_1118 (O_1118,N_9904,N_9893);
xnor UO_1119 (O_1119,N_9976,N_9833);
or UO_1120 (O_1120,N_9835,N_9896);
nor UO_1121 (O_1121,N_9814,N_9989);
and UO_1122 (O_1122,N_9854,N_9857);
nor UO_1123 (O_1123,N_9991,N_9813);
nand UO_1124 (O_1124,N_9891,N_9926);
and UO_1125 (O_1125,N_9942,N_9906);
xnor UO_1126 (O_1126,N_9998,N_9952);
xor UO_1127 (O_1127,N_9911,N_9960);
xor UO_1128 (O_1128,N_9913,N_9961);
and UO_1129 (O_1129,N_9965,N_9960);
or UO_1130 (O_1130,N_9938,N_9956);
xnor UO_1131 (O_1131,N_9845,N_9824);
nand UO_1132 (O_1132,N_9849,N_9861);
or UO_1133 (O_1133,N_9864,N_9925);
or UO_1134 (O_1134,N_9860,N_9883);
and UO_1135 (O_1135,N_9938,N_9902);
and UO_1136 (O_1136,N_9965,N_9936);
and UO_1137 (O_1137,N_9900,N_9905);
or UO_1138 (O_1138,N_9991,N_9833);
or UO_1139 (O_1139,N_9909,N_9850);
xnor UO_1140 (O_1140,N_9997,N_9926);
and UO_1141 (O_1141,N_9846,N_9947);
and UO_1142 (O_1142,N_9941,N_9884);
and UO_1143 (O_1143,N_9931,N_9986);
xnor UO_1144 (O_1144,N_9877,N_9999);
nor UO_1145 (O_1145,N_9837,N_9829);
xor UO_1146 (O_1146,N_9880,N_9993);
xnor UO_1147 (O_1147,N_9989,N_9950);
and UO_1148 (O_1148,N_9833,N_9963);
or UO_1149 (O_1149,N_9873,N_9980);
and UO_1150 (O_1150,N_9986,N_9914);
or UO_1151 (O_1151,N_9922,N_9880);
nand UO_1152 (O_1152,N_9946,N_9893);
or UO_1153 (O_1153,N_9837,N_9853);
xor UO_1154 (O_1154,N_9899,N_9920);
nor UO_1155 (O_1155,N_9805,N_9882);
nand UO_1156 (O_1156,N_9852,N_9971);
and UO_1157 (O_1157,N_9851,N_9842);
nor UO_1158 (O_1158,N_9802,N_9918);
or UO_1159 (O_1159,N_9900,N_9985);
nand UO_1160 (O_1160,N_9914,N_9912);
nand UO_1161 (O_1161,N_9997,N_9927);
xor UO_1162 (O_1162,N_9960,N_9890);
xnor UO_1163 (O_1163,N_9885,N_9809);
or UO_1164 (O_1164,N_9886,N_9952);
nor UO_1165 (O_1165,N_9854,N_9926);
xor UO_1166 (O_1166,N_9991,N_9978);
nor UO_1167 (O_1167,N_9847,N_9898);
or UO_1168 (O_1168,N_9911,N_9811);
or UO_1169 (O_1169,N_9856,N_9803);
xor UO_1170 (O_1170,N_9951,N_9949);
nor UO_1171 (O_1171,N_9930,N_9934);
nand UO_1172 (O_1172,N_9898,N_9875);
nor UO_1173 (O_1173,N_9815,N_9997);
nand UO_1174 (O_1174,N_9883,N_9938);
and UO_1175 (O_1175,N_9933,N_9976);
xor UO_1176 (O_1176,N_9936,N_9850);
nand UO_1177 (O_1177,N_9808,N_9851);
and UO_1178 (O_1178,N_9907,N_9978);
nand UO_1179 (O_1179,N_9843,N_9927);
nor UO_1180 (O_1180,N_9837,N_9908);
or UO_1181 (O_1181,N_9915,N_9914);
nand UO_1182 (O_1182,N_9886,N_9849);
nand UO_1183 (O_1183,N_9995,N_9865);
nand UO_1184 (O_1184,N_9834,N_9956);
and UO_1185 (O_1185,N_9976,N_9801);
xnor UO_1186 (O_1186,N_9935,N_9832);
xnor UO_1187 (O_1187,N_9942,N_9989);
and UO_1188 (O_1188,N_9870,N_9975);
nor UO_1189 (O_1189,N_9921,N_9909);
and UO_1190 (O_1190,N_9978,N_9872);
and UO_1191 (O_1191,N_9845,N_9955);
nand UO_1192 (O_1192,N_9919,N_9961);
xnor UO_1193 (O_1193,N_9946,N_9824);
and UO_1194 (O_1194,N_9822,N_9948);
or UO_1195 (O_1195,N_9889,N_9911);
and UO_1196 (O_1196,N_9837,N_9884);
or UO_1197 (O_1197,N_9862,N_9995);
nand UO_1198 (O_1198,N_9842,N_9930);
and UO_1199 (O_1199,N_9849,N_9913);
nor UO_1200 (O_1200,N_9932,N_9891);
nor UO_1201 (O_1201,N_9954,N_9886);
nor UO_1202 (O_1202,N_9820,N_9834);
or UO_1203 (O_1203,N_9915,N_9895);
nand UO_1204 (O_1204,N_9987,N_9888);
and UO_1205 (O_1205,N_9875,N_9948);
nand UO_1206 (O_1206,N_9862,N_9946);
nor UO_1207 (O_1207,N_9894,N_9986);
xnor UO_1208 (O_1208,N_9922,N_9808);
nor UO_1209 (O_1209,N_9851,N_9903);
nor UO_1210 (O_1210,N_9962,N_9830);
xnor UO_1211 (O_1211,N_9850,N_9806);
xnor UO_1212 (O_1212,N_9861,N_9879);
or UO_1213 (O_1213,N_9894,N_9811);
nand UO_1214 (O_1214,N_9924,N_9846);
xnor UO_1215 (O_1215,N_9871,N_9813);
and UO_1216 (O_1216,N_9877,N_9987);
and UO_1217 (O_1217,N_9822,N_9888);
nand UO_1218 (O_1218,N_9829,N_9940);
nor UO_1219 (O_1219,N_9890,N_9988);
and UO_1220 (O_1220,N_9918,N_9945);
or UO_1221 (O_1221,N_9943,N_9818);
xnor UO_1222 (O_1222,N_9811,N_9964);
or UO_1223 (O_1223,N_9872,N_9928);
nand UO_1224 (O_1224,N_9971,N_9826);
nor UO_1225 (O_1225,N_9876,N_9878);
nor UO_1226 (O_1226,N_9979,N_9912);
and UO_1227 (O_1227,N_9918,N_9865);
nor UO_1228 (O_1228,N_9822,N_9997);
nor UO_1229 (O_1229,N_9816,N_9987);
nand UO_1230 (O_1230,N_9810,N_9902);
and UO_1231 (O_1231,N_9812,N_9846);
xnor UO_1232 (O_1232,N_9879,N_9851);
nor UO_1233 (O_1233,N_9920,N_9911);
nor UO_1234 (O_1234,N_9891,N_9882);
or UO_1235 (O_1235,N_9826,N_9945);
nand UO_1236 (O_1236,N_9866,N_9872);
xor UO_1237 (O_1237,N_9913,N_9996);
nand UO_1238 (O_1238,N_9957,N_9981);
nand UO_1239 (O_1239,N_9969,N_9954);
xnor UO_1240 (O_1240,N_9828,N_9800);
or UO_1241 (O_1241,N_9923,N_9810);
xor UO_1242 (O_1242,N_9836,N_9855);
xor UO_1243 (O_1243,N_9818,N_9998);
xnor UO_1244 (O_1244,N_9825,N_9810);
or UO_1245 (O_1245,N_9950,N_9916);
and UO_1246 (O_1246,N_9891,N_9901);
and UO_1247 (O_1247,N_9982,N_9807);
xnor UO_1248 (O_1248,N_9962,N_9906);
xnor UO_1249 (O_1249,N_9876,N_9885);
and UO_1250 (O_1250,N_9905,N_9836);
and UO_1251 (O_1251,N_9935,N_9903);
nand UO_1252 (O_1252,N_9958,N_9943);
nor UO_1253 (O_1253,N_9997,N_9878);
or UO_1254 (O_1254,N_9915,N_9802);
and UO_1255 (O_1255,N_9967,N_9816);
and UO_1256 (O_1256,N_9892,N_9874);
nand UO_1257 (O_1257,N_9914,N_9917);
and UO_1258 (O_1258,N_9806,N_9949);
nor UO_1259 (O_1259,N_9896,N_9900);
and UO_1260 (O_1260,N_9897,N_9872);
or UO_1261 (O_1261,N_9951,N_9954);
and UO_1262 (O_1262,N_9821,N_9933);
or UO_1263 (O_1263,N_9932,N_9996);
nor UO_1264 (O_1264,N_9842,N_9821);
nor UO_1265 (O_1265,N_9990,N_9883);
xor UO_1266 (O_1266,N_9810,N_9837);
xor UO_1267 (O_1267,N_9812,N_9914);
and UO_1268 (O_1268,N_9973,N_9968);
xnor UO_1269 (O_1269,N_9974,N_9882);
nor UO_1270 (O_1270,N_9902,N_9909);
nand UO_1271 (O_1271,N_9945,N_9895);
nand UO_1272 (O_1272,N_9874,N_9982);
and UO_1273 (O_1273,N_9980,N_9953);
xor UO_1274 (O_1274,N_9958,N_9997);
nand UO_1275 (O_1275,N_9815,N_9847);
or UO_1276 (O_1276,N_9930,N_9926);
or UO_1277 (O_1277,N_9931,N_9991);
and UO_1278 (O_1278,N_9873,N_9834);
nor UO_1279 (O_1279,N_9994,N_9906);
nand UO_1280 (O_1280,N_9957,N_9881);
nand UO_1281 (O_1281,N_9864,N_9943);
nor UO_1282 (O_1282,N_9987,N_9914);
or UO_1283 (O_1283,N_9918,N_9984);
or UO_1284 (O_1284,N_9964,N_9915);
and UO_1285 (O_1285,N_9953,N_9844);
xor UO_1286 (O_1286,N_9930,N_9836);
nand UO_1287 (O_1287,N_9968,N_9964);
and UO_1288 (O_1288,N_9850,N_9853);
nor UO_1289 (O_1289,N_9953,N_9872);
and UO_1290 (O_1290,N_9820,N_9807);
nor UO_1291 (O_1291,N_9947,N_9931);
or UO_1292 (O_1292,N_9957,N_9997);
nand UO_1293 (O_1293,N_9980,N_9845);
nor UO_1294 (O_1294,N_9853,N_9934);
nand UO_1295 (O_1295,N_9880,N_9857);
nand UO_1296 (O_1296,N_9822,N_9957);
and UO_1297 (O_1297,N_9937,N_9924);
and UO_1298 (O_1298,N_9803,N_9895);
xnor UO_1299 (O_1299,N_9967,N_9968);
nand UO_1300 (O_1300,N_9887,N_9861);
nor UO_1301 (O_1301,N_9983,N_9950);
nor UO_1302 (O_1302,N_9938,N_9977);
nand UO_1303 (O_1303,N_9862,N_9818);
and UO_1304 (O_1304,N_9935,N_9836);
or UO_1305 (O_1305,N_9802,N_9900);
nor UO_1306 (O_1306,N_9805,N_9918);
nand UO_1307 (O_1307,N_9815,N_9920);
and UO_1308 (O_1308,N_9973,N_9871);
xnor UO_1309 (O_1309,N_9973,N_9873);
xor UO_1310 (O_1310,N_9802,N_9980);
xor UO_1311 (O_1311,N_9942,N_9876);
xnor UO_1312 (O_1312,N_9859,N_9982);
nor UO_1313 (O_1313,N_9981,N_9940);
nand UO_1314 (O_1314,N_9815,N_9959);
nor UO_1315 (O_1315,N_9964,N_9807);
or UO_1316 (O_1316,N_9924,N_9975);
xnor UO_1317 (O_1317,N_9992,N_9912);
and UO_1318 (O_1318,N_9962,N_9981);
xnor UO_1319 (O_1319,N_9871,N_9879);
nand UO_1320 (O_1320,N_9879,N_9888);
nand UO_1321 (O_1321,N_9951,N_9840);
xnor UO_1322 (O_1322,N_9842,N_9854);
and UO_1323 (O_1323,N_9984,N_9894);
and UO_1324 (O_1324,N_9913,N_9899);
and UO_1325 (O_1325,N_9907,N_9949);
and UO_1326 (O_1326,N_9849,N_9979);
nand UO_1327 (O_1327,N_9951,N_9912);
and UO_1328 (O_1328,N_9842,N_9976);
nand UO_1329 (O_1329,N_9939,N_9910);
and UO_1330 (O_1330,N_9969,N_9928);
or UO_1331 (O_1331,N_9951,N_9817);
and UO_1332 (O_1332,N_9812,N_9824);
nor UO_1333 (O_1333,N_9916,N_9957);
and UO_1334 (O_1334,N_9895,N_9972);
and UO_1335 (O_1335,N_9972,N_9816);
nor UO_1336 (O_1336,N_9902,N_9847);
nand UO_1337 (O_1337,N_9868,N_9821);
nor UO_1338 (O_1338,N_9855,N_9965);
or UO_1339 (O_1339,N_9967,N_9990);
nand UO_1340 (O_1340,N_9920,N_9854);
or UO_1341 (O_1341,N_9939,N_9980);
and UO_1342 (O_1342,N_9826,N_9860);
or UO_1343 (O_1343,N_9856,N_9902);
nand UO_1344 (O_1344,N_9800,N_9930);
nand UO_1345 (O_1345,N_9848,N_9908);
nor UO_1346 (O_1346,N_9894,N_9856);
nor UO_1347 (O_1347,N_9878,N_9910);
or UO_1348 (O_1348,N_9962,N_9857);
xnor UO_1349 (O_1349,N_9899,N_9963);
and UO_1350 (O_1350,N_9908,N_9855);
xnor UO_1351 (O_1351,N_9842,N_9903);
nor UO_1352 (O_1352,N_9888,N_9974);
xnor UO_1353 (O_1353,N_9895,N_9864);
nor UO_1354 (O_1354,N_9805,N_9947);
or UO_1355 (O_1355,N_9918,N_9873);
nand UO_1356 (O_1356,N_9944,N_9891);
and UO_1357 (O_1357,N_9927,N_9996);
nor UO_1358 (O_1358,N_9893,N_9918);
nand UO_1359 (O_1359,N_9984,N_9983);
nor UO_1360 (O_1360,N_9865,N_9846);
nor UO_1361 (O_1361,N_9910,N_9920);
or UO_1362 (O_1362,N_9971,N_9892);
and UO_1363 (O_1363,N_9872,N_9849);
nor UO_1364 (O_1364,N_9938,N_9803);
nand UO_1365 (O_1365,N_9836,N_9901);
and UO_1366 (O_1366,N_9955,N_9880);
and UO_1367 (O_1367,N_9897,N_9849);
nor UO_1368 (O_1368,N_9915,N_9873);
nand UO_1369 (O_1369,N_9916,N_9956);
xor UO_1370 (O_1370,N_9911,N_9822);
and UO_1371 (O_1371,N_9823,N_9822);
nand UO_1372 (O_1372,N_9864,N_9854);
nor UO_1373 (O_1373,N_9987,N_9851);
nor UO_1374 (O_1374,N_9806,N_9990);
xnor UO_1375 (O_1375,N_9961,N_9959);
nand UO_1376 (O_1376,N_9876,N_9944);
nor UO_1377 (O_1377,N_9919,N_9841);
nor UO_1378 (O_1378,N_9875,N_9985);
nand UO_1379 (O_1379,N_9852,N_9990);
nor UO_1380 (O_1380,N_9910,N_9837);
and UO_1381 (O_1381,N_9966,N_9817);
nand UO_1382 (O_1382,N_9826,N_9939);
and UO_1383 (O_1383,N_9817,N_9802);
nor UO_1384 (O_1384,N_9831,N_9866);
nand UO_1385 (O_1385,N_9893,N_9853);
or UO_1386 (O_1386,N_9872,N_9973);
nand UO_1387 (O_1387,N_9968,N_9909);
nand UO_1388 (O_1388,N_9932,N_9928);
nand UO_1389 (O_1389,N_9958,N_9887);
and UO_1390 (O_1390,N_9856,N_9824);
nand UO_1391 (O_1391,N_9839,N_9991);
and UO_1392 (O_1392,N_9811,N_9834);
and UO_1393 (O_1393,N_9849,N_9997);
nor UO_1394 (O_1394,N_9810,N_9848);
xnor UO_1395 (O_1395,N_9902,N_9890);
xor UO_1396 (O_1396,N_9867,N_9897);
and UO_1397 (O_1397,N_9805,N_9952);
and UO_1398 (O_1398,N_9861,N_9899);
and UO_1399 (O_1399,N_9962,N_9943);
or UO_1400 (O_1400,N_9855,N_9887);
nor UO_1401 (O_1401,N_9892,N_9825);
or UO_1402 (O_1402,N_9995,N_9934);
nand UO_1403 (O_1403,N_9849,N_9863);
xor UO_1404 (O_1404,N_9884,N_9894);
nor UO_1405 (O_1405,N_9896,N_9904);
xor UO_1406 (O_1406,N_9801,N_9838);
nor UO_1407 (O_1407,N_9864,N_9934);
xnor UO_1408 (O_1408,N_9898,N_9914);
nand UO_1409 (O_1409,N_9907,N_9902);
nand UO_1410 (O_1410,N_9850,N_9863);
and UO_1411 (O_1411,N_9998,N_9867);
nor UO_1412 (O_1412,N_9852,N_9966);
xor UO_1413 (O_1413,N_9829,N_9836);
or UO_1414 (O_1414,N_9895,N_9811);
and UO_1415 (O_1415,N_9941,N_9982);
or UO_1416 (O_1416,N_9978,N_9869);
or UO_1417 (O_1417,N_9887,N_9809);
or UO_1418 (O_1418,N_9915,N_9948);
xor UO_1419 (O_1419,N_9871,N_9930);
nor UO_1420 (O_1420,N_9957,N_9879);
or UO_1421 (O_1421,N_9861,N_9834);
nor UO_1422 (O_1422,N_9960,N_9808);
nand UO_1423 (O_1423,N_9813,N_9931);
nand UO_1424 (O_1424,N_9980,N_9919);
and UO_1425 (O_1425,N_9862,N_9936);
xor UO_1426 (O_1426,N_9868,N_9893);
nand UO_1427 (O_1427,N_9830,N_9996);
or UO_1428 (O_1428,N_9809,N_9826);
and UO_1429 (O_1429,N_9871,N_9892);
and UO_1430 (O_1430,N_9895,N_9958);
or UO_1431 (O_1431,N_9940,N_9804);
xor UO_1432 (O_1432,N_9868,N_9840);
or UO_1433 (O_1433,N_9897,N_9805);
xnor UO_1434 (O_1434,N_9877,N_9960);
or UO_1435 (O_1435,N_9827,N_9866);
xor UO_1436 (O_1436,N_9923,N_9880);
xor UO_1437 (O_1437,N_9803,N_9973);
nand UO_1438 (O_1438,N_9847,N_9961);
xor UO_1439 (O_1439,N_9985,N_9947);
and UO_1440 (O_1440,N_9978,N_9846);
nor UO_1441 (O_1441,N_9932,N_9906);
and UO_1442 (O_1442,N_9860,N_9898);
and UO_1443 (O_1443,N_9934,N_9809);
xnor UO_1444 (O_1444,N_9938,N_9860);
nor UO_1445 (O_1445,N_9981,N_9886);
nand UO_1446 (O_1446,N_9855,N_9906);
or UO_1447 (O_1447,N_9988,N_9886);
or UO_1448 (O_1448,N_9965,N_9827);
and UO_1449 (O_1449,N_9871,N_9901);
nor UO_1450 (O_1450,N_9908,N_9927);
xor UO_1451 (O_1451,N_9888,N_9973);
or UO_1452 (O_1452,N_9999,N_9913);
nand UO_1453 (O_1453,N_9944,N_9963);
nand UO_1454 (O_1454,N_9862,N_9925);
and UO_1455 (O_1455,N_9946,N_9854);
and UO_1456 (O_1456,N_9867,N_9946);
nand UO_1457 (O_1457,N_9841,N_9832);
xor UO_1458 (O_1458,N_9998,N_9834);
nand UO_1459 (O_1459,N_9922,N_9862);
nand UO_1460 (O_1460,N_9869,N_9860);
nand UO_1461 (O_1461,N_9895,N_9814);
nand UO_1462 (O_1462,N_9900,N_9904);
and UO_1463 (O_1463,N_9913,N_9974);
nor UO_1464 (O_1464,N_9957,N_9906);
xor UO_1465 (O_1465,N_9952,N_9853);
or UO_1466 (O_1466,N_9884,N_9954);
nor UO_1467 (O_1467,N_9917,N_9876);
nand UO_1468 (O_1468,N_9967,N_9947);
nand UO_1469 (O_1469,N_9897,N_9845);
and UO_1470 (O_1470,N_9839,N_9935);
nor UO_1471 (O_1471,N_9921,N_9945);
and UO_1472 (O_1472,N_9897,N_9868);
nor UO_1473 (O_1473,N_9860,N_9927);
xnor UO_1474 (O_1474,N_9937,N_9986);
and UO_1475 (O_1475,N_9826,N_9891);
nand UO_1476 (O_1476,N_9852,N_9916);
xnor UO_1477 (O_1477,N_9995,N_9973);
xor UO_1478 (O_1478,N_9856,N_9892);
and UO_1479 (O_1479,N_9812,N_9887);
nor UO_1480 (O_1480,N_9986,N_9990);
nor UO_1481 (O_1481,N_9877,N_9996);
xor UO_1482 (O_1482,N_9867,N_9964);
nor UO_1483 (O_1483,N_9877,N_9932);
nor UO_1484 (O_1484,N_9869,N_9866);
or UO_1485 (O_1485,N_9927,N_9844);
nand UO_1486 (O_1486,N_9863,N_9934);
xnor UO_1487 (O_1487,N_9807,N_9869);
or UO_1488 (O_1488,N_9839,N_9945);
nand UO_1489 (O_1489,N_9803,N_9843);
nor UO_1490 (O_1490,N_9944,N_9850);
nand UO_1491 (O_1491,N_9923,N_9937);
and UO_1492 (O_1492,N_9966,N_9823);
nand UO_1493 (O_1493,N_9847,N_9841);
xnor UO_1494 (O_1494,N_9912,N_9935);
nor UO_1495 (O_1495,N_9887,N_9832);
and UO_1496 (O_1496,N_9978,N_9875);
and UO_1497 (O_1497,N_9892,N_9960);
and UO_1498 (O_1498,N_9859,N_9883);
or UO_1499 (O_1499,N_9985,N_9891);
endmodule