module basic_2000_20000_2500_40_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
or U0 (N_0,In_1426,In_139);
xor U1 (N_1,In_1364,In_1370);
xor U2 (N_2,In_1732,In_754);
or U3 (N_3,In_677,In_214);
nand U4 (N_4,In_1022,In_1693);
nor U5 (N_5,In_1915,In_1388);
or U6 (N_6,In_380,In_1583);
nor U7 (N_7,In_892,In_1139);
and U8 (N_8,In_1104,In_982);
nor U9 (N_9,In_596,In_1911);
nand U10 (N_10,In_226,In_104);
nand U11 (N_11,In_827,In_1475);
or U12 (N_12,In_1895,In_366);
or U13 (N_13,In_1562,In_419);
xor U14 (N_14,In_1770,In_1215);
xor U15 (N_15,In_692,In_1571);
nor U16 (N_16,In_1170,In_926);
or U17 (N_17,In_1643,In_937);
nand U18 (N_18,In_415,In_1821);
or U19 (N_19,In_1203,In_138);
xnor U20 (N_20,In_1691,In_1406);
nor U21 (N_21,In_963,In_1809);
and U22 (N_22,In_164,In_494);
and U23 (N_23,In_1570,In_433);
xor U24 (N_24,In_432,In_1260);
nor U25 (N_25,In_1673,In_134);
nor U26 (N_26,In_1187,In_64);
xor U27 (N_27,In_377,In_72);
nor U28 (N_28,In_1578,In_1630);
nor U29 (N_29,In_1354,In_1361);
nor U30 (N_30,In_1748,In_1652);
nor U31 (N_31,In_1950,In_1917);
or U32 (N_32,In_94,In_1649);
nor U33 (N_33,In_956,In_365);
xor U34 (N_34,In_586,In_811);
and U35 (N_35,In_1700,In_817);
and U36 (N_36,In_866,In_255);
or U37 (N_37,In_1306,In_1900);
xnor U38 (N_38,In_1541,In_1112);
nor U39 (N_39,In_1314,In_1898);
nand U40 (N_40,In_587,In_24);
nor U41 (N_41,In_1269,In_742);
or U42 (N_42,In_1471,In_1461);
or U43 (N_43,In_1702,In_1101);
nand U44 (N_44,In_1189,In_324);
or U45 (N_45,In_484,In_1538);
nor U46 (N_46,In_805,In_1865);
xor U47 (N_47,In_514,In_573);
and U48 (N_48,In_1252,In_1226);
and U49 (N_49,In_1177,In_710);
nor U50 (N_50,In_397,In_37);
or U51 (N_51,In_853,In_644);
xnor U52 (N_52,In_160,In_1337);
or U53 (N_53,In_1443,In_1543);
or U54 (N_54,In_229,In_1517);
xor U55 (N_55,In_1592,In_1730);
nand U56 (N_56,In_442,In_955);
nor U57 (N_57,In_1333,In_1676);
xnor U58 (N_58,In_1131,In_1457);
nor U59 (N_59,In_1942,In_1540);
nand U60 (N_60,In_1885,In_1612);
nor U61 (N_61,In_1875,In_527);
xnor U62 (N_62,In_962,In_1175);
or U63 (N_63,In_815,In_364);
and U64 (N_64,In_1497,In_1739);
and U65 (N_65,In_253,In_283);
and U66 (N_66,In_1125,In_1546);
nand U67 (N_67,In_1358,In_1587);
nand U68 (N_68,In_719,In_763);
or U69 (N_69,In_554,In_1931);
nor U70 (N_70,In_947,In_1986);
nor U71 (N_71,In_1282,In_661);
nor U72 (N_72,In_562,In_907);
nor U73 (N_73,In_898,In_1347);
and U74 (N_74,In_839,In_1514);
nor U75 (N_75,In_1864,In_1644);
nand U76 (N_76,In_553,In_1262);
or U77 (N_77,In_949,In_1647);
and U78 (N_78,In_784,In_462);
nand U79 (N_79,In_86,In_518);
xnor U80 (N_80,In_1007,In_1486);
xnor U81 (N_81,In_1180,In_1281);
and U82 (N_82,In_1901,In_870);
nand U83 (N_83,In_471,In_1965);
nor U84 (N_84,In_1648,In_589);
or U85 (N_85,In_943,In_1925);
nor U86 (N_86,In_837,In_1631);
xnor U87 (N_87,In_542,In_356);
nor U88 (N_88,In_808,In_1485);
or U89 (N_89,In_656,In_549);
nand U90 (N_90,In_1329,In_386);
xnor U91 (N_91,In_1808,In_888);
or U92 (N_92,In_939,In_1929);
nor U93 (N_93,In_1659,In_938);
nand U94 (N_94,In_1529,In_1653);
xnor U95 (N_95,In_909,In_1696);
and U96 (N_96,In_1431,In_1108);
nand U97 (N_97,In_87,In_1709);
and U98 (N_98,In_1382,In_1615);
xor U99 (N_99,In_1403,In_1103);
or U100 (N_100,In_1427,In_1919);
and U101 (N_101,In_479,In_18);
xor U102 (N_102,In_544,In_502);
xor U103 (N_103,In_1147,In_1816);
nor U104 (N_104,In_1316,In_806);
nand U105 (N_105,In_819,In_388);
nor U106 (N_106,In_1122,In_584);
nand U107 (N_107,In_749,In_338);
and U108 (N_108,In_1502,In_1760);
nor U109 (N_109,In_5,In_1729);
nand U110 (N_110,In_1810,In_1544);
or U111 (N_111,In_1555,In_721);
nor U112 (N_112,In_1725,In_1014);
nand U113 (N_113,In_192,In_1);
xor U114 (N_114,In_895,In_883);
nor U115 (N_115,In_740,In_430);
nand U116 (N_116,In_1363,In_531);
nand U117 (N_117,In_1060,In_1258);
nand U118 (N_118,In_1871,In_1671);
nor U119 (N_119,In_1876,In_1339);
nand U120 (N_120,In_950,In_1073);
or U121 (N_121,In_941,In_410);
or U122 (N_122,In_1505,In_1684);
nand U123 (N_123,In_463,In_492);
or U124 (N_124,In_1241,In_1307);
nand U125 (N_125,In_1407,In_1928);
or U126 (N_126,In_290,In_1651);
xor U127 (N_127,In_363,In_355);
xnor U128 (N_128,In_450,In_602);
or U129 (N_129,In_280,In_1656);
nor U130 (N_130,In_474,In_1952);
nor U131 (N_131,In_731,In_796);
xnor U132 (N_132,In_1920,In_137);
xnor U133 (N_133,In_15,In_1657);
nor U134 (N_134,In_1229,In_1195);
or U135 (N_135,In_143,In_406);
nand U136 (N_136,In_1371,In_12);
and U137 (N_137,In_1141,In_159);
or U138 (N_138,In_974,In_1528);
nand U139 (N_139,In_966,In_1111);
nor U140 (N_140,In_268,In_1254);
nand U141 (N_141,In_1133,In_257);
xnor U142 (N_142,In_294,In_1736);
nand U143 (N_143,In_1313,In_1698);
or U144 (N_144,In_1627,In_1588);
nor U145 (N_145,In_263,In_1510);
nand U146 (N_146,In_597,In_1897);
and U147 (N_147,In_653,In_1123);
nor U148 (N_148,In_1896,In_266);
nor U149 (N_149,In_1604,In_551);
nor U150 (N_150,In_1420,In_720);
or U151 (N_151,In_900,In_1397);
nor U152 (N_152,In_1172,In_389);
nor U153 (N_153,In_110,In_967);
xnor U154 (N_154,In_1513,In_603);
and U155 (N_155,In_336,In_795);
nand U156 (N_156,In_1597,In_67);
or U157 (N_157,In_858,In_121);
xnor U158 (N_158,In_964,In_1899);
nand U159 (N_159,In_716,In_1609);
nor U160 (N_160,In_1550,In_256);
nor U161 (N_161,In_337,In_1413);
and U162 (N_162,In_912,In_733);
nand U163 (N_163,In_384,In_609);
and U164 (N_164,In_1954,In_1688);
xnor U165 (N_165,In_605,In_1704);
xor U166 (N_166,In_833,In_1741);
nand U167 (N_167,In_759,In_113);
nor U168 (N_168,In_198,In_259);
nand U169 (N_169,In_1309,In_427);
or U170 (N_170,In_1018,In_534);
and U171 (N_171,In_1381,In_1573);
or U172 (N_172,In_1466,In_1994);
nor U173 (N_173,In_730,In_1048);
and U174 (N_174,In_1375,In_131);
xnor U175 (N_175,In_770,In_243);
xor U176 (N_176,In_155,In_92);
or U177 (N_177,In_150,In_1474);
or U178 (N_178,In_979,In_1149);
nand U179 (N_179,In_687,In_845);
and U180 (N_180,In_439,In_1489);
xor U181 (N_181,In_1107,In_1763);
or U182 (N_182,In_101,In_1146);
or U183 (N_183,In_1166,In_1286);
nor U184 (N_184,In_1839,In_798);
xnor U185 (N_185,In_572,In_591);
and U186 (N_186,In_488,In_1065);
nand U187 (N_187,In_1368,In_1251);
xor U188 (N_188,In_1212,In_1710);
or U189 (N_189,In_1047,In_297);
nand U190 (N_190,In_1798,In_1357);
or U191 (N_191,In_1490,In_1789);
and U192 (N_192,In_655,In_623);
or U193 (N_193,In_1178,In_832);
nor U194 (N_194,In_915,In_404);
xor U195 (N_195,In_485,In_1584);
xor U196 (N_196,In_891,In_750);
xnor U197 (N_197,In_1345,In_1914);
nor U198 (N_198,In_1625,In_1138);
nand U199 (N_199,In_896,In_714);
xnor U200 (N_200,In_1677,In_411);
nand U201 (N_201,In_3,In_456);
nor U202 (N_202,In_1465,In_1365);
nor U203 (N_203,In_287,In_882);
and U204 (N_204,In_1311,In_1767);
and U205 (N_205,In_1995,In_973);
nand U206 (N_206,In_1744,In_1522);
or U207 (N_207,In_535,In_508);
xor U208 (N_208,In_1015,In_868);
nand U209 (N_209,In_1068,In_333);
xor U210 (N_210,In_948,In_807);
or U211 (N_211,In_1072,In_1854);
nor U212 (N_212,In_1479,In_913);
and U213 (N_213,In_1790,In_1873);
or U214 (N_214,In_599,In_1967);
and U215 (N_215,In_959,In_1672);
nor U216 (N_216,In_1569,In_1038);
nand U217 (N_217,In_100,In_580);
xor U218 (N_218,In_1416,In_1932);
and U219 (N_219,In_1784,In_1830);
or U220 (N_220,In_626,In_393);
xor U221 (N_221,In_855,In_1011);
nor U222 (N_222,In_395,In_678);
nand U223 (N_223,In_1738,In_1705);
and U224 (N_224,In_1781,In_1992);
nand U225 (N_225,In_620,In_1591);
nor U226 (N_226,In_398,In_762);
xor U227 (N_227,In_1987,In_307);
or U228 (N_228,In_842,In_1442);
nor U229 (N_229,In_249,In_322);
nand U230 (N_230,In_1655,In_771);
nand U231 (N_231,In_1728,In_1113);
xnor U232 (N_232,In_107,In_1859);
or U233 (N_233,In_169,In_1521);
xnor U234 (N_234,In_1988,In_1835);
nand U235 (N_235,In_616,In_1795);
and U236 (N_236,In_752,In_505);
xnor U237 (N_237,In_594,In_1083);
nand U238 (N_238,In_1678,In_766);
nand U239 (N_239,In_765,In_1266);
or U240 (N_240,In_934,In_717);
and U241 (N_241,In_315,In_124);
nor U242 (N_242,In_1686,In_1318);
nor U243 (N_243,In_1059,In_940);
and U244 (N_244,In_1091,In_1878);
and U245 (N_245,In_1579,In_417);
xnor U246 (N_246,In_455,In_1006);
and U247 (N_247,In_1974,In_1126);
xor U248 (N_248,In_1613,In_1747);
or U249 (N_249,In_1405,In_1848);
or U250 (N_250,In_308,In_179);
and U251 (N_251,In_1909,In_99);
nor U252 (N_252,In_206,In_1893);
nand U253 (N_253,In_516,In_1323);
nor U254 (N_254,In_666,In_250);
nand U255 (N_255,In_914,In_1167);
xnor U256 (N_256,In_558,In_787);
and U257 (N_257,In_1850,In_1445);
or U258 (N_258,In_1908,In_1500);
nand U259 (N_259,In_1356,In_693);
and U260 (N_260,In_1483,In_1844);
nand U261 (N_261,In_515,In_241);
xnor U262 (N_262,In_303,In_1979);
xnor U263 (N_263,In_1906,In_1135);
nand U264 (N_264,In_1636,In_1774);
or U265 (N_265,In_537,In_1983);
and U266 (N_266,In_886,In_123);
xor U267 (N_267,In_1183,In_295);
and U268 (N_268,In_557,In_202);
nor U269 (N_269,In_208,In_781);
and U270 (N_270,In_893,In_1089);
nor U271 (N_271,In_353,In_985);
xor U272 (N_272,In_1496,In_185);
and U273 (N_273,In_854,In_1826);
or U274 (N_274,In_1359,In_60);
or U275 (N_275,In_451,In_1937);
nand U276 (N_276,In_1157,In_1423);
and U277 (N_277,In_718,In_1338);
nor U278 (N_278,In_1837,In_1295);
nor U279 (N_279,In_1595,In_538);
nand U280 (N_280,In_1629,In_1322);
and U281 (N_281,In_239,In_1076);
and U282 (N_282,In_16,In_1594);
nand U283 (N_283,In_1294,In_713);
or U284 (N_284,In_1945,In_680);
or U285 (N_285,In_1412,In_299);
xnor U286 (N_286,In_1163,In_1953);
nand U287 (N_287,In_828,In_1803);
nor U288 (N_288,In_316,In_1196);
xor U289 (N_289,In_988,In_1634);
nor U290 (N_290,In_1389,In_55);
nand U291 (N_291,In_651,In_585);
nand U292 (N_292,In_1030,In_1096);
nor U293 (N_293,In_311,In_598);
nor U294 (N_294,In_35,In_1255);
or U295 (N_295,In_513,In_1581);
and U296 (N_296,In_1504,In_401);
nand U297 (N_297,In_1956,In_1161);
nand U298 (N_298,In_23,In_180);
or U299 (N_299,In_1280,In_1831);
xnor U300 (N_300,In_894,In_1793);
nor U301 (N_301,In_235,In_446);
or U302 (N_302,In_77,In_1086);
nand U303 (N_303,In_997,In_1626);
nand U304 (N_304,In_1257,In_753);
xor U305 (N_305,In_1754,In_768);
nand U306 (N_306,In_1981,In_1088);
or U307 (N_307,In_119,In_744);
nor U308 (N_308,In_650,In_1780);
nand U309 (N_309,In_539,In_619);
xnor U310 (N_310,In_617,In_234);
or U311 (N_311,In_1300,In_1176);
and U312 (N_312,In_359,In_989);
and U313 (N_313,In_588,In_218);
nor U314 (N_314,In_1058,In_1114);
nor U315 (N_315,In_747,In_1317);
and U316 (N_316,In_385,In_4);
and U317 (N_317,In_1436,In_372);
or U318 (N_318,In_1325,In_178);
and U319 (N_319,In_1775,In_812);
and U320 (N_320,In_1127,In_458);
nor U321 (N_321,In_1327,In_1548);
or U322 (N_322,In_167,In_1978);
nor U323 (N_323,In_1998,In_1777);
or U324 (N_324,In_1033,In_1962);
xnor U325 (N_325,In_304,In_1828);
xor U326 (N_326,In_1236,In_1005);
nand U327 (N_327,In_210,In_567);
nand U328 (N_328,In_1616,In_1886);
or U329 (N_329,In_215,In_1075);
xor U330 (N_330,In_40,In_431);
nand U331 (N_331,In_1418,In_1002);
and U332 (N_332,In_1285,In_88);
nand U333 (N_333,In_165,In_1223);
and U334 (N_334,In_1745,In_200);
nand U335 (N_335,In_1063,In_157);
xor U336 (N_336,In_672,In_1256);
nand U337 (N_337,In_663,In_1969);
or U338 (N_338,In_769,In_457);
or U339 (N_339,In_277,In_1824);
nand U340 (N_340,In_258,In_1362);
nand U341 (N_341,In_1145,In_305);
xor U342 (N_342,In_1439,In_1444);
xnor U343 (N_343,In_212,In_646);
xnor U344 (N_344,In_822,In_32);
and U345 (N_345,In_135,In_595);
xnor U346 (N_346,In_657,In_449);
xor U347 (N_347,In_296,In_203);
nor U348 (N_348,In_1348,In_1605);
nor U349 (N_349,In_1235,In_1305);
xnor U350 (N_350,In_1207,In_608);
xor U351 (N_351,In_1585,In_418);
and U352 (N_352,In_830,In_47);
nor U353 (N_353,In_376,In_1293);
nand U354 (N_354,In_1185,In_615);
or U355 (N_355,In_1851,In_50);
nand U356 (N_356,In_379,In_618);
nor U357 (N_357,In_470,In_1438);
nand U358 (N_358,In_130,In_635);
nor U359 (N_359,In_8,In_1695);
or U360 (N_360,In_510,In_1391);
xor U361 (N_361,In_676,In_865);
or U362 (N_362,In_96,In_901);
nor U363 (N_363,In_671,In_1124);
or U364 (N_364,In_739,In_785);
xnor U365 (N_365,In_320,In_1913);
nand U366 (N_366,In_1884,In_1755);
nand U367 (N_367,In_319,In_1572);
and U368 (N_368,In_339,In_1128);
xor U369 (N_369,In_629,In_496);
nor U370 (N_370,In_1949,In_70);
nor U371 (N_371,In_276,In_1031);
nor U372 (N_372,In_1610,In_610);
nand U373 (N_373,In_141,In_1542);
xor U374 (N_374,In_1624,In_1353);
and U375 (N_375,In_1188,In_1503);
nand U376 (N_376,In_1301,In_528);
nor U377 (N_377,In_1319,In_699);
nand U378 (N_378,In_1401,In_84);
or U379 (N_379,In_1843,In_467);
xnor U380 (N_380,In_162,In_1296);
or U381 (N_381,In_1246,In_935);
nor U382 (N_382,In_148,In_525);
and U383 (N_383,In_285,In_550);
nand U384 (N_384,In_1202,In_1463);
or U385 (N_385,In_1586,In_387);
or U386 (N_386,In_1669,In_1882);
nand U387 (N_387,In_1692,In_1726);
xnor U388 (N_388,In_1742,In_1263);
nor U389 (N_389,In_523,In_209);
xor U390 (N_390,In_59,In_1576);
or U391 (N_391,In_354,In_607);
and U392 (N_392,In_936,In_1057);
nor U393 (N_393,In_899,In_278);
and U394 (N_394,In_1452,In_1746);
nor U395 (N_395,In_122,In_105);
and U396 (N_396,In_975,In_66);
and U397 (N_397,In_1193,In_682);
nand U398 (N_398,In_480,In_62);
or U399 (N_399,In_1640,In_1298);
and U400 (N_400,In_1240,In_1469);
xor U401 (N_401,In_13,In_816);
and U402 (N_402,In_673,In_1087);
nand U403 (N_403,In_1666,In_1055);
or U404 (N_404,In_1043,In_1472);
and U405 (N_405,In_1972,In_1819);
and U406 (N_406,In_746,In_264);
and U407 (N_407,In_625,In_503);
xnor U408 (N_408,In_288,In_1476);
nand U409 (N_409,In_686,In_660);
or U410 (N_410,In_340,In_1756);
nor U411 (N_411,In_325,In_244);
xor U412 (N_412,In_1247,In_772);
and U413 (N_413,In_126,In_1303);
or U414 (N_414,In_1239,In_1010);
or U415 (N_415,In_1923,In_97);
and U416 (N_416,In_1097,In_345);
and U417 (N_417,In_1737,In_1182);
nor U418 (N_418,In_1130,In_1102);
nand U419 (N_419,In_761,In_1894);
and U420 (N_420,In_791,In_343);
and U421 (N_421,In_1703,In_1567);
and U422 (N_422,In_521,In_1551);
xnor U423 (N_423,In_91,In_413);
nor U424 (N_424,In_48,In_1685);
xnor U425 (N_425,In_1797,In_1140);
and U426 (N_426,In_22,In_416);
xor U427 (N_427,In_946,In_78);
and U428 (N_428,In_929,In_6);
or U429 (N_429,In_1155,In_631);
nand U430 (N_430,In_568,In_383);
nor U431 (N_431,In_1706,In_1200);
nand U432 (N_432,In_932,In_927);
nand U433 (N_433,In_1811,In_1186);
nor U434 (N_434,In_1874,In_944);
xnor U435 (N_435,In_593,In_1424);
or U436 (N_436,In_1951,In_374);
nand U437 (N_437,In_1233,In_1197);
or U438 (N_438,In_1532,In_1805);
and U439 (N_439,In_640,In_1759);
nand U440 (N_440,In_286,In_1017);
xnor U441 (N_441,In_1042,In_1752);
and U442 (N_442,In_228,In_151);
nand U443 (N_443,In_1454,In_1171);
nor U444 (N_444,In_1034,In_756);
and U445 (N_445,In_1430,In_403);
nand U446 (N_446,In_1079,In_662);
or U447 (N_447,In_1715,In_889);
nor U448 (N_448,In_1720,In_79);
nor U449 (N_449,In_426,In_689);
xor U450 (N_450,In_146,In_1536);
and U451 (N_451,In_543,In_261);
nor U452 (N_452,In_63,In_362);
or U453 (N_453,In_1531,In_1001);
or U454 (N_454,In_1515,In_39);
nand U455 (N_455,In_399,In_1922);
and U456 (N_456,In_1066,In_1115);
nand U457 (N_457,In_924,In_1619);
xor U458 (N_458,In_1813,In_98);
nand U459 (N_459,In_983,In_641);
and U460 (N_460,In_466,In_1734);
xor U461 (N_461,In_1907,In_1404);
nand U462 (N_462,In_852,In_1159);
and U463 (N_463,In_802,In_957);
xnor U464 (N_464,In_1971,In_1267);
and U465 (N_465,In_1132,In_792);
xor U466 (N_466,In_1872,In_1053);
nor U467 (N_467,In_1862,In_1376);
nor U468 (N_468,In_701,In_1346);
nor U469 (N_469,In_443,In_272);
nand U470 (N_470,In_1209,In_1456);
xor U471 (N_471,In_487,In_321);
nand U472 (N_472,In_27,In_1041);
nand U473 (N_473,In_1930,In_201);
nand U474 (N_474,In_563,In_350);
or U475 (N_475,In_423,In_526);
nor U476 (N_476,In_846,In_1451);
or U477 (N_477,In_887,In_820);
nand U478 (N_478,In_506,In_1230);
nor U479 (N_479,In_1330,In_880);
nand U480 (N_480,In_1462,In_1153);
nor U481 (N_481,In_1121,In_1259);
xnor U482 (N_482,In_1682,In_996);
and U483 (N_483,In_1411,In_1284);
xnor U484 (N_484,In_724,In_65);
nand U485 (N_485,In_1535,In_1044);
nor U486 (N_486,In_483,In_630);
nor U487 (N_487,In_1966,In_1563);
xor U488 (N_488,In_81,In_981);
and U489 (N_489,In_778,In_703);
nand U490 (N_490,In_1869,In_327);
and U491 (N_491,In_1557,In_194);
nand U492 (N_492,In_237,In_1482);
and U493 (N_493,In_738,In_1796);
xnor U494 (N_494,In_574,In_649);
nand U495 (N_495,In_783,In_1310);
nor U496 (N_496,In_1632,In_1735);
nand U497 (N_497,In_1164,In_755);
nand U498 (N_498,In_1879,In_972);
xor U499 (N_499,In_519,In_1350);
xnor U500 (N_500,In_153,In_369);
or U501 (N_501,In_472,In_933);
nand U502 (N_502,In_1812,In_44);
or U503 (N_503,In_357,In_1028);
nor U504 (N_504,In_378,In_848);
and U505 (N_505,In_844,In_1665);
nor U506 (N_506,N_205,In_1437);
nand U507 (N_507,N_50,In_166);
nor U508 (N_508,In_1109,N_112);
and U509 (N_509,N_270,In_1880);
nand U510 (N_510,In_1667,N_34);
nand U511 (N_511,In_547,In_1464);
xor U512 (N_512,N_232,In_637);
xor U513 (N_513,In_1392,In_190);
or U514 (N_514,In_1921,N_369);
or U515 (N_515,N_370,In_1600);
xnor U516 (N_516,In_529,In_628);
nand U517 (N_517,In_829,In_1650);
xnor U518 (N_518,In_634,In_33);
xnor U519 (N_519,N_374,N_215);
nor U520 (N_520,In_329,In_309);
nor U521 (N_521,In_438,In_232);
nand U522 (N_522,In_632,In_1094);
and U523 (N_523,In_1646,In_590);
and U524 (N_524,In_1184,In_332);
nor U525 (N_525,N_365,In_112);
nor U526 (N_526,In_1023,In_1621);
nor U527 (N_527,In_368,In_1846);
nor U528 (N_528,In_878,N_161);
xnor U529 (N_529,In_1589,In_511);
nor U530 (N_530,In_318,In_1518);
and U531 (N_531,N_28,In_1237);
or U532 (N_532,In_144,In_1393);
xor U533 (N_533,In_1198,N_354);
and U534 (N_534,In_548,N_337);
nand U535 (N_535,In_712,N_52);
and U536 (N_536,In_220,N_21);
xor U537 (N_537,In_961,In_1941);
or U538 (N_538,In_1421,In_1334);
nor U539 (N_539,In_1783,In_421);
nor U540 (N_540,N_158,N_139);
xor U541 (N_541,In_1008,In_1792);
nand U542 (N_542,In_1487,In_1045);
nand U543 (N_543,N_170,In_1374);
xor U544 (N_544,In_330,In_1387);
xor U545 (N_545,In_1225,N_96);
xnor U546 (N_546,N_144,In_1106);
nand U547 (N_547,N_276,N_193);
or U548 (N_548,N_198,In_813);
nand U549 (N_549,N_203,In_270);
and U550 (N_550,In_1989,In_1516);
xnor U551 (N_551,In_556,In_265);
nand U552 (N_552,In_642,In_1355);
nor U553 (N_553,N_388,In_1287);
or U554 (N_554,In_358,N_136);
xnor U555 (N_555,N_62,In_1787);
nor U556 (N_556,In_1208,In_1369);
or U557 (N_557,In_262,In_1993);
and U558 (N_558,N_49,In_953);
nor U559 (N_559,N_386,In_1757);
and U560 (N_560,In_1867,In_1292);
nor U561 (N_561,In_582,N_449);
nand U562 (N_562,N_48,In_1332);
or U563 (N_563,In_1791,In_500);
nor U564 (N_564,In_873,In_1838);
and U565 (N_565,In_1856,In_306);
xnor U566 (N_566,N_95,In_434);
or U567 (N_567,N_404,In_810);
xnor U568 (N_568,In_776,In_1156);
nand U569 (N_569,In_1224,In_903);
nand U570 (N_570,In_1249,N_181);
or U571 (N_571,In_1694,In_1519);
nand U572 (N_572,In_847,N_478);
nand U573 (N_573,In_1933,N_182);
or U574 (N_574,N_429,N_145);
nor U575 (N_575,N_406,N_255);
nand U576 (N_576,In_1806,In_1003);
or U577 (N_577,In_669,In_1771);
and U578 (N_578,N_278,N_290);
or U579 (N_579,In_902,In_25);
xnor U580 (N_580,N_20,In_1385);
nor U581 (N_581,In_1642,In_11);
xnor U582 (N_582,N_173,N_243);
or U583 (N_583,N_338,In_1577);
nand U584 (N_584,N_199,In_1414);
xor U585 (N_585,In_222,In_1975);
xor U586 (N_586,In_561,In_1165);
nand U587 (N_587,In_181,N_26);
nor U588 (N_588,N_77,In_274);
and U589 (N_589,In_1491,N_111);
or U590 (N_590,In_723,N_272);
or U591 (N_591,In_1459,In_93);
and U592 (N_592,In_726,N_367);
nor U593 (N_593,N_314,N_344);
nand U594 (N_594,In_1093,N_230);
nand U595 (N_595,In_61,In_1935);
nand U596 (N_596,N_175,N_47);
and U597 (N_597,In_251,In_424);
and U598 (N_598,In_874,In_1151);
nor U599 (N_599,In_835,In_136);
nor U600 (N_600,N_30,N_328);
or U601 (N_601,N_489,In_1384);
nand U602 (N_602,N_248,In_774);
or U603 (N_603,In_1697,N_398);
or U604 (N_604,In_1608,In_1912);
nor U605 (N_605,In_317,In_698);
nor U606 (N_606,N_474,In_622);
xor U607 (N_607,In_344,In_334);
nor U608 (N_608,N_437,N_363);
nor U609 (N_609,In_1481,In_1940);
xnor U610 (N_610,N_4,In_977);
xnor U611 (N_611,In_1032,In_1714);
nand U612 (N_612,In_734,In_117);
nor U613 (N_613,N_409,In_1080);
and U614 (N_614,N_343,In_1150);
and U615 (N_615,In_127,In_1144);
xor U616 (N_616,In_367,In_1877);
xnor U617 (N_617,In_1349,N_178);
nor U618 (N_618,In_1534,In_1372);
and U619 (N_619,N_41,In_118);
and U620 (N_620,In_1335,In_51);
nor U621 (N_621,In_1679,N_128);
or U622 (N_622,In_1985,N_357);
nor U623 (N_623,In_1553,N_479);
nor U624 (N_624,In_555,N_219);
xnor U625 (N_625,In_1558,N_339);
nor U626 (N_626,In_881,N_397);
nor U627 (N_627,In_1085,N_179);
or U628 (N_628,In_1035,N_281);
xnor U629 (N_629,N_375,In_400);
or U630 (N_630,In_879,In_1549);
or U631 (N_631,In_1964,N_275);
nand U632 (N_632,In_1717,In_1680);
and U633 (N_633,In_444,N_133);
nand U634 (N_634,In_930,In_1440);
or U635 (N_635,In_396,In_954);
nor U636 (N_636,In_1525,In_1415);
or U637 (N_637,In_1959,In_1711);
nor U638 (N_638,In_481,N_108);
nor U639 (N_639,N_149,In_1611);
nor U640 (N_640,N_110,N_250);
and U641 (N_641,In_453,N_5);
xnor U642 (N_642,In_1799,N_242);
nor U643 (N_643,In_1495,In_818);
or U644 (N_644,In_757,In_328);
nor U645 (N_645,N_56,N_499);
xor U646 (N_646,In_1868,In_779);
nor U647 (N_647,In_1204,In_1433);
and U648 (N_648,In_1845,In_1243);
xnor U649 (N_649,In_452,In_1825);
nor U650 (N_650,In_722,In_1276);
nand U651 (N_651,In_187,In_639);
xnor U652 (N_652,N_292,In_583);
or U653 (N_653,In_645,N_491);
xor U654 (N_654,In_1957,In_31);
or U655 (N_655,In_441,In_420);
xnor U656 (N_656,N_115,N_66);
nand U657 (N_657,In_801,In_826);
nand U658 (N_658,N_176,In_298);
and U659 (N_659,N_326,N_231);
and U660 (N_660,N_84,In_1564);
nand U661 (N_661,N_311,In_238);
nand U662 (N_662,In_30,N_361);
nand U663 (N_663,In_188,In_1980);
xor U664 (N_664,N_459,In_1883);
nor U665 (N_665,N_470,N_39);
or U666 (N_666,N_389,N_316);
and U667 (N_667,In_1523,In_1801);
nor U668 (N_668,In_1277,In_872);
and U669 (N_669,N_273,In_925);
nor U670 (N_670,N_377,In_1708);
xnor U671 (N_671,N_410,In_302);
or U672 (N_672,In_352,N_296);
nor U673 (N_673,In_1782,In_1090);
xnor U674 (N_674,In_1026,In_1077);
or U675 (N_675,In_1419,N_423);
nor U676 (N_676,In_1435,N_373);
xnor U677 (N_677,In_133,In_922);
and U678 (N_678,In_1654,In_1219);
nor U679 (N_679,In_681,N_288);
nand U680 (N_680,N_498,In_764);
nor U681 (N_681,In_675,In_428);
xnor U682 (N_682,In_273,In_240);
nand U683 (N_683,N_261,N_253);
xnor U684 (N_684,In_1341,N_426);
or U685 (N_685,N_279,In_942);
and U686 (N_686,In_28,N_14);
xnor U687 (N_687,N_317,In_184);
and U688 (N_688,In_54,N_94);
nand U689 (N_689,In_83,In_1707);
nand U690 (N_690,In_1100,In_1997);
xor U691 (N_691,In_1559,In_1448);
xor U692 (N_692,N_280,N_120);
nor U693 (N_693,N_436,In_841);
nor U694 (N_694,In_34,N_213);
and U695 (N_695,In_291,N_55);
nor U696 (N_696,N_141,N_356);
or U697 (N_697,N_135,N_40);
nor U698 (N_698,In_1834,In_1105);
and U699 (N_699,N_355,In_1750);
or U700 (N_700,N_411,In_1841);
and U701 (N_701,In_1661,N_100);
nor U702 (N_702,N_222,N_448);
and U703 (N_703,In_1719,N_194);
or U704 (N_704,In_1823,N_297);
or U705 (N_705,In_1064,In_552);
nor U706 (N_706,In_1765,N_114);
and U707 (N_707,In_247,In_1289);
nand U708 (N_708,In_565,In_435);
nor U709 (N_709,N_43,N_480);
and U710 (N_710,N_214,In_313);
nor U711 (N_711,N_75,In_897);
nor U712 (N_712,N_61,In_729);
and U713 (N_713,In_1614,In_643);
and U714 (N_714,In_1539,In_690);
nand U715 (N_715,In_706,In_1639);
and U716 (N_716,N_484,N_267);
nand U717 (N_717,N_238,N_15);
nor U718 (N_718,N_446,N_315);
nand U719 (N_719,In_1227,N_400);
or U720 (N_720,N_425,N_172);
and U721 (N_721,In_600,In_1331);
or U722 (N_722,In_524,N_482);
nand U723 (N_723,In_168,N_209);
xor U724 (N_724,In_1453,In_803);
and U725 (N_725,In_1213,In_73);
or U726 (N_726,In_998,In_1924);
nor U727 (N_727,In_1948,N_165);
xor U728 (N_728,In_1683,In_116);
and U729 (N_729,In_743,N_71);
or U730 (N_730,In_1488,In_1829);
and U731 (N_731,In_1009,In_293);
or U732 (N_732,In_1723,In_928);
and U733 (N_733,N_22,In_41);
nand U734 (N_734,In_1052,In_592);
nand U735 (N_735,In_211,N_83);
and U736 (N_736,N_432,In_838);
nor U737 (N_737,In_1429,In_654);
or U738 (N_738,In_578,N_119);
and U739 (N_739,In_1379,In_850);
xor U740 (N_740,N_266,N_366);
nand U741 (N_741,In_1264,N_463);
xor U742 (N_742,In_132,In_1499);
nor U743 (N_743,In_170,In_75);
and U744 (N_744,In_242,In_1507);
and U745 (N_745,In_695,In_715);
or U746 (N_746,In_409,N_117);
xnor U747 (N_747,In_1336,N_228);
xor U748 (N_748,In_871,In_517);
xnor U749 (N_749,N_87,In_414);
xnor U750 (N_750,In_1367,In_347);
or U751 (N_751,In_1772,N_415);
and U752 (N_752,In_464,In_1866);
or U753 (N_753,N_57,In_860);
nor U754 (N_754,In_857,In_1904);
nand U755 (N_755,In_824,In_1910);
and U756 (N_756,N_318,In_1432);
xor U757 (N_757,In_489,N_109);
or U758 (N_758,N_137,N_31);
nor U759 (N_759,N_73,N_190);
or U760 (N_760,N_438,N_486);
and U761 (N_761,In_1468,In_1458);
nand U762 (N_762,N_159,In_1822);
and U763 (N_763,In_478,In_799);
xor U764 (N_764,In_213,In_797);
nand U765 (N_765,In_331,In_624);
xnor U766 (N_766,In_1039,N_217);
xor U767 (N_767,In_370,In_20);
nor U768 (N_768,In_53,N_252);
or U769 (N_769,N_229,N_223);
xnor U770 (N_770,In_727,N_147);
xor U771 (N_771,In_1599,N_116);
xnor U772 (N_772,N_483,In_1390);
and U773 (N_773,In_965,N_306);
nor U774 (N_774,In_1179,In_825);
or U775 (N_775,N_191,In_275);
or U776 (N_776,In_636,In_737);
or U777 (N_777,N_481,N_378);
nor U778 (N_778,In_794,In_193);
nand U779 (N_779,In_1377,N_372);
and U780 (N_780,In_1396,N_312);
nand U781 (N_781,In_751,In_1261);
and U782 (N_782,In_1927,In_1395);
nand U783 (N_783,N_472,In_659);
xor U784 (N_784,In_292,N_259);
nand U785 (N_785,In_1242,In_1271);
and U786 (N_786,In_1618,In_856);
xnor U787 (N_787,In_1291,In_708);
xor U788 (N_788,In_507,N_300);
nor U789 (N_789,In_1727,In_541);
nand U790 (N_790,In_1288,N_65);
or U791 (N_791,In_960,N_186);
xnor U792 (N_792,N_91,In_191);
xor U793 (N_793,In_102,In_728);
nor U794 (N_794,N_274,N_254);
nor U795 (N_795,In_1344,In_1556);
nor U796 (N_796,In_459,In_207);
and U797 (N_797,In_559,In_314);
nand U798 (N_798,In_454,In_346);
nand U799 (N_799,In_1351,In_1633);
or U800 (N_800,N_310,N_291);
or U801 (N_801,N_0,In_1380);
xor U802 (N_802,N_78,In_1977);
nor U803 (N_803,In_1205,N_469);
nand U804 (N_804,In_1054,In_1552);
xnor U805 (N_805,N_271,In_217);
xor U806 (N_806,In_1099,In_1820);
nand U807 (N_807,N_460,In_1070);
nor U808 (N_808,In_9,In_195);
xnor U809 (N_809,In_612,In_606);
nand U810 (N_810,In_987,In_142);
or U811 (N_811,In_282,In_103);
and U812 (N_812,In_1449,N_439);
or U813 (N_813,In_1450,N_129);
or U814 (N_814,In_1299,In_683);
nor U815 (N_815,In_1849,N_347);
and U816 (N_816,N_227,In_1976);
nand U817 (N_817,In_231,N_126);
nand U818 (N_818,N_82,In_497);
and U819 (N_819,In_1118,In_154);
xnor U820 (N_820,In_532,In_1713);
nand U821 (N_821,In_1400,In_42);
nand U822 (N_822,In_1455,N_476);
xnor U823 (N_823,N_258,In_1162);
and U824 (N_824,In_341,N_402);
or U825 (N_825,N_257,In_910);
nor U826 (N_826,In_1250,In_475);
and U827 (N_827,In_1724,N_156);
nand U828 (N_828,In_7,N_473);
xor U829 (N_829,In_1918,N_395);
nor U830 (N_830,In_1012,In_1852);
and U831 (N_831,In_469,In_1493);
or U832 (N_832,N_8,N_249);
xor U833 (N_833,In_1326,In_498);
and U834 (N_834,In_906,N_351);
nor U835 (N_835,In_1598,In_522);
or U836 (N_836,In_1037,In_1641);
nor U837 (N_837,N_462,In_1231);
nand U838 (N_838,In_1520,In_114);
and U839 (N_839,N_468,In_809);
nand U840 (N_840,In_1383,In_777);
nor U841 (N_841,In_1574,In_700);
or U842 (N_842,N_81,In_611);
xor U843 (N_843,In_233,In_540);
xnor U844 (N_844,N_188,In_986);
xnor U845 (N_845,In_1409,N_331);
xor U846 (N_846,In_1484,In_978);
nor U847 (N_847,N_346,In_1191);
nor U848 (N_848,In_533,N_35);
and U849 (N_849,In_995,N_342);
or U850 (N_850,N_485,N_121);
nor U851 (N_851,In_108,N_148);
nor U852 (N_852,N_309,N_330);
or U853 (N_853,In_1062,In_821);
nand U854 (N_854,In_69,N_340);
or U855 (N_855,In_1302,In_1056);
nand U856 (N_856,In_1174,In_849);
nor U857 (N_857,In_670,N_399);
nor U858 (N_858,N_106,N_146);
and U859 (N_859,N_445,In_1232);
xor U860 (N_860,N_236,N_60);
or U861 (N_861,N_224,N_225);
or U862 (N_862,In_1328,In_980);
xor U863 (N_863,In_1891,In_1881);
nand U864 (N_864,In_405,N_447);
xnor U865 (N_865,In_509,In_1938);
and U866 (N_866,In_348,N_132);
nor U867 (N_867,In_1689,N_192);
and U868 (N_868,N_103,N_334);
xnor U869 (N_869,N_327,In_1214);
and U870 (N_870,In_95,In_1253);
or U871 (N_871,N_32,In_183);
xor U872 (N_872,In_1352,In_884);
and U873 (N_873,In_668,In_836);
or U874 (N_874,N_237,In_1842);
or U875 (N_875,In_1120,N_79);
or U876 (N_876,In_1733,In_696);
nand U877 (N_877,In_1622,In_1360);
nor U878 (N_878,N_283,In_1773);
and U879 (N_879,In_725,In_1814);
and U880 (N_880,N_413,N_401);
or U881 (N_881,In_1142,In_1947);
xor U882 (N_882,N_262,N_245);
and U883 (N_883,In_1343,N_263);
nor U884 (N_884,In_1273,In_1802);
xor U885 (N_885,N_200,In_1761);
or U886 (N_886,N_184,In_1117);
nor U887 (N_887,In_1422,In_1658);
xor U888 (N_888,In_1982,N_368);
and U889 (N_889,In_674,In_908);
xnor U890 (N_890,In_863,N_325);
and U891 (N_891,N_58,N_7);
and U892 (N_892,In_495,N_303);
xor U893 (N_893,In_1082,In_735);
nand U894 (N_894,In_1441,In_991);
and U895 (N_895,In_1478,N_392);
nand U896 (N_896,In_1378,N_424);
nand U897 (N_897,In_461,In_1019);
nand U898 (N_898,N_307,In_1498);
and U899 (N_899,N_321,In_1533);
nor U900 (N_900,N_269,In_1575);
xor U901 (N_901,N_414,In_1137);
nor U902 (N_902,N_371,In_546);
or U903 (N_903,In_679,In_402);
or U904 (N_904,In_172,In_360);
nand U905 (N_905,In_1807,N_475);
or U906 (N_906,N_430,In_1545);
or U907 (N_907,N_207,In_476);
or U908 (N_908,N_268,In_575);
or U909 (N_909,In_1749,N_130);
and U910 (N_910,In_736,In_877);
nand U911 (N_911,N_335,In_1148);
nand U912 (N_912,In_1818,In_1861);
nand U913 (N_913,In_919,N_69);
or U914 (N_914,N_256,N_285);
nand U915 (N_915,In_916,In_1216);
nand U916 (N_916,In_289,N_461);
or U917 (N_917,N_134,In_1492);
and U918 (N_918,In_1013,In_236);
xnor U919 (N_919,In_1786,N_113);
nand U920 (N_920,N_234,In_312);
nor U921 (N_921,In_90,N_162);
nor U922 (N_922,N_138,In_1968);
and U923 (N_923,In_705,In_140);
and U924 (N_924,In_800,In_269);
nand U925 (N_925,In_1218,In_468);
nor U926 (N_926,In_252,In_976);
nor U927 (N_927,In_758,In_613);
nor U928 (N_928,In_875,N_488);
nor U929 (N_929,In_196,N_412);
nand U930 (N_930,In_460,In_1607);
xnor U931 (N_931,In_1386,In_1228);
xor U932 (N_932,In_990,In_323);
xnor U933 (N_933,In_182,N_54);
and U934 (N_934,In_923,In_691);
nor U935 (N_935,In_1036,In_71);
nand U936 (N_936,In_1800,N_360);
nand U937 (N_937,In_1168,In_447);
and U938 (N_938,N_226,N_102);
or U939 (N_939,In_1690,In_0);
or U940 (N_940,In_504,In_905);
xnor U941 (N_941,In_1833,N_59);
xor U942 (N_942,In_225,In_1081);
nor U943 (N_943,In_301,In_1991);
and U944 (N_944,In_1234,In_1434);
and U945 (N_945,N_305,In_448);
or U946 (N_946,N_160,In_1222);
xnor U947 (N_947,In_604,In_1129);
nand U948 (N_948,In_576,In_1902);
and U949 (N_949,N_11,N_324);
or U950 (N_950,In_1662,In_1785);
xor U951 (N_951,N_464,N_10);
or U952 (N_952,N_185,In_890);
or U953 (N_953,N_177,In_125);
xnor U954 (N_954,In_106,In_790);
nand U955 (N_955,In_186,In_1916);
and U956 (N_956,In_831,N_118);
nand U957 (N_957,N_68,N_353);
xnor U958 (N_958,In_1903,N_376);
nand U959 (N_959,N_246,In_1961);
or U960 (N_960,N_150,N_308);
xor U961 (N_961,In_1304,In_149);
nor U962 (N_962,In_1061,In_1398);
nor U963 (N_963,In_375,N_319);
nand U964 (N_964,In_545,In_1999);
xnor U965 (N_965,N_90,In_685);
xor U966 (N_966,In_1593,In_199);
xnor U967 (N_967,N_380,N_1);
and U968 (N_968,N_298,N_171);
nor U969 (N_969,In_1511,In_145);
nor U970 (N_970,In_437,In_694);
and U971 (N_971,In_1628,In_436);
xnor U972 (N_972,N_72,N_16);
nor U973 (N_973,N_211,N_201);
nand U974 (N_974,In_709,In_1278);
xor U975 (N_975,In_1602,In_281);
or U976 (N_976,N_487,In_1758);
nor U977 (N_977,N_383,In_1721);
xnor U978 (N_978,In_1526,N_416);
nor U979 (N_979,In_1887,In_361);
or U980 (N_980,In_931,In_412);
and U981 (N_981,In_1173,In_1815);
nor U982 (N_982,In_571,N_183);
nor U983 (N_983,In_1764,In_1731);
nor U984 (N_984,In_970,In_1892);
nand U985 (N_985,In_1394,In_1870);
nand U986 (N_986,In_1857,In_851);
nor U987 (N_987,In_1027,In_1681);
nand U988 (N_988,In_702,N_493);
nand U989 (N_989,In_1660,In_43);
nor U990 (N_990,In_1554,In_984);
and U991 (N_991,In_147,In_1668);
xor U992 (N_992,N_240,In_373);
and U993 (N_993,In_429,N_167);
nor U994 (N_994,In_1722,In_1926);
nand U995 (N_995,N_23,In_1315);
xnor U996 (N_996,N_216,N_456);
and U997 (N_997,N_197,In_1324);
or U998 (N_998,N_329,In_560);
xnor U999 (N_999,In_391,In_1320);
xnor U1000 (N_1000,N_667,N_123);
xnor U1001 (N_1001,In_1847,In_161);
nand U1002 (N_1002,In_1074,N_928);
and U1003 (N_1003,N_504,In_1084);
and U1004 (N_1004,N_289,In_1425);
or U1005 (N_1005,N_492,N_626);
nand U1006 (N_1006,In_260,In_732);
xor U1007 (N_1007,N_212,N_690);
nor U1008 (N_1008,In_1804,In_1154);
xnor U1009 (N_1009,In_408,N_859);
nand U1010 (N_1010,In_1561,N_998);
nand U1011 (N_1011,N_733,N_727);
nand U1012 (N_1012,N_169,In_440);
xnor U1013 (N_1013,In_1016,N_442);
nand U1014 (N_1014,N_594,N_900);
nand U1015 (N_1015,N_909,N_961);
or U1016 (N_1016,N_920,N_584);
or U1017 (N_1017,In_1210,N_251);
nand U1018 (N_1018,In_371,N_393);
or U1019 (N_1019,N_965,N_997);
or U1020 (N_1020,N_662,N_875);
nor U1021 (N_1021,In_1939,N_688);
nand U1022 (N_1022,In_971,N_505);
nand U1023 (N_1023,N_511,In_38);
and U1024 (N_1024,In_176,In_499);
xnor U1025 (N_1025,N_671,N_323);
nand U1026 (N_1026,In_1265,N_12);
or U1027 (N_1027,N_163,In_1092);
or U1028 (N_1028,N_679,N_739);
nand U1029 (N_1029,N_613,N_921);
and U1030 (N_1030,In_156,N_708);
xor U1031 (N_1031,N_615,N_546);
nor U1032 (N_1032,In_921,N_532);
nand U1033 (N_1033,N_725,N_906);
and U1034 (N_1034,N_812,In_351);
or U1035 (N_1035,N_573,In_425);
or U1036 (N_1036,N_362,N_852);
nor U1037 (N_1037,In_786,N_872);
and U1038 (N_1038,In_1194,N_814);
xor U1039 (N_1039,In_57,N_629);
or U1040 (N_1040,N_549,N_140);
nor U1041 (N_1041,N_706,N_907);
and U1042 (N_1042,N_76,In_869);
and U1043 (N_1043,In_310,N_967);
nor U1044 (N_1044,In_1776,N_883);
xnor U1045 (N_1045,N_164,N_574);
nand U1046 (N_1046,N_726,In_120);
nand U1047 (N_1047,N_780,N_101);
xnor U1048 (N_1048,In_1158,N_548);
nor U1049 (N_1049,N_518,N_990);
nor U1050 (N_1050,In_390,In_223);
and U1051 (N_1051,N_454,N_443);
nor U1052 (N_1052,N_945,N_689);
nor U1053 (N_1053,In_945,N_915);
or U1054 (N_1054,N_382,N_19);
and U1055 (N_1055,N_822,In_876);
and U1056 (N_1056,N_534,N_957);
or U1057 (N_1057,In_1095,N_320);
and U1058 (N_1058,N_698,N_806);
and U1059 (N_1059,N_614,N_966);
nand U1060 (N_1060,N_729,N_897);
xnor U1061 (N_1061,N_25,N_743);
xor U1062 (N_1062,N_912,In_1366);
or U1063 (N_1063,In_773,N_685);
or U1064 (N_1064,N_809,In_1617);
nand U1065 (N_1065,N_564,In_129);
and U1066 (N_1066,N_828,In_1620);
or U1067 (N_1067,N_678,N_752);
nor U1068 (N_1068,N_844,N_892);
and U1069 (N_1069,In_482,N_665);
and U1070 (N_1070,N_746,In_21);
and U1071 (N_1071,In_1905,In_1275);
nand U1072 (N_1072,N_742,N_958);
and U1073 (N_1073,In_1944,N_465);
nor U1074 (N_1074,In_904,In_445);
nor U1075 (N_1075,N_450,In_861);
and U1076 (N_1076,N_36,N_854);
nand U1077 (N_1077,In_175,In_1000);
or U1078 (N_1078,N_540,N_790);
nand U1079 (N_1079,In_840,In_1004);
or U1080 (N_1080,N_981,N_798);
xnor U1081 (N_1081,N_526,N_580);
and U1082 (N_1082,In_1638,In_667);
xor U1083 (N_1083,N_841,In_1410);
nor U1084 (N_1084,N_98,N_587);
or U1085 (N_1085,N_836,In_1778);
and U1086 (N_1086,In_227,N_876);
or U1087 (N_1087,N_623,N_994);
or U1088 (N_1088,N_293,N_507);
nor U1089 (N_1089,In_1199,N_984);
nor U1090 (N_1090,In_633,N_865);
xnor U1091 (N_1091,In_1623,In_1480);
nand U1092 (N_1092,In_174,N_407);
and U1093 (N_1093,In_1863,N_861);
xor U1094 (N_1094,N_599,N_683);
nor U1095 (N_1095,In_68,In_477);
or U1096 (N_1096,N_648,In_115);
or U1097 (N_1097,In_205,N_466);
nand U1098 (N_1098,N_931,N_607);
nor U1099 (N_1099,N_660,N_808);
nor U1100 (N_1100,N_694,In_46);
nor U1101 (N_1101,N_919,N_533);
nand U1102 (N_1102,N_884,In_1025);
and U1103 (N_1103,N_716,In_1836);
and U1104 (N_1104,N_830,N_583);
nor U1105 (N_1105,In_14,N_956);
and U1106 (N_1106,N_44,In_969);
xnor U1107 (N_1107,N_544,N_829);
nand U1108 (N_1108,N_105,N_97);
nor U1109 (N_1109,In_1788,N_929);
nor U1110 (N_1110,N_863,In_248);
or U1111 (N_1111,N_969,N_642);
xnor U1112 (N_1112,N_771,N_952);
xor U1113 (N_1113,N_444,N_239);
xor U1114 (N_1114,In_1768,N_630);
nand U1115 (N_1115,In_109,N_500);
xnor U1116 (N_1116,N_517,N_831);
nor U1117 (N_1117,In_1740,N_650);
xor U1118 (N_1118,N_433,N_800);
nor U1119 (N_1119,N_821,N_911);
or U1120 (N_1120,N_88,N_979);
and U1121 (N_1121,N_51,In_1402);
nor U1122 (N_1122,N_772,In_1958);
nand U1123 (N_1123,N_799,In_1603);
or U1124 (N_1124,In_224,N_85);
xnor U1125 (N_1125,N_46,N_781);
nand U1126 (N_1126,N_882,N_441);
nor U1127 (N_1127,N_348,N_576);
or U1128 (N_1128,N_37,N_817);
or U1129 (N_1129,In_128,In_917);
and U1130 (N_1130,N_490,N_616);
and U1131 (N_1131,In_1160,N_537);
xor U1132 (N_1132,In_1568,N_295);
or U1133 (N_1133,N_513,In_993);
nand U1134 (N_1134,N_871,In_1098);
nor U1135 (N_1135,N_552,In_1268);
and U1136 (N_1136,N_950,In_1936);
nor U1137 (N_1137,In_823,In_486);
xor U1138 (N_1138,N_536,N_757);
xnor U1139 (N_1139,In_1769,In_1050);
and U1140 (N_1140,N_837,N_696);
xnor U1141 (N_1141,In_1537,In_1283);
nor U1142 (N_1142,In_1399,N_477);
nand U1143 (N_1143,N_92,In_834);
xor U1144 (N_1144,N_918,N_948);
or U1145 (N_1145,In_300,In_1110);
or U1146 (N_1146,N_714,In_1408);
nor U1147 (N_1147,In_920,N_637);
nor U1148 (N_1148,N_503,N_811);
or U1149 (N_1149,N_592,N_265);
nand U1150 (N_1150,N_24,N_74);
or U1151 (N_1151,N_453,In_782);
and U1152 (N_1152,N_196,In_45);
and U1153 (N_1153,N_313,N_602);
and U1154 (N_1154,N_840,In_1297);
nor U1155 (N_1155,In_1342,N_776);
or U1156 (N_1156,N_804,N_955);
or U1157 (N_1157,N_612,In_1701);
and U1158 (N_1158,N_455,N_515);
and U1159 (N_1159,N_428,In_1645);
or U1160 (N_1160,In_867,N_510);
xnor U1161 (N_1161,N_604,N_827);
nand U1162 (N_1162,N_666,In_1029);
or U1163 (N_1163,N_38,N_260);
xor U1164 (N_1164,N_962,In_382);
or U1165 (N_1165,N_512,N_759);
nor U1166 (N_1166,In_1477,In_1566);
and U1167 (N_1167,In_804,N_624);
and U1168 (N_1168,N_595,In_158);
nor U1169 (N_1169,N_349,N_693);
nand U1170 (N_1170,N_204,In_85);
and U1171 (N_1171,In_1290,N_913);
nor U1172 (N_1172,N_558,N_632);
or U1173 (N_1173,In_10,N_881);
xnor U1174 (N_1174,N_301,N_417);
and U1175 (N_1175,N_67,N_641);
nor U1176 (N_1176,N_795,N_560);
xor U1177 (N_1177,In_80,N_601);
nor U1178 (N_1178,N_736,N_673);
nand U1179 (N_1179,N_235,N_802);
or U1180 (N_1180,N_577,In_501);
nand U1181 (N_1181,N_735,N_762);
xnor U1182 (N_1182,In_1446,N_420);
nor U1183 (N_1183,N_658,N_33);
and U1184 (N_1184,N_963,N_755);
xnor U1185 (N_1185,In_1447,In_1470);
nand U1186 (N_1186,In_219,N_991);
nor U1187 (N_1187,N_718,N_568);
and U1188 (N_1188,In_1270,N_784);
and U1189 (N_1189,In_958,N_745);
and U1190 (N_1190,N_86,In_36);
or U1191 (N_1191,In_1670,N_959);
or U1192 (N_1192,N_639,N_396);
and U1193 (N_1193,N_717,In_1664);
nand U1194 (N_1194,In_284,N_125);
and U1195 (N_1195,N_701,In_1817);
nor U1196 (N_1196,N_652,In_1889);
and U1197 (N_1197,In_163,In_569);
nand U1198 (N_1198,N_302,N_677);
xor U1199 (N_1199,N_27,In_862);
xor U1200 (N_1200,In_1190,N_341);
nor U1201 (N_1201,In_1181,N_894);
or U1202 (N_1202,N_647,N_538);
or U1203 (N_1203,In_1508,N_825);
nor U1204 (N_1204,N_509,In_1743);
xnor U1205 (N_1205,N_857,N_704);
and U1206 (N_1206,N_390,N_45);
nor U1207 (N_1207,N_770,N_885);
xnor U1208 (N_1208,In_1766,N_942);
and U1209 (N_1209,In_1606,N_527);
nand U1210 (N_1210,N_946,N_421);
or U1211 (N_1211,In_1244,In_267);
nand U1212 (N_1212,N_29,N_670);
or U1213 (N_1213,N_940,N_778);
or U1214 (N_1214,N_646,In_864);
and U1215 (N_1215,N_107,N_970);
xnor U1216 (N_1216,N_682,N_530);
nand U1217 (N_1217,In_89,N_535);
nand U1218 (N_1218,In_19,N_675);
or U1219 (N_1219,N_332,N_996);
or U1220 (N_1220,N_870,N_864);
nor U1221 (N_1221,In_271,In_775);
nand U1222 (N_1222,N_987,N_767);
nor U1223 (N_1223,N_610,In_29);
nor U1224 (N_1224,N_17,N_555);
nand U1225 (N_1225,N_801,N_972);
nor U1226 (N_1226,In_1687,N_394);
nand U1227 (N_1227,N_794,N_157);
or U1228 (N_1228,N_709,N_422);
nand U1229 (N_1229,N_839,N_989);
nand U1230 (N_1230,N_923,N_853);
xnor U1231 (N_1231,In_999,N_649);
and U1232 (N_1232,N_786,N_758);
nand U1233 (N_1233,N_333,N_886);
nand U1234 (N_1234,N_598,N_600);
nand U1235 (N_1235,In_254,N_585);
or U1236 (N_1236,N_638,N_849);
nand U1237 (N_1237,N_902,N_788);
xnor U1238 (N_1238,N_627,In_1637);
or U1239 (N_1239,In_245,N_152);
nor U1240 (N_1240,N_651,In_1751);
xnor U1241 (N_1241,N_521,In_1217);
and U1242 (N_1242,N_796,N_927);
nor U1243 (N_1243,N_703,N_964);
xor U1244 (N_1244,N_571,N_528);
nor U1245 (N_1245,In_859,In_1580);
or U1246 (N_1246,In_204,N_345);
or U1247 (N_1247,N_519,N_572);
and U1248 (N_1248,In_1560,N_954);
xor U1249 (N_1249,N_299,N_605);
xor U1250 (N_1250,In_1635,N_643);
nor U1251 (N_1251,N_496,In_473);
nor U1252 (N_1252,N_589,In_1565);
nand U1253 (N_1253,In_564,N_350);
xnor U1254 (N_1254,N_663,N_988);
nand U1255 (N_1255,In_1046,N_661);
nor U1256 (N_1256,N_980,N_155);
or U1257 (N_1257,N_789,N_760);
nand U1258 (N_1258,N_3,N_352);
or U1259 (N_1259,N_938,In_1860);
nor U1260 (N_1260,N_766,N_13);
xor U1261 (N_1261,N_553,N_233);
and U1262 (N_1262,N_634,In_711);
nor U1263 (N_1263,N_761,N_131);
nand U1264 (N_1264,N_815,In_82);
or U1265 (N_1265,N_824,N_935);
nand U1266 (N_1266,N_699,In_1460);
xor U1267 (N_1267,In_1245,In_407);
or U1268 (N_1268,N_960,N_569);
nor U1269 (N_1269,N_834,N_932);
and U1270 (N_1270,N_70,N_974);
or U1271 (N_1271,In_520,N_654);
and U1272 (N_1272,In_1853,N_563);
nand U1273 (N_1273,In_1832,In_968);
xnor U1274 (N_1274,N_896,In_342);
or U1275 (N_1275,In_1428,N_993);
xnor U1276 (N_1276,N_914,N_951);
and U1277 (N_1277,In_1206,N_713);
and U1278 (N_1278,N_810,N_554);
nand U1279 (N_1279,In_1116,In_1143);
or U1280 (N_1280,In_326,In_1674);
and U1281 (N_1281,N_550,In_760);
and U1282 (N_1282,N_702,N_151);
or U1283 (N_1283,N_586,N_764);
or U1284 (N_1284,N_851,N_561);
xor U1285 (N_1285,N_566,In_1524);
and U1286 (N_1286,N_692,N_656);
nor U1287 (N_1287,In_665,In_49);
and U1288 (N_1288,In_1051,In_1220);
and U1289 (N_1289,N_893,In_1340);
nand U1290 (N_1290,N_730,In_58);
xor U1291 (N_1291,In_1890,In_17);
or U1292 (N_1292,N_823,N_868);
and U1293 (N_1293,N_724,In_1530);
or U1294 (N_1294,N_543,In_664);
nand U1295 (N_1295,In_392,N_835);
or U1296 (N_1296,N_846,In_952);
nor U1297 (N_1297,N_506,In_647);
nand U1298 (N_1298,In_1762,In_1827);
xor U1299 (N_1299,N_9,N_779);
xor U1300 (N_1300,N_797,N_842);
xor U1301 (N_1301,N_408,N_731);
or U1302 (N_1302,N_793,N_953);
nand U1303 (N_1303,N_887,N_791);
nand U1304 (N_1304,In_748,N_895);
or U1305 (N_1305,N_628,N_562);
nand U1306 (N_1306,N_581,N_832);
and U1307 (N_1307,In_1494,In_1718);
and U1308 (N_1308,N_6,N_53);
or U1309 (N_1309,N_419,In_152);
xnor U1310 (N_1310,N_621,N_856);
or U1311 (N_1311,N_879,N_684);
nand U1312 (N_1312,N_686,N_986);
nor U1313 (N_1313,N_452,N_588);
or U1314 (N_1314,In_788,N_947);
nand U1315 (N_1315,In_1373,In_1527);
xnor U1316 (N_1316,In_74,In_621);
xnor U1317 (N_1317,In_76,N_153);
xor U1318 (N_1318,In_614,N_934);
and U1319 (N_1319,In_1020,In_707);
nor U1320 (N_1320,In_1675,N_403);
and U1321 (N_1321,N_977,N_187);
and U1322 (N_1322,In_741,In_648);
nor U1323 (N_1323,In_601,N_732);
xor U1324 (N_1324,N_925,In_1169);
or U1325 (N_1325,N_495,N_559);
nor U1326 (N_1326,N_785,N_287);
and U1327 (N_1327,N_653,In_1467);
nand U1328 (N_1328,N_633,N_195);
or U1329 (N_1329,N_978,In_843);
and U1330 (N_1330,N_220,In_1308);
xor U1331 (N_1331,N_691,N_2);
and U1332 (N_1332,In_1753,N_202);
or U1333 (N_1333,In_1136,In_1312);
or U1334 (N_1334,N_304,In_177);
nand U1335 (N_1335,N_244,N_597);
xor U1336 (N_1336,In_1501,N_578);
and U1337 (N_1337,N_18,N_845);
or U1338 (N_1338,N_924,N_753);
nand U1339 (N_1339,In_688,In_52);
and U1340 (N_1340,N_608,N_567);
nor U1341 (N_1341,In_1021,In_1590);
xor U1342 (N_1342,N_750,In_171);
or U1343 (N_1343,N_104,N_734);
xor U1344 (N_1344,N_286,N_860);
nand U1345 (N_1345,N_208,N_777);
or U1346 (N_1346,N_763,In_951);
nand U1347 (N_1347,N_609,N_619);
or U1348 (N_1348,N_221,N_710);
and U1349 (N_1349,N_596,In_814);
or U1350 (N_1350,N_282,N_611);
and U1351 (N_1351,N_494,In_1984);
and U1352 (N_1352,In_1858,N_531);
or U1353 (N_1353,N_659,N_582);
and U1354 (N_1354,In_918,In_221);
and U1355 (N_1355,N_862,N_922);
or U1356 (N_1356,N_142,In_767);
and U1357 (N_1357,N_754,N_976);
xnor U1358 (N_1358,In_1049,N_944);
and U1359 (N_1359,In_1279,In_1943);
and U1360 (N_1360,In_1596,N_154);
nor U1361 (N_1361,N_218,N_431);
and U1362 (N_1362,In_1152,N_565);
nand U1363 (N_1363,N_42,In_1078);
or U1364 (N_1364,N_803,N_434);
or U1365 (N_1365,In_1221,In_465);
xor U1366 (N_1366,N_277,N_937);
nor U1367 (N_1367,N_756,N_381);
xnor U1368 (N_1368,N_99,N_644);
nor U1369 (N_1369,N_728,In_1888);
nor U1370 (N_1370,N_387,In_652);
xnor U1371 (N_1371,N_910,N_631);
or U1372 (N_1372,N_384,In_1211);
and U1373 (N_1373,N_774,N_591);
or U1374 (N_1374,N_617,In_1712);
and U1375 (N_1375,N_880,In_536);
nand U1376 (N_1376,N_992,In_1069);
nand U1377 (N_1377,N_636,In_279);
or U1378 (N_1378,N_189,In_1934);
and U1379 (N_1379,N_805,N_635);
nand U1380 (N_1380,In_992,N_949);
or U1381 (N_1381,In_1321,In_885);
or U1382 (N_1382,In_789,N_707);
nand U1383 (N_1383,N_792,N_697);
and U1384 (N_1384,N_869,N_904);
xnor U1385 (N_1385,N_622,N_737);
nand U1386 (N_1386,In_1071,In_1955);
xor U1387 (N_1387,N_680,N_529);
and U1388 (N_1388,N_440,In_1990);
nand U1389 (N_1389,N_80,In_1970);
nor U1390 (N_1390,N_542,N_983);
nand U1391 (N_1391,In_246,In_26);
xnor U1392 (N_1392,N_556,N_941);
and U1393 (N_1393,N_525,N_874);
nor U1394 (N_1394,In_1201,N_833);
nor U1395 (N_1395,In_1716,N_514);
nand U1396 (N_1396,N_787,N_818);
and U1397 (N_1397,N_664,N_749);
and U1398 (N_1398,In_381,N_681);
and U1399 (N_1399,In_394,In_1192);
nor U1400 (N_1400,N_551,N_850);
or U1401 (N_1401,In_684,N_712);
nand U1402 (N_1402,N_890,N_738);
nor U1403 (N_1403,In_1238,N_593);
or U1404 (N_1404,N_174,N_816);
nor U1405 (N_1405,N_63,In_491);
and U1406 (N_1406,In_1960,N_926);
or U1407 (N_1407,In_780,N_206);
and U1408 (N_1408,N_982,In_577);
and U1409 (N_1409,N_502,N_847);
xnor U1410 (N_1410,N_606,N_975);
xnor U1411 (N_1411,N_640,N_557);
and U1412 (N_1412,N_522,In_335);
nand U1413 (N_1413,N_379,In_216);
nand U1414 (N_1414,N_768,In_1473);
or U1415 (N_1415,N_723,In_1699);
or U1416 (N_1416,N_775,In_1779);
or U1417 (N_1417,N_657,N_547);
and U1418 (N_1418,N_524,N_705);
nor U1419 (N_1419,In_111,In_638);
xor U1420 (N_1420,N_210,N_501);
xor U1421 (N_1421,N_166,N_916);
or U1422 (N_1422,N_359,N_933);
and U1423 (N_1423,In_1794,N_720);
or U1424 (N_1424,In_1547,N_873);
xnor U1425 (N_1425,N_570,N_722);
nor U1426 (N_1426,N_180,N_858);
or U1427 (N_1427,N_508,N_898);
xnor U1428 (N_1428,N_322,N_127);
nor U1429 (N_1429,N_64,N_747);
or U1430 (N_1430,N_676,In_490);
nor U1431 (N_1431,N_539,N_939);
and U1432 (N_1432,N_284,N_936);
nor U1433 (N_1433,In_2,In_704);
nand U1434 (N_1434,N_751,In_1946);
nand U1435 (N_1435,N_973,N_855);
and U1436 (N_1436,In_579,In_1024);
and U1437 (N_1437,In_1272,N_669);
nor U1438 (N_1438,N_467,In_422);
xnor U1439 (N_1439,In_570,N_807);
or U1440 (N_1440,In_1973,N_497);
or U1441 (N_1441,In_627,In_1509);
and U1442 (N_1442,In_745,In_1040);
nor U1443 (N_1443,In_1840,N_995);
and U1444 (N_1444,N_471,N_620);
or U1445 (N_1445,N_999,In_1417);
and U1446 (N_1446,N_674,N_247);
or U1447 (N_1447,In_56,N_740);
xor U1448 (N_1448,N_336,N_866);
nor U1449 (N_1449,N_451,N_905);
or U1450 (N_1450,N_741,N_943);
nor U1451 (N_1451,N_748,In_658);
xor U1452 (N_1452,N_917,N_603);
nand U1453 (N_1453,N_458,N_930);
nand U1454 (N_1454,N_819,N_655);
or U1455 (N_1455,N_391,N_241);
nand U1456 (N_1456,N_838,In_1855);
nor U1457 (N_1457,In_1248,N_719);
or U1458 (N_1458,In_566,N_124);
xnor U1459 (N_1459,N_901,N_687);
xor U1460 (N_1460,N_888,N_418);
and U1461 (N_1461,N_668,N_695);
or U1462 (N_1462,N_889,N_782);
xor U1463 (N_1463,In_697,N_813);
and U1464 (N_1464,In_349,N_405);
or U1465 (N_1465,N_769,N_457);
nand U1466 (N_1466,N_385,N_516);
xor U1467 (N_1467,N_908,N_358);
or U1468 (N_1468,N_579,In_1274);
or U1469 (N_1469,N_843,In_493);
nand U1470 (N_1470,N_826,N_700);
xnor U1471 (N_1471,In_1601,N_168);
nand U1472 (N_1472,In_1582,N_541);
and U1473 (N_1473,In_530,N_89);
and U1474 (N_1474,In_1067,N_878);
nand U1475 (N_1475,N_711,N_968);
nand U1476 (N_1476,N_427,In_1119);
or U1477 (N_1477,N_820,In_793);
or U1478 (N_1478,N_985,N_590);
xnor U1479 (N_1479,N_575,N_867);
nand U1480 (N_1480,In_1506,In_173);
and U1481 (N_1481,N_523,N_364);
nand U1482 (N_1482,N_520,N_435);
and U1483 (N_1483,N_971,In_230);
nand U1484 (N_1484,N_891,N_618);
and U1485 (N_1485,N_765,N_715);
xnor U1486 (N_1486,N_264,In_189);
or U1487 (N_1487,In_911,N_773);
nor U1488 (N_1488,N_877,N_903);
and U1489 (N_1489,N_625,N_122);
xor U1490 (N_1490,N_783,In_512);
nand U1491 (N_1491,In_1663,In_581);
and U1492 (N_1492,In_1512,N_899);
xnor U1493 (N_1493,In_1996,N_744);
xor U1494 (N_1494,N_848,In_1134);
and U1495 (N_1495,N_721,N_294);
or U1496 (N_1496,N_645,N_143);
nand U1497 (N_1497,In_1963,N_93);
xor U1498 (N_1498,In_197,N_672);
and U1499 (N_1499,N_545,In_994);
or U1500 (N_1500,N_1413,N_1486);
or U1501 (N_1501,N_1176,N_1476);
or U1502 (N_1502,N_1110,N_1237);
xor U1503 (N_1503,N_1179,N_1243);
and U1504 (N_1504,N_1496,N_1226);
xnor U1505 (N_1505,N_1040,N_1172);
or U1506 (N_1506,N_1274,N_1078);
xor U1507 (N_1507,N_1264,N_1364);
xor U1508 (N_1508,N_1156,N_1347);
nand U1509 (N_1509,N_1444,N_1059);
or U1510 (N_1510,N_1038,N_1021);
or U1511 (N_1511,N_1007,N_1152);
nand U1512 (N_1512,N_1448,N_1189);
xnor U1513 (N_1513,N_1390,N_1341);
and U1514 (N_1514,N_1279,N_1062);
and U1515 (N_1515,N_1100,N_1463);
xnor U1516 (N_1516,N_1026,N_1308);
xnor U1517 (N_1517,N_1309,N_1254);
xor U1518 (N_1518,N_1103,N_1468);
or U1519 (N_1519,N_1410,N_1113);
or U1520 (N_1520,N_1003,N_1075);
nor U1521 (N_1521,N_1415,N_1092);
nand U1522 (N_1522,N_1411,N_1198);
and U1523 (N_1523,N_1029,N_1174);
nand U1524 (N_1524,N_1348,N_1057);
nor U1525 (N_1525,N_1447,N_1249);
and U1526 (N_1526,N_1036,N_1474);
or U1527 (N_1527,N_1127,N_1073);
nand U1528 (N_1528,N_1091,N_1184);
xnor U1529 (N_1529,N_1282,N_1423);
or U1530 (N_1530,N_1183,N_1216);
or U1531 (N_1531,N_1193,N_1461);
xor U1532 (N_1532,N_1061,N_1495);
xor U1533 (N_1533,N_1464,N_1039);
nand U1534 (N_1534,N_1335,N_1303);
or U1535 (N_1535,N_1241,N_1289);
nand U1536 (N_1536,N_1440,N_1164);
and U1537 (N_1537,N_1295,N_1351);
nand U1538 (N_1538,N_1436,N_1281);
and U1539 (N_1539,N_1354,N_1380);
nor U1540 (N_1540,N_1227,N_1481);
or U1541 (N_1541,N_1359,N_1235);
nor U1542 (N_1542,N_1162,N_1318);
and U1543 (N_1543,N_1201,N_1446);
and U1544 (N_1544,N_1072,N_1311);
and U1545 (N_1545,N_1493,N_1480);
nand U1546 (N_1546,N_1037,N_1370);
xor U1547 (N_1547,N_1208,N_1365);
and U1548 (N_1548,N_1117,N_1181);
xnor U1549 (N_1549,N_1104,N_1221);
and U1550 (N_1550,N_1171,N_1366);
xnor U1551 (N_1551,N_1149,N_1321);
and U1552 (N_1552,N_1324,N_1150);
xor U1553 (N_1553,N_1132,N_1025);
xnor U1554 (N_1554,N_1345,N_1420);
nor U1555 (N_1555,N_1031,N_1197);
and U1556 (N_1556,N_1097,N_1041);
and U1557 (N_1557,N_1027,N_1294);
or U1558 (N_1558,N_1369,N_1098);
nor U1559 (N_1559,N_1070,N_1261);
nor U1560 (N_1560,N_1142,N_1238);
nand U1561 (N_1561,N_1185,N_1044);
xor U1562 (N_1562,N_1310,N_1112);
and U1563 (N_1563,N_1213,N_1144);
xor U1564 (N_1564,N_1114,N_1232);
nor U1565 (N_1565,N_1192,N_1123);
nand U1566 (N_1566,N_1166,N_1450);
nor U1567 (N_1567,N_1313,N_1373);
nor U1568 (N_1568,N_1343,N_1256);
nor U1569 (N_1569,N_1383,N_1161);
xnor U1570 (N_1570,N_1317,N_1022);
nand U1571 (N_1571,N_1304,N_1405);
or U1572 (N_1572,N_1432,N_1404);
or U1573 (N_1573,N_1374,N_1377);
nor U1574 (N_1574,N_1401,N_1322);
nand U1575 (N_1575,N_1403,N_1080);
nand U1576 (N_1576,N_1290,N_1280);
nand U1577 (N_1577,N_1454,N_1427);
or U1578 (N_1578,N_1332,N_1473);
or U1579 (N_1579,N_1008,N_1252);
nand U1580 (N_1580,N_1260,N_1225);
or U1581 (N_1581,N_1387,N_1336);
or U1582 (N_1582,N_1167,N_1002);
nand U1583 (N_1583,N_1067,N_1083);
nand U1584 (N_1584,N_1076,N_1456);
nor U1585 (N_1585,N_1048,N_1023);
xnor U1586 (N_1586,N_1458,N_1173);
nor U1587 (N_1587,N_1168,N_1465);
nor U1588 (N_1588,N_1084,N_1485);
xor U1589 (N_1589,N_1498,N_1055);
nor U1590 (N_1590,N_1207,N_1269);
nor U1591 (N_1591,N_1270,N_1305);
nor U1592 (N_1592,N_1466,N_1094);
or U1593 (N_1593,N_1169,N_1014);
xnor U1594 (N_1594,N_1133,N_1071);
and U1595 (N_1595,N_1491,N_1268);
nand U1596 (N_1596,N_1375,N_1135);
nor U1597 (N_1597,N_1233,N_1372);
nor U1598 (N_1598,N_1439,N_1180);
nor U1599 (N_1599,N_1319,N_1276);
nand U1600 (N_1600,N_1064,N_1175);
nor U1601 (N_1601,N_1066,N_1312);
nor U1602 (N_1602,N_1361,N_1217);
or U1603 (N_1603,N_1384,N_1273);
xnor U1604 (N_1604,N_1316,N_1120);
or U1605 (N_1605,N_1222,N_1090);
xor U1606 (N_1606,N_1130,N_1326);
or U1607 (N_1607,N_1329,N_1340);
nor U1608 (N_1608,N_1015,N_1299);
nand U1609 (N_1609,N_1253,N_1125);
or U1610 (N_1610,N_1000,N_1388);
and U1611 (N_1611,N_1391,N_1407);
nor U1612 (N_1612,N_1054,N_1457);
nand U1613 (N_1613,N_1255,N_1490);
or U1614 (N_1614,N_1477,N_1460);
xnor U1615 (N_1615,N_1005,N_1393);
nand U1616 (N_1616,N_1052,N_1060);
nand U1617 (N_1617,N_1194,N_1355);
nand U1618 (N_1618,N_1165,N_1096);
and U1619 (N_1619,N_1042,N_1306);
xnor U1620 (N_1620,N_1385,N_1471);
nor U1621 (N_1621,N_1020,N_1275);
or U1622 (N_1622,N_1362,N_1065);
and U1623 (N_1623,N_1246,N_1399);
and U1624 (N_1624,N_1215,N_1497);
nor U1625 (N_1625,N_1089,N_1129);
xnor U1626 (N_1626,N_1445,N_1333);
nand U1627 (N_1627,N_1400,N_1344);
xnor U1628 (N_1628,N_1251,N_1301);
xor U1629 (N_1629,N_1224,N_1286);
nand U1630 (N_1630,N_1484,N_1105);
and U1631 (N_1631,N_1487,N_1392);
nor U1632 (N_1632,N_1155,N_1160);
nor U1633 (N_1633,N_1131,N_1302);
or U1634 (N_1634,N_1187,N_1267);
nand U1635 (N_1635,N_1479,N_1236);
nor U1636 (N_1636,N_1438,N_1019);
or U1637 (N_1637,N_1158,N_1297);
and U1638 (N_1638,N_1107,N_1462);
nor U1639 (N_1639,N_1430,N_1489);
or U1640 (N_1640,N_1240,N_1408);
nor U1641 (N_1641,N_1272,N_1327);
nand U1642 (N_1642,N_1367,N_1093);
and U1643 (N_1643,N_1102,N_1234);
or U1644 (N_1644,N_1209,N_1188);
or U1645 (N_1645,N_1368,N_1292);
or U1646 (N_1646,N_1079,N_1353);
or U1647 (N_1647,N_1121,N_1382);
nand U1648 (N_1648,N_1459,N_1013);
and U1649 (N_1649,N_1219,N_1146);
nand U1650 (N_1650,N_1032,N_1017);
nand U1651 (N_1651,N_1009,N_1035);
xnor U1652 (N_1652,N_1205,N_1346);
and U1653 (N_1653,N_1350,N_1196);
and U1654 (N_1654,N_1159,N_1378);
nand U1655 (N_1655,N_1425,N_1126);
nor U1656 (N_1656,N_1177,N_1379);
and U1657 (N_1657,N_1050,N_1074);
nand U1658 (N_1658,N_1431,N_1239);
nor U1659 (N_1659,N_1053,N_1056);
nand U1660 (N_1660,N_1178,N_1043);
and U1661 (N_1661,N_1470,N_1195);
xor U1662 (N_1662,N_1266,N_1262);
xor U1663 (N_1663,N_1394,N_1101);
xnor U1664 (N_1664,N_1320,N_1331);
or U1665 (N_1665,N_1141,N_1452);
nand U1666 (N_1666,N_1298,N_1287);
or U1667 (N_1667,N_1360,N_1030);
and U1668 (N_1668,N_1140,N_1284);
or U1669 (N_1669,N_1263,N_1277);
and U1670 (N_1670,N_1386,N_1285);
nand U1671 (N_1671,N_1069,N_1455);
or U1672 (N_1672,N_1244,N_1402);
and U1673 (N_1673,N_1492,N_1356);
xor U1674 (N_1674,N_1325,N_1218);
nor U1675 (N_1675,N_1242,N_1397);
and U1676 (N_1676,N_1106,N_1339);
nor U1677 (N_1677,N_1124,N_1257);
xor U1678 (N_1678,N_1398,N_1211);
nor U1679 (N_1679,N_1488,N_1229);
nor U1680 (N_1680,N_1451,N_1472);
and U1681 (N_1681,N_1191,N_1396);
nor U1682 (N_1682,N_1109,N_1006);
or U1683 (N_1683,N_1342,N_1422);
or U1684 (N_1684,N_1151,N_1139);
and U1685 (N_1685,N_1307,N_1338);
and U1686 (N_1686,N_1182,N_1190);
and U1687 (N_1687,N_1424,N_1300);
nor U1688 (N_1688,N_1001,N_1435);
nand U1689 (N_1689,N_1437,N_1247);
nor U1690 (N_1690,N_1482,N_1494);
and U1691 (N_1691,N_1330,N_1046);
nor U1692 (N_1692,N_1296,N_1137);
or U1693 (N_1693,N_1077,N_1442);
or U1694 (N_1694,N_1028,N_1063);
nor U1695 (N_1695,N_1337,N_1134);
nand U1696 (N_1696,N_1204,N_1047);
xnor U1697 (N_1697,N_1145,N_1115);
and U1698 (N_1698,N_1228,N_1418);
or U1699 (N_1699,N_1434,N_1004);
nor U1700 (N_1700,N_1406,N_1467);
nand U1701 (N_1701,N_1441,N_1250);
xnor U1702 (N_1702,N_1389,N_1163);
xnor U1703 (N_1703,N_1265,N_1118);
nor U1704 (N_1704,N_1016,N_1358);
nor U1705 (N_1705,N_1409,N_1099);
or U1706 (N_1706,N_1199,N_1010);
or U1707 (N_1707,N_1323,N_1315);
xor U1708 (N_1708,N_1412,N_1111);
nor U1709 (N_1709,N_1414,N_1283);
and U1710 (N_1710,N_1085,N_1258);
xor U1711 (N_1711,N_1186,N_1314);
xor U1712 (N_1712,N_1024,N_1475);
nand U1713 (N_1713,N_1148,N_1449);
xor U1714 (N_1714,N_1088,N_1352);
xor U1715 (N_1715,N_1011,N_1081);
nand U1716 (N_1716,N_1433,N_1453);
nand U1717 (N_1717,N_1293,N_1328);
xnor U1718 (N_1718,N_1428,N_1214);
and U1719 (N_1719,N_1245,N_1051);
and U1720 (N_1720,N_1202,N_1138);
nor U1721 (N_1721,N_1058,N_1483);
nand U1722 (N_1722,N_1068,N_1376);
and U1723 (N_1723,N_1095,N_1381);
or U1724 (N_1724,N_1116,N_1334);
xor U1725 (N_1725,N_1395,N_1012);
nor U1726 (N_1726,N_1018,N_1478);
nor U1727 (N_1727,N_1278,N_1154);
nand U1728 (N_1728,N_1033,N_1212);
and U1729 (N_1729,N_1421,N_1416);
xnor U1730 (N_1730,N_1170,N_1049);
nor U1731 (N_1731,N_1363,N_1417);
nand U1732 (N_1732,N_1371,N_1419);
xor U1733 (N_1733,N_1143,N_1119);
or U1734 (N_1734,N_1499,N_1157);
and U1735 (N_1735,N_1206,N_1248);
and U1736 (N_1736,N_1122,N_1136);
or U1737 (N_1737,N_1128,N_1223);
nor U1738 (N_1738,N_1357,N_1203);
nor U1739 (N_1739,N_1288,N_1147);
xor U1740 (N_1740,N_1469,N_1082);
or U1741 (N_1741,N_1349,N_1087);
xnor U1742 (N_1742,N_1153,N_1210);
and U1743 (N_1743,N_1034,N_1086);
nand U1744 (N_1744,N_1259,N_1443);
and U1745 (N_1745,N_1200,N_1429);
nor U1746 (N_1746,N_1271,N_1108);
nor U1747 (N_1747,N_1291,N_1231);
or U1748 (N_1748,N_1220,N_1045);
nor U1749 (N_1749,N_1230,N_1426);
and U1750 (N_1750,N_1073,N_1224);
nor U1751 (N_1751,N_1020,N_1351);
nor U1752 (N_1752,N_1399,N_1408);
xnor U1753 (N_1753,N_1183,N_1096);
nand U1754 (N_1754,N_1394,N_1424);
nor U1755 (N_1755,N_1310,N_1388);
xnor U1756 (N_1756,N_1107,N_1054);
nand U1757 (N_1757,N_1136,N_1356);
nor U1758 (N_1758,N_1218,N_1329);
or U1759 (N_1759,N_1206,N_1096);
or U1760 (N_1760,N_1300,N_1026);
nor U1761 (N_1761,N_1183,N_1415);
and U1762 (N_1762,N_1450,N_1237);
nand U1763 (N_1763,N_1450,N_1113);
or U1764 (N_1764,N_1091,N_1290);
nor U1765 (N_1765,N_1384,N_1014);
or U1766 (N_1766,N_1263,N_1444);
xor U1767 (N_1767,N_1218,N_1355);
or U1768 (N_1768,N_1121,N_1024);
or U1769 (N_1769,N_1356,N_1363);
nor U1770 (N_1770,N_1333,N_1230);
and U1771 (N_1771,N_1448,N_1251);
xnor U1772 (N_1772,N_1447,N_1363);
or U1773 (N_1773,N_1378,N_1333);
nor U1774 (N_1774,N_1215,N_1266);
nand U1775 (N_1775,N_1396,N_1056);
xnor U1776 (N_1776,N_1357,N_1317);
xnor U1777 (N_1777,N_1156,N_1146);
nor U1778 (N_1778,N_1240,N_1326);
nor U1779 (N_1779,N_1207,N_1359);
xor U1780 (N_1780,N_1018,N_1264);
nand U1781 (N_1781,N_1134,N_1256);
and U1782 (N_1782,N_1127,N_1202);
and U1783 (N_1783,N_1237,N_1285);
nand U1784 (N_1784,N_1121,N_1415);
or U1785 (N_1785,N_1028,N_1301);
nor U1786 (N_1786,N_1041,N_1370);
xor U1787 (N_1787,N_1097,N_1146);
xor U1788 (N_1788,N_1083,N_1454);
or U1789 (N_1789,N_1378,N_1183);
nand U1790 (N_1790,N_1466,N_1006);
xor U1791 (N_1791,N_1028,N_1341);
xnor U1792 (N_1792,N_1301,N_1372);
or U1793 (N_1793,N_1489,N_1236);
xnor U1794 (N_1794,N_1006,N_1078);
nor U1795 (N_1795,N_1185,N_1371);
nand U1796 (N_1796,N_1269,N_1487);
nor U1797 (N_1797,N_1404,N_1086);
and U1798 (N_1798,N_1041,N_1145);
nor U1799 (N_1799,N_1090,N_1406);
nand U1800 (N_1800,N_1196,N_1347);
and U1801 (N_1801,N_1012,N_1457);
xnor U1802 (N_1802,N_1094,N_1152);
xor U1803 (N_1803,N_1227,N_1247);
xor U1804 (N_1804,N_1376,N_1065);
and U1805 (N_1805,N_1258,N_1322);
nor U1806 (N_1806,N_1266,N_1149);
xor U1807 (N_1807,N_1287,N_1442);
or U1808 (N_1808,N_1068,N_1462);
and U1809 (N_1809,N_1187,N_1307);
nand U1810 (N_1810,N_1090,N_1316);
nor U1811 (N_1811,N_1154,N_1104);
or U1812 (N_1812,N_1486,N_1005);
nand U1813 (N_1813,N_1268,N_1167);
xor U1814 (N_1814,N_1480,N_1157);
and U1815 (N_1815,N_1295,N_1071);
or U1816 (N_1816,N_1428,N_1026);
nor U1817 (N_1817,N_1262,N_1302);
or U1818 (N_1818,N_1248,N_1048);
xnor U1819 (N_1819,N_1235,N_1290);
nor U1820 (N_1820,N_1400,N_1259);
and U1821 (N_1821,N_1322,N_1303);
nor U1822 (N_1822,N_1083,N_1262);
nand U1823 (N_1823,N_1072,N_1402);
nand U1824 (N_1824,N_1476,N_1168);
xnor U1825 (N_1825,N_1208,N_1154);
nand U1826 (N_1826,N_1313,N_1231);
and U1827 (N_1827,N_1289,N_1254);
nor U1828 (N_1828,N_1339,N_1419);
and U1829 (N_1829,N_1363,N_1145);
or U1830 (N_1830,N_1488,N_1057);
nor U1831 (N_1831,N_1198,N_1149);
nor U1832 (N_1832,N_1289,N_1474);
xnor U1833 (N_1833,N_1047,N_1002);
nand U1834 (N_1834,N_1473,N_1135);
and U1835 (N_1835,N_1222,N_1268);
nor U1836 (N_1836,N_1359,N_1401);
xnor U1837 (N_1837,N_1444,N_1403);
nor U1838 (N_1838,N_1320,N_1176);
and U1839 (N_1839,N_1341,N_1340);
nor U1840 (N_1840,N_1415,N_1205);
xor U1841 (N_1841,N_1269,N_1345);
or U1842 (N_1842,N_1165,N_1088);
nor U1843 (N_1843,N_1256,N_1168);
xor U1844 (N_1844,N_1354,N_1337);
nand U1845 (N_1845,N_1477,N_1254);
nand U1846 (N_1846,N_1083,N_1366);
and U1847 (N_1847,N_1159,N_1143);
or U1848 (N_1848,N_1431,N_1162);
and U1849 (N_1849,N_1000,N_1392);
or U1850 (N_1850,N_1190,N_1472);
nand U1851 (N_1851,N_1230,N_1346);
nand U1852 (N_1852,N_1052,N_1408);
or U1853 (N_1853,N_1499,N_1280);
or U1854 (N_1854,N_1014,N_1326);
xnor U1855 (N_1855,N_1089,N_1316);
or U1856 (N_1856,N_1162,N_1488);
nor U1857 (N_1857,N_1320,N_1039);
or U1858 (N_1858,N_1138,N_1080);
xor U1859 (N_1859,N_1341,N_1385);
nand U1860 (N_1860,N_1070,N_1045);
nor U1861 (N_1861,N_1156,N_1417);
xor U1862 (N_1862,N_1320,N_1268);
and U1863 (N_1863,N_1499,N_1310);
xor U1864 (N_1864,N_1328,N_1399);
nor U1865 (N_1865,N_1103,N_1318);
and U1866 (N_1866,N_1436,N_1315);
and U1867 (N_1867,N_1205,N_1095);
xor U1868 (N_1868,N_1295,N_1047);
or U1869 (N_1869,N_1210,N_1179);
or U1870 (N_1870,N_1211,N_1057);
and U1871 (N_1871,N_1184,N_1223);
and U1872 (N_1872,N_1009,N_1172);
xor U1873 (N_1873,N_1142,N_1135);
nor U1874 (N_1874,N_1123,N_1329);
or U1875 (N_1875,N_1193,N_1264);
xor U1876 (N_1876,N_1141,N_1001);
or U1877 (N_1877,N_1467,N_1082);
nand U1878 (N_1878,N_1453,N_1213);
and U1879 (N_1879,N_1314,N_1173);
nand U1880 (N_1880,N_1188,N_1030);
nand U1881 (N_1881,N_1016,N_1116);
nor U1882 (N_1882,N_1404,N_1111);
or U1883 (N_1883,N_1302,N_1330);
and U1884 (N_1884,N_1187,N_1252);
xor U1885 (N_1885,N_1416,N_1408);
nand U1886 (N_1886,N_1209,N_1229);
or U1887 (N_1887,N_1345,N_1168);
nand U1888 (N_1888,N_1415,N_1058);
xor U1889 (N_1889,N_1162,N_1198);
nand U1890 (N_1890,N_1455,N_1092);
nand U1891 (N_1891,N_1274,N_1150);
and U1892 (N_1892,N_1070,N_1400);
or U1893 (N_1893,N_1364,N_1498);
nor U1894 (N_1894,N_1393,N_1201);
nor U1895 (N_1895,N_1436,N_1152);
nor U1896 (N_1896,N_1325,N_1151);
xor U1897 (N_1897,N_1046,N_1203);
nor U1898 (N_1898,N_1007,N_1426);
nor U1899 (N_1899,N_1390,N_1303);
or U1900 (N_1900,N_1283,N_1319);
and U1901 (N_1901,N_1496,N_1472);
or U1902 (N_1902,N_1174,N_1033);
and U1903 (N_1903,N_1005,N_1389);
and U1904 (N_1904,N_1190,N_1401);
or U1905 (N_1905,N_1276,N_1030);
nand U1906 (N_1906,N_1401,N_1309);
or U1907 (N_1907,N_1196,N_1273);
nor U1908 (N_1908,N_1077,N_1090);
nand U1909 (N_1909,N_1121,N_1274);
nor U1910 (N_1910,N_1479,N_1298);
and U1911 (N_1911,N_1127,N_1108);
or U1912 (N_1912,N_1315,N_1485);
nor U1913 (N_1913,N_1088,N_1034);
xnor U1914 (N_1914,N_1413,N_1048);
and U1915 (N_1915,N_1277,N_1312);
nor U1916 (N_1916,N_1114,N_1493);
nand U1917 (N_1917,N_1251,N_1343);
nand U1918 (N_1918,N_1486,N_1409);
nand U1919 (N_1919,N_1013,N_1487);
or U1920 (N_1920,N_1208,N_1485);
or U1921 (N_1921,N_1113,N_1310);
xnor U1922 (N_1922,N_1321,N_1473);
xor U1923 (N_1923,N_1022,N_1223);
nor U1924 (N_1924,N_1353,N_1497);
nand U1925 (N_1925,N_1152,N_1463);
and U1926 (N_1926,N_1154,N_1389);
or U1927 (N_1927,N_1143,N_1391);
nand U1928 (N_1928,N_1038,N_1331);
xnor U1929 (N_1929,N_1090,N_1424);
nor U1930 (N_1930,N_1345,N_1424);
or U1931 (N_1931,N_1146,N_1397);
nand U1932 (N_1932,N_1411,N_1322);
xor U1933 (N_1933,N_1400,N_1047);
nor U1934 (N_1934,N_1417,N_1061);
nor U1935 (N_1935,N_1269,N_1095);
and U1936 (N_1936,N_1288,N_1278);
nor U1937 (N_1937,N_1499,N_1082);
nand U1938 (N_1938,N_1488,N_1278);
xnor U1939 (N_1939,N_1262,N_1132);
and U1940 (N_1940,N_1063,N_1212);
nand U1941 (N_1941,N_1300,N_1032);
and U1942 (N_1942,N_1058,N_1439);
or U1943 (N_1943,N_1382,N_1015);
xor U1944 (N_1944,N_1123,N_1006);
and U1945 (N_1945,N_1483,N_1258);
nand U1946 (N_1946,N_1246,N_1433);
or U1947 (N_1947,N_1137,N_1484);
or U1948 (N_1948,N_1388,N_1117);
or U1949 (N_1949,N_1143,N_1074);
or U1950 (N_1950,N_1159,N_1148);
and U1951 (N_1951,N_1157,N_1004);
and U1952 (N_1952,N_1244,N_1391);
and U1953 (N_1953,N_1110,N_1171);
and U1954 (N_1954,N_1067,N_1087);
xnor U1955 (N_1955,N_1341,N_1458);
or U1956 (N_1956,N_1048,N_1424);
xor U1957 (N_1957,N_1436,N_1335);
nand U1958 (N_1958,N_1385,N_1354);
and U1959 (N_1959,N_1213,N_1208);
nor U1960 (N_1960,N_1051,N_1054);
xnor U1961 (N_1961,N_1073,N_1077);
or U1962 (N_1962,N_1051,N_1006);
nand U1963 (N_1963,N_1319,N_1171);
or U1964 (N_1964,N_1227,N_1319);
nor U1965 (N_1965,N_1277,N_1396);
nand U1966 (N_1966,N_1007,N_1200);
nor U1967 (N_1967,N_1206,N_1183);
xor U1968 (N_1968,N_1381,N_1463);
xor U1969 (N_1969,N_1499,N_1031);
nor U1970 (N_1970,N_1354,N_1122);
xnor U1971 (N_1971,N_1454,N_1164);
and U1972 (N_1972,N_1142,N_1456);
and U1973 (N_1973,N_1277,N_1476);
nor U1974 (N_1974,N_1414,N_1483);
and U1975 (N_1975,N_1223,N_1451);
and U1976 (N_1976,N_1111,N_1155);
nand U1977 (N_1977,N_1241,N_1150);
xor U1978 (N_1978,N_1024,N_1003);
and U1979 (N_1979,N_1430,N_1358);
xor U1980 (N_1980,N_1275,N_1131);
nor U1981 (N_1981,N_1424,N_1287);
nor U1982 (N_1982,N_1205,N_1142);
or U1983 (N_1983,N_1017,N_1231);
and U1984 (N_1984,N_1005,N_1301);
or U1985 (N_1985,N_1431,N_1376);
nor U1986 (N_1986,N_1254,N_1259);
nand U1987 (N_1987,N_1390,N_1209);
nor U1988 (N_1988,N_1225,N_1406);
and U1989 (N_1989,N_1048,N_1092);
nor U1990 (N_1990,N_1116,N_1043);
nor U1991 (N_1991,N_1244,N_1020);
xnor U1992 (N_1992,N_1236,N_1008);
or U1993 (N_1993,N_1449,N_1067);
and U1994 (N_1994,N_1475,N_1389);
nor U1995 (N_1995,N_1457,N_1226);
xor U1996 (N_1996,N_1220,N_1359);
xnor U1997 (N_1997,N_1499,N_1129);
nor U1998 (N_1998,N_1287,N_1279);
nand U1999 (N_1999,N_1333,N_1467);
xnor U2000 (N_2000,N_1658,N_1643);
xor U2001 (N_2001,N_1539,N_1743);
and U2002 (N_2002,N_1890,N_1669);
nand U2003 (N_2003,N_1969,N_1674);
or U2004 (N_2004,N_1550,N_1945);
or U2005 (N_2005,N_1659,N_1966);
xor U2006 (N_2006,N_1955,N_1730);
or U2007 (N_2007,N_1874,N_1508);
nand U2008 (N_2008,N_1719,N_1615);
xor U2009 (N_2009,N_1897,N_1849);
or U2010 (N_2010,N_1698,N_1833);
and U2011 (N_2011,N_1650,N_1984);
and U2012 (N_2012,N_1645,N_1841);
xnor U2013 (N_2013,N_1559,N_1635);
nand U2014 (N_2014,N_1510,N_1552);
nor U2015 (N_2015,N_1830,N_1921);
and U2016 (N_2016,N_1706,N_1678);
or U2017 (N_2017,N_1912,N_1987);
and U2018 (N_2018,N_1600,N_1954);
xor U2019 (N_2019,N_1710,N_1862);
or U2020 (N_2020,N_1977,N_1699);
and U2021 (N_2021,N_1957,N_1813);
nor U2022 (N_2022,N_1863,N_1625);
nor U2023 (N_2023,N_1958,N_1622);
nand U2024 (N_2024,N_1795,N_1522);
and U2025 (N_2025,N_1629,N_1994);
xor U2026 (N_2026,N_1656,N_1758);
xor U2027 (N_2027,N_1762,N_1964);
or U2028 (N_2028,N_1616,N_1821);
xor U2029 (N_2029,N_1558,N_1648);
or U2030 (N_2030,N_1720,N_1634);
and U2031 (N_2031,N_1537,N_1940);
xnor U2032 (N_2032,N_1501,N_1746);
or U2033 (N_2033,N_1544,N_1968);
xnor U2034 (N_2034,N_1599,N_1823);
xor U2035 (N_2035,N_1563,N_1541);
nand U2036 (N_2036,N_1668,N_1651);
nor U2037 (N_2037,N_1690,N_1763);
nor U2038 (N_2038,N_1785,N_1637);
or U2039 (N_2039,N_1889,N_1827);
or U2040 (N_2040,N_1584,N_1524);
or U2041 (N_2041,N_1619,N_1594);
or U2042 (N_2042,N_1859,N_1775);
nor U2043 (N_2043,N_1755,N_1998);
nor U2044 (N_2044,N_1799,N_1923);
xnor U2045 (N_2045,N_1511,N_1893);
xnor U2046 (N_2046,N_1655,N_1902);
xor U2047 (N_2047,N_1670,N_1687);
nor U2048 (N_2048,N_1523,N_1515);
nand U2049 (N_2049,N_1694,N_1995);
and U2050 (N_2050,N_1744,N_1811);
or U2051 (N_2051,N_1514,N_1817);
and U2052 (N_2052,N_1895,N_1961);
or U2053 (N_2053,N_1723,N_1586);
or U2054 (N_2054,N_1748,N_1759);
nor U2055 (N_2055,N_1892,N_1636);
or U2056 (N_2056,N_1884,N_1596);
or U2057 (N_2057,N_1938,N_1567);
nand U2058 (N_2058,N_1836,N_1781);
or U2059 (N_2059,N_1916,N_1891);
or U2060 (N_2060,N_1920,N_1808);
and U2061 (N_2061,N_1624,N_1732);
nand U2062 (N_2062,N_1948,N_1547);
nand U2063 (N_2063,N_1734,N_1903);
xor U2064 (N_2064,N_1516,N_1826);
nand U2065 (N_2065,N_1975,N_1639);
or U2066 (N_2066,N_1810,N_1695);
nand U2067 (N_2067,N_1745,N_1926);
and U2068 (N_2068,N_1882,N_1803);
nand U2069 (N_2069,N_1804,N_1708);
and U2070 (N_2070,N_1500,N_1798);
nand U2071 (N_2071,N_1820,N_1854);
nand U2072 (N_2072,N_1910,N_1702);
or U2073 (N_2073,N_1992,N_1993);
nand U2074 (N_2074,N_1942,N_1953);
nor U2075 (N_2075,N_1727,N_1872);
nor U2076 (N_2076,N_1822,N_1664);
xnor U2077 (N_2077,N_1579,N_1780);
xnor U2078 (N_2078,N_1535,N_1856);
xnor U2079 (N_2079,N_1574,N_1869);
nor U2080 (N_2080,N_1649,N_1561);
and U2081 (N_2081,N_1627,N_1580);
nor U2082 (N_2082,N_1877,N_1517);
or U2083 (N_2083,N_1972,N_1828);
xnor U2084 (N_2084,N_1991,N_1733);
xor U2085 (N_2085,N_1838,N_1739);
or U2086 (N_2086,N_1576,N_1794);
nand U2087 (N_2087,N_1875,N_1566);
xor U2088 (N_2088,N_1887,N_1899);
or U2089 (N_2089,N_1800,N_1963);
and U2090 (N_2090,N_1617,N_1684);
or U2091 (N_2091,N_1738,N_1860);
and U2092 (N_2092,N_1531,N_1568);
and U2093 (N_2093,N_1513,N_1960);
and U2094 (N_2094,N_1852,N_1685);
xor U2095 (N_2095,N_1931,N_1604);
or U2096 (N_2096,N_1789,N_1693);
nor U2097 (N_2097,N_1613,N_1703);
or U2098 (N_2098,N_1638,N_1740);
nand U2099 (N_2099,N_1666,N_1512);
and U2100 (N_2100,N_1881,N_1915);
xor U2101 (N_2101,N_1707,N_1614);
and U2102 (N_2102,N_1598,N_1937);
or U2103 (N_2103,N_1952,N_1667);
nand U2104 (N_2104,N_1644,N_1592);
nand U2105 (N_2105,N_1990,N_1959);
nand U2106 (N_2106,N_1564,N_1533);
or U2107 (N_2107,N_1737,N_1979);
nand U2108 (N_2108,N_1560,N_1529);
or U2109 (N_2109,N_1878,N_1855);
nand U2110 (N_2110,N_1770,N_1816);
xor U2111 (N_2111,N_1769,N_1765);
nand U2112 (N_2112,N_1595,N_1534);
nand U2113 (N_2113,N_1741,N_1905);
and U2114 (N_2114,N_1831,N_1605);
or U2115 (N_2115,N_1686,N_1840);
nand U2116 (N_2116,N_1754,N_1705);
nor U2117 (N_2117,N_1851,N_1628);
xor U2118 (N_2118,N_1587,N_1936);
or U2119 (N_2119,N_1802,N_1502);
nor U2120 (N_2120,N_1554,N_1787);
xor U2121 (N_2121,N_1527,N_1725);
xor U2122 (N_2122,N_1988,N_1809);
and U2123 (N_2123,N_1825,N_1724);
nand U2124 (N_2124,N_1853,N_1562);
xor U2125 (N_2125,N_1914,N_1868);
or U2126 (N_2126,N_1601,N_1776);
or U2127 (N_2127,N_1525,N_1918);
nand U2128 (N_2128,N_1528,N_1555);
nand U2129 (N_2129,N_1908,N_1679);
nor U2130 (N_2130,N_1962,N_1578);
xnor U2131 (N_2131,N_1919,N_1760);
nand U2132 (N_2132,N_1753,N_1714);
and U2133 (N_2133,N_1997,N_1973);
or U2134 (N_2134,N_1581,N_1682);
and U2135 (N_2135,N_1929,N_1927);
nor U2136 (N_2136,N_1783,N_1688);
nor U2137 (N_2137,N_1689,N_1761);
and U2138 (N_2138,N_1711,N_1771);
xnor U2139 (N_2139,N_1640,N_1965);
xor U2140 (N_2140,N_1812,N_1607);
nand U2141 (N_2141,N_1848,N_1786);
or U2142 (N_2142,N_1709,N_1553);
xnor U2143 (N_2143,N_1548,N_1873);
xnor U2144 (N_2144,N_1538,N_1888);
or U2145 (N_2145,N_1967,N_1999);
nor U2146 (N_2146,N_1949,N_1835);
nand U2147 (N_2147,N_1571,N_1612);
xnor U2148 (N_2148,N_1509,N_1520);
or U2149 (N_2149,N_1925,N_1700);
xor U2150 (N_2150,N_1911,N_1844);
nand U2151 (N_2151,N_1526,N_1665);
xnor U2152 (N_2152,N_1570,N_1729);
or U2153 (N_2153,N_1573,N_1597);
or U2154 (N_2154,N_1909,N_1819);
xnor U2155 (N_2155,N_1557,N_1663);
nand U2156 (N_2156,N_1653,N_1657);
or U2157 (N_2157,N_1676,N_1536);
or U2158 (N_2158,N_1591,N_1671);
and U2159 (N_2159,N_1626,N_1660);
nand U2160 (N_2160,N_1572,N_1623);
or U2161 (N_2161,N_1867,N_1583);
or U2162 (N_2162,N_1503,N_1989);
or U2163 (N_2163,N_1641,N_1834);
xnor U2164 (N_2164,N_1716,N_1970);
nand U2165 (N_2165,N_1982,N_1519);
or U2166 (N_2166,N_1662,N_1824);
and U2167 (N_2167,N_1642,N_1551);
nor U2168 (N_2168,N_1815,N_1588);
nor U2169 (N_2169,N_1871,N_1589);
nor U2170 (N_2170,N_1749,N_1611);
or U2171 (N_2171,N_1784,N_1779);
and U2172 (N_2172,N_1506,N_1713);
xor U2173 (N_2173,N_1933,N_1518);
nor U2174 (N_2174,N_1843,N_1842);
or U2175 (N_2175,N_1565,N_1829);
xor U2176 (N_2176,N_1906,N_1778);
nand U2177 (N_2177,N_1752,N_1876);
and U2178 (N_2178,N_1814,N_1672);
and U2179 (N_2179,N_1864,N_1947);
nor U2180 (N_2180,N_1593,N_1898);
nor U2181 (N_2181,N_1850,N_1845);
xor U2182 (N_2182,N_1673,N_1807);
and U2183 (N_2183,N_1880,N_1545);
nand U2184 (N_2184,N_1913,N_1704);
nand U2185 (N_2185,N_1904,N_1943);
xnor U2186 (N_2186,N_1791,N_1652);
and U2187 (N_2187,N_1788,N_1900);
and U2188 (N_2188,N_1505,N_1736);
nand U2189 (N_2189,N_1722,N_1757);
nand U2190 (N_2190,N_1546,N_1974);
nor U2191 (N_2191,N_1896,N_1782);
and U2192 (N_2192,N_1647,N_1606);
nor U2193 (N_2193,N_1777,N_1712);
nand U2194 (N_2194,N_1901,N_1654);
and U2195 (N_2195,N_1944,N_1886);
or U2196 (N_2196,N_1747,N_1633);
and U2197 (N_2197,N_1774,N_1932);
xor U2198 (N_2198,N_1922,N_1806);
nor U2199 (N_2199,N_1618,N_1620);
xor U2200 (N_2200,N_1631,N_1773);
and U2201 (N_2201,N_1575,N_1728);
nand U2202 (N_2202,N_1764,N_1818);
and U2203 (N_2203,N_1677,N_1569);
and U2204 (N_2204,N_1696,N_1907);
and U2205 (N_2205,N_1832,N_1742);
nor U2206 (N_2206,N_1930,N_1766);
xnor U2207 (N_2207,N_1950,N_1585);
nor U2208 (N_2208,N_1981,N_1951);
xor U2209 (N_2209,N_1610,N_1885);
or U2210 (N_2210,N_1701,N_1879);
and U2211 (N_2211,N_1646,N_1680);
or U2212 (N_2212,N_1837,N_1621);
or U2213 (N_2213,N_1976,N_1796);
nor U2214 (N_2214,N_1590,N_1790);
or U2215 (N_2215,N_1630,N_1692);
nand U2216 (N_2216,N_1731,N_1756);
nand U2217 (N_2217,N_1996,N_1768);
xnor U2218 (N_2218,N_1521,N_1956);
and U2219 (N_2219,N_1939,N_1772);
nand U2220 (N_2220,N_1507,N_1717);
and U2221 (N_2221,N_1793,N_1532);
nand U2222 (N_2222,N_1540,N_1928);
and U2223 (N_2223,N_1917,N_1846);
and U2224 (N_2224,N_1847,N_1935);
xnor U2225 (N_2225,N_1697,N_1632);
and U2226 (N_2226,N_1735,N_1983);
xnor U2227 (N_2227,N_1675,N_1504);
xnor U2228 (N_2228,N_1602,N_1870);
nand U2229 (N_2229,N_1530,N_1718);
or U2230 (N_2230,N_1978,N_1985);
nand U2231 (N_2231,N_1894,N_1549);
and U2232 (N_2232,N_1858,N_1980);
or U2233 (N_2233,N_1866,N_1726);
nand U2234 (N_2234,N_1577,N_1805);
xnor U2235 (N_2235,N_1582,N_1556);
or U2236 (N_2236,N_1603,N_1934);
or U2237 (N_2237,N_1542,N_1751);
or U2238 (N_2238,N_1883,N_1721);
nor U2239 (N_2239,N_1683,N_1797);
and U2240 (N_2240,N_1865,N_1857);
or U2241 (N_2241,N_1661,N_1750);
or U2242 (N_2242,N_1767,N_1543);
nor U2243 (N_2243,N_1924,N_1839);
xnor U2244 (N_2244,N_1946,N_1691);
nand U2245 (N_2245,N_1681,N_1941);
or U2246 (N_2246,N_1971,N_1986);
or U2247 (N_2247,N_1792,N_1801);
nor U2248 (N_2248,N_1861,N_1608);
nand U2249 (N_2249,N_1609,N_1715);
nand U2250 (N_2250,N_1574,N_1737);
xor U2251 (N_2251,N_1579,N_1582);
nand U2252 (N_2252,N_1867,N_1659);
nor U2253 (N_2253,N_1687,N_1799);
nand U2254 (N_2254,N_1980,N_1591);
nand U2255 (N_2255,N_1979,N_1714);
nor U2256 (N_2256,N_1604,N_1881);
nand U2257 (N_2257,N_1651,N_1778);
and U2258 (N_2258,N_1648,N_1890);
and U2259 (N_2259,N_1733,N_1925);
and U2260 (N_2260,N_1725,N_1532);
and U2261 (N_2261,N_1801,N_1955);
or U2262 (N_2262,N_1567,N_1774);
xor U2263 (N_2263,N_1614,N_1569);
and U2264 (N_2264,N_1637,N_1522);
or U2265 (N_2265,N_1527,N_1649);
nand U2266 (N_2266,N_1890,N_1980);
nand U2267 (N_2267,N_1653,N_1576);
and U2268 (N_2268,N_1990,N_1613);
or U2269 (N_2269,N_1896,N_1808);
xnor U2270 (N_2270,N_1635,N_1855);
or U2271 (N_2271,N_1685,N_1968);
and U2272 (N_2272,N_1640,N_1962);
or U2273 (N_2273,N_1932,N_1872);
nor U2274 (N_2274,N_1600,N_1500);
nand U2275 (N_2275,N_1962,N_1644);
nor U2276 (N_2276,N_1786,N_1552);
nand U2277 (N_2277,N_1727,N_1928);
and U2278 (N_2278,N_1586,N_1791);
nand U2279 (N_2279,N_1684,N_1611);
nand U2280 (N_2280,N_1536,N_1926);
nor U2281 (N_2281,N_1685,N_1818);
nand U2282 (N_2282,N_1760,N_1610);
and U2283 (N_2283,N_1843,N_1920);
and U2284 (N_2284,N_1904,N_1514);
and U2285 (N_2285,N_1746,N_1945);
xor U2286 (N_2286,N_1950,N_1644);
xnor U2287 (N_2287,N_1663,N_1893);
xor U2288 (N_2288,N_1749,N_1573);
nand U2289 (N_2289,N_1873,N_1564);
xor U2290 (N_2290,N_1666,N_1899);
and U2291 (N_2291,N_1955,N_1862);
nand U2292 (N_2292,N_1587,N_1830);
nand U2293 (N_2293,N_1876,N_1554);
nand U2294 (N_2294,N_1708,N_1765);
xnor U2295 (N_2295,N_1560,N_1612);
and U2296 (N_2296,N_1658,N_1949);
or U2297 (N_2297,N_1655,N_1782);
nor U2298 (N_2298,N_1793,N_1894);
or U2299 (N_2299,N_1716,N_1710);
xor U2300 (N_2300,N_1929,N_1794);
xor U2301 (N_2301,N_1918,N_1531);
nor U2302 (N_2302,N_1940,N_1974);
or U2303 (N_2303,N_1622,N_1731);
nor U2304 (N_2304,N_1600,N_1961);
xnor U2305 (N_2305,N_1506,N_1787);
nor U2306 (N_2306,N_1537,N_1927);
nand U2307 (N_2307,N_1783,N_1880);
and U2308 (N_2308,N_1971,N_1627);
nor U2309 (N_2309,N_1693,N_1628);
and U2310 (N_2310,N_1912,N_1696);
nor U2311 (N_2311,N_1604,N_1812);
and U2312 (N_2312,N_1537,N_1949);
xor U2313 (N_2313,N_1594,N_1864);
xor U2314 (N_2314,N_1682,N_1864);
nor U2315 (N_2315,N_1552,N_1690);
and U2316 (N_2316,N_1679,N_1789);
nor U2317 (N_2317,N_1651,N_1542);
xnor U2318 (N_2318,N_1716,N_1637);
xnor U2319 (N_2319,N_1939,N_1713);
xor U2320 (N_2320,N_1892,N_1555);
nor U2321 (N_2321,N_1544,N_1528);
nor U2322 (N_2322,N_1759,N_1918);
xor U2323 (N_2323,N_1638,N_1703);
xnor U2324 (N_2324,N_1513,N_1872);
or U2325 (N_2325,N_1670,N_1828);
and U2326 (N_2326,N_1809,N_1734);
xor U2327 (N_2327,N_1937,N_1925);
and U2328 (N_2328,N_1501,N_1504);
nor U2329 (N_2329,N_1853,N_1867);
and U2330 (N_2330,N_1774,N_1792);
nor U2331 (N_2331,N_1525,N_1648);
and U2332 (N_2332,N_1921,N_1537);
xnor U2333 (N_2333,N_1846,N_1992);
nand U2334 (N_2334,N_1961,N_1646);
or U2335 (N_2335,N_1569,N_1658);
nor U2336 (N_2336,N_1801,N_1768);
and U2337 (N_2337,N_1541,N_1854);
xnor U2338 (N_2338,N_1677,N_1594);
and U2339 (N_2339,N_1739,N_1915);
xor U2340 (N_2340,N_1974,N_1680);
xor U2341 (N_2341,N_1865,N_1823);
or U2342 (N_2342,N_1818,N_1961);
and U2343 (N_2343,N_1703,N_1599);
and U2344 (N_2344,N_1979,N_1973);
xor U2345 (N_2345,N_1820,N_1880);
or U2346 (N_2346,N_1616,N_1615);
nand U2347 (N_2347,N_1721,N_1868);
xor U2348 (N_2348,N_1677,N_1835);
nand U2349 (N_2349,N_1640,N_1614);
or U2350 (N_2350,N_1537,N_1588);
or U2351 (N_2351,N_1522,N_1748);
or U2352 (N_2352,N_1829,N_1952);
and U2353 (N_2353,N_1995,N_1889);
nor U2354 (N_2354,N_1775,N_1747);
and U2355 (N_2355,N_1927,N_1989);
xor U2356 (N_2356,N_1927,N_1894);
and U2357 (N_2357,N_1745,N_1800);
nor U2358 (N_2358,N_1525,N_1915);
nand U2359 (N_2359,N_1746,N_1656);
nor U2360 (N_2360,N_1774,N_1815);
nand U2361 (N_2361,N_1500,N_1979);
or U2362 (N_2362,N_1959,N_1572);
or U2363 (N_2363,N_1545,N_1673);
or U2364 (N_2364,N_1583,N_1921);
and U2365 (N_2365,N_1529,N_1841);
xnor U2366 (N_2366,N_1897,N_1949);
nand U2367 (N_2367,N_1851,N_1874);
xor U2368 (N_2368,N_1528,N_1770);
or U2369 (N_2369,N_1920,N_1521);
xnor U2370 (N_2370,N_1924,N_1571);
xor U2371 (N_2371,N_1876,N_1946);
nor U2372 (N_2372,N_1567,N_1513);
and U2373 (N_2373,N_1685,N_1929);
nor U2374 (N_2374,N_1639,N_1856);
and U2375 (N_2375,N_1890,N_1941);
nor U2376 (N_2376,N_1823,N_1968);
or U2377 (N_2377,N_1740,N_1759);
or U2378 (N_2378,N_1802,N_1680);
and U2379 (N_2379,N_1899,N_1657);
nor U2380 (N_2380,N_1983,N_1913);
and U2381 (N_2381,N_1978,N_1521);
nor U2382 (N_2382,N_1530,N_1941);
xnor U2383 (N_2383,N_1686,N_1961);
xnor U2384 (N_2384,N_1981,N_1683);
nor U2385 (N_2385,N_1685,N_1840);
nand U2386 (N_2386,N_1551,N_1742);
and U2387 (N_2387,N_1611,N_1887);
and U2388 (N_2388,N_1679,N_1724);
or U2389 (N_2389,N_1900,N_1754);
xnor U2390 (N_2390,N_1924,N_1572);
xor U2391 (N_2391,N_1951,N_1527);
nand U2392 (N_2392,N_1751,N_1624);
xnor U2393 (N_2393,N_1608,N_1728);
nand U2394 (N_2394,N_1650,N_1689);
xor U2395 (N_2395,N_1744,N_1719);
and U2396 (N_2396,N_1727,N_1970);
nor U2397 (N_2397,N_1794,N_1820);
and U2398 (N_2398,N_1942,N_1543);
nand U2399 (N_2399,N_1813,N_1870);
and U2400 (N_2400,N_1587,N_1556);
and U2401 (N_2401,N_1670,N_1730);
or U2402 (N_2402,N_1608,N_1875);
or U2403 (N_2403,N_1536,N_1696);
nor U2404 (N_2404,N_1690,N_1743);
nor U2405 (N_2405,N_1608,N_1884);
xor U2406 (N_2406,N_1928,N_1940);
and U2407 (N_2407,N_1509,N_1901);
nor U2408 (N_2408,N_1784,N_1988);
xor U2409 (N_2409,N_1516,N_1794);
or U2410 (N_2410,N_1892,N_1982);
xnor U2411 (N_2411,N_1692,N_1640);
nand U2412 (N_2412,N_1664,N_1669);
xnor U2413 (N_2413,N_1502,N_1614);
nand U2414 (N_2414,N_1585,N_1855);
xnor U2415 (N_2415,N_1852,N_1920);
nand U2416 (N_2416,N_1799,N_1812);
nor U2417 (N_2417,N_1756,N_1767);
nand U2418 (N_2418,N_1625,N_1784);
xnor U2419 (N_2419,N_1899,N_1727);
and U2420 (N_2420,N_1828,N_1776);
xnor U2421 (N_2421,N_1540,N_1509);
or U2422 (N_2422,N_1639,N_1823);
and U2423 (N_2423,N_1704,N_1596);
and U2424 (N_2424,N_1701,N_1947);
and U2425 (N_2425,N_1571,N_1645);
nor U2426 (N_2426,N_1943,N_1877);
or U2427 (N_2427,N_1798,N_1825);
xnor U2428 (N_2428,N_1698,N_1515);
xnor U2429 (N_2429,N_1750,N_1545);
nand U2430 (N_2430,N_1655,N_1868);
or U2431 (N_2431,N_1682,N_1508);
xnor U2432 (N_2432,N_1888,N_1692);
nand U2433 (N_2433,N_1784,N_1832);
or U2434 (N_2434,N_1952,N_1725);
xnor U2435 (N_2435,N_1940,N_1767);
nand U2436 (N_2436,N_1534,N_1668);
or U2437 (N_2437,N_1930,N_1687);
xor U2438 (N_2438,N_1995,N_1862);
nor U2439 (N_2439,N_1805,N_1959);
and U2440 (N_2440,N_1924,N_1579);
and U2441 (N_2441,N_1503,N_1540);
and U2442 (N_2442,N_1756,N_1522);
nor U2443 (N_2443,N_1593,N_1737);
xnor U2444 (N_2444,N_1800,N_1545);
nor U2445 (N_2445,N_1934,N_1984);
xnor U2446 (N_2446,N_1804,N_1516);
nor U2447 (N_2447,N_1851,N_1770);
or U2448 (N_2448,N_1875,N_1501);
xor U2449 (N_2449,N_1780,N_1723);
nor U2450 (N_2450,N_1783,N_1943);
or U2451 (N_2451,N_1596,N_1795);
or U2452 (N_2452,N_1886,N_1707);
and U2453 (N_2453,N_1723,N_1968);
nor U2454 (N_2454,N_1553,N_1842);
or U2455 (N_2455,N_1698,N_1554);
nor U2456 (N_2456,N_1819,N_1648);
nand U2457 (N_2457,N_1765,N_1776);
or U2458 (N_2458,N_1599,N_1934);
or U2459 (N_2459,N_1880,N_1835);
xor U2460 (N_2460,N_1759,N_1684);
nor U2461 (N_2461,N_1856,N_1755);
nand U2462 (N_2462,N_1745,N_1731);
or U2463 (N_2463,N_1728,N_1983);
nand U2464 (N_2464,N_1695,N_1648);
nand U2465 (N_2465,N_1865,N_1817);
xnor U2466 (N_2466,N_1553,N_1948);
nand U2467 (N_2467,N_1734,N_1917);
nand U2468 (N_2468,N_1559,N_1550);
and U2469 (N_2469,N_1937,N_1523);
xnor U2470 (N_2470,N_1777,N_1995);
xnor U2471 (N_2471,N_1525,N_1991);
or U2472 (N_2472,N_1624,N_1833);
and U2473 (N_2473,N_1836,N_1728);
nor U2474 (N_2474,N_1980,N_1985);
and U2475 (N_2475,N_1776,N_1901);
or U2476 (N_2476,N_1801,N_1745);
nor U2477 (N_2477,N_1623,N_1664);
or U2478 (N_2478,N_1924,N_1545);
nor U2479 (N_2479,N_1541,N_1520);
or U2480 (N_2480,N_1783,N_1892);
or U2481 (N_2481,N_1724,N_1916);
nor U2482 (N_2482,N_1575,N_1566);
nor U2483 (N_2483,N_1778,N_1967);
and U2484 (N_2484,N_1752,N_1583);
or U2485 (N_2485,N_1522,N_1776);
xor U2486 (N_2486,N_1785,N_1828);
nand U2487 (N_2487,N_1790,N_1534);
xnor U2488 (N_2488,N_1979,N_1691);
nand U2489 (N_2489,N_1718,N_1746);
nand U2490 (N_2490,N_1912,N_1903);
xnor U2491 (N_2491,N_1535,N_1539);
and U2492 (N_2492,N_1959,N_1999);
or U2493 (N_2493,N_1664,N_1567);
xor U2494 (N_2494,N_1871,N_1677);
and U2495 (N_2495,N_1534,N_1917);
xnor U2496 (N_2496,N_1664,N_1960);
nor U2497 (N_2497,N_1504,N_1795);
nand U2498 (N_2498,N_1626,N_1558);
nor U2499 (N_2499,N_1714,N_1911);
nor U2500 (N_2500,N_2021,N_2156);
nor U2501 (N_2501,N_2121,N_2274);
or U2502 (N_2502,N_2016,N_2051);
or U2503 (N_2503,N_2480,N_2026);
nor U2504 (N_2504,N_2487,N_2437);
nor U2505 (N_2505,N_2246,N_2090);
or U2506 (N_2506,N_2429,N_2425);
xnor U2507 (N_2507,N_2332,N_2102);
and U2508 (N_2508,N_2066,N_2019);
nand U2509 (N_2509,N_2368,N_2142);
nor U2510 (N_2510,N_2493,N_2385);
nand U2511 (N_2511,N_2128,N_2290);
nor U2512 (N_2512,N_2123,N_2056);
nor U2513 (N_2513,N_2189,N_2285);
xor U2514 (N_2514,N_2125,N_2101);
xnor U2515 (N_2515,N_2243,N_2150);
nor U2516 (N_2516,N_2039,N_2229);
nor U2517 (N_2517,N_2457,N_2439);
or U2518 (N_2518,N_2009,N_2103);
and U2519 (N_2519,N_2374,N_2273);
nor U2520 (N_2520,N_2499,N_2052);
nor U2521 (N_2521,N_2436,N_2376);
nand U2522 (N_2522,N_2395,N_2187);
or U2523 (N_2523,N_2448,N_2244);
and U2524 (N_2524,N_2111,N_2108);
or U2525 (N_2525,N_2268,N_2151);
nor U2526 (N_2526,N_2441,N_2209);
nand U2527 (N_2527,N_2276,N_2269);
xnor U2528 (N_2528,N_2261,N_2099);
nor U2529 (N_2529,N_2232,N_2015);
nor U2530 (N_2530,N_2037,N_2221);
xnor U2531 (N_2531,N_2062,N_2422);
and U2532 (N_2532,N_2020,N_2494);
nor U2533 (N_2533,N_2396,N_2278);
nand U2534 (N_2534,N_2392,N_2450);
and U2535 (N_2535,N_2074,N_2069);
or U2536 (N_2536,N_2314,N_2418);
and U2537 (N_2537,N_2067,N_2444);
and U2538 (N_2538,N_2239,N_2098);
xnor U2539 (N_2539,N_2149,N_2137);
xor U2540 (N_2540,N_2033,N_2050);
nand U2541 (N_2541,N_2322,N_2479);
nor U2542 (N_2542,N_2485,N_2434);
and U2543 (N_2543,N_2346,N_2220);
and U2544 (N_2544,N_2207,N_2451);
nand U2545 (N_2545,N_2250,N_2370);
or U2546 (N_2546,N_2405,N_2011);
and U2547 (N_2547,N_2177,N_2400);
and U2548 (N_2548,N_2394,N_2185);
nand U2549 (N_2549,N_2198,N_2148);
nor U2550 (N_2550,N_2327,N_2204);
nand U2551 (N_2551,N_2159,N_2364);
or U2552 (N_2552,N_2470,N_2331);
nand U2553 (N_2553,N_2100,N_2416);
or U2554 (N_2554,N_2134,N_2265);
and U2555 (N_2555,N_2218,N_2203);
nor U2556 (N_2556,N_2191,N_2311);
nand U2557 (N_2557,N_2248,N_2296);
nand U2558 (N_2558,N_2180,N_2312);
nand U2559 (N_2559,N_2288,N_2181);
or U2560 (N_2560,N_2133,N_2300);
or U2561 (N_2561,N_2294,N_2302);
nand U2562 (N_2562,N_2162,N_2000);
and U2563 (N_2563,N_2379,N_2305);
nand U2564 (N_2564,N_2028,N_2393);
or U2565 (N_2565,N_2467,N_2030);
and U2566 (N_2566,N_2006,N_2138);
nand U2567 (N_2567,N_2184,N_2168);
or U2568 (N_2568,N_2275,N_2061);
or U2569 (N_2569,N_2462,N_2147);
xor U2570 (N_2570,N_2118,N_2017);
nor U2571 (N_2571,N_2064,N_2043);
and U2572 (N_2572,N_2366,N_2386);
nor U2573 (N_2573,N_2131,N_2365);
nor U2574 (N_2574,N_2266,N_2035);
xnor U2575 (N_2575,N_2421,N_2157);
nor U2576 (N_2576,N_2308,N_2389);
and U2577 (N_2577,N_2072,N_2349);
xor U2578 (N_2578,N_2027,N_2235);
and U2579 (N_2579,N_2415,N_2040);
nor U2580 (N_2580,N_2330,N_2258);
nand U2581 (N_2581,N_2486,N_2446);
nor U2582 (N_2582,N_2110,N_2169);
nor U2583 (N_2583,N_2424,N_2048);
nor U2584 (N_2584,N_2292,N_2183);
xor U2585 (N_2585,N_2371,N_2438);
nand U2586 (N_2586,N_2497,N_2054);
nor U2587 (N_2587,N_2233,N_2245);
nand U2588 (N_2588,N_2242,N_2076);
and U2589 (N_2589,N_2464,N_2155);
and U2590 (N_2590,N_2046,N_2139);
nor U2591 (N_2591,N_2409,N_2193);
xnor U2592 (N_2592,N_2211,N_2080);
nor U2593 (N_2593,N_2075,N_2401);
nor U2594 (N_2594,N_2283,N_2380);
xnor U2595 (N_2595,N_2321,N_2045);
or U2596 (N_2596,N_2141,N_2445);
and U2597 (N_2597,N_2166,N_2483);
xnor U2598 (N_2598,N_2031,N_2154);
nand U2599 (N_2599,N_2260,N_2105);
nor U2600 (N_2600,N_2022,N_2124);
nor U2601 (N_2601,N_2328,N_2354);
nor U2602 (N_2602,N_2230,N_2489);
nor U2603 (N_2603,N_2025,N_2143);
xnor U2604 (N_2604,N_2454,N_2014);
or U2605 (N_2605,N_2295,N_2478);
nor U2606 (N_2606,N_2092,N_2406);
nand U2607 (N_2607,N_2091,N_2329);
or U2608 (N_2608,N_2362,N_2315);
and U2609 (N_2609,N_2176,N_2058);
and U2610 (N_2610,N_2114,N_2428);
or U2611 (N_2611,N_2231,N_2469);
nand U2612 (N_2612,N_2047,N_2381);
nor U2613 (N_2613,N_2281,N_2414);
nor U2614 (N_2614,N_2316,N_2094);
xor U2615 (N_2615,N_2456,N_2347);
xnor U2616 (N_2616,N_2299,N_2471);
xnor U2617 (N_2617,N_2303,N_2431);
nor U2618 (N_2618,N_2356,N_2367);
nor U2619 (N_2619,N_2034,N_2144);
or U2620 (N_2620,N_2167,N_2267);
xnor U2621 (N_2621,N_2065,N_2241);
nand U2622 (N_2622,N_2213,N_2369);
and U2623 (N_2623,N_2093,N_2490);
nor U2624 (N_2624,N_2112,N_2382);
and U2625 (N_2625,N_2289,N_2391);
nor U2626 (N_2626,N_2357,N_2145);
xor U2627 (N_2627,N_2284,N_2277);
and U2628 (N_2628,N_2481,N_2287);
nand U2629 (N_2629,N_2097,N_2377);
nor U2630 (N_2630,N_2440,N_2461);
nor U2631 (N_2631,N_2326,N_2498);
and U2632 (N_2632,N_2003,N_2082);
or U2633 (N_2633,N_2373,N_2247);
xor U2634 (N_2634,N_2307,N_2126);
xnor U2635 (N_2635,N_2472,N_2200);
and U2636 (N_2636,N_2443,N_2004);
or U2637 (N_2637,N_2104,N_2345);
and U2638 (N_2638,N_2175,N_2343);
nor U2639 (N_2639,N_2334,N_2317);
nor U2640 (N_2640,N_2419,N_2130);
nand U2641 (N_2641,N_2106,N_2081);
and U2642 (N_2642,N_2383,N_2353);
nand U2643 (N_2643,N_2412,N_2073);
nand U2644 (N_2644,N_2163,N_2029);
xor U2645 (N_2645,N_2205,N_2227);
nor U2646 (N_2646,N_2442,N_2199);
or U2647 (N_2647,N_2378,N_2077);
xor U2648 (N_2648,N_2358,N_2254);
or U2649 (N_2649,N_2182,N_2466);
nor U2650 (N_2650,N_2279,N_2234);
nand U2651 (N_2651,N_2397,N_2116);
xor U2652 (N_2652,N_2161,N_2088);
xnor U2653 (N_2653,N_2060,N_2018);
nor U2654 (N_2654,N_2120,N_2049);
or U2655 (N_2655,N_2070,N_2262);
and U2656 (N_2656,N_2482,N_2172);
nand U2657 (N_2657,N_2463,N_2236);
xor U2658 (N_2658,N_2491,N_2348);
nand U2659 (N_2659,N_2320,N_2053);
nand U2660 (N_2660,N_2170,N_2360);
nand U2661 (N_2661,N_2132,N_2055);
xor U2662 (N_2662,N_2251,N_2257);
nand U2663 (N_2663,N_2350,N_2372);
nor U2664 (N_2664,N_2410,N_2044);
xnor U2665 (N_2665,N_2146,N_2324);
or U2666 (N_2666,N_2336,N_2313);
or U2667 (N_2667,N_2115,N_2340);
xor U2668 (N_2668,N_2224,N_2476);
or U2669 (N_2669,N_2122,N_2083);
or U2670 (N_2670,N_2012,N_2459);
xnor U2671 (N_2671,N_2192,N_2452);
xor U2672 (N_2672,N_2086,N_2407);
xnor U2673 (N_2673,N_2351,N_2319);
nand U2674 (N_2674,N_2223,N_2335);
nor U2675 (N_2675,N_2024,N_2488);
nor U2676 (N_2676,N_2399,N_2007);
nor U2677 (N_2677,N_2252,N_2363);
xor U2678 (N_2678,N_2474,N_2013);
nand U2679 (N_2679,N_2484,N_2071);
nand U2680 (N_2680,N_2270,N_2427);
or U2681 (N_2681,N_2085,N_2129);
nand U2682 (N_2682,N_2460,N_2160);
nand U2683 (N_2683,N_2352,N_2339);
or U2684 (N_2684,N_2178,N_2453);
nand U2685 (N_2685,N_2008,N_2465);
nand U2686 (N_2686,N_2206,N_2164);
xor U2687 (N_2687,N_2318,N_2310);
and U2688 (N_2688,N_2225,N_2256);
nand U2689 (N_2689,N_2002,N_2238);
or U2690 (N_2690,N_2195,N_2495);
xor U2691 (N_2691,N_2304,N_2286);
nand U2692 (N_2692,N_2216,N_2113);
xnor U2693 (N_2693,N_2153,N_2387);
or U2694 (N_2694,N_2240,N_2344);
and U2695 (N_2695,N_2001,N_2194);
and U2696 (N_2696,N_2219,N_2468);
nand U2697 (N_2697,N_2190,N_2117);
xnor U2698 (N_2698,N_2271,N_2398);
and U2699 (N_2699,N_2068,N_2402);
xor U2700 (N_2700,N_2388,N_2447);
or U2701 (N_2701,N_2165,N_2095);
or U2702 (N_2702,N_2323,N_2403);
xnor U2703 (N_2703,N_2337,N_2127);
or U2704 (N_2704,N_2084,N_2210);
nor U2705 (N_2705,N_2171,N_2449);
nand U2706 (N_2706,N_2222,N_2038);
xor U2707 (N_2707,N_2023,N_2306);
nand U2708 (N_2708,N_2384,N_2390);
nor U2709 (N_2709,N_2263,N_2215);
and U2710 (N_2710,N_2433,N_2423);
and U2711 (N_2711,N_2041,N_2059);
and U2712 (N_2712,N_2341,N_2087);
nor U2713 (N_2713,N_2492,N_2355);
and U2714 (N_2714,N_2136,N_2253);
or U2715 (N_2715,N_2036,N_2455);
or U2716 (N_2716,N_2214,N_2338);
xor U2717 (N_2717,N_2107,N_2226);
and U2718 (N_2718,N_2140,N_2197);
or U2719 (N_2719,N_2359,N_2426);
and U2720 (N_2720,N_2411,N_2473);
nor U2721 (N_2721,N_2417,N_2096);
nand U2722 (N_2722,N_2089,N_2158);
or U2723 (N_2723,N_2293,N_2301);
nor U2724 (N_2724,N_2063,N_2196);
nor U2725 (N_2725,N_2430,N_2217);
or U2726 (N_2726,N_2325,N_2435);
xnor U2727 (N_2727,N_2282,N_2475);
nor U2728 (N_2728,N_2259,N_2135);
nand U2729 (N_2729,N_2408,N_2309);
nor U2730 (N_2730,N_2208,N_2010);
and U2731 (N_2731,N_2477,N_2202);
or U2732 (N_2732,N_2255,N_2079);
or U2733 (N_2733,N_2057,N_2174);
nand U2734 (N_2734,N_2298,N_2032);
xor U2735 (N_2735,N_2375,N_2264);
nor U2736 (N_2736,N_2297,N_2361);
nor U2737 (N_2737,N_2272,N_2458);
nand U2738 (N_2738,N_2342,N_2420);
nor U2739 (N_2739,N_2413,N_2291);
xor U2740 (N_2740,N_2237,N_2173);
xor U2741 (N_2741,N_2201,N_2119);
xor U2742 (N_2742,N_2432,N_2188);
nor U2743 (N_2743,N_2078,N_2005);
xnor U2744 (N_2744,N_2186,N_2280);
or U2745 (N_2745,N_2179,N_2212);
nor U2746 (N_2746,N_2109,N_2249);
and U2747 (N_2747,N_2152,N_2228);
xnor U2748 (N_2748,N_2404,N_2333);
xor U2749 (N_2749,N_2042,N_2496);
or U2750 (N_2750,N_2377,N_2160);
and U2751 (N_2751,N_2104,N_2146);
nor U2752 (N_2752,N_2098,N_2471);
or U2753 (N_2753,N_2303,N_2152);
nor U2754 (N_2754,N_2037,N_2050);
and U2755 (N_2755,N_2276,N_2110);
xnor U2756 (N_2756,N_2441,N_2374);
nand U2757 (N_2757,N_2387,N_2272);
nand U2758 (N_2758,N_2320,N_2314);
nand U2759 (N_2759,N_2400,N_2097);
or U2760 (N_2760,N_2147,N_2471);
xor U2761 (N_2761,N_2200,N_2104);
xnor U2762 (N_2762,N_2230,N_2452);
and U2763 (N_2763,N_2043,N_2307);
nand U2764 (N_2764,N_2033,N_2299);
nor U2765 (N_2765,N_2081,N_2026);
nor U2766 (N_2766,N_2055,N_2285);
nand U2767 (N_2767,N_2363,N_2178);
nand U2768 (N_2768,N_2108,N_2345);
nand U2769 (N_2769,N_2469,N_2036);
xnor U2770 (N_2770,N_2294,N_2117);
nor U2771 (N_2771,N_2182,N_2428);
nand U2772 (N_2772,N_2090,N_2191);
xnor U2773 (N_2773,N_2344,N_2407);
xnor U2774 (N_2774,N_2211,N_2008);
or U2775 (N_2775,N_2367,N_2477);
nor U2776 (N_2776,N_2427,N_2117);
nor U2777 (N_2777,N_2494,N_2117);
xor U2778 (N_2778,N_2149,N_2251);
nor U2779 (N_2779,N_2163,N_2015);
nand U2780 (N_2780,N_2292,N_2333);
xor U2781 (N_2781,N_2195,N_2362);
or U2782 (N_2782,N_2422,N_2328);
or U2783 (N_2783,N_2255,N_2055);
nor U2784 (N_2784,N_2380,N_2051);
nor U2785 (N_2785,N_2015,N_2220);
xnor U2786 (N_2786,N_2198,N_2331);
xor U2787 (N_2787,N_2259,N_2371);
xor U2788 (N_2788,N_2314,N_2374);
nor U2789 (N_2789,N_2071,N_2180);
nor U2790 (N_2790,N_2476,N_2022);
nor U2791 (N_2791,N_2248,N_2221);
and U2792 (N_2792,N_2470,N_2094);
nand U2793 (N_2793,N_2112,N_2029);
nand U2794 (N_2794,N_2300,N_2009);
nor U2795 (N_2795,N_2064,N_2314);
nand U2796 (N_2796,N_2127,N_2136);
xnor U2797 (N_2797,N_2039,N_2369);
nand U2798 (N_2798,N_2125,N_2290);
nand U2799 (N_2799,N_2485,N_2307);
xnor U2800 (N_2800,N_2495,N_2358);
or U2801 (N_2801,N_2447,N_2027);
or U2802 (N_2802,N_2064,N_2026);
nor U2803 (N_2803,N_2332,N_2128);
and U2804 (N_2804,N_2328,N_2180);
nor U2805 (N_2805,N_2388,N_2463);
xnor U2806 (N_2806,N_2101,N_2029);
xor U2807 (N_2807,N_2424,N_2140);
xnor U2808 (N_2808,N_2498,N_2439);
xor U2809 (N_2809,N_2005,N_2339);
nor U2810 (N_2810,N_2172,N_2124);
nand U2811 (N_2811,N_2272,N_2244);
xor U2812 (N_2812,N_2007,N_2445);
and U2813 (N_2813,N_2493,N_2423);
nor U2814 (N_2814,N_2488,N_2010);
or U2815 (N_2815,N_2120,N_2103);
nor U2816 (N_2816,N_2165,N_2489);
or U2817 (N_2817,N_2034,N_2419);
and U2818 (N_2818,N_2271,N_2043);
xor U2819 (N_2819,N_2385,N_2145);
nor U2820 (N_2820,N_2339,N_2073);
xor U2821 (N_2821,N_2089,N_2106);
nand U2822 (N_2822,N_2372,N_2313);
xor U2823 (N_2823,N_2298,N_2029);
nand U2824 (N_2824,N_2099,N_2422);
nor U2825 (N_2825,N_2255,N_2172);
xor U2826 (N_2826,N_2232,N_2484);
nand U2827 (N_2827,N_2230,N_2226);
and U2828 (N_2828,N_2439,N_2074);
nor U2829 (N_2829,N_2266,N_2221);
or U2830 (N_2830,N_2388,N_2053);
nor U2831 (N_2831,N_2447,N_2137);
nand U2832 (N_2832,N_2162,N_2454);
nand U2833 (N_2833,N_2349,N_2291);
or U2834 (N_2834,N_2302,N_2415);
nand U2835 (N_2835,N_2389,N_2316);
xnor U2836 (N_2836,N_2320,N_2034);
xnor U2837 (N_2837,N_2028,N_2410);
and U2838 (N_2838,N_2193,N_2240);
and U2839 (N_2839,N_2044,N_2178);
and U2840 (N_2840,N_2106,N_2174);
and U2841 (N_2841,N_2007,N_2292);
and U2842 (N_2842,N_2430,N_2181);
nand U2843 (N_2843,N_2280,N_2388);
and U2844 (N_2844,N_2145,N_2120);
xnor U2845 (N_2845,N_2455,N_2217);
or U2846 (N_2846,N_2484,N_2046);
xor U2847 (N_2847,N_2376,N_2263);
xor U2848 (N_2848,N_2479,N_2028);
and U2849 (N_2849,N_2186,N_2260);
or U2850 (N_2850,N_2180,N_2066);
nand U2851 (N_2851,N_2282,N_2404);
or U2852 (N_2852,N_2288,N_2434);
nor U2853 (N_2853,N_2449,N_2384);
and U2854 (N_2854,N_2308,N_2490);
or U2855 (N_2855,N_2371,N_2275);
nand U2856 (N_2856,N_2440,N_2103);
xnor U2857 (N_2857,N_2287,N_2115);
and U2858 (N_2858,N_2165,N_2082);
or U2859 (N_2859,N_2360,N_2160);
nand U2860 (N_2860,N_2394,N_2487);
or U2861 (N_2861,N_2421,N_2101);
xnor U2862 (N_2862,N_2078,N_2171);
nand U2863 (N_2863,N_2275,N_2464);
or U2864 (N_2864,N_2103,N_2322);
nor U2865 (N_2865,N_2273,N_2364);
nor U2866 (N_2866,N_2295,N_2290);
nor U2867 (N_2867,N_2101,N_2188);
and U2868 (N_2868,N_2059,N_2264);
xor U2869 (N_2869,N_2328,N_2375);
or U2870 (N_2870,N_2409,N_2391);
nand U2871 (N_2871,N_2095,N_2317);
or U2872 (N_2872,N_2436,N_2292);
xor U2873 (N_2873,N_2048,N_2198);
nor U2874 (N_2874,N_2402,N_2261);
nand U2875 (N_2875,N_2128,N_2083);
xor U2876 (N_2876,N_2051,N_2019);
nand U2877 (N_2877,N_2057,N_2155);
or U2878 (N_2878,N_2475,N_2291);
xnor U2879 (N_2879,N_2316,N_2001);
nor U2880 (N_2880,N_2390,N_2163);
or U2881 (N_2881,N_2022,N_2038);
and U2882 (N_2882,N_2066,N_2398);
nand U2883 (N_2883,N_2183,N_2115);
and U2884 (N_2884,N_2019,N_2119);
and U2885 (N_2885,N_2247,N_2128);
xnor U2886 (N_2886,N_2362,N_2139);
nand U2887 (N_2887,N_2288,N_2207);
and U2888 (N_2888,N_2342,N_2170);
xor U2889 (N_2889,N_2159,N_2304);
nor U2890 (N_2890,N_2317,N_2185);
or U2891 (N_2891,N_2091,N_2133);
or U2892 (N_2892,N_2207,N_2117);
or U2893 (N_2893,N_2188,N_2139);
and U2894 (N_2894,N_2357,N_2271);
and U2895 (N_2895,N_2129,N_2150);
and U2896 (N_2896,N_2310,N_2262);
or U2897 (N_2897,N_2045,N_2229);
nor U2898 (N_2898,N_2117,N_2236);
and U2899 (N_2899,N_2194,N_2461);
nand U2900 (N_2900,N_2066,N_2298);
xnor U2901 (N_2901,N_2051,N_2059);
nand U2902 (N_2902,N_2452,N_2283);
xor U2903 (N_2903,N_2050,N_2134);
nor U2904 (N_2904,N_2014,N_2295);
or U2905 (N_2905,N_2047,N_2481);
nor U2906 (N_2906,N_2151,N_2235);
nand U2907 (N_2907,N_2171,N_2486);
xnor U2908 (N_2908,N_2298,N_2479);
or U2909 (N_2909,N_2261,N_2165);
and U2910 (N_2910,N_2396,N_2326);
and U2911 (N_2911,N_2130,N_2451);
xor U2912 (N_2912,N_2124,N_2402);
and U2913 (N_2913,N_2431,N_2193);
or U2914 (N_2914,N_2332,N_2424);
xor U2915 (N_2915,N_2258,N_2238);
xor U2916 (N_2916,N_2353,N_2182);
and U2917 (N_2917,N_2022,N_2490);
xnor U2918 (N_2918,N_2454,N_2231);
and U2919 (N_2919,N_2291,N_2465);
nand U2920 (N_2920,N_2333,N_2037);
nand U2921 (N_2921,N_2073,N_2029);
nor U2922 (N_2922,N_2025,N_2186);
xor U2923 (N_2923,N_2098,N_2235);
or U2924 (N_2924,N_2460,N_2052);
nand U2925 (N_2925,N_2229,N_2496);
and U2926 (N_2926,N_2432,N_2490);
nor U2927 (N_2927,N_2206,N_2035);
or U2928 (N_2928,N_2417,N_2274);
and U2929 (N_2929,N_2004,N_2307);
nand U2930 (N_2930,N_2227,N_2427);
and U2931 (N_2931,N_2084,N_2285);
and U2932 (N_2932,N_2144,N_2153);
nand U2933 (N_2933,N_2387,N_2474);
nand U2934 (N_2934,N_2444,N_2363);
nand U2935 (N_2935,N_2269,N_2362);
and U2936 (N_2936,N_2292,N_2413);
nand U2937 (N_2937,N_2087,N_2226);
xor U2938 (N_2938,N_2373,N_2139);
nor U2939 (N_2939,N_2331,N_2454);
xnor U2940 (N_2940,N_2068,N_2434);
or U2941 (N_2941,N_2225,N_2116);
and U2942 (N_2942,N_2477,N_2349);
xor U2943 (N_2943,N_2354,N_2302);
xor U2944 (N_2944,N_2024,N_2008);
and U2945 (N_2945,N_2455,N_2049);
and U2946 (N_2946,N_2085,N_2430);
and U2947 (N_2947,N_2302,N_2471);
xnor U2948 (N_2948,N_2269,N_2207);
or U2949 (N_2949,N_2224,N_2176);
xnor U2950 (N_2950,N_2199,N_2290);
nand U2951 (N_2951,N_2466,N_2382);
nand U2952 (N_2952,N_2374,N_2464);
nor U2953 (N_2953,N_2031,N_2298);
xor U2954 (N_2954,N_2440,N_2023);
nor U2955 (N_2955,N_2257,N_2268);
or U2956 (N_2956,N_2460,N_2448);
xor U2957 (N_2957,N_2181,N_2403);
xor U2958 (N_2958,N_2164,N_2065);
nor U2959 (N_2959,N_2045,N_2424);
and U2960 (N_2960,N_2359,N_2238);
nor U2961 (N_2961,N_2348,N_2368);
and U2962 (N_2962,N_2494,N_2200);
nor U2963 (N_2963,N_2214,N_2368);
or U2964 (N_2964,N_2119,N_2348);
or U2965 (N_2965,N_2183,N_2332);
and U2966 (N_2966,N_2142,N_2056);
or U2967 (N_2967,N_2482,N_2194);
xor U2968 (N_2968,N_2200,N_2016);
nand U2969 (N_2969,N_2026,N_2405);
or U2970 (N_2970,N_2137,N_2396);
and U2971 (N_2971,N_2143,N_2488);
xnor U2972 (N_2972,N_2342,N_2057);
or U2973 (N_2973,N_2328,N_2353);
and U2974 (N_2974,N_2281,N_2154);
or U2975 (N_2975,N_2209,N_2331);
xor U2976 (N_2976,N_2461,N_2363);
nor U2977 (N_2977,N_2473,N_2102);
nand U2978 (N_2978,N_2162,N_2080);
and U2979 (N_2979,N_2047,N_2044);
xor U2980 (N_2980,N_2422,N_2221);
xnor U2981 (N_2981,N_2152,N_2048);
or U2982 (N_2982,N_2071,N_2367);
nand U2983 (N_2983,N_2447,N_2124);
and U2984 (N_2984,N_2093,N_2394);
xor U2985 (N_2985,N_2197,N_2027);
or U2986 (N_2986,N_2084,N_2439);
xnor U2987 (N_2987,N_2217,N_2182);
nand U2988 (N_2988,N_2192,N_2031);
nor U2989 (N_2989,N_2152,N_2160);
or U2990 (N_2990,N_2104,N_2312);
and U2991 (N_2991,N_2107,N_2327);
xor U2992 (N_2992,N_2428,N_2226);
xor U2993 (N_2993,N_2042,N_2211);
xnor U2994 (N_2994,N_2491,N_2072);
nor U2995 (N_2995,N_2101,N_2446);
nor U2996 (N_2996,N_2034,N_2232);
or U2997 (N_2997,N_2018,N_2210);
nand U2998 (N_2998,N_2104,N_2247);
nand U2999 (N_2999,N_2131,N_2000);
nor U3000 (N_3000,N_2543,N_2742);
nand U3001 (N_3001,N_2991,N_2998);
nor U3002 (N_3002,N_2519,N_2695);
xor U3003 (N_3003,N_2608,N_2567);
xor U3004 (N_3004,N_2732,N_2734);
nand U3005 (N_3005,N_2805,N_2525);
nor U3006 (N_3006,N_2673,N_2807);
xor U3007 (N_3007,N_2554,N_2802);
nor U3008 (N_3008,N_2876,N_2728);
xor U3009 (N_3009,N_2796,N_2665);
xnor U3010 (N_3010,N_2677,N_2671);
xnor U3011 (N_3011,N_2992,N_2588);
and U3012 (N_3012,N_2682,N_2566);
and U3013 (N_3013,N_2598,N_2620);
and U3014 (N_3014,N_2771,N_2971);
nor U3015 (N_3015,N_2655,N_2885);
nand U3016 (N_3016,N_2947,N_2662);
nor U3017 (N_3017,N_2630,N_2999);
and U3018 (N_3018,N_2663,N_2723);
and U3019 (N_3019,N_2714,N_2846);
xor U3020 (N_3020,N_2793,N_2816);
and U3021 (N_3021,N_2821,N_2739);
nand U3022 (N_3022,N_2894,N_2975);
nor U3023 (N_3023,N_2617,N_2657);
nand U3024 (N_3024,N_2965,N_2518);
nand U3025 (N_3025,N_2571,N_2904);
nor U3026 (N_3026,N_2704,N_2718);
and U3027 (N_3027,N_2862,N_2854);
nor U3028 (N_3028,N_2563,N_2969);
xnor U3029 (N_3029,N_2605,N_2836);
or U3030 (N_3030,N_2936,N_2843);
and U3031 (N_3031,N_2908,N_2613);
nor U3032 (N_3032,N_2906,N_2831);
or U3033 (N_3033,N_2957,N_2985);
and U3034 (N_3034,N_2648,N_2698);
nor U3035 (N_3035,N_2596,N_2614);
and U3036 (N_3036,N_2790,N_2694);
and U3037 (N_3037,N_2607,N_2735);
nand U3038 (N_3038,N_2818,N_2763);
and U3039 (N_3039,N_2747,N_2559);
and U3040 (N_3040,N_2560,N_2562);
or U3041 (N_3041,N_2510,N_2949);
nand U3042 (N_3042,N_2645,N_2515);
nor U3043 (N_3043,N_2882,N_2811);
or U3044 (N_3044,N_2661,N_2606);
or U3045 (N_3045,N_2956,N_2886);
or U3046 (N_3046,N_2578,N_2691);
and U3047 (N_3047,N_2819,N_2856);
nor U3048 (N_3048,N_2675,N_2979);
or U3049 (N_3049,N_2600,N_2887);
and U3050 (N_3050,N_2914,N_2909);
nor U3051 (N_3051,N_2919,N_2597);
nand U3052 (N_3052,N_2869,N_2859);
xnor U3053 (N_3053,N_2641,N_2916);
nor U3054 (N_3054,N_2801,N_2551);
and U3055 (N_3055,N_2676,N_2511);
nor U3056 (N_3056,N_2656,N_2706);
nor U3057 (N_3057,N_2794,N_2789);
nor U3058 (N_3058,N_2660,N_2729);
nor U3059 (N_3059,N_2824,N_2644);
or U3060 (N_3060,N_2674,N_2669);
and U3061 (N_3061,N_2603,N_2604);
and U3062 (N_3062,N_2950,N_2736);
xor U3063 (N_3063,N_2530,N_2888);
xor U3064 (N_3064,N_2526,N_2637);
nor U3065 (N_3065,N_2837,N_2590);
and U3066 (N_3066,N_2754,N_2690);
and U3067 (N_3067,N_2780,N_2829);
xnor U3068 (N_3068,N_2533,N_2785);
and U3069 (N_3069,N_2595,N_2795);
and U3070 (N_3070,N_2582,N_2528);
nor U3071 (N_3071,N_2863,N_2642);
nand U3072 (N_3072,N_2594,N_2726);
and U3073 (N_3073,N_2941,N_2777);
nand U3074 (N_3074,N_2502,N_2800);
and U3075 (N_3075,N_2685,N_2911);
and U3076 (N_3076,N_2589,N_2577);
nor U3077 (N_3077,N_2834,N_2918);
nor U3078 (N_3078,N_2759,N_2939);
xnor U3079 (N_3079,N_2974,N_2967);
xor U3080 (N_3080,N_2501,N_2897);
xor U3081 (N_3081,N_2953,N_2550);
nor U3082 (N_3082,N_2568,N_2858);
nor U3083 (N_3083,N_2988,N_2973);
nand U3084 (N_3084,N_2782,N_2527);
or U3085 (N_3085,N_2961,N_2653);
nor U3086 (N_3086,N_2922,N_2875);
or U3087 (N_3087,N_2764,N_2631);
and U3088 (N_3088,N_2583,N_2715);
nor U3089 (N_3089,N_2776,N_2505);
nand U3090 (N_3090,N_2743,N_2730);
and U3091 (N_3091,N_2640,N_2522);
nor U3092 (N_3092,N_2970,N_2748);
xnor U3093 (N_3093,N_2866,N_2556);
or U3094 (N_3094,N_2822,N_2737);
and U3095 (N_3095,N_2927,N_2907);
nor U3096 (N_3096,N_2788,N_2878);
xnor U3097 (N_3097,N_2855,N_2937);
and U3098 (N_3098,N_2902,N_2930);
nor U3099 (N_3099,N_2622,N_2591);
xnor U3100 (N_3100,N_2632,N_2980);
or U3101 (N_3101,N_2751,N_2972);
xnor U3102 (N_3102,N_2891,N_2963);
nand U3103 (N_3103,N_2636,N_2835);
xor U3104 (N_3104,N_2996,N_2851);
nor U3105 (N_3105,N_2757,N_2848);
nand U3106 (N_3106,N_2761,N_2981);
nand U3107 (N_3107,N_2845,N_2978);
nor U3108 (N_3108,N_2865,N_2534);
or U3109 (N_3109,N_2841,N_2731);
or U3110 (N_3110,N_2699,N_2868);
nand U3111 (N_3111,N_2544,N_2575);
xnor U3112 (N_3112,N_2516,N_2758);
or U3113 (N_3113,N_2820,N_2667);
nand U3114 (N_3114,N_2532,N_2633);
nor U3115 (N_3115,N_2768,N_2808);
or U3116 (N_3116,N_2553,N_2716);
nand U3117 (N_3117,N_2925,N_2599);
nand U3118 (N_3118,N_2787,N_2923);
or U3119 (N_3119,N_2746,N_2549);
and U3120 (N_3120,N_2627,N_2592);
and U3121 (N_3121,N_2546,N_2744);
and U3122 (N_3122,N_2700,N_2727);
nor U3123 (N_3123,N_2773,N_2889);
and U3124 (N_3124,N_2586,N_2781);
nor U3125 (N_3125,N_2733,N_2572);
or U3126 (N_3126,N_2569,N_2537);
nor U3127 (N_3127,N_2982,N_2760);
nand U3128 (N_3128,N_2539,N_2680);
xnor U3129 (N_3129,N_2721,N_2839);
nor U3130 (N_3130,N_2647,N_2809);
and U3131 (N_3131,N_2994,N_2799);
nor U3132 (N_3132,N_2585,N_2755);
or U3133 (N_3133,N_2709,N_2587);
and U3134 (N_3134,N_2725,N_2752);
xnor U3135 (N_3135,N_2946,N_2703);
and U3136 (N_3136,N_2626,N_2581);
or U3137 (N_3137,N_2536,N_2954);
nand U3138 (N_3138,N_2649,N_2625);
and U3139 (N_3139,N_2535,N_2769);
and U3140 (N_3140,N_2508,N_2666);
or U3141 (N_3141,N_2783,N_2984);
nor U3142 (N_3142,N_2995,N_2864);
nand U3143 (N_3143,N_2684,N_2903);
nor U3144 (N_3144,N_2616,N_2683);
nor U3145 (N_3145,N_2654,N_2881);
and U3146 (N_3146,N_2986,N_2940);
and U3147 (N_3147,N_2584,N_2926);
xor U3148 (N_3148,N_2514,N_2942);
or U3149 (N_3149,N_2542,N_2920);
xnor U3150 (N_3150,N_2696,N_2652);
nor U3151 (N_3151,N_2929,N_2883);
nand U3152 (N_3152,N_2558,N_2833);
nor U3153 (N_3153,N_2870,N_2933);
xor U3154 (N_3154,N_2803,N_2798);
and U3155 (N_3155,N_2860,N_2893);
or U3156 (N_3156,N_2749,N_2651);
and U3157 (N_3157,N_2917,N_2555);
or U3158 (N_3158,N_2951,N_2852);
xnor U3159 (N_3159,N_2989,N_2952);
nand U3160 (N_3160,N_2576,N_2720);
nand U3161 (N_3161,N_2838,N_2968);
nor U3162 (N_3162,N_2997,N_2692);
xnor U3163 (N_3163,N_2830,N_2842);
xnor U3164 (N_3164,N_2915,N_2712);
xor U3165 (N_3165,N_2570,N_2976);
nor U3166 (N_3166,N_2959,N_2810);
and U3167 (N_3167,N_2948,N_2847);
xor U3168 (N_3168,N_2681,N_2503);
nand U3169 (N_3169,N_2541,N_2879);
or U3170 (N_3170,N_2900,N_2705);
or U3171 (N_3171,N_2964,N_2877);
or U3172 (N_3172,N_2987,N_2552);
and U3173 (N_3173,N_2701,N_2618);
xnor U3174 (N_3174,N_2643,N_2924);
xor U3175 (N_3175,N_2849,N_2774);
nand U3176 (N_3176,N_2874,N_2500);
nand U3177 (N_3177,N_2990,N_2766);
nor U3178 (N_3178,N_2504,N_2786);
or U3179 (N_3179,N_2668,N_2901);
nand U3180 (N_3180,N_2797,N_2791);
nand U3181 (N_3181,N_2612,N_2628);
or U3182 (N_3182,N_2813,N_2619);
nand U3183 (N_3183,N_2659,N_2910);
nor U3184 (N_3184,N_2650,N_2825);
and U3185 (N_3185,N_2966,N_2639);
or U3186 (N_3186,N_2804,N_2523);
nor U3187 (N_3187,N_2890,N_2512);
nor U3188 (N_3188,N_2688,N_2601);
nand U3189 (N_3189,N_2962,N_2686);
or U3190 (N_3190,N_2713,N_2812);
nand U3191 (N_3191,N_2767,N_2853);
nand U3192 (N_3192,N_2531,N_2934);
nand U3193 (N_3193,N_2778,N_2564);
and U3194 (N_3194,N_2689,N_2658);
nand U3195 (N_3195,N_2944,N_2529);
and U3196 (N_3196,N_2679,N_2943);
nor U3197 (N_3197,N_2557,N_2753);
or U3198 (N_3198,N_2707,N_2850);
and U3199 (N_3199,N_2827,N_2521);
nand U3200 (N_3200,N_2895,N_2823);
nor U3201 (N_3201,N_2765,N_2872);
or U3202 (N_3202,N_2517,N_2921);
nor U3203 (N_3203,N_2702,N_2506);
nand U3204 (N_3204,N_2779,N_2932);
xnor U3205 (N_3205,N_2857,N_2670);
xnor U3206 (N_3206,N_2960,N_2770);
or U3207 (N_3207,N_2621,N_2724);
xor U3208 (N_3208,N_2815,N_2896);
or U3209 (N_3209,N_2693,N_2548);
xor U3210 (N_3210,N_2762,N_2638);
nand U3211 (N_3211,N_2624,N_2928);
nand U3212 (N_3212,N_2861,N_2738);
nor U3213 (N_3213,N_2871,N_2898);
xor U3214 (N_3214,N_2672,N_2905);
nand U3215 (N_3215,N_2873,N_2678);
nand U3216 (N_3216,N_2772,N_2775);
nor U3217 (N_3217,N_2756,N_2817);
xor U3218 (N_3218,N_2561,N_2806);
xor U3219 (N_3219,N_2513,N_2832);
nor U3220 (N_3220,N_2828,N_2880);
nor U3221 (N_3221,N_2892,N_2722);
nand U3222 (N_3222,N_2580,N_2687);
and U3223 (N_3223,N_2750,N_2711);
or U3224 (N_3224,N_2545,N_2912);
nor U3225 (N_3225,N_2565,N_2538);
nand U3226 (N_3226,N_2977,N_2708);
nand U3227 (N_3227,N_2945,N_2814);
nor U3228 (N_3228,N_2524,N_2547);
and U3229 (N_3229,N_2938,N_2602);
xor U3230 (N_3230,N_2792,N_2983);
nor U3231 (N_3231,N_2579,N_2664);
or U3232 (N_3232,N_2958,N_2719);
or U3233 (N_3233,N_2615,N_2574);
nand U3234 (N_3234,N_2573,N_2741);
nand U3235 (N_3235,N_2509,N_2913);
or U3236 (N_3236,N_2507,N_2935);
or U3237 (N_3237,N_2899,N_2635);
nand U3238 (N_3238,N_2717,N_2710);
xnor U3239 (N_3239,N_2609,N_2520);
nand U3240 (N_3240,N_2993,N_2629);
nand U3241 (N_3241,N_2611,N_2634);
or U3242 (N_3242,N_2540,N_2745);
nor U3243 (N_3243,N_2884,N_2867);
nand U3244 (N_3244,N_2931,N_2697);
or U3245 (N_3245,N_2844,N_2955);
nand U3246 (N_3246,N_2623,N_2646);
xnor U3247 (N_3247,N_2826,N_2593);
nand U3248 (N_3248,N_2784,N_2740);
nor U3249 (N_3249,N_2840,N_2610);
nor U3250 (N_3250,N_2507,N_2805);
nand U3251 (N_3251,N_2872,N_2539);
nor U3252 (N_3252,N_2633,N_2809);
xor U3253 (N_3253,N_2911,N_2934);
and U3254 (N_3254,N_2808,N_2835);
xnor U3255 (N_3255,N_2745,N_2657);
xor U3256 (N_3256,N_2646,N_2567);
or U3257 (N_3257,N_2847,N_2914);
and U3258 (N_3258,N_2685,N_2895);
nor U3259 (N_3259,N_2739,N_2529);
xnor U3260 (N_3260,N_2733,N_2680);
nor U3261 (N_3261,N_2508,N_2921);
xnor U3262 (N_3262,N_2719,N_2512);
and U3263 (N_3263,N_2705,N_2798);
or U3264 (N_3264,N_2555,N_2718);
and U3265 (N_3265,N_2671,N_2590);
nand U3266 (N_3266,N_2851,N_2733);
or U3267 (N_3267,N_2631,N_2854);
or U3268 (N_3268,N_2976,N_2711);
xor U3269 (N_3269,N_2553,N_2676);
or U3270 (N_3270,N_2663,N_2970);
nor U3271 (N_3271,N_2500,N_2914);
or U3272 (N_3272,N_2838,N_2911);
nor U3273 (N_3273,N_2607,N_2693);
nand U3274 (N_3274,N_2612,N_2992);
nor U3275 (N_3275,N_2777,N_2568);
and U3276 (N_3276,N_2864,N_2918);
or U3277 (N_3277,N_2608,N_2842);
nor U3278 (N_3278,N_2807,N_2830);
xor U3279 (N_3279,N_2845,N_2772);
nor U3280 (N_3280,N_2600,N_2851);
nor U3281 (N_3281,N_2913,N_2756);
xor U3282 (N_3282,N_2535,N_2622);
nand U3283 (N_3283,N_2791,N_2751);
xnor U3284 (N_3284,N_2530,N_2916);
and U3285 (N_3285,N_2555,N_2713);
xor U3286 (N_3286,N_2622,N_2621);
xor U3287 (N_3287,N_2525,N_2785);
nand U3288 (N_3288,N_2700,N_2606);
xor U3289 (N_3289,N_2593,N_2681);
and U3290 (N_3290,N_2621,N_2642);
nand U3291 (N_3291,N_2576,N_2561);
or U3292 (N_3292,N_2539,N_2765);
nand U3293 (N_3293,N_2513,N_2755);
nor U3294 (N_3294,N_2654,N_2996);
nand U3295 (N_3295,N_2655,N_2841);
and U3296 (N_3296,N_2740,N_2974);
and U3297 (N_3297,N_2993,N_2553);
nor U3298 (N_3298,N_2794,N_2741);
xnor U3299 (N_3299,N_2532,N_2845);
nor U3300 (N_3300,N_2749,N_2948);
nor U3301 (N_3301,N_2910,N_2711);
nand U3302 (N_3302,N_2900,N_2625);
xor U3303 (N_3303,N_2910,N_2845);
and U3304 (N_3304,N_2529,N_2869);
nand U3305 (N_3305,N_2937,N_2858);
nand U3306 (N_3306,N_2758,N_2680);
and U3307 (N_3307,N_2869,N_2820);
and U3308 (N_3308,N_2542,N_2603);
nand U3309 (N_3309,N_2556,N_2773);
nand U3310 (N_3310,N_2831,N_2919);
and U3311 (N_3311,N_2600,N_2949);
xnor U3312 (N_3312,N_2705,N_2971);
xnor U3313 (N_3313,N_2789,N_2864);
nand U3314 (N_3314,N_2505,N_2552);
xnor U3315 (N_3315,N_2863,N_2942);
or U3316 (N_3316,N_2516,N_2566);
nand U3317 (N_3317,N_2782,N_2876);
nand U3318 (N_3318,N_2675,N_2621);
nand U3319 (N_3319,N_2518,N_2724);
nor U3320 (N_3320,N_2806,N_2909);
nand U3321 (N_3321,N_2514,N_2711);
nor U3322 (N_3322,N_2789,N_2707);
or U3323 (N_3323,N_2995,N_2538);
and U3324 (N_3324,N_2760,N_2728);
nor U3325 (N_3325,N_2543,N_2778);
xnor U3326 (N_3326,N_2796,N_2578);
xnor U3327 (N_3327,N_2762,N_2790);
or U3328 (N_3328,N_2976,N_2766);
xor U3329 (N_3329,N_2698,N_2971);
xnor U3330 (N_3330,N_2916,N_2539);
or U3331 (N_3331,N_2735,N_2604);
xor U3332 (N_3332,N_2793,N_2517);
nor U3333 (N_3333,N_2501,N_2758);
xor U3334 (N_3334,N_2769,N_2857);
or U3335 (N_3335,N_2521,N_2668);
and U3336 (N_3336,N_2559,N_2818);
and U3337 (N_3337,N_2849,N_2583);
and U3338 (N_3338,N_2735,N_2991);
and U3339 (N_3339,N_2586,N_2828);
nor U3340 (N_3340,N_2601,N_2944);
nor U3341 (N_3341,N_2809,N_2965);
nand U3342 (N_3342,N_2761,N_2658);
xnor U3343 (N_3343,N_2620,N_2786);
xor U3344 (N_3344,N_2712,N_2569);
nor U3345 (N_3345,N_2672,N_2954);
or U3346 (N_3346,N_2919,N_2697);
or U3347 (N_3347,N_2675,N_2772);
xor U3348 (N_3348,N_2556,N_2535);
nor U3349 (N_3349,N_2961,N_2934);
or U3350 (N_3350,N_2943,N_2647);
nand U3351 (N_3351,N_2679,N_2531);
and U3352 (N_3352,N_2726,N_2731);
xor U3353 (N_3353,N_2705,N_2678);
and U3354 (N_3354,N_2785,N_2985);
or U3355 (N_3355,N_2881,N_2660);
xor U3356 (N_3356,N_2671,N_2579);
or U3357 (N_3357,N_2912,N_2957);
or U3358 (N_3358,N_2534,N_2655);
and U3359 (N_3359,N_2700,N_2529);
and U3360 (N_3360,N_2723,N_2645);
or U3361 (N_3361,N_2519,N_2726);
nor U3362 (N_3362,N_2753,N_2994);
nand U3363 (N_3363,N_2691,N_2851);
or U3364 (N_3364,N_2956,N_2963);
or U3365 (N_3365,N_2699,N_2879);
and U3366 (N_3366,N_2741,N_2607);
nand U3367 (N_3367,N_2937,N_2712);
xnor U3368 (N_3368,N_2759,N_2964);
nor U3369 (N_3369,N_2567,N_2589);
xor U3370 (N_3370,N_2600,N_2607);
nor U3371 (N_3371,N_2870,N_2613);
xnor U3372 (N_3372,N_2835,N_2990);
xnor U3373 (N_3373,N_2932,N_2830);
or U3374 (N_3374,N_2777,N_2976);
and U3375 (N_3375,N_2726,N_2670);
xor U3376 (N_3376,N_2856,N_2503);
xor U3377 (N_3377,N_2961,N_2573);
or U3378 (N_3378,N_2708,N_2791);
or U3379 (N_3379,N_2971,N_2642);
nand U3380 (N_3380,N_2825,N_2642);
and U3381 (N_3381,N_2578,N_2921);
nor U3382 (N_3382,N_2568,N_2727);
xnor U3383 (N_3383,N_2998,N_2640);
xnor U3384 (N_3384,N_2607,N_2804);
nand U3385 (N_3385,N_2750,N_2617);
nand U3386 (N_3386,N_2617,N_2725);
or U3387 (N_3387,N_2678,N_2871);
xnor U3388 (N_3388,N_2592,N_2731);
nand U3389 (N_3389,N_2923,N_2544);
xor U3390 (N_3390,N_2679,N_2727);
nor U3391 (N_3391,N_2822,N_2818);
xor U3392 (N_3392,N_2673,N_2789);
or U3393 (N_3393,N_2763,N_2744);
nand U3394 (N_3394,N_2878,N_2765);
nor U3395 (N_3395,N_2886,N_2585);
xor U3396 (N_3396,N_2747,N_2655);
nand U3397 (N_3397,N_2637,N_2940);
nor U3398 (N_3398,N_2546,N_2730);
nor U3399 (N_3399,N_2775,N_2725);
nand U3400 (N_3400,N_2914,N_2603);
nor U3401 (N_3401,N_2842,N_2643);
or U3402 (N_3402,N_2709,N_2750);
and U3403 (N_3403,N_2562,N_2767);
nand U3404 (N_3404,N_2742,N_2897);
nor U3405 (N_3405,N_2508,N_2696);
and U3406 (N_3406,N_2594,N_2745);
and U3407 (N_3407,N_2959,N_2923);
nor U3408 (N_3408,N_2708,N_2529);
or U3409 (N_3409,N_2807,N_2670);
nand U3410 (N_3410,N_2876,N_2985);
nor U3411 (N_3411,N_2761,N_2945);
and U3412 (N_3412,N_2880,N_2939);
nor U3413 (N_3413,N_2891,N_2625);
xnor U3414 (N_3414,N_2901,N_2539);
and U3415 (N_3415,N_2955,N_2936);
xor U3416 (N_3416,N_2553,N_2987);
nor U3417 (N_3417,N_2741,N_2848);
or U3418 (N_3418,N_2534,N_2727);
and U3419 (N_3419,N_2945,N_2608);
or U3420 (N_3420,N_2606,N_2911);
or U3421 (N_3421,N_2714,N_2645);
and U3422 (N_3422,N_2853,N_2894);
xor U3423 (N_3423,N_2555,N_2863);
or U3424 (N_3424,N_2783,N_2995);
nand U3425 (N_3425,N_2688,N_2817);
and U3426 (N_3426,N_2590,N_2712);
nor U3427 (N_3427,N_2961,N_2511);
or U3428 (N_3428,N_2944,N_2564);
or U3429 (N_3429,N_2953,N_2811);
xnor U3430 (N_3430,N_2963,N_2659);
nor U3431 (N_3431,N_2897,N_2841);
nand U3432 (N_3432,N_2857,N_2633);
or U3433 (N_3433,N_2879,N_2616);
nand U3434 (N_3434,N_2897,N_2811);
xnor U3435 (N_3435,N_2621,N_2665);
or U3436 (N_3436,N_2807,N_2544);
nor U3437 (N_3437,N_2938,N_2526);
xnor U3438 (N_3438,N_2769,N_2797);
xnor U3439 (N_3439,N_2706,N_2612);
or U3440 (N_3440,N_2715,N_2536);
nor U3441 (N_3441,N_2589,N_2941);
nor U3442 (N_3442,N_2988,N_2940);
nand U3443 (N_3443,N_2978,N_2997);
and U3444 (N_3444,N_2522,N_2878);
nor U3445 (N_3445,N_2931,N_2642);
nor U3446 (N_3446,N_2918,N_2691);
or U3447 (N_3447,N_2997,N_2968);
nand U3448 (N_3448,N_2644,N_2702);
or U3449 (N_3449,N_2817,N_2654);
nor U3450 (N_3450,N_2559,N_2725);
and U3451 (N_3451,N_2616,N_2654);
or U3452 (N_3452,N_2951,N_2705);
and U3453 (N_3453,N_2890,N_2548);
nand U3454 (N_3454,N_2959,N_2768);
nor U3455 (N_3455,N_2988,N_2953);
or U3456 (N_3456,N_2929,N_2693);
and U3457 (N_3457,N_2974,N_2970);
xor U3458 (N_3458,N_2856,N_2686);
and U3459 (N_3459,N_2892,N_2801);
xnor U3460 (N_3460,N_2992,N_2948);
or U3461 (N_3461,N_2999,N_2939);
or U3462 (N_3462,N_2845,N_2959);
nor U3463 (N_3463,N_2556,N_2877);
nor U3464 (N_3464,N_2939,N_2972);
and U3465 (N_3465,N_2580,N_2807);
nand U3466 (N_3466,N_2773,N_2838);
and U3467 (N_3467,N_2624,N_2878);
xnor U3468 (N_3468,N_2893,N_2756);
nand U3469 (N_3469,N_2778,N_2557);
or U3470 (N_3470,N_2836,N_2973);
nor U3471 (N_3471,N_2959,N_2937);
and U3472 (N_3472,N_2680,N_2798);
nor U3473 (N_3473,N_2837,N_2975);
nand U3474 (N_3474,N_2516,N_2817);
xor U3475 (N_3475,N_2688,N_2874);
xor U3476 (N_3476,N_2657,N_2986);
and U3477 (N_3477,N_2838,N_2777);
xnor U3478 (N_3478,N_2566,N_2641);
nand U3479 (N_3479,N_2964,N_2635);
nor U3480 (N_3480,N_2524,N_2857);
nand U3481 (N_3481,N_2740,N_2919);
nand U3482 (N_3482,N_2626,N_2653);
nand U3483 (N_3483,N_2830,N_2707);
nor U3484 (N_3484,N_2769,N_2900);
xor U3485 (N_3485,N_2733,N_2918);
xor U3486 (N_3486,N_2830,N_2998);
nor U3487 (N_3487,N_2671,N_2687);
nor U3488 (N_3488,N_2603,N_2870);
nor U3489 (N_3489,N_2504,N_2870);
or U3490 (N_3490,N_2993,N_2522);
nand U3491 (N_3491,N_2682,N_2768);
nand U3492 (N_3492,N_2865,N_2894);
and U3493 (N_3493,N_2540,N_2589);
nor U3494 (N_3494,N_2864,N_2641);
and U3495 (N_3495,N_2729,N_2996);
and U3496 (N_3496,N_2511,N_2993);
nand U3497 (N_3497,N_2897,N_2651);
or U3498 (N_3498,N_2614,N_2607);
or U3499 (N_3499,N_2704,N_2790);
and U3500 (N_3500,N_3298,N_3326);
xor U3501 (N_3501,N_3257,N_3267);
nand U3502 (N_3502,N_3055,N_3442);
or U3503 (N_3503,N_3303,N_3026);
nor U3504 (N_3504,N_3333,N_3205);
nor U3505 (N_3505,N_3066,N_3388);
and U3506 (N_3506,N_3287,N_3317);
or U3507 (N_3507,N_3063,N_3186);
nand U3508 (N_3508,N_3289,N_3010);
xnor U3509 (N_3509,N_3188,N_3421);
and U3510 (N_3510,N_3212,N_3369);
nand U3511 (N_3511,N_3008,N_3274);
and U3512 (N_3512,N_3254,N_3223);
nor U3513 (N_3513,N_3194,N_3418);
xor U3514 (N_3514,N_3004,N_3094);
nand U3515 (N_3515,N_3099,N_3276);
xor U3516 (N_3516,N_3376,N_3422);
or U3517 (N_3517,N_3312,N_3323);
nand U3518 (N_3518,N_3451,N_3320);
and U3519 (N_3519,N_3414,N_3357);
and U3520 (N_3520,N_3042,N_3358);
nor U3521 (N_3521,N_3490,N_3306);
nand U3522 (N_3522,N_3169,N_3109);
xor U3523 (N_3523,N_3086,N_3144);
xor U3524 (N_3524,N_3469,N_3404);
nor U3525 (N_3525,N_3208,N_3371);
xor U3526 (N_3526,N_3077,N_3210);
nor U3527 (N_3527,N_3219,N_3350);
nor U3528 (N_3528,N_3222,N_3083);
xor U3529 (N_3529,N_3344,N_3220);
xor U3530 (N_3530,N_3088,N_3059);
nor U3531 (N_3531,N_3087,N_3439);
nand U3532 (N_3532,N_3262,N_3382);
and U3533 (N_3533,N_3031,N_3394);
nand U3534 (N_3534,N_3495,N_3067);
nor U3535 (N_3535,N_3492,N_3161);
and U3536 (N_3536,N_3060,N_3441);
xor U3537 (N_3537,N_3329,N_3201);
xnor U3538 (N_3538,N_3191,N_3244);
xnor U3539 (N_3539,N_3124,N_3266);
nor U3540 (N_3540,N_3258,N_3061);
nand U3541 (N_3541,N_3227,N_3221);
xor U3542 (N_3542,N_3453,N_3057);
and U3543 (N_3543,N_3102,N_3330);
xor U3544 (N_3544,N_3431,N_3494);
nor U3545 (N_3545,N_3468,N_3082);
nor U3546 (N_3546,N_3052,N_3435);
nand U3547 (N_3547,N_3167,N_3229);
and U3548 (N_3548,N_3447,N_3268);
or U3549 (N_3549,N_3147,N_3401);
or U3550 (N_3550,N_3377,N_3296);
xor U3551 (N_3551,N_3148,N_3051);
or U3552 (N_3552,N_3024,N_3381);
or U3553 (N_3553,N_3036,N_3118);
nor U3554 (N_3554,N_3001,N_3458);
nor U3555 (N_3555,N_3277,N_3236);
and U3556 (N_3556,N_3297,N_3246);
or U3557 (N_3557,N_3065,N_3231);
xor U3558 (N_3558,N_3311,N_3396);
and U3559 (N_3559,N_3180,N_3362);
nor U3560 (N_3560,N_3319,N_3101);
xor U3561 (N_3561,N_3135,N_3470);
or U3562 (N_3562,N_3259,N_3255);
or U3563 (N_3563,N_3175,N_3264);
nand U3564 (N_3564,N_3378,N_3355);
nand U3565 (N_3565,N_3058,N_3069);
nor U3566 (N_3566,N_3288,N_3410);
xnor U3567 (N_3567,N_3429,N_3260);
nand U3568 (N_3568,N_3129,N_3073);
nor U3569 (N_3569,N_3419,N_3136);
or U3570 (N_3570,N_3375,N_3482);
or U3571 (N_3571,N_3301,N_3183);
xor U3572 (N_3572,N_3016,N_3325);
or U3573 (N_3573,N_3361,N_3199);
xnor U3574 (N_3574,N_3143,N_3206);
and U3575 (N_3575,N_3075,N_3146);
nor U3576 (N_3576,N_3462,N_3145);
nor U3577 (N_3577,N_3335,N_3444);
nand U3578 (N_3578,N_3017,N_3006);
or U3579 (N_3579,N_3153,N_3339);
and U3580 (N_3580,N_3243,N_3480);
and U3581 (N_3581,N_3193,N_3202);
and U3582 (N_3582,N_3224,N_3228);
nand U3583 (N_3583,N_3280,N_3190);
and U3584 (N_3584,N_3198,N_3211);
nand U3585 (N_3585,N_3126,N_3238);
xnor U3586 (N_3586,N_3397,N_3033);
xor U3587 (N_3587,N_3484,N_3040);
and U3588 (N_3588,N_3415,N_3345);
xor U3589 (N_3589,N_3034,N_3430);
nand U3590 (N_3590,N_3411,N_3125);
xnor U3591 (N_3591,N_3425,N_3286);
nand U3592 (N_3592,N_3253,N_3428);
or U3593 (N_3593,N_3437,N_3474);
nand U3594 (N_3594,N_3030,N_3283);
or U3595 (N_3595,N_3467,N_3292);
or U3596 (N_3596,N_3291,N_3389);
and U3597 (N_3597,N_3426,N_3113);
or U3598 (N_3598,N_3157,N_3155);
xor U3599 (N_3599,N_3047,N_3078);
nor U3600 (N_3600,N_3491,N_3440);
nand U3601 (N_3601,N_3110,N_3218);
and U3602 (N_3602,N_3304,N_3424);
or U3603 (N_3603,N_3035,N_3460);
nand U3604 (N_3604,N_3332,N_3089);
and U3605 (N_3605,N_3300,N_3107);
or U3606 (N_3606,N_3115,N_3295);
xnor U3607 (N_3607,N_3393,N_3189);
and U3608 (N_3608,N_3408,N_3173);
or U3609 (N_3609,N_3261,N_3200);
xor U3610 (N_3610,N_3321,N_3331);
or U3611 (N_3611,N_3354,N_3241);
nor U3612 (N_3612,N_3207,N_3130);
or U3613 (N_3613,N_3009,N_3204);
or U3614 (N_3614,N_3380,N_3475);
nor U3615 (N_3615,N_3497,N_3203);
and U3616 (N_3616,N_3316,N_3449);
nand U3617 (N_3617,N_3402,N_3456);
nor U3618 (N_3618,N_3463,N_3248);
nand U3619 (N_3619,N_3093,N_3464);
and U3620 (N_3620,N_3049,N_3434);
nand U3621 (N_3621,N_3454,N_3233);
xnor U3622 (N_3622,N_3364,N_3108);
nand U3623 (N_3623,N_3092,N_3348);
and U3624 (N_3624,N_3164,N_3363);
nor U3625 (N_3625,N_3485,N_3247);
xnor U3626 (N_3626,N_3085,N_3400);
xnor U3627 (N_3627,N_3347,N_3406);
and U3628 (N_3628,N_3112,N_3056);
xnor U3629 (N_3629,N_3405,N_3154);
nor U3630 (N_3630,N_3322,N_3021);
nor U3631 (N_3631,N_3471,N_3028);
or U3632 (N_3632,N_3174,N_3139);
and U3633 (N_3633,N_3372,N_3476);
xnor U3634 (N_3634,N_3346,N_3318);
nand U3635 (N_3635,N_3466,N_3324);
or U3636 (N_3636,N_3072,N_3003);
or U3637 (N_3637,N_3279,N_3217);
nor U3638 (N_3638,N_3080,N_3216);
nor U3639 (N_3639,N_3379,N_3436);
xnor U3640 (N_3640,N_3237,N_3366);
xor U3641 (N_3641,N_3064,N_3472);
nor U3642 (N_3642,N_3493,N_3281);
xor U3643 (N_3643,N_3041,N_3070);
nand U3644 (N_3644,N_3473,N_3448);
nor U3645 (N_3645,N_3023,N_3095);
nor U3646 (N_3646,N_3019,N_3062);
or U3647 (N_3647,N_3018,N_3168);
and U3648 (N_3648,N_3116,N_3373);
nand U3649 (N_3649,N_3097,N_3170);
xor U3650 (N_3650,N_3461,N_3310);
nand U3651 (N_3651,N_3487,N_3142);
nor U3652 (N_3652,N_3048,N_3427);
nor U3653 (N_3653,N_3103,N_3235);
or U3654 (N_3654,N_3334,N_3360);
xnor U3655 (N_3655,N_3446,N_3012);
and U3656 (N_3656,N_3341,N_3141);
xnor U3657 (N_3657,N_3081,N_3140);
or U3658 (N_3658,N_3119,N_3315);
nor U3659 (N_3659,N_3071,N_3328);
and U3660 (N_3660,N_3340,N_3152);
nand U3661 (N_3661,N_3284,N_3163);
nand U3662 (N_3662,N_3007,N_3225);
nand U3663 (N_3663,N_3486,N_3015);
xor U3664 (N_3664,N_3137,N_3150);
or U3665 (N_3665,N_3242,N_3054);
nor U3666 (N_3666,N_3213,N_3162);
or U3667 (N_3667,N_3053,N_3002);
xnor U3668 (N_3668,N_3412,N_3403);
and U3669 (N_3669,N_3477,N_3395);
xor U3670 (N_3670,N_3383,N_3230);
and U3671 (N_3671,N_3293,N_3044);
nor U3672 (N_3672,N_3478,N_3443);
xnor U3673 (N_3673,N_3353,N_3285);
and U3674 (N_3674,N_3417,N_3166);
xnor U3675 (N_3675,N_3215,N_3457);
nand U3676 (N_3676,N_3171,N_3005);
nand U3677 (N_3677,N_3336,N_3309);
nor U3678 (N_3678,N_3359,N_3131);
or U3679 (N_3679,N_3367,N_3249);
xor U3680 (N_3680,N_3197,N_3313);
nand U3681 (N_3681,N_3032,N_3263);
nor U3682 (N_3682,N_3273,N_3134);
or U3683 (N_3683,N_3374,N_3352);
and U3684 (N_3684,N_3098,N_3299);
nor U3685 (N_3685,N_3384,N_3182);
xnor U3686 (N_3686,N_3278,N_3122);
nor U3687 (N_3687,N_3481,N_3327);
or U3688 (N_3688,N_3305,N_3416);
nand U3689 (N_3689,N_3117,N_3176);
nor U3690 (N_3690,N_3120,N_3250);
nand U3691 (N_3691,N_3160,N_3488);
and U3692 (N_3692,N_3132,N_3029);
nor U3693 (N_3693,N_3181,N_3165);
nand U3694 (N_3694,N_3011,N_3014);
and U3695 (N_3695,N_3184,N_3351);
xnor U3696 (N_3696,N_3079,N_3156);
nor U3697 (N_3697,N_3251,N_3365);
and U3698 (N_3698,N_3432,N_3096);
or U3699 (N_3699,N_3209,N_3423);
xor U3700 (N_3700,N_3172,N_3149);
xor U3701 (N_3701,N_3282,N_3046);
nand U3702 (N_3702,N_3226,N_3127);
nor U3703 (N_3703,N_3391,N_3270);
and U3704 (N_3704,N_3106,N_3294);
xnor U3705 (N_3705,N_3158,N_3138);
nor U3706 (N_3706,N_3271,N_3256);
or U3707 (N_3707,N_3038,N_3465);
nor U3708 (N_3708,N_3370,N_3133);
xor U3709 (N_3709,N_3496,N_3045);
and U3710 (N_3710,N_3192,N_3177);
and U3711 (N_3711,N_3104,N_3314);
xnor U3712 (N_3712,N_3068,N_3269);
or U3713 (N_3713,N_3399,N_3076);
and U3714 (N_3714,N_3091,N_3123);
or U3715 (N_3715,N_3022,N_3234);
xnor U3716 (N_3716,N_3498,N_3185);
nor U3717 (N_3717,N_3179,N_3390);
and U3718 (N_3718,N_3187,N_3343);
nor U3719 (N_3719,N_3452,N_3265);
nor U3720 (N_3720,N_3105,N_3385);
and U3721 (N_3721,N_3114,N_3499);
and U3722 (N_3722,N_3037,N_3455);
xor U3723 (N_3723,N_3387,N_3392);
nand U3724 (N_3724,N_3438,N_3338);
and U3725 (N_3725,N_3356,N_3349);
nor U3726 (N_3726,N_3027,N_3420);
nand U3727 (N_3727,N_3013,N_3074);
nand U3728 (N_3728,N_3398,N_3239);
or U3729 (N_3729,N_3084,N_3025);
and U3730 (N_3730,N_3290,N_3240);
nand U3731 (N_3731,N_3111,N_3489);
nand U3732 (N_3732,N_3245,N_3043);
xnor U3733 (N_3733,N_3407,N_3000);
xnor U3734 (N_3734,N_3450,N_3178);
or U3735 (N_3735,N_3386,N_3214);
nor U3736 (N_3736,N_3121,N_3433);
xor U3737 (N_3737,N_3020,N_3337);
or U3738 (N_3738,N_3159,N_3252);
and U3739 (N_3739,N_3368,N_3090);
and U3740 (N_3740,N_3459,N_3302);
xnor U3741 (N_3741,N_3128,N_3050);
xor U3742 (N_3742,N_3413,N_3483);
xnor U3743 (N_3743,N_3479,N_3039);
or U3744 (N_3744,N_3409,N_3232);
or U3745 (N_3745,N_3100,N_3275);
and U3746 (N_3746,N_3308,N_3151);
xor U3747 (N_3747,N_3196,N_3195);
or U3748 (N_3748,N_3342,N_3307);
xor U3749 (N_3749,N_3272,N_3445);
or U3750 (N_3750,N_3457,N_3302);
xnor U3751 (N_3751,N_3424,N_3163);
or U3752 (N_3752,N_3124,N_3411);
and U3753 (N_3753,N_3118,N_3241);
xor U3754 (N_3754,N_3139,N_3420);
and U3755 (N_3755,N_3456,N_3034);
nand U3756 (N_3756,N_3231,N_3313);
nand U3757 (N_3757,N_3202,N_3040);
nand U3758 (N_3758,N_3246,N_3348);
xor U3759 (N_3759,N_3419,N_3394);
or U3760 (N_3760,N_3334,N_3356);
and U3761 (N_3761,N_3191,N_3250);
nor U3762 (N_3762,N_3064,N_3219);
xnor U3763 (N_3763,N_3082,N_3151);
nor U3764 (N_3764,N_3393,N_3206);
or U3765 (N_3765,N_3233,N_3013);
xor U3766 (N_3766,N_3168,N_3195);
nor U3767 (N_3767,N_3060,N_3073);
and U3768 (N_3768,N_3187,N_3165);
nand U3769 (N_3769,N_3235,N_3046);
and U3770 (N_3770,N_3165,N_3337);
and U3771 (N_3771,N_3377,N_3244);
nor U3772 (N_3772,N_3189,N_3241);
nor U3773 (N_3773,N_3007,N_3440);
xnor U3774 (N_3774,N_3448,N_3088);
and U3775 (N_3775,N_3125,N_3276);
nor U3776 (N_3776,N_3237,N_3402);
and U3777 (N_3777,N_3038,N_3347);
nand U3778 (N_3778,N_3189,N_3423);
and U3779 (N_3779,N_3046,N_3110);
xnor U3780 (N_3780,N_3498,N_3016);
xnor U3781 (N_3781,N_3394,N_3034);
nand U3782 (N_3782,N_3252,N_3239);
nand U3783 (N_3783,N_3396,N_3302);
xor U3784 (N_3784,N_3375,N_3266);
xnor U3785 (N_3785,N_3063,N_3201);
xnor U3786 (N_3786,N_3413,N_3293);
nor U3787 (N_3787,N_3234,N_3171);
nand U3788 (N_3788,N_3219,N_3197);
nand U3789 (N_3789,N_3475,N_3218);
nor U3790 (N_3790,N_3199,N_3046);
or U3791 (N_3791,N_3204,N_3089);
nand U3792 (N_3792,N_3280,N_3020);
nor U3793 (N_3793,N_3386,N_3404);
or U3794 (N_3794,N_3387,N_3030);
or U3795 (N_3795,N_3481,N_3491);
nor U3796 (N_3796,N_3030,N_3175);
xor U3797 (N_3797,N_3398,N_3450);
nor U3798 (N_3798,N_3159,N_3460);
xnor U3799 (N_3799,N_3197,N_3015);
nand U3800 (N_3800,N_3289,N_3341);
xnor U3801 (N_3801,N_3345,N_3072);
nor U3802 (N_3802,N_3492,N_3256);
or U3803 (N_3803,N_3073,N_3377);
nor U3804 (N_3804,N_3149,N_3131);
xnor U3805 (N_3805,N_3442,N_3025);
xor U3806 (N_3806,N_3449,N_3266);
xnor U3807 (N_3807,N_3303,N_3233);
nor U3808 (N_3808,N_3197,N_3029);
nor U3809 (N_3809,N_3346,N_3381);
and U3810 (N_3810,N_3192,N_3302);
or U3811 (N_3811,N_3370,N_3157);
and U3812 (N_3812,N_3024,N_3457);
nand U3813 (N_3813,N_3442,N_3389);
nand U3814 (N_3814,N_3274,N_3390);
or U3815 (N_3815,N_3237,N_3053);
nor U3816 (N_3816,N_3166,N_3174);
xnor U3817 (N_3817,N_3012,N_3097);
nor U3818 (N_3818,N_3386,N_3168);
nand U3819 (N_3819,N_3160,N_3135);
nand U3820 (N_3820,N_3225,N_3034);
nor U3821 (N_3821,N_3332,N_3021);
xor U3822 (N_3822,N_3027,N_3346);
or U3823 (N_3823,N_3274,N_3120);
or U3824 (N_3824,N_3219,N_3254);
and U3825 (N_3825,N_3401,N_3413);
or U3826 (N_3826,N_3158,N_3479);
and U3827 (N_3827,N_3206,N_3277);
nor U3828 (N_3828,N_3363,N_3128);
xor U3829 (N_3829,N_3456,N_3184);
and U3830 (N_3830,N_3231,N_3409);
or U3831 (N_3831,N_3447,N_3035);
nor U3832 (N_3832,N_3083,N_3063);
xnor U3833 (N_3833,N_3104,N_3394);
and U3834 (N_3834,N_3261,N_3458);
nor U3835 (N_3835,N_3123,N_3283);
or U3836 (N_3836,N_3474,N_3427);
xor U3837 (N_3837,N_3063,N_3044);
and U3838 (N_3838,N_3338,N_3353);
and U3839 (N_3839,N_3237,N_3441);
nand U3840 (N_3840,N_3084,N_3312);
nor U3841 (N_3841,N_3499,N_3292);
or U3842 (N_3842,N_3356,N_3210);
nand U3843 (N_3843,N_3396,N_3480);
nand U3844 (N_3844,N_3371,N_3479);
and U3845 (N_3845,N_3444,N_3468);
nand U3846 (N_3846,N_3390,N_3067);
or U3847 (N_3847,N_3276,N_3222);
or U3848 (N_3848,N_3129,N_3441);
xor U3849 (N_3849,N_3034,N_3356);
xor U3850 (N_3850,N_3447,N_3285);
and U3851 (N_3851,N_3251,N_3164);
xor U3852 (N_3852,N_3453,N_3028);
and U3853 (N_3853,N_3048,N_3366);
xnor U3854 (N_3854,N_3291,N_3422);
xnor U3855 (N_3855,N_3370,N_3060);
xor U3856 (N_3856,N_3277,N_3273);
or U3857 (N_3857,N_3366,N_3043);
or U3858 (N_3858,N_3459,N_3011);
nor U3859 (N_3859,N_3220,N_3161);
nor U3860 (N_3860,N_3289,N_3108);
nor U3861 (N_3861,N_3400,N_3197);
nor U3862 (N_3862,N_3198,N_3433);
xnor U3863 (N_3863,N_3429,N_3057);
and U3864 (N_3864,N_3193,N_3284);
and U3865 (N_3865,N_3419,N_3421);
xor U3866 (N_3866,N_3144,N_3216);
nand U3867 (N_3867,N_3042,N_3331);
and U3868 (N_3868,N_3289,N_3062);
nor U3869 (N_3869,N_3142,N_3073);
and U3870 (N_3870,N_3220,N_3431);
nor U3871 (N_3871,N_3294,N_3324);
or U3872 (N_3872,N_3173,N_3413);
and U3873 (N_3873,N_3131,N_3159);
nor U3874 (N_3874,N_3297,N_3084);
xnor U3875 (N_3875,N_3022,N_3031);
or U3876 (N_3876,N_3277,N_3477);
nand U3877 (N_3877,N_3210,N_3046);
xor U3878 (N_3878,N_3022,N_3277);
nand U3879 (N_3879,N_3190,N_3237);
nand U3880 (N_3880,N_3119,N_3410);
and U3881 (N_3881,N_3158,N_3156);
nor U3882 (N_3882,N_3091,N_3015);
and U3883 (N_3883,N_3441,N_3291);
nor U3884 (N_3884,N_3166,N_3195);
and U3885 (N_3885,N_3406,N_3299);
nand U3886 (N_3886,N_3390,N_3447);
or U3887 (N_3887,N_3183,N_3129);
or U3888 (N_3888,N_3128,N_3437);
nor U3889 (N_3889,N_3346,N_3268);
nand U3890 (N_3890,N_3345,N_3159);
nor U3891 (N_3891,N_3298,N_3193);
and U3892 (N_3892,N_3015,N_3161);
and U3893 (N_3893,N_3016,N_3278);
or U3894 (N_3894,N_3041,N_3287);
xnor U3895 (N_3895,N_3378,N_3496);
and U3896 (N_3896,N_3372,N_3411);
nand U3897 (N_3897,N_3251,N_3245);
xor U3898 (N_3898,N_3013,N_3322);
nor U3899 (N_3899,N_3064,N_3422);
nor U3900 (N_3900,N_3132,N_3225);
xor U3901 (N_3901,N_3121,N_3056);
nand U3902 (N_3902,N_3427,N_3252);
or U3903 (N_3903,N_3389,N_3204);
or U3904 (N_3904,N_3379,N_3165);
or U3905 (N_3905,N_3191,N_3497);
and U3906 (N_3906,N_3336,N_3470);
xor U3907 (N_3907,N_3346,N_3178);
and U3908 (N_3908,N_3407,N_3141);
xnor U3909 (N_3909,N_3003,N_3111);
nor U3910 (N_3910,N_3083,N_3006);
or U3911 (N_3911,N_3492,N_3361);
nor U3912 (N_3912,N_3432,N_3227);
and U3913 (N_3913,N_3390,N_3224);
or U3914 (N_3914,N_3321,N_3145);
nand U3915 (N_3915,N_3099,N_3405);
or U3916 (N_3916,N_3198,N_3078);
nand U3917 (N_3917,N_3433,N_3008);
nand U3918 (N_3918,N_3055,N_3221);
nor U3919 (N_3919,N_3218,N_3258);
xnor U3920 (N_3920,N_3451,N_3314);
xnor U3921 (N_3921,N_3050,N_3105);
and U3922 (N_3922,N_3023,N_3210);
or U3923 (N_3923,N_3035,N_3234);
or U3924 (N_3924,N_3483,N_3244);
or U3925 (N_3925,N_3184,N_3152);
nand U3926 (N_3926,N_3090,N_3369);
and U3927 (N_3927,N_3114,N_3169);
nor U3928 (N_3928,N_3131,N_3090);
nor U3929 (N_3929,N_3499,N_3378);
nor U3930 (N_3930,N_3007,N_3372);
xor U3931 (N_3931,N_3111,N_3412);
and U3932 (N_3932,N_3304,N_3494);
and U3933 (N_3933,N_3237,N_3173);
and U3934 (N_3934,N_3004,N_3363);
xnor U3935 (N_3935,N_3493,N_3387);
xor U3936 (N_3936,N_3210,N_3490);
nand U3937 (N_3937,N_3373,N_3193);
nand U3938 (N_3938,N_3453,N_3053);
xor U3939 (N_3939,N_3249,N_3215);
nand U3940 (N_3940,N_3434,N_3315);
and U3941 (N_3941,N_3210,N_3274);
nand U3942 (N_3942,N_3016,N_3339);
nand U3943 (N_3943,N_3154,N_3143);
xor U3944 (N_3944,N_3311,N_3231);
xnor U3945 (N_3945,N_3386,N_3208);
and U3946 (N_3946,N_3097,N_3415);
nor U3947 (N_3947,N_3497,N_3184);
or U3948 (N_3948,N_3078,N_3297);
nor U3949 (N_3949,N_3086,N_3283);
or U3950 (N_3950,N_3291,N_3333);
nor U3951 (N_3951,N_3078,N_3169);
nand U3952 (N_3952,N_3141,N_3437);
xnor U3953 (N_3953,N_3119,N_3346);
nand U3954 (N_3954,N_3370,N_3489);
nor U3955 (N_3955,N_3003,N_3280);
and U3956 (N_3956,N_3159,N_3134);
xor U3957 (N_3957,N_3264,N_3067);
nor U3958 (N_3958,N_3002,N_3258);
or U3959 (N_3959,N_3092,N_3200);
nand U3960 (N_3960,N_3120,N_3074);
or U3961 (N_3961,N_3196,N_3399);
xor U3962 (N_3962,N_3342,N_3315);
nand U3963 (N_3963,N_3125,N_3275);
nor U3964 (N_3964,N_3478,N_3139);
and U3965 (N_3965,N_3030,N_3190);
or U3966 (N_3966,N_3284,N_3031);
nor U3967 (N_3967,N_3189,N_3456);
or U3968 (N_3968,N_3151,N_3018);
nor U3969 (N_3969,N_3306,N_3428);
and U3970 (N_3970,N_3175,N_3199);
or U3971 (N_3971,N_3375,N_3333);
nor U3972 (N_3972,N_3123,N_3095);
or U3973 (N_3973,N_3116,N_3189);
nand U3974 (N_3974,N_3095,N_3341);
nand U3975 (N_3975,N_3124,N_3468);
nand U3976 (N_3976,N_3018,N_3038);
xnor U3977 (N_3977,N_3018,N_3126);
xnor U3978 (N_3978,N_3068,N_3039);
or U3979 (N_3979,N_3078,N_3374);
and U3980 (N_3980,N_3236,N_3424);
nand U3981 (N_3981,N_3391,N_3419);
nand U3982 (N_3982,N_3062,N_3415);
xnor U3983 (N_3983,N_3068,N_3271);
xnor U3984 (N_3984,N_3245,N_3371);
nand U3985 (N_3985,N_3055,N_3355);
nand U3986 (N_3986,N_3046,N_3345);
or U3987 (N_3987,N_3466,N_3426);
or U3988 (N_3988,N_3121,N_3169);
or U3989 (N_3989,N_3014,N_3382);
or U3990 (N_3990,N_3126,N_3288);
xnor U3991 (N_3991,N_3448,N_3125);
and U3992 (N_3992,N_3425,N_3028);
xor U3993 (N_3993,N_3184,N_3252);
nand U3994 (N_3994,N_3208,N_3352);
and U3995 (N_3995,N_3254,N_3087);
nor U3996 (N_3996,N_3449,N_3481);
xnor U3997 (N_3997,N_3145,N_3165);
nor U3998 (N_3998,N_3430,N_3253);
nor U3999 (N_3999,N_3080,N_3184);
nand U4000 (N_4000,N_3812,N_3608);
and U4001 (N_4001,N_3753,N_3726);
nand U4002 (N_4002,N_3627,N_3752);
nor U4003 (N_4003,N_3574,N_3859);
and U4004 (N_4004,N_3618,N_3768);
and U4005 (N_4005,N_3815,N_3534);
or U4006 (N_4006,N_3542,N_3703);
and U4007 (N_4007,N_3502,N_3868);
and U4008 (N_4008,N_3748,N_3723);
xnor U4009 (N_4009,N_3702,N_3897);
xor U4010 (N_4010,N_3934,N_3952);
nor U4011 (N_4011,N_3580,N_3631);
and U4012 (N_4012,N_3509,N_3557);
nand U4013 (N_4013,N_3535,N_3654);
nand U4014 (N_4014,N_3544,N_3762);
nand U4015 (N_4015,N_3829,N_3609);
nand U4016 (N_4016,N_3983,N_3782);
xnor U4017 (N_4017,N_3927,N_3976);
nand U4018 (N_4018,N_3882,N_3994);
or U4019 (N_4019,N_3809,N_3643);
or U4020 (N_4020,N_3827,N_3770);
xnor U4021 (N_4021,N_3811,N_3675);
or U4022 (N_4022,N_3517,N_3584);
or U4023 (N_4023,N_3792,N_3958);
xor U4024 (N_4024,N_3657,N_3674);
and U4025 (N_4025,N_3599,N_3521);
nand U4026 (N_4026,N_3567,N_3971);
nand U4027 (N_4027,N_3781,N_3734);
nand U4028 (N_4028,N_3755,N_3601);
and U4029 (N_4029,N_3769,N_3602);
nor U4030 (N_4030,N_3975,N_3805);
nand U4031 (N_4031,N_3759,N_3767);
nor U4032 (N_4032,N_3772,N_3801);
xnor U4033 (N_4033,N_3948,N_3757);
nor U4034 (N_4034,N_3523,N_3932);
xnor U4035 (N_4035,N_3662,N_3735);
xor U4036 (N_4036,N_3854,N_3558);
or U4037 (N_4037,N_3501,N_3559);
or U4038 (N_4038,N_3921,N_3705);
nand U4039 (N_4039,N_3611,N_3615);
nand U4040 (N_4040,N_3655,N_3540);
xnor U4041 (N_4041,N_3986,N_3573);
nand U4042 (N_4042,N_3904,N_3933);
nor U4043 (N_4043,N_3585,N_3865);
or U4044 (N_4044,N_3862,N_3879);
xor U4045 (N_4045,N_3589,N_3842);
nand U4046 (N_4046,N_3858,N_3708);
nand U4047 (N_4047,N_3813,N_3784);
and U4048 (N_4048,N_3953,N_3505);
xnor U4049 (N_4049,N_3852,N_3909);
or U4050 (N_4050,N_3733,N_3962);
nand U4051 (N_4051,N_3890,N_3777);
xor U4052 (N_4052,N_3612,N_3774);
or U4053 (N_4053,N_3543,N_3889);
xor U4054 (N_4054,N_3530,N_3623);
and U4055 (N_4055,N_3649,N_3990);
and U4056 (N_4056,N_3931,N_3595);
and U4057 (N_4057,N_3626,N_3873);
and U4058 (N_4058,N_3856,N_3711);
xor U4059 (N_4059,N_3853,N_3714);
xor U4060 (N_4060,N_3709,N_3637);
nor U4061 (N_4061,N_3959,N_3855);
nor U4062 (N_4062,N_3713,N_3866);
and U4063 (N_4063,N_3681,N_3785);
or U4064 (N_4064,N_3954,N_3569);
nor U4065 (N_4065,N_3577,N_3652);
xor U4066 (N_4066,N_3835,N_3506);
xor U4067 (N_4067,N_3894,N_3957);
and U4068 (N_4068,N_3791,N_3514);
xor U4069 (N_4069,N_3686,N_3666);
xnor U4070 (N_4070,N_3508,N_3836);
and U4071 (N_4071,N_3789,N_3729);
and U4072 (N_4072,N_3997,N_3669);
or U4073 (N_4073,N_3594,N_3556);
nand U4074 (N_4074,N_3843,N_3683);
or U4075 (N_4075,N_3925,N_3749);
or U4076 (N_4076,N_3989,N_3916);
or U4077 (N_4077,N_3878,N_3846);
nand U4078 (N_4078,N_3597,N_3507);
and U4079 (N_4079,N_3562,N_3522);
nor U4080 (N_4080,N_3832,N_3533);
nor U4081 (N_4081,N_3511,N_3906);
or U4082 (N_4082,N_3902,N_3691);
or U4083 (N_4083,N_3678,N_3680);
and U4084 (N_4084,N_3717,N_3642);
xnor U4085 (N_4085,N_3775,N_3718);
or U4086 (N_4086,N_3780,N_3740);
or U4087 (N_4087,N_3870,N_3677);
or U4088 (N_4088,N_3564,N_3621);
nand U4089 (N_4089,N_3650,N_3788);
nand U4090 (N_4090,N_3583,N_3531);
nand U4091 (N_4091,N_3941,N_3880);
and U4092 (N_4092,N_3515,N_3869);
xor U4093 (N_4093,N_3824,N_3929);
nand U4094 (N_4094,N_3696,N_3992);
and U4095 (N_4095,N_3571,N_3946);
nor U4096 (N_4096,N_3687,N_3503);
nor U4097 (N_4097,N_3923,N_3742);
and U4098 (N_4098,N_3945,N_3779);
xnor U4099 (N_4099,N_3526,N_3908);
and U4100 (N_4100,N_3937,N_3978);
xnor U4101 (N_4101,N_3638,N_3525);
and U4102 (N_4102,N_3625,N_3797);
and U4103 (N_4103,N_3624,N_3684);
and U4104 (N_4104,N_3689,N_3539);
and U4105 (N_4105,N_3758,N_3529);
and U4106 (N_4106,N_3861,N_3596);
xor U4107 (N_4107,N_3950,N_3910);
nand U4108 (N_4108,N_3695,N_3560);
xnor U4109 (N_4109,N_3730,N_3587);
nor U4110 (N_4110,N_3619,N_3914);
nand U4111 (N_4111,N_3743,N_3613);
nor U4112 (N_4112,N_3776,N_3973);
nand U4113 (N_4113,N_3907,N_3938);
nand U4114 (N_4114,N_3722,N_3510);
xor U4115 (N_4115,N_3872,N_3874);
xnor U4116 (N_4116,N_3547,N_3598);
xnor U4117 (N_4117,N_3765,N_3831);
or U4118 (N_4118,N_3839,N_3693);
and U4119 (N_4119,N_3988,N_3548);
or U4120 (N_4120,N_3851,N_3778);
nand U4121 (N_4121,N_3817,N_3793);
nor U4122 (N_4122,N_3926,N_3947);
or U4123 (N_4123,N_3754,N_3712);
and U4124 (N_4124,N_3640,N_3924);
or U4125 (N_4125,N_3731,N_3935);
nor U4126 (N_4126,N_3885,N_3513);
nor U4127 (N_4127,N_3512,N_3527);
xor U4128 (N_4128,N_3578,N_3900);
nor U4129 (N_4129,N_3970,N_3636);
xor U4130 (N_4130,N_3773,N_3803);
or U4131 (N_4131,N_3984,N_3532);
or U4132 (N_4132,N_3746,N_3646);
nor U4133 (N_4133,N_3576,N_3998);
xnor U4134 (N_4134,N_3668,N_3566);
or U4135 (N_4135,N_3600,N_3982);
nor U4136 (N_4136,N_3592,N_3673);
or U4137 (N_4137,N_3806,N_3790);
or U4138 (N_4138,N_3555,N_3688);
nor U4139 (N_4139,N_3800,N_3896);
nor U4140 (N_4140,N_3725,N_3912);
nand U4141 (N_4141,N_3930,N_3710);
xnor U4142 (N_4142,N_3698,N_3605);
or U4143 (N_4143,N_3500,N_3645);
nand U4144 (N_4144,N_3991,N_3891);
xor U4145 (N_4145,N_3917,N_3575);
nor U4146 (N_4146,N_3802,N_3699);
xnor U4147 (N_4147,N_3922,N_3568);
xor U4148 (N_4148,N_3849,N_3732);
and U4149 (N_4149,N_3553,N_3750);
or U4150 (N_4150,N_3738,N_3648);
nor U4151 (N_4151,N_3617,N_3565);
xnor U4152 (N_4152,N_3760,N_3644);
nand U4153 (N_4153,N_3672,N_3951);
nand U4154 (N_4154,N_3972,N_3963);
nand U4155 (N_4155,N_3588,N_3647);
and U4156 (N_4156,N_3724,N_3867);
or U4157 (N_4157,N_3898,N_3787);
or U4158 (N_4158,N_3728,N_3814);
nand U4159 (N_4159,N_3936,N_3823);
nor U4160 (N_4160,N_3524,N_3996);
nand U4161 (N_4161,N_3821,N_3819);
nand U4162 (N_4162,N_3520,N_3629);
xnor U4163 (N_4163,N_3628,N_3993);
or U4164 (N_4164,N_3940,N_3607);
nand U4165 (N_4165,N_3545,N_3876);
xnor U4166 (N_4166,N_3561,N_3721);
and U4167 (N_4167,N_3603,N_3961);
xor U4168 (N_4168,N_3804,N_3579);
xnor U4169 (N_4169,N_3536,N_3707);
and U4170 (N_4170,N_3816,N_3664);
xor U4171 (N_4171,N_3554,N_3719);
or U4172 (N_4172,N_3877,N_3563);
nand U4173 (N_4173,N_3679,N_3883);
and U4174 (N_4174,N_3736,N_3670);
nor U4175 (N_4175,N_3949,N_3822);
or U4176 (N_4176,N_3622,N_3519);
xor U4177 (N_4177,N_3969,N_3895);
nor U4178 (N_4178,N_3786,N_3987);
xnor U4179 (N_4179,N_3834,N_3630);
nand U4180 (N_4180,N_3911,N_3960);
and U4181 (N_4181,N_3682,N_3651);
nor U4182 (N_4182,N_3838,N_3863);
and U4183 (N_4183,N_3999,N_3905);
nand U4184 (N_4184,N_3884,N_3604);
or U4185 (N_4185,N_3761,N_3860);
nand U4186 (N_4186,N_3826,N_3593);
nor U4187 (N_4187,N_3572,N_3632);
nand U4188 (N_4188,N_3541,N_3964);
nor U4189 (N_4189,N_3528,N_3901);
nor U4190 (N_4190,N_3979,N_3968);
xor U4191 (N_4191,N_3701,N_3704);
xor U4192 (N_4192,N_3844,N_3537);
xor U4193 (N_4193,N_3766,N_3985);
nand U4194 (N_4194,N_3659,N_3538);
and U4195 (N_4195,N_3833,N_3771);
or U4196 (N_4196,N_3614,N_3639);
nor U4197 (N_4197,N_3763,N_3837);
and U4198 (N_4198,N_3518,N_3706);
xnor U4199 (N_4199,N_3516,N_3915);
xnor U4200 (N_4200,N_3825,N_3848);
xor U4201 (N_4201,N_3549,N_3918);
and U4202 (N_4202,N_3692,N_3658);
and U4203 (N_4203,N_3810,N_3606);
xnor U4204 (N_4204,N_3751,N_3840);
nor U4205 (N_4205,N_3665,N_3956);
nand U4206 (N_4206,N_3697,N_3888);
xnor U4207 (N_4207,N_3995,N_3764);
and U4208 (N_4208,N_3828,N_3570);
xnor U4209 (N_4209,N_3955,N_3716);
xnor U4210 (N_4210,N_3841,N_3620);
nand U4211 (N_4211,N_3974,N_3820);
xor U4212 (N_4212,N_3980,N_3756);
and U4213 (N_4213,N_3667,N_3794);
nor U4214 (N_4214,N_3807,N_3641);
and U4215 (N_4215,N_3942,N_3818);
nor U4216 (N_4216,N_3864,N_3977);
or U4217 (N_4217,N_3944,N_3965);
nand U4218 (N_4218,N_3634,N_3913);
nand U4219 (N_4219,N_3700,N_3887);
nor U4220 (N_4220,N_3967,N_3720);
xor U4221 (N_4221,N_3727,N_3656);
or U4222 (N_4222,N_3881,N_3830);
nand U4223 (N_4223,N_3671,N_3783);
or U4224 (N_4224,N_3660,N_3850);
or U4225 (N_4225,N_3808,N_3581);
and U4226 (N_4226,N_3920,N_3610);
nor U4227 (N_4227,N_3899,N_3893);
xnor U4228 (N_4228,N_3616,N_3676);
and U4229 (N_4229,N_3847,N_3795);
nand U4230 (N_4230,N_3966,N_3745);
and U4231 (N_4231,N_3892,N_3737);
nand U4232 (N_4232,N_3744,N_3635);
xnor U4233 (N_4233,N_3939,N_3591);
or U4234 (N_4234,N_3690,N_3633);
xnor U4235 (N_4235,N_3715,N_3875);
and U4236 (N_4236,N_3871,N_3582);
nand U4237 (N_4237,N_3694,N_3504);
nor U4238 (N_4238,N_3685,N_3590);
nand U4239 (N_4239,N_3546,N_3796);
or U4240 (N_4240,N_3747,N_3552);
nand U4241 (N_4241,N_3903,N_3550);
nor U4242 (N_4242,N_3739,N_3845);
nor U4243 (N_4243,N_3981,N_3919);
and U4244 (N_4244,N_3798,N_3663);
xor U4245 (N_4245,N_3799,N_3586);
or U4246 (N_4246,N_3857,N_3928);
nand U4247 (N_4247,N_3741,N_3886);
xor U4248 (N_4248,N_3551,N_3661);
and U4249 (N_4249,N_3653,N_3943);
xor U4250 (N_4250,N_3734,N_3724);
nor U4251 (N_4251,N_3925,N_3666);
or U4252 (N_4252,N_3839,N_3911);
and U4253 (N_4253,N_3756,N_3848);
xnor U4254 (N_4254,N_3622,N_3557);
xor U4255 (N_4255,N_3956,N_3687);
xnor U4256 (N_4256,N_3883,N_3874);
nor U4257 (N_4257,N_3716,N_3679);
xnor U4258 (N_4258,N_3933,N_3992);
nor U4259 (N_4259,N_3648,N_3890);
nand U4260 (N_4260,N_3514,N_3740);
nor U4261 (N_4261,N_3888,N_3770);
nor U4262 (N_4262,N_3507,N_3720);
xor U4263 (N_4263,N_3619,N_3560);
xor U4264 (N_4264,N_3831,N_3651);
xor U4265 (N_4265,N_3957,N_3866);
nand U4266 (N_4266,N_3509,N_3680);
and U4267 (N_4267,N_3584,N_3877);
nor U4268 (N_4268,N_3525,N_3645);
xnor U4269 (N_4269,N_3740,N_3788);
nor U4270 (N_4270,N_3628,N_3873);
xnor U4271 (N_4271,N_3560,N_3919);
and U4272 (N_4272,N_3511,N_3694);
or U4273 (N_4273,N_3632,N_3511);
or U4274 (N_4274,N_3840,N_3838);
or U4275 (N_4275,N_3939,N_3567);
xor U4276 (N_4276,N_3835,N_3809);
or U4277 (N_4277,N_3923,N_3980);
xor U4278 (N_4278,N_3648,N_3543);
nor U4279 (N_4279,N_3524,N_3629);
and U4280 (N_4280,N_3928,N_3604);
or U4281 (N_4281,N_3832,N_3602);
nand U4282 (N_4282,N_3910,N_3723);
nand U4283 (N_4283,N_3994,N_3666);
or U4284 (N_4284,N_3528,N_3956);
nor U4285 (N_4285,N_3962,N_3869);
or U4286 (N_4286,N_3614,N_3755);
and U4287 (N_4287,N_3644,N_3694);
and U4288 (N_4288,N_3988,N_3981);
or U4289 (N_4289,N_3799,N_3617);
nor U4290 (N_4290,N_3640,N_3785);
or U4291 (N_4291,N_3750,N_3716);
nand U4292 (N_4292,N_3775,N_3837);
nand U4293 (N_4293,N_3526,N_3990);
nand U4294 (N_4294,N_3751,N_3564);
and U4295 (N_4295,N_3841,N_3742);
nand U4296 (N_4296,N_3735,N_3568);
or U4297 (N_4297,N_3678,N_3744);
or U4298 (N_4298,N_3639,N_3653);
nand U4299 (N_4299,N_3709,N_3847);
nor U4300 (N_4300,N_3537,N_3883);
xor U4301 (N_4301,N_3660,N_3552);
or U4302 (N_4302,N_3927,N_3517);
nand U4303 (N_4303,N_3911,N_3986);
nand U4304 (N_4304,N_3812,N_3999);
and U4305 (N_4305,N_3592,N_3978);
nor U4306 (N_4306,N_3640,N_3580);
xnor U4307 (N_4307,N_3642,N_3920);
and U4308 (N_4308,N_3779,N_3738);
or U4309 (N_4309,N_3741,N_3896);
nor U4310 (N_4310,N_3504,N_3620);
and U4311 (N_4311,N_3684,N_3685);
xor U4312 (N_4312,N_3682,N_3587);
xor U4313 (N_4313,N_3830,N_3769);
and U4314 (N_4314,N_3763,N_3944);
or U4315 (N_4315,N_3696,N_3506);
nand U4316 (N_4316,N_3559,N_3647);
nand U4317 (N_4317,N_3518,N_3924);
xnor U4318 (N_4318,N_3959,N_3799);
nand U4319 (N_4319,N_3612,N_3989);
nor U4320 (N_4320,N_3824,N_3951);
nor U4321 (N_4321,N_3963,N_3767);
nor U4322 (N_4322,N_3596,N_3586);
or U4323 (N_4323,N_3966,N_3778);
or U4324 (N_4324,N_3766,N_3909);
and U4325 (N_4325,N_3815,N_3633);
nor U4326 (N_4326,N_3911,N_3774);
or U4327 (N_4327,N_3968,N_3771);
or U4328 (N_4328,N_3670,N_3923);
xor U4329 (N_4329,N_3758,N_3941);
nand U4330 (N_4330,N_3933,N_3694);
and U4331 (N_4331,N_3969,N_3760);
or U4332 (N_4332,N_3779,N_3812);
xor U4333 (N_4333,N_3934,N_3516);
nor U4334 (N_4334,N_3557,N_3922);
and U4335 (N_4335,N_3544,N_3508);
xor U4336 (N_4336,N_3547,N_3656);
nand U4337 (N_4337,N_3656,N_3575);
or U4338 (N_4338,N_3662,N_3837);
nand U4339 (N_4339,N_3919,N_3789);
nor U4340 (N_4340,N_3704,N_3979);
and U4341 (N_4341,N_3766,N_3908);
nor U4342 (N_4342,N_3714,N_3625);
nor U4343 (N_4343,N_3993,N_3789);
nand U4344 (N_4344,N_3616,N_3758);
and U4345 (N_4345,N_3887,N_3619);
or U4346 (N_4346,N_3743,N_3596);
nor U4347 (N_4347,N_3934,N_3792);
nor U4348 (N_4348,N_3683,N_3773);
nand U4349 (N_4349,N_3764,N_3997);
xnor U4350 (N_4350,N_3648,N_3761);
xor U4351 (N_4351,N_3891,N_3560);
or U4352 (N_4352,N_3616,N_3784);
xnor U4353 (N_4353,N_3812,N_3738);
or U4354 (N_4354,N_3838,N_3980);
nand U4355 (N_4355,N_3698,N_3550);
nor U4356 (N_4356,N_3839,N_3943);
nand U4357 (N_4357,N_3583,N_3882);
or U4358 (N_4358,N_3617,N_3629);
nor U4359 (N_4359,N_3762,N_3764);
xnor U4360 (N_4360,N_3533,N_3827);
nor U4361 (N_4361,N_3947,N_3621);
xor U4362 (N_4362,N_3591,N_3561);
nand U4363 (N_4363,N_3894,N_3994);
xor U4364 (N_4364,N_3503,N_3897);
nand U4365 (N_4365,N_3776,N_3839);
nand U4366 (N_4366,N_3831,N_3682);
and U4367 (N_4367,N_3725,N_3693);
or U4368 (N_4368,N_3531,N_3669);
or U4369 (N_4369,N_3645,N_3560);
xor U4370 (N_4370,N_3648,N_3694);
and U4371 (N_4371,N_3957,N_3571);
nor U4372 (N_4372,N_3560,N_3842);
or U4373 (N_4373,N_3688,N_3890);
nor U4374 (N_4374,N_3953,N_3908);
and U4375 (N_4375,N_3707,N_3963);
nand U4376 (N_4376,N_3913,N_3942);
or U4377 (N_4377,N_3932,N_3507);
nand U4378 (N_4378,N_3987,N_3671);
nand U4379 (N_4379,N_3687,N_3949);
nor U4380 (N_4380,N_3530,N_3817);
nor U4381 (N_4381,N_3762,N_3980);
nand U4382 (N_4382,N_3510,N_3614);
xor U4383 (N_4383,N_3526,N_3975);
or U4384 (N_4384,N_3674,N_3897);
xnor U4385 (N_4385,N_3776,N_3773);
and U4386 (N_4386,N_3966,N_3712);
nor U4387 (N_4387,N_3537,N_3889);
nand U4388 (N_4388,N_3957,N_3738);
xor U4389 (N_4389,N_3823,N_3667);
xor U4390 (N_4390,N_3957,N_3703);
or U4391 (N_4391,N_3654,N_3505);
xor U4392 (N_4392,N_3762,N_3821);
or U4393 (N_4393,N_3762,N_3625);
and U4394 (N_4394,N_3959,N_3985);
nand U4395 (N_4395,N_3837,N_3684);
nor U4396 (N_4396,N_3908,N_3781);
nor U4397 (N_4397,N_3580,N_3540);
and U4398 (N_4398,N_3815,N_3971);
and U4399 (N_4399,N_3585,N_3599);
and U4400 (N_4400,N_3849,N_3794);
or U4401 (N_4401,N_3686,N_3921);
nand U4402 (N_4402,N_3727,N_3929);
xnor U4403 (N_4403,N_3752,N_3509);
nor U4404 (N_4404,N_3727,N_3984);
nand U4405 (N_4405,N_3847,N_3652);
or U4406 (N_4406,N_3932,N_3500);
and U4407 (N_4407,N_3912,N_3858);
and U4408 (N_4408,N_3699,N_3940);
xor U4409 (N_4409,N_3828,N_3652);
nand U4410 (N_4410,N_3679,N_3595);
nand U4411 (N_4411,N_3766,N_3914);
xnor U4412 (N_4412,N_3761,N_3810);
nor U4413 (N_4413,N_3687,N_3881);
and U4414 (N_4414,N_3542,N_3958);
xor U4415 (N_4415,N_3891,N_3688);
and U4416 (N_4416,N_3963,N_3817);
or U4417 (N_4417,N_3969,N_3684);
xor U4418 (N_4418,N_3769,N_3656);
xnor U4419 (N_4419,N_3855,N_3970);
nor U4420 (N_4420,N_3837,N_3853);
or U4421 (N_4421,N_3970,N_3856);
nand U4422 (N_4422,N_3553,N_3821);
and U4423 (N_4423,N_3855,N_3933);
nand U4424 (N_4424,N_3603,N_3879);
nor U4425 (N_4425,N_3616,N_3829);
nand U4426 (N_4426,N_3732,N_3713);
xnor U4427 (N_4427,N_3855,N_3771);
nor U4428 (N_4428,N_3768,N_3993);
nor U4429 (N_4429,N_3547,N_3702);
xnor U4430 (N_4430,N_3572,N_3867);
nand U4431 (N_4431,N_3525,N_3654);
nor U4432 (N_4432,N_3923,N_3834);
and U4433 (N_4433,N_3601,N_3988);
nor U4434 (N_4434,N_3620,N_3524);
and U4435 (N_4435,N_3694,N_3955);
xnor U4436 (N_4436,N_3870,N_3800);
and U4437 (N_4437,N_3754,N_3622);
nor U4438 (N_4438,N_3541,N_3554);
or U4439 (N_4439,N_3668,N_3612);
nand U4440 (N_4440,N_3929,N_3956);
nand U4441 (N_4441,N_3546,N_3971);
nor U4442 (N_4442,N_3750,N_3920);
and U4443 (N_4443,N_3551,N_3598);
or U4444 (N_4444,N_3542,N_3821);
xor U4445 (N_4445,N_3657,N_3527);
or U4446 (N_4446,N_3795,N_3906);
nand U4447 (N_4447,N_3898,N_3552);
nand U4448 (N_4448,N_3945,N_3673);
nand U4449 (N_4449,N_3539,N_3877);
and U4450 (N_4450,N_3661,N_3544);
and U4451 (N_4451,N_3555,N_3835);
nand U4452 (N_4452,N_3548,N_3832);
nor U4453 (N_4453,N_3989,N_3677);
nand U4454 (N_4454,N_3949,N_3852);
nand U4455 (N_4455,N_3580,N_3791);
or U4456 (N_4456,N_3583,N_3962);
nand U4457 (N_4457,N_3911,N_3982);
nor U4458 (N_4458,N_3827,N_3576);
or U4459 (N_4459,N_3641,N_3992);
xor U4460 (N_4460,N_3904,N_3986);
xnor U4461 (N_4461,N_3691,N_3980);
xor U4462 (N_4462,N_3582,N_3878);
nand U4463 (N_4463,N_3657,N_3873);
nand U4464 (N_4464,N_3883,N_3520);
or U4465 (N_4465,N_3624,N_3766);
nor U4466 (N_4466,N_3784,N_3852);
or U4467 (N_4467,N_3967,N_3857);
nor U4468 (N_4468,N_3937,N_3783);
nand U4469 (N_4469,N_3611,N_3746);
nand U4470 (N_4470,N_3759,N_3755);
or U4471 (N_4471,N_3877,N_3594);
nor U4472 (N_4472,N_3633,N_3538);
xnor U4473 (N_4473,N_3527,N_3858);
nor U4474 (N_4474,N_3676,N_3683);
and U4475 (N_4475,N_3962,N_3739);
xnor U4476 (N_4476,N_3612,N_3976);
nor U4477 (N_4477,N_3660,N_3876);
nor U4478 (N_4478,N_3975,N_3928);
nor U4479 (N_4479,N_3982,N_3903);
or U4480 (N_4480,N_3606,N_3876);
nor U4481 (N_4481,N_3920,N_3632);
nor U4482 (N_4482,N_3627,N_3690);
and U4483 (N_4483,N_3672,N_3794);
nand U4484 (N_4484,N_3956,N_3899);
xnor U4485 (N_4485,N_3866,N_3637);
and U4486 (N_4486,N_3579,N_3728);
xor U4487 (N_4487,N_3958,N_3718);
xnor U4488 (N_4488,N_3520,N_3719);
nand U4489 (N_4489,N_3521,N_3917);
and U4490 (N_4490,N_3665,N_3846);
or U4491 (N_4491,N_3951,N_3665);
xnor U4492 (N_4492,N_3610,N_3707);
nand U4493 (N_4493,N_3953,N_3618);
and U4494 (N_4494,N_3561,N_3951);
nand U4495 (N_4495,N_3630,N_3560);
nand U4496 (N_4496,N_3860,N_3886);
and U4497 (N_4497,N_3686,N_3612);
and U4498 (N_4498,N_3509,N_3600);
xor U4499 (N_4499,N_3763,N_3543);
xnor U4500 (N_4500,N_4105,N_4259);
or U4501 (N_4501,N_4121,N_4173);
and U4502 (N_4502,N_4056,N_4260);
or U4503 (N_4503,N_4469,N_4099);
or U4504 (N_4504,N_4077,N_4395);
and U4505 (N_4505,N_4083,N_4413);
xor U4506 (N_4506,N_4135,N_4000);
or U4507 (N_4507,N_4347,N_4479);
and U4508 (N_4508,N_4127,N_4404);
nand U4509 (N_4509,N_4444,N_4346);
or U4510 (N_4510,N_4217,N_4033);
nor U4511 (N_4511,N_4451,N_4115);
nand U4512 (N_4512,N_4351,N_4252);
nand U4513 (N_4513,N_4380,N_4468);
xor U4514 (N_4514,N_4063,N_4234);
nand U4515 (N_4515,N_4097,N_4279);
or U4516 (N_4516,N_4406,N_4455);
nor U4517 (N_4517,N_4006,N_4074);
and U4518 (N_4518,N_4283,N_4141);
xor U4519 (N_4519,N_4303,N_4355);
xor U4520 (N_4520,N_4409,N_4493);
or U4521 (N_4521,N_4086,N_4071);
xor U4522 (N_4522,N_4136,N_4463);
or U4523 (N_4523,N_4341,N_4179);
xor U4524 (N_4524,N_4453,N_4011);
and U4525 (N_4525,N_4288,N_4114);
xor U4526 (N_4526,N_4198,N_4315);
nor U4527 (N_4527,N_4297,N_4250);
xnor U4528 (N_4528,N_4045,N_4080);
nor U4529 (N_4529,N_4075,N_4160);
nand U4530 (N_4530,N_4427,N_4344);
and U4531 (N_4531,N_4372,N_4123);
nor U4532 (N_4532,N_4428,N_4248);
nand U4533 (N_4533,N_4254,N_4324);
nor U4534 (N_4534,N_4014,N_4354);
nand U4535 (N_4535,N_4214,N_4246);
xnor U4536 (N_4536,N_4041,N_4102);
xor U4537 (N_4537,N_4161,N_4447);
xor U4538 (N_4538,N_4226,N_4300);
nand U4539 (N_4539,N_4302,N_4025);
or U4540 (N_4540,N_4332,N_4164);
nand U4541 (N_4541,N_4122,N_4239);
or U4542 (N_4542,N_4190,N_4233);
xnor U4543 (N_4543,N_4415,N_4094);
nand U4544 (N_4544,N_4058,N_4130);
nand U4545 (N_4545,N_4282,N_4062);
and U4546 (N_4546,N_4081,N_4445);
or U4547 (N_4547,N_4399,N_4436);
or U4548 (N_4548,N_4256,N_4112);
nand U4549 (N_4549,N_4417,N_4365);
and U4550 (N_4550,N_4481,N_4392);
and U4551 (N_4551,N_4047,N_4118);
xor U4552 (N_4552,N_4318,N_4496);
xor U4553 (N_4553,N_4420,N_4472);
xor U4554 (N_4554,N_4319,N_4325);
nand U4555 (N_4555,N_4187,N_4188);
and U4556 (N_4556,N_4433,N_4322);
and U4557 (N_4557,N_4040,N_4490);
nor U4558 (N_4558,N_4360,N_4036);
nor U4559 (N_4559,N_4208,N_4009);
nand U4560 (N_4560,N_4206,N_4059);
and U4561 (N_4561,N_4383,N_4305);
xor U4562 (N_4562,N_4416,N_4317);
and U4563 (N_4563,N_4342,N_4480);
xor U4564 (N_4564,N_4149,N_4159);
nor U4565 (N_4565,N_4477,N_4065);
xor U4566 (N_4566,N_4350,N_4263);
or U4567 (N_4567,N_4334,N_4143);
or U4568 (N_4568,N_4189,N_4138);
xnor U4569 (N_4569,N_4157,N_4090);
xnor U4570 (N_4570,N_4343,N_4264);
nor U4571 (N_4571,N_4061,N_4460);
xor U4572 (N_4572,N_4113,N_4398);
nand U4573 (N_4573,N_4269,N_4464);
and U4574 (N_4574,N_4111,N_4128);
xnor U4575 (N_4575,N_4396,N_4022);
xnor U4576 (N_4576,N_4265,N_4275);
xnor U4577 (N_4577,N_4196,N_4170);
xnor U4578 (N_4578,N_4418,N_4280);
or U4579 (N_4579,N_4311,N_4219);
xor U4580 (N_4580,N_4296,N_4287);
nor U4581 (N_4581,N_4085,N_4032);
or U4582 (N_4582,N_4419,N_4229);
nand U4583 (N_4583,N_4457,N_4154);
and U4584 (N_4584,N_4374,N_4235);
nor U4585 (N_4585,N_4446,N_4377);
or U4586 (N_4586,N_4211,N_4262);
and U4587 (N_4587,N_4035,N_4495);
xnor U4588 (N_4588,N_4001,N_4470);
nor U4589 (N_4589,N_4004,N_4096);
xor U4590 (N_4590,N_4371,N_4023);
nand U4591 (N_4591,N_4176,N_4438);
xor U4592 (N_4592,N_4203,N_4223);
or U4593 (N_4593,N_4289,N_4379);
and U4594 (N_4594,N_4232,N_4320);
xnor U4595 (N_4595,N_4313,N_4168);
or U4596 (N_4596,N_4078,N_4201);
nand U4597 (N_4597,N_4192,N_4244);
nand U4598 (N_4598,N_4057,N_4349);
and U4599 (N_4599,N_4142,N_4278);
nand U4600 (N_4600,N_4104,N_4020);
and U4601 (N_4601,N_4156,N_4465);
nand U4602 (N_4602,N_4301,N_4434);
or U4603 (N_4603,N_4286,N_4306);
or U4604 (N_4604,N_4100,N_4166);
nand U4605 (N_4605,N_4281,N_4184);
nor U4606 (N_4606,N_4145,N_4109);
nor U4607 (N_4607,N_4304,N_4027);
nor U4608 (N_4608,N_4221,N_4255);
xnor U4609 (N_4609,N_4017,N_4437);
and U4610 (N_4610,N_4331,N_4373);
nor U4611 (N_4611,N_4378,N_4044);
or U4612 (N_4612,N_4243,N_4180);
and U4613 (N_4613,N_4454,N_4367);
and U4614 (N_4614,N_4362,N_4107);
nor U4615 (N_4615,N_4284,N_4034);
and U4616 (N_4616,N_4340,N_4258);
nand U4617 (N_4617,N_4484,N_4019);
nand U4618 (N_4618,N_4220,N_4067);
or U4619 (N_4619,N_4052,N_4150);
or U4620 (N_4620,N_4273,N_4467);
xor U4621 (N_4621,N_4345,N_4125);
nand U4622 (N_4622,N_4441,N_4240);
nor U4623 (N_4623,N_4440,N_4016);
and U4624 (N_4624,N_4224,N_4400);
nor U4625 (N_4625,N_4298,N_4162);
and U4626 (N_4626,N_4394,N_4316);
or U4627 (N_4627,N_4486,N_4257);
or U4628 (N_4628,N_4386,N_4294);
nand U4629 (N_4629,N_4266,N_4356);
nor U4630 (N_4630,N_4018,N_4411);
or U4631 (N_4631,N_4382,N_4124);
or U4632 (N_4632,N_4483,N_4402);
and U4633 (N_4633,N_4106,N_4195);
or U4634 (N_4634,N_4155,N_4238);
nor U4635 (N_4635,N_4326,N_4485);
xnor U4636 (N_4636,N_4348,N_4171);
and U4637 (N_4637,N_4426,N_4037);
xor U4638 (N_4638,N_4291,N_4271);
nor U4639 (N_4639,N_4132,N_4012);
nand U4640 (N_4640,N_4497,N_4225);
nor U4641 (N_4641,N_4309,N_4335);
nor U4642 (N_4642,N_4439,N_4144);
or U4643 (N_4643,N_4376,N_4274);
nor U4644 (N_4644,N_4370,N_4007);
and U4645 (N_4645,N_4277,N_4227);
xnor U4646 (N_4646,N_4448,N_4363);
and U4647 (N_4647,N_4388,N_4393);
nor U4648 (N_4648,N_4352,N_4423);
and U4649 (N_4649,N_4055,N_4381);
and U4650 (N_4650,N_4333,N_4270);
or U4651 (N_4651,N_4177,N_4401);
xor U4652 (N_4652,N_4131,N_4133);
nand U4653 (N_4653,N_4222,N_4432);
nor U4654 (N_4654,N_4048,N_4200);
nand U4655 (N_4655,N_4163,N_4053);
nand U4656 (N_4656,N_4169,N_4435);
xor U4657 (N_4657,N_4430,N_4307);
or U4658 (N_4658,N_4153,N_4207);
xor U4659 (N_4659,N_4414,N_4199);
xnor U4660 (N_4660,N_4236,N_4237);
and U4661 (N_4661,N_4231,N_4389);
xnor U4662 (N_4662,N_4029,N_4049);
nand U4663 (N_4663,N_4116,N_4405);
nor U4664 (N_4664,N_4272,N_4101);
and U4665 (N_4665,N_4013,N_4174);
xnor U4666 (N_4666,N_4499,N_4494);
nor U4667 (N_4667,N_4197,N_4407);
and U4668 (N_4668,N_4152,N_4043);
or U4669 (N_4669,N_4194,N_4060);
nand U4670 (N_4670,N_4292,N_4475);
nand U4671 (N_4671,N_4148,N_4218);
nor U4672 (N_4672,N_4366,N_4321);
or U4673 (N_4673,N_4461,N_4146);
nand U4674 (N_4674,N_4183,N_4204);
xnor U4675 (N_4675,N_4073,N_4165);
nand U4676 (N_4676,N_4488,N_4357);
nand U4677 (N_4677,N_4491,N_4005);
or U4678 (N_4678,N_4103,N_4337);
xnor U4679 (N_4679,N_4425,N_4253);
nor U4680 (N_4680,N_4230,N_4158);
nand U4681 (N_4681,N_4046,N_4110);
nor U4682 (N_4682,N_4482,N_4421);
nand U4683 (N_4683,N_4329,N_4242);
xor U4684 (N_4684,N_4087,N_4247);
and U4685 (N_4685,N_4010,N_4205);
xnor U4686 (N_4686,N_4353,N_4129);
or U4687 (N_4687,N_4456,N_4471);
xor U4688 (N_4688,N_4098,N_4368);
nor U4689 (N_4689,N_4002,N_4095);
nand U4690 (N_4690,N_4068,N_4361);
xor U4691 (N_4691,N_4391,N_4358);
nor U4692 (N_4692,N_4290,N_4185);
xnor U4693 (N_4693,N_4069,N_4450);
nor U4694 (N_4694,N_4338,N_4431);
xnor U4695 (N_4695,N_4030,N_4015);
nand U4696 (N_4696,N_4108,N_4092);
and U4697 (N_4697,N_4228,N_4178);
and U4698 (N_4698,N_4093,N_4251);
and U4699 (N_4699,N_4091,N_4193);
or U4700 (N_4700,N_4139,N_4167);
or U4701 (N_4701,N_4498,N_4489);
nor U4702 (N_4702,N_4210,N_4385);
or U4703 (N_4703,N_4293,N_4397);
nand U4704 (N_4704,N_4449,N_4462);
nor U4705 (N_4705,N_4314,N_4212);
and U4706 (N_4706,N_4323,N_4089);
xor U4707 (N_4707,N_4117,N_4299);
or U4708 (N_4708,N_4175,N_4459);
xor U4709 (N_4709,N_4458,N_4492);
or U4710 (N_4710,N_4051,N_4245);
nand U4711 (N_4711,N_4137,N_4066);
or U4712 (N_4712,N_4126,N_4327);
nand U4713 (N_4713,N_4072,N_4120);
nor U4714 (N_4714,N_4364,N_4215);
xnor U4715 (N_4715,N_4186,N_4267);
nand U4716 (N_4716,N_4369,N_4202);
nand U4717 (N_4717,N_4330,N_4261);
or U4718 (N_4718,N_4336,N_4308);
and U4719 (N_4719,N_4042,N_4410);
and U4720 (N_4720,N_4429,N_4424);
or U4721 (N_4721,N_4249,N_4403);
or U4722 (N_4722,N_4375,N_4172);
nand U4723 (N_4723,N_4339,N_4408);
and U4724 (N_4724,N_4079,N_4310);
xnor U4725 (N_4725,N_4359,N_4054);
nand U4726 (N_4726,N_4021,N_4241);
and U4727 (N_4727,N_4487,N_4084);
nor U4728 (N_4728,N_4276,N_4076);
and U4729 (N_4729,N_4390,N_4312);
and U4730 (N_4730,N_4119,N_4442);
nand U4731 (N_4731,N_4140,N_4328);
nor U4732 (N_4732,N_4384,N_4387);
and U4733 (N_4733,N_4050,N_4082);
xnor U4734 (N_4734,N_4466,N_4209);
nor U4735 (N_4735,N_4064,N_4268);
xnor U4736 (N_4736,N_4182,N_4422);
nand U4737 (N_4737,N_4452,N_4134);
nand U4738 (N_4738,N_4412,N_4039);
nand U4739 (N_4739,N_4295,N_4026);
or U4740 (N_4740,N_4181,N_4038);
and U4741 (N_4741,N_4474,N_4147);
nor U4742 (N_4742,N_4031,N_4151);
or U4743 (N_4743,N_4003,N_4216);
nor U4744 (N_4744,N_4213,N_4473);
xor U4745 (N_4745,N_4443,N_4285);
nand U4746 (N_4746,N_4024,N_4008);
xor U4747 (N_4747,N_4070,N_4478);
xor U4748 (N_4748,N_4191,N_4476);
and U4749 (N_4749,N_4088,N_4028);
xor U4750 (N_4750,N_4441,N_4034);
nand U4751 (N_4751,N_4402,N_4101);
nor U4752 (N_4752,N_4297,N_4092);
nor U4753 (N_4753,N_4021,N_4467);
nand U4754 (N_4754,N_4361,N_4031);
or U4755 (N_4755,N_4124,N_4498);
or U4756 (N_4756,N_4345,N_4445);
xnor U4757 (N_4757,N_4342,N_4263);
or U4758 (N_4758,N_4276,N_4244);
xnor U4759 (N_4759,N_4476,N_4447);
or U4760 (N_4760,N_4082,N_4203);
and U4761 (N_4761,N_4343,N_4184);
nor U4762 (N_4762,N_4287,N_4451);
and U4763 (N_4763,N_4422,N_4029);
or U4764 (N_4764,N_4001,N_4297);
nor U4765 (N_4765,N_4060,N_4016);
or U4766 (N_4766,N_4452,N_4206);
nor U4767 (N_4767,N_4406,N_4294);
or U4768 (N_4768,N_4212,N_4023);
nand U4769 (N_4769,N_4392,N_4327);
nand U4770 (N_4770,N_4185,N_4207);
nor U4771 (N_4771,N_4432,N_4358);
nor U4772 (N_4772,N_4004,N_4285);
nand U4773 (N_4773,N_4117,N_4228);
nand U4774 (N_4774,N_4380,N_4260);
or U4775 (N_4775,N_4199,N_4369);
nor U4776 (N_4776,N_4313,N_4055);
nand U4777 (N_4777,N_4008,N_4159);
nor U4778 (N_4778,N_4143,N_4313);
xor U4779 (N_4779,N_4141,N_4312);
xnor U4780 (N_4780,N_4174,N_4159);
and U4781 (N_4781,N_4026,N_4117);
nor U4782 (N_4782,N_4071,N_4038);
nor U4783 (N_4783,N_4233,N_4034);
xor U4784 (N_4784,N_4242,N_4124);
nand U4785 (N_4785,N_4463,N_4491);
and U4786 (N_4786,N_4248,N_4140);
nand U4787 (N_4787,N_4204,N_4400);
xnor U4788 (N_4788,N_4437,N_4233);
or U4789 (N_4789,N_4138,N_4013);
and U4790 (N_4790,N_4204,N_4261);
nand U4791 (N_4791,N_4130,N_4163);
or U4792 (N_4792,N_4350,N_4161);
nand U4793 (N_4793,N_4259,N_4457);
and U4794 (N_4794,N_4056,N_4316);
and U4795 (N_4795,N_4411,N_4326);
and U4796 (N_4796,N_4035,N_4376);
xor U4797 (N_4797,N_4158,N_4077);
nand U4798 (N_4798,N_4282,N_4254);
or U4799 (N_4799,N_4092,N_4089);
nor U4800 (N_4800,N_4102,N_4251);
or U4801 (N_4801,N_4295,N_4485);
nand U4802 (N_4802,N_4353,N_4085);
and U4803 (N_4803,N_4304,N_4437);
xor U4804 (N_4804,N_4074,N_4261);
nand U4805 (N_4805,N_4389,N_4468);
nand U4806 (N_4806,N_4375,N_4092);
nand U4807 (N_4807,N_4416,N_4438);
and U4808 (N_4808,N_4237,N_4199);
nor U4809 (N_4809,N_4118,N_4130);
or U4810 (N_4810,N_4181,N_4020);
xnor U4811 (N_4811,N_4028,N_4317);
or U4812 (N_4812,N_4332,N_4480);
xor U4813 (N_4813,N_4464,N_4129);
xor U4814 (N_4814,N_4105,N_4027);
or U4815 (N_4815,N_4190,N_4367);
xnor U4816 (N_4816,N_4197,N_4403);
xnor U4817 (N_4817,N_4129,N_4418);
and U4818 (N_4818,N_4492,N_4425);
and U4819 (N_4819,N_4247,N_4081);
and U4820 (N_4820,N_4277,N_4110);
nand U4821 (N_4821,N_4125,N_4356);
nor U4822 (N_4822,N_4096,N_4415);
or U4823 (N_4823,N_4447,N_4259);
and U4824 (N_4824,N_4091,N_4043);
or U4825 (N_4825,N_4354,N_4003);
xnor U4826 (N_4826,N_4392,N_4247);
nor U4827 (N_4827,N_4391,N_4067);
nand U4828 (N_4828,N_4347,N_4474);
nor U4829 (N_4829,N_4279,N_4353);
nor U4830 (N_4830,N_4114,N_4343);
and U4831 (N_4831,N_4282,N_4192);
and U4832 (N_4832,N_4350,N_4356);
and U4833 (N_4833,N_4008,N_4396);
nand U4834 (N_4834,N_4015,N_4208);
and U4835 (N_4835,N_4443,N_4301);
xnor U4836 (N_4836,N_4445,N_4084);
or U4837 (N_4837,N_4476,N_4152);
and U4838 (N_4838,N_4463,N_4214);
xnor U4839 (N_4839,N_4025,N_4261);
nand U4840 (N_4840,N_4031,N_4052);
nor U4841 (N_4841,N_4096,N_4423);
nor U4842 (N_4842,N_4008,N_4454);
xor U4843 (N_4843,N_4008,N_4490);
xor U4844 (N_4844,N_4127,N_4224);
nand U4845 (N_4845,N_4223,N_4194);
xnor U4846 (N_4846,N_4360,N_4262);
xor U4847 (N_4847,N_4362,N_4465);
xnor U4848 (N_4848,N_4324,N_4085);
nand U4849 (N_4849,N_4092,N_4218);
nand U4850 (N_4850,N_4491,N_4328);
nor U4851 (N_4851,N_4408,N_4306);
nor U4852 (N_4852,N_4095,N_4487);
and U4853 (N_4853,N_4195,N_4277);
xnor U4854 (N_4854,N_4182,N_4364);
nand U4855 (N_4855,N_4271,N_4004);
nor U4856 (N_4856,N_4034,N_4446);
nand U4857 (N_4857,N_4264,N_4246);
nand U4858 (N_4858,N_4355,N_4313);
xnor U4859 (N_4859,N_4465,N_4137);
xnor U4860 (N_4860,N_4016,N_4406);
nor U4861 (N_4861,N_4356,N_4401);
nand U4862 (N_4862,N_4406,N_4385);
xor U4863 (N_4863,N_4337,N_4324);
xor U4864 (N_4864,N_4068,N_4326);
nor U4865 (N_4865,N_4080,N_4090);
nor U4866 (N_4866,N_4371,N_4497);
nor U4867 (N_4867,N_4277,N_4472);
nand U4868 (N_4868,N_4317,N_4060);
xnor U4869 (N_4869,N_4028,N_4360);
xor U4870 (N_4870,N_4117,N_4351);
xor U4871 (N_4871,N_4432,N_4240);
xor U4872 (N_4872,N_4221,N_4411);
or U4873 (N_4873,N_4319,N_4208);
and U4874 (N_4874,N_4211,N_4151);
and U4875 (N_4875,N_4034,N_4372);
nor U4876 (N_4876,N_4208,N_4030);
xnor U4877 (N_4877,N_4073,N_4484);
and U4878 (N_4878,N_4176,N_4018);
nor U4879 (N_4879,N_4484,N_4466);
nor U4880 (N_4880,N_4292,N_4086);
xor U4881 (N_4881,N_4346,N_4138);
and U4882 (N_4882,N_4104,N_4223);
nand U4883 (N_4883,N_4021,N_4254);
xnor U4884 (N_4884,N_4036,N_4019);
or U4885 (N_4885,N_4145,N_4108);
or U4886 (N_4886,N_4186,N_4183);
or U4887 (N_4887,N_4296,N_4089);
xnor U4888 (N_4888,N_4279,N_4058);
or U4889 (N_4889,N_4092,N_4184);
and U4890 (N_4890,N_4383,N_4240);
and U4891 (N_4891,N_4468,N_4142);
xnor U4892 (N_4892,N_4317,N_4091);
or U4893 (N_4893,N_4188,N_4168);
nand U4894 (N_4894,N_4343,N_4353);
nand U4895 (N_4895,N_4094,N_4243);
or U4896 (N_4896,N_4125,N_4057);
and U4897 (N_4897,N_4086,N_4352);
nand U4898 (N_4898,N_4148,N_4464);
and U4899 (N_4899,N_4159,N_4391);
xor U4900 (N_4900,N_4201,N_4052);
and U4901 (N_4901,N_4097,N_4010);
nor U4902 (N_4902,N_4287,N_4080);
or U4903 (N_4903,N_4124,N_4138);
xor U4904 (N_4904,N_4268,N_4205);
nand U4905 (N_4905,N_4078,N_4210);
nand U4906 (N_4906,N_4104,N_4264);
nand U4907 (N_4907,N_4084,N_4077);
xor U4908 (N_4908,N_4132,N_4207);
nor U4909 (N_4909,N_4466,N_4020);
or U4910 (N_4910,N_4006,N_4284);
and U4911 (N_4911,N_4381,N_4025);
xnor U4912 (N_4912,N_4215,N_4407);
xor U4913 (N_4913,N_4358,N_4229);
or U4914 (N_4914,N_4257,N_4289);
or U4915 (N_4915,N_4095,N_4039);
and U4916 (N_4916,N_4206,N_4097);
and U4917 (N_4917,N_4427,N_4406);
xnor U4918 (N_4918,N_4131,N_4235);
and U4919 (N_4919,N_4381,N_4082);
or U4920 (N_4920,N_4338,N_4441);
nor U4921 (N_4921,N_4220,N_4100);
or U4922 (N_4922,N_4184,N_4445);
nand U4923 (N_4923,N_4226,N_4100);
xor U4924 (N_4924,N_4486,N_4423);
nand U4925 (N_4925,N_4115,N_4114);
nand U4926 (N_4926,N_4417,N_4308);
and U4927 (N_4927,N_4239,N_4260);
nand U4928 (N_4928,N_4497,N_4232);
xor U4929 (N_4929,N_4162,N_4352);
nor U4930 (N_4930,N_4295,N_4389);
nor U4931 (N_4931,N_4035,N_4248);
or U4932 (N_4932,N_4018,N_4038);
or U4933 (N_4933,N_4095,N_4126);
nand U4934 (N_4934,N_4147,N_4121);
and U4935 (N_4935,N_4311,N_4238);
or U4936 (N_4936,N_4490,N_4318);
nor U4937 (N_4937,N_4147,N_4227);
nor U4938 (N_4938,N_4213,N_4284);
nand U4939 (N_4939,N_4296,N_4120);
or U4940 (N_4940,N_4140,N_4304);
nor U4941 (N_4941,N_4396,N_4287);
nand U4942 (N_4942,N_4172,N_4057);
nand U4943 (N_4943,N_4439,N_4421);
xor U4944 (N_4944,N_4289,N_4422);
and U4945 (N_4945,N_4130,N_4478);
and U4946 (N_4946,N_4004,N_4133);
nand U4947 (N_4947,N_4228,N_4297);
nand U4948 (N_4948,N_4185,N_4220);
xnor U4949 (N_4949,N_4020,N_4404);
and U4950 (N_4950,N_4094,N_4256);
nand U4951 (N_4951,N_4497,N_4174);
nor U4952 (N_4952,N_4074,N_4119);
nor U4953 (N_4953,N_4481,N_4403);
xnor U4954 (N_4954,N_4322,N_4130);
or U4955 (N_4955,N_4196,N_4100);
or U4956 (N_4956,N_4271,N_4220);
or U4957 (N_4957,N_4487,N_4012);
or U4958 (N_4958,N_4459,N_4383);
nor U4959 (N_4959,N_4015,N_4290);
nand U4960 (N_4960,N_4449,N_4153);
and U4961 (N_4961,N_4001,N_4049);
nand U4962 (N_4962,N_4183,N_4220);
nand U4963 (N_4963,N_4131,N_4006);
or U4964 (N_4964,N_4217,N_4467);
nand U4965 (N_4965,N_4073,N_4191);
nand U4966 (N_4966,N_4187,N_4149);
nor U4967 (N_4967,N_4086,N_4420);
or U4968 (N_4968,N_4498,N_4253);
nand U4969 (N_4969,N_4462,N_4417);
nor U4970 (N_4970,N_4188,N_4175);
or U4971 (N_4971,N_4189,N_4471);
xnor U4972 (N_4972,N_4125,N_4272);
or U4973 (N_4973,N_4268,N_4117);
nor U4974 (N_4974,N_4490,N_4338);
xnor U4975 (N_4975,N_4324,N_4023);
or U4976 (N_4976,N_4002,N_4325);
xor U4977 (N_4977,N_4329,N_4116);
or U4978 (N_4978,N_4429,N_4362);
or U4979 (N_4979,N_4429,N_4048);
xor U4980 (N_4980,N_4094,N_4302);
and U4981 (N_4981,N_4129,N_4415);
or U4982 (N_4982,N_4472,N_4257);
nor U4983 (N_4983,N_4044,N_4098);
nor U4984 (N_4984,N_4105,N_4397);
xnor U4985 (N_4985,N_4445,N_4261);
xor U4986 (N_4986,N_4097,N_4143);
nor U4987 (N_4987,N_4331,N_4071);
xor U4988 (N_4988,N_4482,N_4267);
nand U4989 (N_4989,N_4285,N_4049);
nor U4990 (N_4990,N_4494,N_4158);
and U4991 (N_4991,N_4206,N_4430);
nand U4992 (N_4992,N_4335,N_4086);
nor U4993 (N_4993,N_4447,N_4008);
or U4994 (N_4994,N_4499,N_4341);
xnor U4995 (N_4995,N_4197,N_4363);
nand U4996 (N_4996,N_4206,N_4117);
or U4997 (N_4997,N_4090,N_4020);
or U4998 (N_4998,N_4424,N_4359);
xnor U4999 (N_4999,N_4117,N_4243);
nand U5000 (N_5000,N_4726,N_4543);
xor U5001 (N_5001,N_4926,N_4928);
or U5002 (N_5002,N_4605,N_4606);
xnor U5003 (N_5003,N_4554,N_4702);
nor U5004 (N_5004,N_4738,N_4569);
and U5005 (N_5005,N_4986,N_4960);
and U5006 (N_5006,N_4627,N_4896);
nand U5007 (N_5007,N_4954,N_4913);
xnor U5008 (N_5008,N_4745,N_4618);
nor U5009 (N_5009,N_4515,N_4837);
nand U5010 (N_5010,N_4899,N_4904);
nor U5011 (N_5011,N_4530,N_4885);
nor U5012 (N_5012,N_4967,N_4567);
xnor U5013 (N_5013,N_4512,N_4843);
nand U5014 (N_5014,N_4563,N_4719);
and U5015 (N_5015,N_4548,N_4908);
nor U5016 (N_5016,N_4560,N_4656);
and U5017 (N_5017,N_4735,N_4792);
and U5018 (N_5018,N_4920,N_4739);
nor U5019 (N_5019,N_4999,N_4815);
or U5020 (N_5020,N_4900,N_4626);
and U5021 (N_5021,N_4944,N_4844);
or U5022 (N_5022,N_4955,N_4595);
or U5023 (N_5023,N_4581,N_4624);
xnor U5024 (N_5024,N_4615,N_4951);
nand U5025 (N_5025,N_4612,N_4639);
nor U5026 (N_5026,N_4832,N_4813);
nor U5027 (N_5027,N_4818,N_4685);
nor U5028 (N_5028,N_4974,N_4614);
xnor U5029 (N_5029,N_4748,N_4891);
or U5030 (N_5030,N_4943,N_4580);
or U5031 (N_5031,N_4524,N_4776);
or U5032 (N_5032,N_4695,N_4816);
nor U5033 (N_5033,N_4947,N_4787);
nand U5034 (N_5034,N_4831,N_4736);
or U5035 (N_5035,N_4852,N_4609);
nand U5036 (N_5036,N_4602,N_4987);
or U5037 (N_5037,N_4935,N_4874);
nand U5038 (N_5038,N_4888,N_4805);
xnor U5039 (N_5039,N_4687,N_4691);
xnor U5040 (N_5040,N_4665,N_4725);
xnor U5041 (N_5041,N_4866,N_4703);
and U5042 (N_5042,N_4948,N_4946);
or U5043 (N_5043,N_4504,N_4829);
and U5044 (N_5044,N_4793,N_4517);
and U5045 (N_5045,N_4522,N_4724);
or U5046 (N_5046,N_4718,N_4962);
nand U5047 (N_5047,N_4868,N_4903);
nor U5048 (N_5048,N_4768,N_4757);
xor U5049 (N_5049,N_4766,N_4763);
and U5050 (N_5050,N_4549,N_4810);
or U5051 (N_5051,N_4635,N_4769);
nor U5052 (N_5052,N_4648,N_4939);
or U5053 (N_5053,N_4911,N_4909);
nand U5054 (N_5054,N_4586,N_4856);
nor U5055 (N_5055,N_4835,N_4647);
nand U5056 (N_5056,N_4644,N_4881);
xor U5057 (N_5057,N_4929,N_4995);
or U5058 (N_5058,N_4544,N_4712);
nand U5059 (N_5059,N_4916,N_4848);
or U5060 (N_5060,N_4621,N_4541);
nor U5061 (N_5061,N_4681,N_4661);
or U5062 (N_5062,N_4864,N_4662);
or U5063 (N_5063,N_4616,N_4906);
and U5064 (N_5064,N_4737,N_4631);
and U5065 (N_5065,N_4603,N_4696);
nor U5066 (N_5066,N_4956,N_4789);
nor U5067 (N_5067,N_4657,N_4600);
or U5068 (N_5068,N_4788,N_4781);
xor U5069 (N_5069,N_4568,N_4806);
nor U5070 (N_5070,N_4550,N_4887);
or U5071 (N_5071,N_4531,N_4985);
xnor U5072 (N_5072,N_4804,N_4773);
and U5073 (N_5073,N_4537,N_4927);
and U5074 (N_5074,N_4976,N_4690);
or U5075 (N_5075,N_4824,N_4750);
and U5076 (N_5076,N_4870,N_4684);
nor U5077 (N_5077,N_4895,N_4667);
xor U5078 (N_5078,N_4535,N_4716);
nor U5079 (N_5079,N_4774,N_4886);
and U5080 (N_5080,N_4525,N_4630);
nor U5081 (N_5081,N_4564,N_4982);
nor U5082 (N_5082,N_4693,N_4758);
and U5083 (N_5083,N_4664,N_4611);
xor U5084 (N_5084,N_4534,N_4589);
nand U5085 (N_5085,N_4968,N_4973);
and U5086 (N_5086,N_4625,N_4936);
or U5087 (N_5087,N_4780,N_4540);
and U5088 (N_5088,N_4526,N_4989);
nor U5089 (N_5089,N_4532,N_4593);
nand U5090 (N_5090,N_4650,N_4889);
nand U5091 (N_5091,N_4752,N_4882);
nand U5092 (N_5092,N_4833,N_4686);
nand U5093 (N_5093,N_4520,N_4849);
or U5094 (N_5094,N_4527,N_4797);
and U5095 (N_5095,N_4777,N_4762);
and U5096 (N_5096,N_4972,N_4673);
or U5097 (N_5097,N_4964,N_4507);
and U5098 (N_5098,N_4508,N_4628);
nand U5099 (N_5099,N_4884,N_4597);
nor U5100 (N_5100,N_4798,N_4596);
nand U5101 (N_5101,N_4692,N_4847);
and U5102 (N_5102,N_4901,N_4915);
or U5103 (N_5103,N_4683,N_4670);
or U5104 (N_5104,N_4853,N_4933);
or U5105 (N_5105,N_4997,N_4717);
or U5106 (N_5106,N_4706,N_4723);
or U5107 (N_5107,N_4655,N_4855);
xnor U5108 (N_5108,N_4809,N_4632);
nand U5109 (N_5109,N_4811,N_4796);
nand U5110 (N_5110,N_4715,N_4820);
nor U5111 (N_5111,N_4511,N_4601);
or U5112 (N_5112,N_4565,N_4858);
or U5113 (N_5113,N_4555,N_4876);
and U5114 (N_5114,N_4937,N_4577);
nand U5115 (N_5115,N_4940,N_4697);
or U5116 (N_5116,N_4764,N_4599);
xor U5117 (N_5117,N_4751,N_4592);
and U5118 (N_5118,N_4642,N_4658);
or U5119 (N_5119,N_4743,N_4679);
xor U5120 (N_5120,N_4710,N_4545);
or U5121 (N_5121,N_4746,N_4689);
and U5122 (N_5122,N_4501,N_4646);
xnor U5123 (N_5123,N_4991,N_4863);
or U5124 (N_5124,N_4506,N_4652);
and U5125 (N_5125,N_4912,N_4910);
xnor U5126 (N_5126,N_4721,N_4790);
and U5127 (N_5127,N_4633,N_4795);
xnor U5128 (N_5128,N_4775,N_4897);
or U5129 (N_5129,N_4699,N_4573);
and U5130 (N_5130,N_4950,N_4975);
xnor U5131 (N_5131,N_4552,N_4572);
xnor U5132 (N_5132,N_4861,N_4701);
and U5133 (N_5133,N_4666,N_4791);
xor U5134 (N_5134,N_4638,N_4669);
xnor U5135 (N_5135,N_4822,N_4519);
nor U5136 (N_5136,N_4807,N_4878);
or U5137 (N_5137,N_4825,N_4588);
and U5138 (N_5138,N_4801,N_4812);
nand U5139 (N_5139,N_4826,N_4629);
or U5140 (N_5140,N_4505,N_4924);
nor U5141 (N_5141,N_4559,N_4959);
nor U5142 (N_5142,N_4918,N_4617);
nand U5143 (N_5143,N_4841,N_4607);
xor U5144 (N_5144,N_4562,N_4518);
nor U5145 (N_5145,N_4539,N_4879);
or U5146 (N_5146,N_4977,N_4732);
nor U5147 (N_5147,N_4556,N_4720);
xor U5148 (N_5148,N_4538,N_4740);
xnor U5149 (N_5149,N_4983,N_4799);
nand U5150 (N_5150,N_4808,N_4575);
xnor U5151 (N_5151,N_4503,N_4965);
and U5152 (N_5152,N_4651,N_4880);
nand U5153 (N_5153,N_4598,N_4574);
nand U5154 (N_5154,N_4707,N_4590);
or U5155 (N_5155,N_4784,N_4523);
nor U5156 (N_5156,N_4640,N_4742);
or U5157 (N_5157,N_4830,N_4902);
nor U5158 (N_5158,N_4753,N_4705);
or U5159 (N_5159,N_4850,N_4620);
nand U5160 (N_5160,N_4747,N_4533);
or U5161 (N_5161,N_4770,N_4838);
nor U5162 (N_5162,N_4694,N_4571);
nor U5163 (N_5163,N_4969,N_4557);
xnor U5164 (N_5164,N_4583,N_4700);
nor U5165 (N_5165,N_4963,N_4988);
nor U5166 (N_5166,N_4898,N_4643);
nor U5167 (N_5167,N_4845,N_4905);
or U5168 (N_5168,N_4942,N_4839);
nor U5169 (N_5169,N_4872,N_4846);
or U5170 (N_5170,N_4698,N_4952);
nor U5171 (N_5171,N_4682,N_4893);
and U5172 (N_5172,N_4677,N_4836);
nand U5173 (N_5173,N_4722,N_4925);
nor U5174 (N_5174,N_4730,N_4553);
or U5175 (N_5175,N_4966,N_4802);
xor U5176 (N_5176,N_4502,N_4949);
or U5177 (N_5177,N_4771,N_4794);
xnor U5178 (N_5178,N_4992,N_4821);
nand U5179 (N_5179,N_4931,N_4984);
or U5180 (N_5180,N_4561,N_4990);
nand U5181 (N_5181,N_4610,N_4783);
or U5182 (N_5182,N_4623,N_4619);
and U5183 (N_5183,N_4923,N_4890);
nor U5184 (N_5184,N_4680,N_4814);
xnor U5185 (N_5185,N_4521,N_4570);
nand U5186 (N_5186,N_4514,N_4529);
xor U5187 (N_5187,N_4819,N_4993);
xor U5188 (N_5188,N_4755,N_4961);
xor U5189 (N_5189,N_4708,N_4981);
xor U5190 (N_5190,N_4765,N_4779);
nand U5191 (N_5191,N_4688,N_4834);
and U5192 (N_5192,N_4772,N_4733);
nor U5193 (N_5193,N_4678,N_4871);
nand U5194 (N_5194,N_4547,N_4786);
and U5195 (N_5195,N_4663,N_4921);
xnor U5196 (N_5196,N_4756,N_4711);
nor U5197 (N_5197,N_4970,N_4536);
xnor U5198 (N_5198,N_4957,N_4576);
xnor U5199 (N_5199,N_4941,N_4613);
or U5200 (N_5200,N_4873,N_4823);
or U5201 (N_5201,N_4637,N_4760);
nor U5202 (N_5202,N_4998,N_4994);
nor U5203 (N_5203,N_4945,N_4587);
nand U5204 (N_5204,N_4729,N_4500);
or U5205 (N_5205,N_4676,N_4907);
nand U5206 (N_5206,N_4542,N_4585);
or U5207 (N_5207,N_4641,N_4857);
nor U5208 (N_5208,N_4660,N_4604);
nand U5209 (N_5209,N_4558,N_4551);
or U5210 (N_5210,N_4649,N_4827);
xor U5211 (N_5211,N_4875,N_4922);
nor U5212 (N_5212,N_4509,N_4767);
nand U5213 (N_5213,N_4914,N_4674);
nor U5214 (N_5214,N_4996,N_4840);
xor U5215 (N_5215,N_4591,N_4727);
and U5216 (N_5216,N_4749,N_4785);
and U5217 (N_5217,N_4579,N_4671);
and U5218 (N_5218,N_4953,N_4582);
nand U5219 (N_5219,N_4851,N_4892);
nor U5220 (N_5220,N_4741,N_4608);
nand U5221 (N_5221,N_4654,N_4653);
nor U5222 (N_5222,N_4584,N_4516);
nor U5223 (N_5223,N_4672,N_4675);
or U5224 (N_5224,N_4894,N_4934);
nand U5225 (N_5225,N_4709,N_4622);
and U5226 (N_5226,N_4594,N_4877);
or U5227 (N_5227,N_4668,N_4842);
nor U5228 (N_5228,N_4744,N_4971);
nand U5229 (N_5229,N_4862,N_4728);
or U5230 (N_5230,N_4714,N_4932);
or U5231 (N_5231,N_4919,N_4782);
or U5232 (N_5232,N_4731,N_4645);
or U5233 (N_5233,N_4803,N_4659);
nand U5234 (N_5234,N_4867,N_4865);
nand U5235 (N_5235,N_4704,N_4734);
nor U5236 (N_5236,N_4854,N_4828);
nand U5237 (N_5237,N_4917,N_4759);
xnor U5238 (N_5238,N_4958,N_4636);
and U5239 (N_5239,N_4528,N_4713);
nor U5240 (N_5240,N_4860,N_4800);
or U5241 (N_5241,N_4859,N_4817);
xor U5242 (N_5242,N_4883,N_4761);
or U5243 (N_5243,N_4546,N_4578);
xor U5244 (N_5244,N_4869,N_4634);
or U5245 (N_5245,N_4566,N_4510);
or U5246 (N_5246,N_4980,N_4938);
and U5247 (N_5247,N_4930,N_4778);
nand U5248 (N_5248,N_4513,N_4754);
nand U5249 (N_5249,N_4978,N_4979);
nand U5250 (N_5250,N_4605,N_4764);
or U5251 (N_5251,N_4667,N_4733);
xnor U5252 (N_5252,N_4800,N_4604);
or U5253 (N_5253,N_4786,N_4828);
nor U5254 (N_5254,N_4774,N_4728);
or U5255 (N_5255,N_4946,N_4790);
or U5256 (N_5256,N_4877,N_4586);
nor U5257 (N_5257,N_4902,N_4511);
nor U5258 (N_5258,N_4787,N_4627);
nor U5259 (N_5259,N_4994,N_4522);
nand U5260 (N_5260,N_4567,N_4814);
or U5261 (N_5261,N_4658,N_4974);
nand U5262 (N_5262,N_4681,N_4654);
xor U5263 (N_5263,N_4963,N_4604);
or U5264 (N_5264,N_4878,N_4864);
and U5265 (N_5265,N_4686,N_4743);
or U5266 (N_5266,N_4972,N_4882);
and U5267 (N_5267,N_4695,N_4503);
and U5268 (N_5268,N_4679,N_4863);
and U5269 (N_5269,N_4750,N_4852);
or U5270 (N_5270,N_4683,N_4509);
nand U5271 (N_5271,N_4593,N_4968);
nand U5272 (N_5272,N_4953,N_4578);
nor U5273 (N_5273,N_4766,N_4832);
or U5274 (N_5274,N_4740,N_4625);
or U5275 (N_5275,N_4687,N_4864);
nor U5276 (N_5276,N_4931,N_4839);
nand U5277 (N_5277,N_4994,N_4883);
and U5278 (N_5278,N_4564,N_4752);
nand U5279 (N_5279,N_4833,N_4900);
nor U5280 (N_5280,N_4814,N_4672);
nor U5281 (N_5281,N_4542,N_4776);
nand U5282 (N_5282,N_4751,N_4890);
nand U5283 (N_5283,N_4532,N_4567);
nand U5284 (N_5284,N_4949,N_4900);
nor U5285 (N_5285,N_4917,N_4692);
and U5286 (N_5286,N_4897,N_4926);
or U5287 (N_5287,N_4822,N_4980);
nor U5288 (N_5288,N_4583,N_4819);
xor U5289 (N_5289,N_4849,N_4968);
nor U5290 (N_5290,N_4945,N_4837);
or U5291 (N_5291,N_4927,N_4727);
nand U5292 (N_5292,N_4549,N_4874);
nor U5293 (N_5293,N_4839,N_4815);
nor U5294 (N_5294,N_4501,N_4727);
or U5295 (N_5295,N_4804,N_4649);
or U5296 (N_5296,N_4873,N_4514);
xor U5297 (N_5297,N_4596,N_4625);
xor U5298 (N_5298,N_4632,N_4966);
and U5299 (N_5299,N_4629,N_4724);
nor U5300 (N_5300,N_4757,N_4618);
nand U5301 (N_5301,N_4661,N_4940);
and U5302 (N_5302,N_4978,N_4573);
xor U5303 (N_5303,N_4675,N_4629);
and U5304 (N_5304,N_4704,N_4813);
nor U5305 (N_5305,N_4518,N_4861);
nor U5306 (N_5306,N_4909,N_4633);
xor U5307 (N_5307,N_4821,N_4605);
nor U5308 (N_5308,N_4931,N_4851);
and U5309 (N_5309,N_4636,N_4501);
nor U5310 (N_5310,N_4556,N_4917);
xor U5311 (N_5311,N_4544,N_4745);
or U5312 (N_5312,N_4940,N_4640);
xor U5313 (N_5313,N_4896,N_4609);
nor U5314 (N_5314,N_4830,N_4640);
or U5315 (N_5315,N_4796,N_4888);
nor U5316 (N_5316,N_4705,N_4544);
nor U5317 (N_5317,N_4847,N_4652);
or U5318 (N_5318,N_4901,N_4514);
xnor U5319 (N_5319,N_4905,N_4856);
nor U5320 (N_5320,N_4704,N_4888);
or U5321 (N_5321,N_4943,N_4773);
or U5322 (N_5322,N_4706,N_4653);
or U5323 (N_5323,N_4963,N_4511);
nand U5324 (N_5324,N_4898,N_4751);
xnor U5325 (N_5325,N_4627,N_4653);
or U5326 (N_5326,N_4945,N_4897);
and U5327 (N_5327,N_4991,N_4575);
and U5328 (N_5328,N_4703,N_4872);
nor U5329 (N_5329,N_4632,N_4833);
nor U5330 (N_5330,N_4909,N_4694);
nor U5331 (N_5331,N_4617,N_4920);
and U5332 (N_5332,N_4702,N_4885);
or U5333 (N_5333,N_4991,N_4815);
nand U5334 (N_5334,N_4877,N_4785);
or U5335 (N_5335,N_4938,N_4772);
nor U5336 (N_5336,N_4745,N_4558);
nand U5337 (N_5337,N_4585,N_4775);
and U5338 (N_5338,N_4867,N_4846);
nor U5339 (N_5339,N_4865,N_4605);
nor U5340 (N_5340,N_4943,N_4643);
and U5341 (N_5341,N_4521,N_4761);
or U5342 (N_5342,N_4941,N_4890);
nor U5343 (N_5343,N_4945,N_4855);
and U5344 (N_5344,N_4647,N_4567);
nor U5345 (N_5345,N_4942,N_4544);
xnor U5346 (N_5346,N_4801,N_4826);
xor U5347 (N_5347,N_4732,N_4800);
nor U5348 (N_5348,N_4581,N_4663);
and U5349 (N_5349,N_4901,N_4587);
xnor U5350 (N_5350,N_4544,N_4554);
or U5351 (N_5351,N_4547,N_4562);
xnor U5352 (N_5352,N_4719,N_4850);
and U5353 (N_5353,N_4660,N_4924);
and U5354 (N_5354,N_4820,N_4657);
or U5355 (N_5355,N_4677,N_4618);
nand U5356 (N_5356,N_4840,N_4734);
nor U5357 (N_5357,N_4987,N_4616);
and U5358 (N_5358,N_4575,N_4663);
nor U5359 (N_5359,N_4860,N_4908);
nand U5360 (N_5360,N_4918,N_4713);
or U5361 (N_5361,N_4744,N_4686);
or U5362 (N_5362,N_4637,N_4791);
or U5363 (N_5363,N_4904,N_4572);
nand U5364 (N_5364,N_4793,N_4802);
and U5365 (N_5365,N_4906,N_4742);
and U5366 (N_5366,N_4938,N_4526);
or U5367 (N_5367,N_4626,N_4776);
and U5368 (N_5368,N_4694,N_4943);
xor U5369 (N_5369,N_4557,N_4831);
nand U5370 (N_5370,N_4974,N_4745);
nor U5371 (N_5371,N_4850,N_4924);
and U5372 (N_5372,N_4867,N_4887);
and U5373 (N_5373,N_4608,N_4985);
nand U5374 (N_5374,N_4846,N_4809);
nand U5375 (N_5375,N_4547,N_4504);
nand U5376 (N_5376,N_4558,N_4597);
or U5377 (N_5377,N_4590,N_4931);
or U5378 (N_5378,N_4662,N_4680);
nand U5379 (N_5379,N_4590,N_4784);
nand U5380 (N_5380,N_4968,N_4615);
or U5381 (N_5381,N_4581,N_4787);
nor U5382 (N_5382,N_4721,N_4714);
or U5383 (N_5383,N_4825,N_4944);
xor U5384 (N_5384,N_4711,N_4712);
or U5385 (N_5385,N_4644,N_4707);
xnor U5386 (N_5386,N_4572,N_4684);
xnor U5387 (N_5387,N_4981,N_4874);
or U5388 (N_5388,N_4502,N_4968);
or U5389 (N_5389,N_4993,N_4970);
or U5390 (N_5390,N_4869,N_4884);
and U5391 (N_5391,N_4926,N_4790);
or U5392 (N_5392,N_4544,N_4742);
nor U5393 (N_5393,N_4751,N_4830);
nor U5394 (N_5394,N_4905,N_4750);
nand U5395 (N_5395,N_4823,N_4736);
nor U5396 (N_5396,N_4542,N_4500);
xnor U5397 (N_5397,N_4750,N_4806);
xnor U5398 (N_5398,N_4652,N_4692);
nor U5399 (N_5399,N_4572,N_4508);
or U5400 (N_5400,N_4828,N_4861);
and U5401 (N_5401,N_4638,N_4651);
and U5402 (N_5402,N_4712,N_4674);
nor U5403 (N_5403,N_4878,N_4677);
xnor U5404 (N_5404,N_4616,N_4800);
xnor U5405 (N_5405,N_4799,N_4521);
or U5406 (N_5406,N_4838,N_4813);
xnor U5407 (N_5407,N_4514,N_4528);
xnor U5408 (N_5408,N_4892,N_4601);
nor U5409 (N_5409,N_4711,N_4629);
nand U5410 (N_5410,N_4840,N_4520);
nor U5411 (N_5411,N_4653,N_4525);
or U5412 (N_5412,N_4599,N_4905);
nor U5413 (N_5413,N_4789,N_4568);
xor U5414 (N_5414,N_4504,N_4725);
nand U5415 (N_5415,N_4692,N_4744);
nor U5416 (N_5416,N_4698,N_4781);
or U5417 (N_5417,N_4580,N_4868);
nor U5418 (N_5418,N_4554,N_4513);
and U5419 (N_5419,N_4835,N_4745);
nand U5420 (N_5420,N_4830,N_4862);
nor U5421 (N_5421,N_4776,N_4772);
or U5422 (N_5422,N_4631,N_4766);
nand U5423 (N_5423,N_4893,N_4834);
nand U5424 (N_5424,N_4746,N_4505);
xnor U5425 (N_5425,N_4651,N_4974);
nor U5426 (N_5426,N_4794,N_4726);
nor U5427 (N_5427,N_4936,N_4559);
nand U5428 (N_5428,N_4836,N_4986);
nand U5429 (N_5429,N_4906,N_4536);
or U5430 (N_5430,N_4594,N_4940);
or U5431 (N_5431,N_4809,N_4902);
nor U5432 (N_5432,N_4838,N_4969);
or U5433 (N_5433,N_4871,N_4510);
nand U5434 (N_5434,N_4740,N_4956);
and U5435 (N_5435,N_4883,N_4673);
nand U5436 (N_5436,N_4902,N_4858);
and U5437 (N_5437,N_4621,N_4669);
nand U5438 (N_5438,N_4956,N_4755);
xnor U5439 (N_5439,N_4653,N_4905);
xnor U5440 (N_5440,N_4778,N_4717);
xnor U5441 (N_5441,N_4980,N_4809);
or U5442 (N_5442,N_4834,N_4745);
nor U5443 (N_5443,N_4594,N_4811);
and U5444 (N_5444,N_4769,N_4848);
nor U5445 (N_5445,N_4634,N_4789);
and U5446 (N_5446,N_4925,N_4503);
or U5447 (N_5447,N_4991,N_4566);
nand U5448 (N_5448,N_4553,N_4887);
or U5449 (N_5449,N_4610,N_4720);
or U5450 (N_5450,N_4620,N_4667);
xnor U5451 (N_5451,N_4670,N_4690);
xnor U5452 (N_5452,N_4727,N_4676);
nand U5453 (N_5453,N_4953,N_4912);
nand U5454 (N_5454,N_4607,N_4518);
xnor U5455 (N_5455,N_4763,N_4574);
xnor U5456 (N_5456,N_4841,N_4589);
and U5457 (N_5457,N_4822,N_4696);
and U5458 (N_5458,N_4802,N_4996);
nor U5459 (N_5459,N_4678,N_4653);
nand U5460 (N_5460,N_4680,N_4735);
or U5461 (N_5461,N_4552,N_4628);
nand U5462 (N_5462,N_4648,N_4581);
nand U5463 (N_5463,N_4918,N_4622);
and U5464 (N_5464,N_4942,N_4581);
nand U5465 (N_5465,N_4691,N_4630);
nor U5466 (N_5466,N_4593,N_4935);
nor U5467 (N_5467,N_4900,N_4609);
nor U5468 (N_5468,N_4835,N_4519);
nor U5469 (N_5469,N_4828,N_4667);
nor U5470 (N_5470,N_4816,N_4654);
or U5471 (N_5471,N_4508,N_4696);
or U5472 (N_5472,N_4581,N_4796);
nand U5473 (N_5473,N_4785,N_4538);
and U5474 (N_5474,N_4979,N_4816);
or U5475 (N_5475,N_4667,N_4953);
and U5476 (N_5476,N_4880,N_4910);
or U5477 (N_5477,N_4944,N_4801);
xor U5478 (N_5478,N_4788,N_4722);
or U5479 (N_5479,N_4778,N_4697);
nor U5480 (N_5480,N_4981,N_4580);
or U5481 (N_5481,N_4555,N_4943);
nor U5482 (N_5482,N_4911,N_4690);
nand U5483 (N_5483,N_4735,N_4798);
nor U5484 (N_5484,N_4694,N_4797);
or U5485 (N_5485,N_4699,N_4672);
nand U5486 (N_5486,N_4717,N_4829);
or U5487 (N_5487,N_4726,N_4520);
nand U5488 (N_5488,N_4577,N_4532);
nor U5489 (N_5489,N_4939,N_4591);
xor U5490 (N_5490,N_4917,N_4621);
nand U5491 (N_5491,N_4931,N_4698);
xnor U5492 (N_5492,N_4881,N_4966);
nand U5493 (N_5493,N_4549,N_4938);
and U5494 (N_5494,N_4618,N_4804);
or U5495 (N_5495,N_4943,N_4711);
nand U5496 (N_5496,N_4976,N_4825);
nand U5497 (N_5497,N_4702,N_4821);
nand U5498 (N_5498,N_4938,N_4757);
xor U5499 (N_5499,N_4566,N_4823);
xor U5500 (N_5500,N_5020,N_5354);
and U5501 (N_5501,N_5279,N_5246);
and U5502 (N_5502,N_5224,N_5332);
xnor U5503 (N_5503,N_5404,N_5449);
and U5504 (N_5504,N_5204,N_5427);
xor U5505 (N_5505,N_5417,N_5406);
nand U5506 (N_5506,N_5353,N_5468);
nor U5507 (N_5507,N_5172,N_5276);
nand U5508 (N_5508,N_5341,N_5208);
or U5509 (N_5509,N_5248,N_5042);
xor U5510 (N_5510,N_5216,N_5037);
xnor U5511 (N_5511,N_5012,N_5373);
or U5512 (N_5512,N_5254,N_5111);
xor U5513 (N_5513,N_5103,N_5402);
nor U5514 (N_5514,N_5307,N_5484);
nand U5515 (N_5515,N_5414,N_5045);
or U5516 (N_5516,N_5145,N_5157);
nand U5517 (N_5517,N_5496,N_5200);
nor U5518 (N_5518,N_5256,N_5375);
xnor U5519 (N_5519,N_5001,N_5244);
nor U5520 (N_5520,N_5053,N_5429);
and U5521 (N_5521,N_5081,N_5228);
nor U5522 (N_5522,N_5051,N_5152);
xnor U5523 (N_5523,N_5359,N_5069);
and U5524 (N_5524,N_5203,N_5362);
and U5525 (N_5525,N_5150,N_5370);
and U5526 (N_5526,N_5030,N_5374);
nand U5527 (N_5527,N_5331,N_5249);
or U5528 (N_5528,N_5304,N_5102);
nand U5529 (N_5529,N_5175,N_5089);
or U5530 (N_5530,N_5445,N_5122);
nor U5531 (N_5531,N_5185,N_5198);
xnor U5532 (N_5532,N_5401,N_5466);
and U5533 (N_5533,N_5367,N_5005);
nor U5534 (N_5534,N_5263,N_5425);
xor U5535 (N_5535,N_5376,N_5132);
or U5536 (N_5536,N_5488,N_5077);
xnor U5537 (N_5537,N_5298,N_5016);
and U5538 (N_5538,N_5292,N_5068);
xnor U5539 (N_5539,N_5194,N_5287);
and U5540 (N_5540,N_5443,N_5312);
and U5541 (N_5541,N_5086,N_5057);
xnor U5542 (N_5542,N_5327,N_5049);
xnor U5543 (N_5543,N_5223,N_5442);
nand U5544 (N_5544,N_5059,N_5105);
nor U5545 (N_5545,N_5014,N_5125);
nor U5546 (N_5546,N_5464,N_5142);
or U5547 (N_5547,N_5120,N_5392);
or U5548 (N_5548,N_5130,N_5044);
nor U5549 (N_5549,N_5078,N_5026);
nand U5550 (N_5550,N_5453,N_5461);
xnor U5551 (N_5551,N_5235,N_5193);
nor U5552 (N_5552,N_5293,N_5237);
or U5553 (N_5553,N_5393,N_5302);
xnor U5554 (N_5554,N_5251,N_5463);
xnor U5555 (N_5555,N_5448,N_5387);
nand U5556 (N_5556,N_5038,N_5064);
and U5557 (N_5557,N_5076,N_5221);
xor U5558 (N_5558,N_5128,N_5270);
nor U5559 (N_5559,N_5188,N_5151);
nor U5560 (N_5560,N_5383,N_5197);
xnor U5561 (N_5561,N_5284,N_5054);
and U5562 (N_5562,N_5211,N_5127);
or U5563 (N_5563,N_5313,N_5169);
and U5564 (N_5564,N_5165,N_5428);
nand U5565 (N_5565,N_5485,N_5305);
nand U5566 (N_5566,N_5478,N_5167);
xnor U5567 (N_5567,N_5195,N_5010);
xnor U5568 (N_5568,N_5029,N_5416);
nor U5569 (N_5569,N_5447,N_5033);
xnor U5570 (N_5570,N_5281,N_5073);
nor U5571 (N_5571,N_5149,N_5368);
nand U5572 (N_5572,N_5098,N_5436);
or U5573 (N_5573,N_5056,N_5477);
and U5574 (N_5574,N_5410,N_5283);
or U5575 (N_5575,N_5498,N_5267);
nor U5576 (N_5576,N_5336,N_5472);
xnor U5577 (N_5577,N_5340,N_5434);
and U5578 (N_5578,N_5280,N_5328);
nor U5579 (N_5579,N_5108,N_5459);
nor U5580 (N_5580,N_5486,N_5024);
nand U5581 (N_5581,N_5239,N_5476);
nand U5582 (N_5582,N_5090,N_5230);
or U5583 (N_5583,N_5201,N_5013);
and U5584 (N_5584,N_5491,N_5225);
xnor U5585 (N_5585,N_5291,N_5273);
nor U5586 (N_5586,N_5371,N_5499);
or U5587 (N_5587,N_5097,N_5344);
nand U5588 (N_5588,N_5389,N_5071);
and U5589 (N_5589,N_5245,N_5063);
nor U5590 (N_5590,N_5300,N_5452);
xnor U5591 (N_5591,N_5382,N_5143);
xnor U5592 (N_5592,N_5092,N_5493);
xor U5593 (N_5593,N_5286,N_5356);
xor U5594 (N_5594,N_5140,N_5243);
and U5595 (N_5595,N_5178,N_5433);
nand U5596 (N_5596,N_5095,N_5317);
xnor U5597 (N_5597,N_5394,N_5288);
and U5598 (N_5598,N_5009,N_5316);
and U5599 (N_5599,N_5358,N_5337);
and U5600 (N_5600,N_5253,N_5289);
and U5601 (N_5601,N_5378,N_5266);
nor U5602 (N_5602,N_5156,N_5413);
xor U5603 (N_5603,N_5310,N_5326);
or U5604 (N_5604,N_5104,N_5171);
or U5605 (N_5605,N_5067,N_5455);
or U5606 (N_5606,N_5096,N_5065);
xor U5607 (N_5607,N_5052,N_5231);
or U5608 (N_5608,N_5047,N_5247);
and U5609 (N_5609,N_5173,N_5349);
nand U5610 (N_5610,N_5347,N_5348);
xnor U5611 (N_5611,N_5023,N_5481);
xor U5612 (N_5612,N_5075,N_5085);
nand U5613 (N_5613,N_5227,N_5421);
or U5614 (N_5614,N_5141,N_5099);
or U5615 (N_5615,N_5207,N_5110);
nor U5616 (N_5616,N_5314,N_5131);
nor U5617 (N_5617,N_5041,N_5192);
and U5618 (N_5618,N_5019,N_5109);
xor U5619 (N_5619,N_5163,N_5384);
or U5620 (N_5620,N_5334,N_5489);
xnor U5621 (N_5621,N_5138,N_5101);
xor U5622 (N_5622,N_5492,N_5240);
and U5623 (N_5623,N_5412,N_5210);
nor U5624 (N_5624,N_5161,N_5351);
nand U5625 (N_5625,N_5366,N_5407);
xnor U5626 (N_5626,N_5028,N_5403);
xnor U5627 (N_5627,N_5206,N_5462);
xor U5628 (N_5628,N_5039,N_5031);
or U5629 (N_5629,N_5218,N_5088);
and U5630 (N_5630,N_5050,N_5058);
nor U5631 (N_5631,N_5220,N_5350);
nand U5632 (N_5632,N_5093,N_5166);
and U5633 (N_5633,N_5055,N_5399);
nand U5634 (N_5634,N_5339,N_5257);
nor U5635 (N_5635,N_5060,N_5277);
nand U5636 (N_5636,N_5315,N_5386);
nand U5637 (N_5637,N_5325,N_5264);
nor U5638 (N_5638,N_5154,N_5074);
nor U5639 (N_5639,N_5318,N_5255);
nand U5640 (N_5640,N_5006,N_5380);
xor U5641 (N_5641,N_5369,N_5061);
and U5642 (N_5642,N_5365,N_5133);
nand U5643 (N_5643,N_5117,N_5397);
and U5644 (N_5644,N_5465,N_5450);
and U5645 (N_5645,N_5377,N_5205);
and U5646 (N_5646,N_5222,N_5182);
or U5647 (N_5647,N_5199,N_5252);
or U5648 (N_5648,N_5311,N_5400);
nor U5649 (N_5649,N_5177,N_5238);
xor U5650 (N_5650,N_5490,N_5144);
nand U5651 (N_5651,N_5112,N_5269);
or U5652 (N_5652,N_5487,N_5431);
and U5653 (N_5653,N_5285,N_5018);
or U5654 (N_5654,N_5209,N_5215);
xor U5655 (N_5655,N_5272,N_5372);
xor U5656 (N_5656,N_5123,N_5242);
nor U5657 (N_5657,N_5419,N_5435);
xor U5658 (N_5658,N_5232,N_5100);
nand U5659 (N_5659,N_5408,N_5438);
nand U5660 (N_5660,N_5441,N_5352);
or U5661 (N_5661,N_5303,N_5008);
nor U5662 (N_5662,N_5148,N_5011);
nor U5663 (N_5663,N_5437,N_5176);
and U5664 (N_5664,N_5473,N_5189);
and U5665 (N_5665,N_5259,N_5034);
and U5666 (N_5666,N_5426,N_5121);
nor U5667 (N_5667,N_5309,N_5274);
and U5668 (N_5668,N_5296,N_5229);
nand U5669 (N_5669,N_5153,N_5226);
nand U5670 (N_5670,N_5391,N_5432);
or U5671 (N_5671,N_5066,N_5282);
nand U5672 (N_5672,N_5470,N_5190);
or U5673 (N_5673,N_5278,N_5233);
and U5674 (N_5674,N_5160,N_5423);
nor U5675 (N_5675,N_5139,N_5381);
xnor U5676 (N_5676,N_5025,N_5361);
xor U5677 (N_5677,N_5196,N_5000);
or U5678 (N_5678,N_5155,N_5213);
nand U5679 (N_5679,N_5258,N_5299);
and U5680 (N_5680,N_5422,N_5364);
xor U5681 (N_5681,N_5043,N_5036);
or U5682 (N_5682,N_5290,N_5457);
xnor U5683 (N_5683,N_5268,N_5191);
nor U5684 (N_5684,N_5342,N_5405);
and U5685 (N_5685,N_5107,N_5079);
and U5686 (N_5686,N_5214,N_5180);
xor U5687 (N_5687,N_5388,N_5396);
and U5688 (N_5688,N_5265,N_5119);
nand U5689 (N_5689,N_5439,N_5308);
nand U5690 (N_5690,N_5135,N_5250);
xor U5691 (N_5691,N_5294,N_5360);
and U5692 (N_5692,N_5343,N_5475);
and U5693 (N_5693,N_5083,N_5480);
nor U5694 (N_5694,N_5219,N_5482);
nor U5695 (N_5695,N_5418,N_5094);
or U5696 (N_5696,N_5116,N_5497);
nor U5697 (N_5697,N_5454,N_5168);
nand U5698 (N_5698,N_5324,N_5467);
nand U5699 (N_5699,N_5474,N_5430);
xnor U5700 (N_5700,N_5321,N_5113);
nor U5701 (N_5701,N_5335,N_5424);
or U5702 (N_5702,N_5297,N_5106);
xnor U5703 (N_5703,N_5084,N_5333);
or U5704 (N_5704,N_5420,N_5015);
nor U5705 (N_5705,N_5091,N_5479);
nand U5706 (N_5706,N_5046,N_5134);
nor U5707 (N_5707,N_5080,N_5346);
or U5708 (N_5708,N_5295,N_5234);
nor U5709 (N_5709,N_5027,N_5184);
or U5710 (N_5710,N_5072,N_5183);
and U5711 (N_5711,N_5040,N_5174);
nor U5712 (N_5712,N_5469,N_5395);
or U5713 (N_5713,N_5241,N_5032);
or U5714 (N_5714,N_5494,N_5379);
xnor U5715 (N_5715,N_5021,N_5390);
xor U5716 (N_5716,N_5070,N_5262);
or U5717 (N_5717,N_5217,N_5017);
xnor U5718 (N_5718,N_5003,N_5271);
nand U5719 (N_5719,N_5471,N_5236);
or U5720 (N_5720,N_5202,N_5458);
nand U5721 (N_5721,N_5147,N_5126);
and U5722 (N_5722,N_5385,N_5301);
nand U5723 (N_5723,N_5320,N_5212);
nor U5724 (N_5724,N_5129,N_5415);
xor U5725 (N_5725,N_5446,N_5146);
nand U5726 (N_5726,N_5260,N_5082);
and U5727 (N_5727,N_5170,N_5363);
and U5728 (N_5728,N_5409,N_5087);
nand U5729 (N_5729,N_5355,N_5398);
nand U5730 (N_5730,N_5062,N_5329);
xor U5731 (N_5731,N_5164,N_5158);
nor U5732 (N_5732,N_5114,N_5179);
nor U5733 (N_5733,N_5181,N_5261);
nor U5734 (N_5734,N_5456,N_5004);
nor U5735 (N_5735,N_5451,N_5136);
nand U5736 (N_5736,N_5323,N_5444);
and U5737 (N_5737,N_5035,N_5159);
and U5738 (N_5738,N_5007,N_5460);
and U5739 (N_5739,N_5022,N_5357);
nand U5740 (N_5740,N_5338,N_5275);
and U5741 (N_5741,N_5162,N_5319);
or U5742 (N_5742,N_5137,N_5048);
nor U5743 (N_5743,N_5187,N_5115);
nor U5744 (N_5744,N_5306,N_5330);
nand U5745 (N_5745,N_5411,N_5345);
nand U5746 (N_5746,N_5322,N_5483);
or U5747 (N_5747,N_5002,N_5495);
nor U5748 (N_5748,N_5440,N_5186);
nand U5749 (N_5749,N_5118,N_5124);
xor U5750 (N_5750,N_5151,N_5471);
or U5751 (N_5751,N_5310,N_5435);
and U5752 (N_5752,N_5274,N_5245);
or U5753 (N_5753,N_5268,N_5411);
or U5754 (N_5754,N_5332,N_5416);
nor U5755 (N_5755,N_5470,N_5348);
and U5756 (N_5756,N_5386,N_5391);
nor U5757 (N_5757,N_5293,N_5158);
xor U5758 (N_5758,N_5378,N_5405);
or U5759 (N_5759,N_5148,N_5203);
nand U5760 (N_5760,N_5433,N_5417);
or U5761 (N_5761,N_5009,N_5460);
and U5762 (N_5762,N_5284,N_5012);
or U5763 (N_5763,N_5316,N_5247);
nand U5764 (N_5764,N_5069,N_5267);
or U5765 (N_5765,N_5140,N_5401);
xnor U5766 (N_5766,N_5414,N_5116);
nand U5767 (N_5767,N_5213,N_5217);
xnor U5768 (N_5768,N_5450,N_5229);
and U5769 (N_5769,N_5456,N_5365);
nor U5770 (N_5770,N_5056,N_5064);
nand U5771 (N_5771,N_5102,N_5457);
nor U5772 (N_5772,N_5155,N_5255);
xor U5773 (N_5773,N_5191,N_5329);
or U5774 (N_5774,N_5369,N_5088);
nand U5775 (N_5775,N_5306,N_5293);
and U5776 (N_5776,N_5460,N_5276);
or U5777 (N_5777,N_5187,N_5335);
nand U5778 (N_5778,N_5111,N_5333);
xor U5779 (N_5779,N_5455,N_5092);
xnor U5780 (N_5780,N_5020,N_5097);
xor U5781 (N_5781,N_5358,N_5059);
and U5782 (N_5782,N_5272,N_5497);
nor U5783 (N_5783,N_5049,N_5336);
xnor U5784 (N_5784,N_5231,N_5036);
nand U5785 (N_5785,N_5406,N_5011);
nand U5786 (N_5786,N_5103,N_5193);
and U5787 (N_5787,N_5494,N_5414);
xor U5788 (N_5788,N_5405,N_5096);
or U5789 (N_5789,N_5388,N_5245);
nand U5790 (N_5790,N_5133,N_5171);
and U5791 (N_5791,N_5399,N_5382);
xnor U5792 (N_5792,N_5374,N_5316);
nand U5793 (N_5793,N_5370,N_5423);
nor U5794 (N_5794,N_5372,N_5008);
nand U5795 (N_5795,N_5075,N_5408);
and U5796 (N_5796,N_5486,N_5104);
xor U5797 (N_5797,N_5479,N_5337);
nor U5798 (N_5798,N_5293,N_5431);
and U5799 (N_5799,N_5046,N_5255);
nand U5800 (N_5800,N_5027,N_5395);
or U5801 (N_5801,N_5288,N_5319);
or U5802 (N_5802,N_5307,N_5159);
xor U5803 (N_5803,N_5167,N_5371);
nor U5804 (N_5804,N_5068,N_5057);
xor U5805 (N_5805,N_5294,N_5017);
and U5806 (N_5806,N_5232,N_5472);
xnor U5807 (N_5807,N_5229,N_5081);
and U5808 (N_5808,N_5208,N_5497);
nor U5809 (N_5809,N_5304,N_5248);
and U5810 (N_5810,N_5319,N_5292);
nor U5811 (N_5811,N_5307,N_5275);
nor U5812 (N_5812,N_5292,N_5300);
xor U5813 (N_5813,N_5190,N_5443);
and U5814 (N_5814,N_5024,N_5367);
xnor U5815 (N_5815,N_5472,N_5481);
nor U5816 (N_5816,N_5201,N_5322);
and U5817 (N_5817,N_5488,N_5368);
nor U5818 (N_5818,N_5076,N_5494);
nand U5819 (N_5819,N_5392,N_5366);
nand U5820 (N_5820,N_5020,N_5060);
nor U5821 (N_5821,N_5286,N_5317);
nor U5822 (N_5822,N_5365,N_5254);
nand U5823 (N_5823,N_5232,N_5044);
nand U5824 (N_5824,N_5286,N_5329);
nand U5825 (N_5825,N_5133,N_5270);
or U5826 (N_5826,N_5003,N_5399);
and U5827 (N_5827,N_5157,N_5124);
xor U5828 (N_5828,N_5030,N_5063);
xnor U5829 (N_5829,N_5087,N_5210);
xnor U5830 (N_5830,N_5058,N_5211);
nand U5831 (N_5831,N_5267,N_5468);
nor U5832 (N_5832,N_5085,N_5168);
xnor U5833 (N_5833,N_5177,N_5396);
nor U5834 (N_5834,N_5215,N_5053);
or U5835 (N_5835,N_5389,N_5404);
nor U5836 (N_5836,N_5499,N_5107);
nand U5837 (N_5837,N_5261,N_5462);
or U5838 (N_5838,N_5290,N_5020);
xnor U5839 (N_5839,N_5203,N_5044);
nor U5840 (N_5840,N_5350,N_5486);
and U5841 (N_5841,N_5017,N_5207);
nand U5842 (N_5842,N_5011,N_5215);
xor U5843 (N_5843,N_5245,N_5292);
nand U5844 (N_5844,N_5167,N_5398);
nand U5845 (N_5845,N_5120,N_5016);
nand U5846 (N_5846,N_5395,N_5281);
and U5847 (N_5847,N_5003,N_5010);
nand U5848 (N_5848,N_5391,N_5049);
xor U5849 (N_5849,N_5128,N_5053);
xor U5850 (N_5850,N_5288,N_5028);
or U5851 (N_5851,N_5364,N_5470);
or U5852 (N_5852,N_5310,N_5062);
and U5853 (N_5853,N_5133,N_5375);
or U5854 (N_5854,N_5154,N_5474);
or U5855 (N_5855,N_5118,N_5096);
nand U5856 (N_5856,N_5496,N_5151);
or U5857 (N_5857,N_5454,N_5055);
and U5858 (N_5858,N_5099,N_5352);
nor U5859 (N_5859,N_5012,N_5347);
or U5860 (N_5860,N_5279,N_5413);
xor U5861 (N_5861,N_5308,N_5133);
xnor U5862 (N_5862,N_5116,N_5094);
or U5863 (N_5863,N_5070,N_5424);
nor U5864 (N_5864,N_5372,N_5134);
xor U5865 (N_5865,N_5202,N_5194);
xnor U5866 (N_5866,N_5184,N_5234);
nand U5867 (N_5867,N_5258,N_5073);
xnor U5868 (N_5868,N_5240,N_5170);
xnor U5869 (N_5869,N_5286,N_5299);
xor U5870 (N_5870,N_5485,N_5340);
nand U5871 (N_5871,N_5156,N_5214);
nand U5872 (N_5872,N_5345,N_5058);
or U5873 (N_5873,N_5077,N_5268);
nor U5874 (N_5874,N_5063,N_5213);
and U5875 (N_5875,N_5045,N_5164);
or U5876 (N_5876,N_5134,N_5287);
nor U5877 (N_5877,N_5165,N_5325);
xor U5878 (N_5878,N_5419,N_5248);
xnor U5879 (N_5879,N_5006,N_5157);
and U5880 (N_5880,N_5336,N_5452);
xor U5881 (N_5881,N_5305,N_5391);
or U5882 (N_5882,N_5101,N_5040);
nor U5883 (N_5883,N_5084,N_5315);
nor U5884 (N_5884,N_5000,N_5359);
or U5885 (N_5885,N_5209,N_5368);
nor U5886 (N_5886,N_5171,N_5298);
nor U5887 (N_5887,N_5054,N_5420);
xnor U5888 (N_5888,N_5075,N_5368);
nand U5889 (N_5889,N_5363,N_5455);
xnor U5890 (N_5890,N_5164,N_5006);
nand U5891 (N_5891,N_5193,N_5434);
nand U5892 (N_5892,N_5095,N_5464);
nor U5893 (N_5893,N_5098,N_5003);
and U5894 (N_5894,N_5414,N_5246);
and U5895 (N_5895,N_5160,N_5112);
nor U5896 (N_5896,N_5486,N_5105);
xnor U5897 (N_5897,N_5011,N_5290);
xnor U5898 (N_5898,N_5182,N_5001);
or U5899 (N_5899,N_5147,N_5164);
or U5900 (N_5900,N_5433,N_5096);
and U5901 (N_5901,N_5355,N_5111);
and U5902 (N_5902,N_5133,N_5231);
or U5903 (N_5903,N_5274,N_5329);
and U5904 (N_5904,N_5305,N_5474);
and U5905 (N_5905,N_5319,N_5336);
xnor U5906 (N_5906,N_5263,N_5321);
nor U5907 (N_5907,N_5397,N_5341);
nand U5908 (N_5908,N_5428,N_5242);
nor U5909 (N_5909,N_5376,N_5413);
or U5910 (N_5910,N_5247,N_5222);
or U5911 (N_5911,N_5465,N_5148);
xnor U5912 (N_5912,N_5388,N_5057);
or U5913 (N_5913,N_5057,N_5450);
and U5914 (N_5914,N_5116,N_5113);
or U5915 (N_5915,N_5094,N_5306);
nand U5916 (N_5916,N_5117,N_5097);
nand U5917 (N_5917,N_5102,N_5169);
xnor U5918 (N_5918,N_5191,N_5174);
or U5919 (N_5919,N_5327,N_5332);
xnor U5920 (N_5920,N_5425,N_5099);
nor U5921 (N_5921,N_5073,N_5322);
xnor U5922 (N_5922,N_5021,N_5068);
nand U5923 (N_5923,N_5260,N_5369);
and U5924 (N_5924,N_5381,N_5311);
or U5925 (N_5925,N_5489,N_5041);
and U5926 (N_5926,N_5192,N_5493);
xnor U5927 (N_5927,N_5300,N_5230);
xor U5928 (N_5928,N_5138,N_5273);
nand U5929 (N_5929,N_5230,N_5101);
xnor U5930 (N_5930,N_5494,N_5079);
xnor U5931 (N_5931,N_5432,N_5253);
and U5932 (N_5932,N_5229,N_5059);
and U5933 (N_5933,N_5044,N_5477);
and U5934 (N_5934,N_5347,N_5300);
or U5935 (N_5935,N_5370,N_5205);
xnor U5936 (N_5936,N_5344,N_5459);
or U5937 (N_5937,N_5234,N_5480);
and U5938 (N_5938,N_5335,N_5239);
xnor U5939 (N_5939,N_5267,N_5030);
and U5940 (N_5940,N_5338,N_5250);
xnor U5941 (N_5941,N_5012,N_5358);
nand U5942 (N_5942,N_5346,N_5102);
and U5943 (N_5943,N_5437,N_5444);
xor U5944 (N_5944,N_5455,N_5274);
xor U5945 (N_5945,N_5409,N_5399);
and U5946 (N_5946,N_5169,N_5396);
xor U5947 (N_5947,N_5320,N_5083);
or U5948 (N_5948,N_5059,N_5252);
nor U5949 (N_5949,N_5153,N_5450);
nor U5950 (N_5950,N_5374,N_5090);
nor U5951 (N_5951,N_5300,N_5350);
xnor U5952 (N_5952,N_5444,N_5337);
nor U5953 (N_5953,N_5267,N_5179);
xnor U5954 (N_5954,N_5241,N_5329);
nand U5955 (N_5955,N_5393,N_5077);
and U5956 (N_5956,N_5034,N_5175);
nand U5957 (N_5957,N_5238,N_5473);
or U5958 (N_5958,N_5437,N_5355);
and U5959 (N_5959,N_5393,N_5120);
nor U5960 (N_5960,N_5366,N_5286);
nand U5961 (N_5961,N_5011,N_5138);
xor U5962 (N_5962,N_5433,N_5354);
nor U5963 (N_5963,N_5037,N_5117);
nor U5964 (N_5964,N_5151,N_5403);
nand U5965 (N_5965,N_5188,N_5404);
nand U5966 (N_5966,N_5169,N_5348);
or U5967 (N_5967,N_5150,N_5340);
nor U5968 (N_5968,N_5099,N_5008);
nand U5969 (N_5969,N_5235,N_5197);
nand U5970 (N_5970,N_5091,N_5418);
and U5971 (N_5971,N_5404,N_5106);
nand U5972 (N_5972,N_5021,N_5498);
or U5973 (N_5973,N_5438,N_5442);
nand U5974 (N_5974,N_5371,N_5498);
nor U5975 (N_5975,N_5077,N_5339);
nand U5976 (N_5976,N_5074,N_5092);
xor U5977 (N_5977,N_5098,N_5063);
nand U5978 (N_5978,N_5077,N_5359);
nor U5979 (N_5979,N_5004,N_5479);
nand U5980 (N_5980,N_5074,N_5098);
and U5981 (N_5981,N_5460,N_5112);
and U5982 (N_5982,N_5212,N_5474);
or U5983 (N_5983,N_5421,N_5363);
or U5984 (N_5984,N_5419,N_5341);
or U5985 (N_5985,N_5042,N_5221);
or U5986 (N_5986,N_5399,N_5087);
nor U5987 (N_5987,N_5131,N_5097);
nor U5988 (N_5988,N_5019,N_5127);
nor U5989 (N_5989,N_5340,N_5209);
and U5990 (N_5990,N_5353,N_5237);
nor U5991 (N_5991,N_5310,N_5123);
nor U5992 (N_5992,N_5260,N_5077);
xor U5993 (N_5993,N_5349,N_5365);
nor U5994 (N_5994,N_5495,N_5276);
or U5995 (N_5995,N_5202,N_5378);
and U5996 (N_5996,N_5223,N_5113);
and U5997 (N_5997,N_5113,N_5032);
xnor U5998 (N_5998,N_5395,N_5476);
nor U5999 (N_5999,N_5357,N_5423);
xnor U6000 (N_6000,N_5652,N_5942);
or U6001 (N_6001,N_5563,N_5705);
or U6002 (N_6002,N_5729,N_5676);
or U6003 (N_6003,N_5742,N_5649);
nor U6004 (N_6004,N_5502,N_5683);
xnor U6005 (N_6005,N_5606,N_5733);
nand U6006 (N_6006,N_5569,N_5710);
xor U6007 (N_6007,N_5909,N_5979);
nand U6008 (N_6008,N_5949,N_5976);
nor U6009 (N_6009,N_5980,N_5720);
nand U6010 (N_6010,N_5646,N_5541);
and U6011 (N_6011,N_5526,N_5878);
nand U6012 (N_6012,N_5828,N_5843);
xnor U6013 (N_6013,N_5616,N_5854);
or U6014 (N_6014,N_5817,N_5774);
or U6015 (N_6015,N_5768,N_5553);
or U6016 (N_6016,N_5713,N_5583);
nand U6017 (N_6017,N_5752,N_5784);
xnor U6018 (N_6018,N_5598,N_5535);
and U6019 (N_6019,N_5723,N_5709);
xnor U6020 (N_6020,N_5617,N_5607);
or U6021 (N_6021,N_5513,N_5807);
nand U6022 (N_6022,N_5995,N_5822);
xnor U6023 (N_6023,N_5687,N_5637);
nand U6024 (N_6024,N_5902,N_5509);
xnor U6025 (N_6025,N_5724,N_5525);
or U6026 (N_6026,N_5930,N_5975);
nor U6027 (N_6027,N_5899,N_5560);
xnor U6028 (N_6028,N_5985,N_5500);
nor U6029 (N_6029,N_5516,N_5791);
nor U6030 (N_6030,N_5593,N_5741);
nand U6031 (N_6031,N_5696,N_5780);
or U6032 (N_6032,N_5934,N_5613);
nand U6033 (N_6033,N_5600,N_5536);
nand U6034 (N_6034,N_5678,N_5658);
or U6035 (N_6035,N_5642,N_5756);
xor U6036 (N_6036,N_5993,N_5505);
xnor U6037 (N_6037,N_5913,N_5944);
and U6038 (N_6038,N_5706,N_5643);
or U6039 (N_6039,N_5892,N_5751);
nor U6040 (N_6040,N_5954,N_5916);
or U6041 (N_6041,N_5827,N_5632);
nor U6042 (N_6042,N_5641,N_5575);
nor U6043 (N_6043,N_5636,N_5801);
nand U6044 (N_6044,N_5818,N_5937);
nor U6045 (N_6045,N_5862,N_5737);
and U6046 (N_6046,N_5883,N_5895);
and U6047 (N_6047,N_5855,N_5701);
nand U6048 (N_6048,N_5625,N_5731);
and U6049 (N_6049,N_5668,N_5840);
and U6050 (N_6050,N_5674,N_5953);
or U6051 (N_6051,N_5823,N_5591);
nand U6052 (N_6052,N_5925,N_5747);
xor U6053 (N_6053,N_5688,N_5689);
nand U6054 (N_6054,N_5787,N_5802);
nand U6055 (N_6055,N_5749,N_5659);
nand U6056 (N_6056,N_5868,N_5578);
nand U6057 (N_6057,N_5721,N_5825);
or U6058 (N_6058,N_5999,N_5962);
or U6059 (N_6059,N_5820,N_5846);
or U6060 (N_6060,N_5859,N_5558);
and U6061 (N_6061,N_5537,N_5857);
nor U6062 (N_6062,N_5933,N_5991);
and U6063 (N_6063,N_5656,N_5750);
or U6064 (N_6064,N_5924,N_5861);
nor U6065 (N_6065,N_5630,N_5703);
nand U6066 (N_6066,N_5865,N_5882);
nand U6067 (N_6067,N_5719,N_5639);
or U6068 (N_6068,N_5549,N_5766);
nor U6069 (N_6069,N_5757,N_5586);
nor U6070 (N_6070,N_5519,N_5534);
and U6071 (N_6071,N_5609,N_5681);
and U6072 (N_6072,N_5811,N_5988);
and U6073 (N_6073,N_5947,N_5810);
nor U6074 (N_6074,N_5596,N_5662);
nand U6075 (N_6075,N_5556,N_5550);
xor U6076 (N_6076,N_5833,N_5884);
nor U6077 (N_6077,N_5615,N_5512);
or U6078 (N_6078,N_5808,N_5671);
and U6079 (N_6079,N_5777,N_5679);
nand U6080 (N_6080,N_5832,N_5798);
and U6081 (N_6081,N_5864,N_5592);
and U6082 (N_6082,N_5917,N_5961);
and U6083 (N_6083,N_5929,N_5858);
and U6084 (N_6084,N_5955,N_5870);
nand U6085 (N_6085,N_5959,N_5809);
and U6086 (N_6086,N_5894,N_5910);
nand U6087 (N_6087,N_5521,N_5973);
nor U6088 (N_6088,N_5812,N_5540);
xor U6089 (N_6089,N_5951,N_5715);
or U6090 (N_6090,N_5634,N_5548);
nor U6091 (N_6091,N_5996,N_5893);
and U6092 (N_6092,N_5717,N_5767);
xor U6093 (N_6093,N_5994,N_5921);
and U6094 (N_6094,N_5901,N_5595);
nand U6095 (N_6095,N_5624,N_5772);
or U6096 (N_6096,N_5667,N_5764);
xnor U6097 (N_6097,N_5898,N_5511);
xor U6098 (N_6098,N_5566,N_5940);
xor U6099 (N_6099,N_5602,N_5522);
or U6100 (N_6100,N_5957,N_5520);
or U6101 (N_6101,N_5806,N_5557);
nand U6102 (N_6102,N_5906,N_5538);
xor U6103 (N_6103,N_5568,N_5844);
xor U6104 (N_6104,N_5783,N_5704);
or U6105 (N_6105,N_5555,N_5869);
or U6106 (N_6106,N_5735,N_5960);
and U6107 (N_6107,N_5956,N_5824);
and U6108 (N_6108,N_5876,N_5506);
and U6109 (N_6109,N_5978,N_5740);
or U6110 (N_6110,N_5997,N_5576);
nor U6111 (N_6111,N_5628,N_5981);
and U6112 (N_6112,N_5837,N_5611);
nand U6113 (N_6113,N_5562,N_5968);
nand U6114 (N_6114,N_5765,N_5793);
xor U6115 (N_6115,N_5559,N_5594);
or U6116 (N_6116,N_5702,N_5773);
nand U6117 (N_6117,N_5836,N_5590);
nand U6118 (N_6118,N_5804,N_5686);
nand U6119 (N_6119,N_5785,N_5904);
nor U6120 (N_6120,N_5838,N_5919);
nor U6121 (N_6121,N_5580,N_5945);
xor U6122 (N_6122,N_5935,N_5946);
and U6123 (N_6123,N_5850,N_5657);
nor U6124 (N_6124,N_5631,N_5873);
xnor U6125 (N_6125,N_5771,N_5915);
and U6126 (N_6126,N_5984,N_5732);
or U6127 (N_6127,N_5603,N_5529);
or U6128 (N_6128,N_5507,N_5531);
xnor U6129 (N_6129,N_5950,N_5938);
xor U6130 (N_6130,N_5788,N_5515);
nor U6131 (N_6131,N_5612,N_5958);
nor U6132 (N_6132,N_5665,N_5573);
xnor U6133 (N_6133,N_5524,N_5527);
and U6134 (N_6134,N_5770,N_5700);
and U6135 (N_6135,N_5663,N_5936);
and U6136 (N_6136,N_5734,N_5746);
or U6137 (N_6137,N_5977,N_5675);
and U6138 (N_6138,N_5651,N_5829);
nor U6139 (N_6139,N_5601,N_5831);
and U6140 (N_6140,N_5670,N_5543);
xnor U6141 (N_6141,N_5508,N_5722);
and U6142 (N_6142,N_5622,N_5896);
nand U6143 (N_6143,N_5875,N_5782);
nand U6144 (N_6144,N_5648,N_5790);
or U6145 (N_6145,N_5677,N_5760);
or U6146 (N_6146,N_5655,N_5755);
or U6147 (N_6147,N_5989,N_5673);
xnor U6148 (N_6148,N_5805,N_5860);
xnor U6149 (N_6149,N_5588,N_5619);
xor U6150 (N_6150,N_5797,N_5718);
and U6151 (N_6151,N_5633,N_5969);
xnor U6152 (N_6152,N_5903,N_5841);
or U6153 (N_6153,N_5927,N_5748);
or U6154 (N_6154,N_5638,N_5738);
nand U6155 (N_6155,N_5964,N_5571);
nand U6156 (N_6156,N_5523,N_5629);
nand U6157 (N_6157,N_5852,N_5775);
xnor U6158 (N_6158,N_5759,N_5839);
and U6159 (N_6159,N_5800,N_5669);
nor U6160 (N_6160,N_5743,N_5672);
nand U6161 (N_6161,N_5694,N_5565);
nand U6162 (N_6162,N_5716,N_5789);
nor U6163 (N_6163,N_5654,N_5684);
nand U6164 (N_6164,N_5943,N_5849);
nor U6165 (N_6165,N_5786,N_5714);
or U6166 (N_6166,N_5708,N_5781);
nor U6167 (N_6167,N_5621,N_5585);
and U6168 (N_6168,N_5547,N_5567);
nand U6169 (N_6169,N_5856,N_5604);
nand U6170 (N_6170,N_5941,N_5645);
or U6171 (N_6171,N_5650,N_5712);
nand U6172 (N_6172,N_5685,N_5666);
nand U6173 (N_6173,N_5584,N_5851);
xor U6174 (N_6174,N_5965,N_5880);
nor U6175 (N_6175,N_5589,N_5819);
nor U6176 (N_6176,N_5900,N_5680);
or U6177 (N_6177,N_5874,N_5504);
nor U6178 (N_6178,N_5660,N_5835);
nand U6179 (N_6179,N_5739,N_5644);
or U6180 (N_6180,N_5830,N_5517);
and U6181 (N_6181,N_5697,N_5577);
or U6182 (N_6182,N_5891,N_5983);
and U6183 (N_6183,N_5779,N_5699);
nand U6184 (N_6184,N_5728,N_5727);
nor U6185 (N_6185,N_5664,N_5542);
nor U6186 (N_6186,N_5982,N_5647);
or U6187 (N_6187,N_5871,N_5769);
nor U6188 (N_6188,N_5610,N_5761);
nand U6189 (N_6189,N_5626,N_5814);
and U6190 (N_6190,N_5758,N_5745);
or U6191 (N_6191,N_5926,N_5762);
nor U6192 (N_6192,N_5753,N_5635);
or U6193 (N_6193,N_5998,N_5581);
nand U6194 (N_6194,N_5693,N_5816);
or U6195 (N_6195,N_5539,N_5778);
nand U6196 (N_6196,N_5897,N_5948);
xor U6197 (N_6197,N_5692,N_5552);
xor U6198 (N_6198,N_5587,N_5914);
or U6199 (N_6199,N_5848,N_5911);
or U6200 (N_6200,N_5928,N_5514);
and U6201 (N_6201,N_5974,N_5564);
or U6202 (N_6202,N_5501,N_5614);
xor U6203 (N_6203,N_5623,N_5923);
xnor U6204 (N_6204,N_5905,N_5796);
nand U6205 (N_6205,N_5726,N_5510);
and U6206 (N_6206,N_5795,N_5561);
nand U6207 (N_6207,N_5826,N_5618);
nand U6208 (N_6208,N_5695,N_5972);
nand U6209 (N_6209,N_5908,N_5690);
xnor U6210 (N_6210,N_5792,N_5885);
nand U6211 (N_6211,N_5834,N_5992);
nand U6212 (N_6212,N_5582,N_5599);
and U6213 (N_6213,N_5863,N_5744);
and U6214 (N_6214,N_5821,N_5640);
nor U6215 (N_6215,N_5952,N_5877);
nor U6216 (N_6216,N_5620,N_5920);
or U6217 (N_6217,N_5932,N_5970);
xnor U6218 (N_6218,N_5963,N_5503);
nor U6219 (N_6219,N_5986,N_5881);
or U6220 (N_6220,N_5888,N_5866);
nand U6221 (N_6221,N_5987,N_5627);
and U6222 (N_6222,N_5853,N_5546);
or U6223 (N_6223,N_5966,N_5551);
nand U6224 (N_6224,N_5813,N_5912);
and U6225 (N_6225,N_5661,N_5554);
xnor U6226 (N_6226,N_5653,N_5872);
xnor U6227 (N_6227,N_5608,N_5545);
nor U6228 (N_6228,N_5528,N_5530);
xnor U6229 (N_6229,N_5815,N_5711);
nand U6230 (N_6230,N_5544,N_5572);
nand U6231 (N_6231,N_5939,N_5967);
and U6232 (N_6232,N_5605,N_5725);
or U6233 (N_6233,N_5707,N_5886);
nor U6234 (N_6234,N_5918,N_5570);
nor U6235 (N_6235,N_5794,N_5730);
or U6236 (N_6236,N_5776,N_5682);
nand U6237 (N_6237,N_5518,N_5907);
xnor U6238 (N_6238,N_5754,N_5691);
or U6239 (N_6239,N_5579,N_5867);
xor U6240 (N_6240,N_5931,N_5845);
nor U6241 (N_6241,N_5890,N_5842);
nand U6242 (N_6242,N_5847,N_5889);
nand U6243 (N_6243,N_5597,N_5971);
xor U6244 (N_6244,N_5532,N_5879);
xnor U6245 (N_6245,N_5698,N_5922);
xnor U6246 (N_6246,N_5799,N_5574);
nand U6247 (N_6247,N_5990,N_5533);
xnor U6248 (N_6248,N_5803,N_5736);
and U6249 (N_6249,N_5887,N_5763);
xnor U6250 (N_6250,N_5662,N_5791);
or U6251 (N_6251,N_5763,N_5965);
and U6252 (N_6252,N_5693,N_5776);
nand U6253 (N_6253,N_5663,N_5779);
or U6254 (N_6254,N_5515,N_5523);
nor U6255 (N_6255,N_5821,N_5932);
nor U6256 (N_6256,N_5744,N_5947);
nor U6257 (N_6257,N_5824,N_5974);
and U6258 (N_6258,N_5894,N_5985);
nor U6259 (N_6259,N_5870,N_5579);
or U6260 (N_6260,N_5942,N_5937);
or U6261 (N_6261,N_5723,N_5513);
nand U6262 (N_6262,N_5988,N_5985);
nand U6263 (N_6263,N_5861,N_5942);
and U6264 (N_6264,N_5848,N_5882);
nand U6265 (N_6265,N_5998,N_5788);
xor U6266 (N_6266,N_5954,N_5589);
or U6267 (N_6267,N_5935,N_5723);
and U6268 (N_6268,N_5576,N_5934);
or U6269 (N_6269,N_5627,N_5559);
xor U6270 (N_6270,N_5954,N_5833);
nand U6271 (N_6271,N_5974,N_5749);
nand U6272 (N_6272,N_5667,N_5720);
xor U6273 (N_6273,N_5653,N_5935);
or U6274 (N_6274,N_5569,N_5864);
or U6275 (N_6275,N_5553,N_5862);
xor U6276 (N_6276,N_5610,N_5580);
nor U6277 (N_6277,N_5799,N_5927);
or U6278 (N_6278,N_5871,N_5898);
nand U6279 (N_6279,N_5678,N_5621);
nand U6280 (N_6280,N_5857,N_5761);
nor U6281 (N_6281,N_5723,N_5516);
and U6282 (N_6282,N_5917,N_5925);
nand U6283 (N_6283,N_5908,N_5809);
or U6284 (N_6284,N_5710,N_5738);
nand U6285 (N_6285,N_5537,N_5675);
nor U6286 (N_6286,N_5585,N_5586);
nand U6287 (N_6287,N_5772,N_5804);
xor U6288 (N_6288,N_5759,N_5749);
or U6289 (N_6289,N_5990,N_5594);
xor U6290 (N_6290,N_5715,N_5716);
and U6291 (N_6291,N_5675,N_5642);
nand U6292 (N_6292,N_5538,N_5729);
xor U6293 (N_6293,N_5726,N_5825);
and U6294 (N_6294,N_5876,N_5674);
nor U6295 (N_6295,N_5519,N_5714);
and U6296 (N_6296,N_5517,N_5589);
or U6297 (N_6297,N_5597,N_5955);
nand U6298 (N_6298,N_5755,N_5672);
and U6299 (N_6299,N_5564,N_5589);
xnor U6300 (N_6300,N_5921,N_5761);
or U6301 (N_6301,N_5921,N_5654);
and U6302 (N_6302,N_5924,N_5990);
xor U6303 (N_6303,N_5814,N_5606);
nor U6304 (N_6304,N_5769,N_5503);
xor U6305 (N_6305,N_5656,N_5895);
nand U6306 (N_6306,N_5628,N_5789);
xnor U6307 (N_6307,N_5979,N_5549);
and U6308 (N_6308,N_5694,N_5599);
nand U6309 (N_6309,N_5943,N_5807);
or U6310 (N_6310,N_5749,N_5646);
nand U6311 (N_6311,N_5671,N_5921);
nor U6312 (N_6312,N_5932,N_5646);
nand U6313 (N_6313,N_5683,N_5658);
nand U6314 (N_6314,N_5570,N_5635);
and U6315 (N_6315,N_5882,N_5635);
xor U6316 (N_6316,N_5713,N_5559);
nor U6317 (N_6317,N_5505,N_5790);
nand U6318 (N_6318,N_5560,N_5608);
nor U6319 (N_6319,N_5729,N_5667);
or U6320 (N_6320,N_5804,N_5746);
xnor U6321 (N_6321,N_5669,N_5651);
nor U6322 (N_6322,N_5569,N_5971);
nand U6323 (N_6323,N_5693,N_5896);
or U6324 (N_6324,N_5640,N_5567);
nand U6325 (N_6325,N_5725,N_5952);
nand U6326 (N_6326,N_5714,N_5731);
xnor U6327 (N_6327,N_5935,N_5797);
or U6328 (N_6328,N_5827,N_5689);
nor U6329 (N_6329,N_5789,N_5718);
or U6330 (N_6330,N_5941,N_5920);
nor U6331 (N_6331,N_5918,N_5957);
or U6332 (N_6332,N_5640,N_5593);
and U6333 (N_6333,N_5548,N_5608);
xnor U6334 (N_6334,N_5601,N_5697);
and U6335 (N_6335,N_5866,N_5683);
or U6336 (N_6336,N_5792,N_5819);
or U6337 (N_6337,N_5771,N_5671);
and U6338 (N_6338,N_5920,N_5561);
or U6339 (N_6339,N_5546,N_5569);
nor U6340 (N_6340,N_5970,N_5593);
or U6341 (N_6341,N_5844,N_5676);
and U6342 (N_6342,N_5628,N_5540);
and U6343 (N_6343,N_5777,N_5736);
nand U6344 (N_6344,N_5727,N_5939);
nand U6345 (N_6345,N_5967,N_5564);
or U6346 (N_6346,N_5799,N_5688);
and U6347 (N_6347,N_5510,N_5669);
nor U6348 (N_6348,N_5583,N_5671);
and U6349 (N_6349,N_5523,N_5760);
xnor U6350 (N_6350,N_5597,N_5838);
and U6351 (N_6351,N_5876,N_5531);
nand U6352 (N_6352,N_5535,N_5619);
xnor U6353 (N_6353,N_5868,N_5651);
xor U6354 (N_6354,N_5885,N_5780);
nand U6355 (N_6355,N_5831,N_5829);
or U6356 (N_6356,N_5678,N_5816);
or U6357 (N_6357,N_5994,N_5785);
nor U6358 (N_6358,N_5615,N_5935);
xnor U6359 (N_6359,N_5786,N_5694);
nor U6360 (N_6360,N_5794,N_5845);
xor U6361 (N_6361,N_5755,N_5610);
nand U6362 (N_6362,N_5777,N_5894);
xor U6363 (N_6363,N_5813,N_5850);
nand U6364 (N_6364,N_5823,N_5931);
and U6365 (N_6365,N_5913,N_5793);
or U6366 (N_6366,N_5797,N_5871);
nor U6367 (N_6367,N_5516,N_5896);
and U6368 (N_6368,N_5869,N_5825);
nand U6369 (N_6369,N_5680,N_5630);
or U6370 (N_6370,N_5585,N_5738);
xnor U6371 (N_6371,N_5722,N_5859);
and U6372 (N_6372,N_5611,N_5624);
or U6373 (N_6373,N_5581,N_5919);
or U6374 (N_6374,N_5771,N_5625);
and U6375 (N_6375,N_5852,N_5575);
or U6376 (N_6376,N_5842,N_5810);
nor U6377 (N_6377,N_5703,N_5862);
nor U6378 (N_6378,N_5862,N_5648);
and U6379 (N_6379,N_5614,N_5714);
nand U6380 (N_6380,N_5736,N_5642);
nand U6381 (N_6381,N_5655,N_5887);
or U6382 (N_6382,N_5605,N_5731);
or U6383 (N_6383,N_5814,N_5708);
nand U6384 (N_6384,N_5731,N_5905);
xnor U6385 (N_6385,N_5763,N_5980);
nor U6386 (N_6386,N_5709,N_5648);
or U6387 (N_6387,N_5888,N_5794);
nor U6388 (N_6388,N_5828,N_5992);
and U6389 (N_6389,N_5819,N_5876);
nor U6390 (N_6390,N_5864,N_5505);
and U6391 (N_6391,N_5664,N_5604);
and U6392 (N_6392,N_5637,N_5520);
xnor U6393 (N_6393,N_5933,N_5550);
and U6394 (N_6394,N_5696,N_5591);
xnor U6395 (N_6395,N_5985,N_5667);
nor U6396 (N_6396,N_5576,N_5984);
and U6397 (N_6397,N_5988,N_5704);
nand U6398 (N_6398,N_5754,N_5876);
and U6399 (N_6399,N_5579,N_5575);
nor U6400 (N_6400,N_5826,N_5963);
and U6401 (N_6401,N_5999,N_5837);
nor U6402 (N_6402,N_5627,N_5682);
xnor U6403 (N_6403,N_5998,N_5991);
nand U6404 (N_6404,N_5658,N_5558);
and U6405 (N_6405,N_5950,N_5545);
nor U6406 (N_6406,N_5580,N_5953);
nor U6407 (N_6407,N_5836,N_5933);
or U6408 (N_6408,N_5882,N_5704);
and U6409 (N_6409,N_5591,N_5755);
xor U6410 (N_6410,N_5885,N_5865);
nor U6411 (N_6411,N_5767,N_5776);
and U6412 (N_6412,N_5751,N_5624);
and U6413 (N_6413,N_5900,N_5824);
or U6414 (N_6414,N_5868,N_5586);
nor U6415 (N_6415,N_5891,N_5524);
nand U6416 (N_6416,N_5928,N_5611);
nand U6417 (N_6417,N_5848,N_5674);
nor U6418 (N_6418,N_5969,N_5589);
nor U6419 (N_6419,N_5943,N_5754);
nand U6420 (N_6420,N_5977,N_5842);
or U6421 (N_6421,N_5674,N_5889);
or U6422 (N_6422,N_5649,N_5652);
xor U6423 (N_6423,N_5917,N_5672);
and U6424 (N_6424,N_5664,N_5677);
nand U6425 (N_6425,N_5996,N_5932);
nor U6426 (N_6426,N_5594,N_5563);
nand U6427 (N_6427,N_5854,N_5894);
and U6428 (N_6428,N_5962,N_5897);
xnor U6429 (N_6429,N_5910,N_5745);
nor U6430 (N_6430,N_5785,N_5569);
nand U6431 (N_6431,N_5623,N_5982);
nor U6432 (N_6432,N_5833,N_5974);
or U6433 (N_6433,N_5575,N_5824);
xnor U6434 (N_6434,N_5536,N_5764);
and U6435 (N_6435,N_5637,N_5943);
and U6436 (N_6436,N_5886,N_5849);
or U6437 (N_6437,N_5742,N_5662);
xnor U6438 (N_6438,N_5838,N_5605);
and U6439 (N_6439,N_5794,N_5837);
nor U6440 (N_6440,N_5541,N_5655);
xnor U6441 (N_6441,N_5690,N_5555);
xnor U6442 (N_6442,N_5796,N_5787);
nor U6443 (N_6443,N_5907,N_5831);
and U6444 (N_6444,N_5813,N_5818);
or U6445 (N_6445,N_5524,N_5890);
or U6446 (N_6446,N_5564,N_5865);
nor U6447 (N_6447,N_5565,N_5578);
nand U6448 (N_6448,N_5599,N_5662);
xnor U6449 (N_6449,N_5781,N_5746);
and U6450 (N_6450,N_5656,N_5793);
nand U6451 (N_6451,N_5850,N_5909);
and U6452 (N_6452,N_5699,N_5955);
and U6453 (N_6453,N_5794,N_5562);
and U6454 (N_6454,N_5594,N_5973);
and U6455 (N_6455,N_5623,N_5961);
nor U6456 (N_6456,N_5930,N_5683);
or U6457 (N_6457,N_5554,N_5975);
nor U6458 (N_6458,N_5834,N_5548);
nand U6459 (N_6459,N_5676,N_5794);
and U6460 (N_6460,N_5575,N_5568);
xor U6461 (N_6461,N_5650,N_5950);
and U6462 (N_6462,N_5825,N_5608);
nand U6463 (N_6463,N_5731,N_5989);
xnor U6464 (N_6464,N_5649,N_5691);
or U6465 (N_6465,N_5951,N_5678);
xor U6466 (N_6466,N_5987,N_5902);
nor U6467 (N_6467,N_5526,N_5695);
and U6468 (N_6468,N_5952,N_5749);
xor U6469 (N_6469,N_5511,N_5564);
or U6470 (N_6470,N_5624,N_5892);
and U6471 (N_6471,N_5857,N_5933);
nor U6472 (N_6472,N_5780,N_5813);
and U6473 (N_6473,N_5537,N_5961);
and U6474 (N_6474,N_5601,N_5871);
xor U6475 (N_6475,N_5905,N_5825);
or U6476 (N_6476,N_5849,N_5882);
xor U6477 (N_6477,N_5647,N_5749);
nand U6478 (N_6478,N_5511,N_5900);
nor U6479 (N_6479,N_5815,N_5774);
and U6480 (N_6480,N_5807,N_5734);
nor U6481 (N_6481,N_5742,N_5713);
nor U6482 (N_6482,N_5978,N_5746);
or U6483 (N_6483,N_5847,N_5953);
nor U6484 (N_6484,N_5844,N_5750);
xor U6485 (N_6485,N_5990,N_5629);
or U6486 (N_6486,N_5661,N_5519);
and U6487 (N_6487,N_5678,N_5859);
xor U6488 (N_6488,N_5883,N_5521);
or U6489 (N_6489,N_5511,N_5897);
nor U6490 (N_6490,N_5618,N_5880);
or U6491 (N_6491,N_5841,N_5847);
and U6492 (N_6492,N_5639,N_5816);
or U6493 (N_6493,N_5505,N_5513);
xor U6494 (N_6494,N_5905,N_5694);
and U6495 (N_6495,N_5604,N_5511);
nand U6496 (N_6496,N_5528,N_5502);
and U6497 (N_6497,N_5769,N_5741);
xor U6498 (N_6498,N_5660,N_5577);
and U6499 (N_6499,N_5591,N_5908);
and U6500 (N_6500,N_6111,N_6266);
and U6501 (N_6501,N_6101,N_6071);
xnor U6502 (N_6502,N_6077,N_6197);
nor U6503 (N_6503,N_6092,N_6464);
xor U6504 (N_6504,N_6063,N_6436);
and U6505 (N_6505,N_6329,N_6315);
xor U6506 (N_6506,N_6350,N_6121);
nor U6507 (N_6507,N_6392,N_6129);
and U6508 (N_6508,N_6496,N_6282);
xnor U6509 (N_6509,N_6478,N_6354);
nand U6510 (N_6510,N_6386,N_6116);
xnor U6511 (N_6511,N_6316,N_6476);
or U6512 (N_6512,N_6135,N_6345);
or U6513 (N_6513,N_6148,N_6061);
nor U6514 (N_6514,N_6170,N_6403);
nor U6515 (N_6515,N_6480,N_6363);
nand U6516 (N_6516,N_6374,N_6455);
xor U6517 (N_6517,N_6167,N_6183);
and U6518 (N_6518,N_6239,N_6078);
xnor U6519 (N_6519,N_6346,N_6497);
or U6520 (N_6520,N_6185,N_6328);
or U6521 (N_6521,N_6140,N_6163);
nand U6522 (N_6522,N_6457,N_6019);
and U6523 (N_6523,N_6380,N_6186);
nand U6524 (N_6524,N_6275,N_6112);
and U6525 (N_6525,N_6371,N_6330);
nand U6526 (N_6526,N_6000,N_6335);
nor U6527 (N_6527,N_6204,N_6168);
xor U6528 (N_6528,N_6070,N_6219);
xor U6529 (N_6529,N_6267,N_6390);
or U6530 (N_6530,N_6094,N_6445);
nand U6531 (N_6531,N_6337,N_6192);
xor U6532 (N_6532,N_6472,N_6288);
or U6533 (N_6533,N_6347,N_6169);
xnor U6534 (N_6534,N_6389,N_6369);
and U6535 (N_6535,N_6110,N_6383);
nand U6536 (N_6536,N_6408,N_6143);
xnor U6537 (N_6537,N_6285,N_6249);
nor U6538 (N_6538,N_6014,N_6271);
or U6539 (N_6539,N_6297,N_6296);
nor U6540 (N_6540,N_6475,N_6032);
nand U6541 (N_6541,N_6470,N_6397);
and U6542 (N_6542,N_6076,N_6366);
xnor U6543 (N_6543,N_6165,N_6274);
or U6544 (N_6544,N_6232,N_6474);
xor U6545 (N_6545,N_6039,N_6115);
nor U6546 (N_6546,N_6171,N_6079);
and U6547 (N_6547,N_6263,N_6352);
nor U6548 (N_6548,N_6237,N_6086);
or U6549 (N_6549,N_6283,N_6405);
and U6550 (N_6550,N_6214,N_6130);
or U6551 (N_6551,N_6359,N_6458);
and U6552 (N_6552,N_6045,N_6294);
xnor U6553 (N_6553,N_6264,N_6291);
nand U6554 (N_6554,N_6377,N_6238);
and U6555 (N_6555,N_6256,N_6339);
xor U6556 (N_6556,N_6479,N_6090);
xnor U6557 (N_6557,N_6320,N_6102);
nand U6558 (N_6558,N_6376,N_6208);
or U6559 (N_6559,N_6146,N_6189);
nand U6560 (N_6560,N_6029,N_6098);
or U6561 (N_6561,N_6492,N_6033);
xnor U6562 (N_6562,N_6428,N_6103);
xnor U6563 (N_6563,N_6338,N_6203);
xnor U6564 (N_6564,N_6318,N_6194);
xnor U6565 (N_6565,N_6388,N_6286);
xor U6566 (N_6566,N_6284,N_6298);
and U6567 (N_6567,N_6051,N_6317);
and U6568 (N_6568,N_6209,N_6424);
nor U6569 (N_6569,N_6401,N_6048);
nor U6570 (N_6570,N_6268,N_6404);
and U6571 (N_6571,N_6097,N_6250);
and U6572 (N_6572,N_6440,N_6336);
nand U6573 (N_6573,N_6423,N_6196);
nand U6574 (N_6574,N_6304,N_6243);
or U6575 (N_6575,N_6142,N_6226);
xor U6576 (N_6576,N_6410,N_6490);
xnor U6577 (N_6577,N_6289,N_6002);
nand U6578 (N_6578,N_6124,N_6152);
xor U6579 (N_6579,N_6444,N_6370);
xnor U6580 (N_6580,N_6295,N_6119);
nand U6581 (N_6581,N_6314,N_6016);
xnor U6582 (N_6582,N_6050,N_6303);
xnor U6583 (N_6583,N_6109,N_6139);
and U6584 (N_6584,N_6198,N_6439);
or U6585 (N_6585,N_6446,N_6481);
and U6586 (N_6586,N_6368,N_6230);
or U6587 (N_6587,N_6413,N_6447);
xnor U6588 (N_6588,N_6128,N_6195);
and U6589 (N_6589,N_6173,N_6099);
or U6590 (N_6590,N_6340,N_6035);
nand U6591 (N_6591,N_6281,N_6027);
nand U6592 (N_6592,N_6151,N_6058);
nor U6593 (N_6593,N_6123,N_6387);
and U6594 (N_6594,N_6187,N_6161);
nand U6595 (N_6595,N_6093,N_6062);
or U6596 (N_6596,N_6017,N_6469);
xnor U6597 (N_6597,N_6415,N_6391);
xnor U6598 (N_6598,N_6085,N_6133);
xnor U6599 (N_6599,N_6269,N_6011);
or U6600 (N_6600,N_6227,N_6299);
xor U6601 (N_6601,N_6026,N_6084);
and U6602 (N_6602,N_6036,N_6348);
nor U6603 (N_6603,N_6435,N_6118);
and U6604 (N_6604,N_6427,N_6212);
nor U6605 (N_6605,N_6041,N_6433);
nand U6606 (N_6606,N_6324,N_6095);
or U6607 (N_6607,N_6057,N_6015);
nor U6608 (N_6608,N_6012,N_6040);
nand U6609 (N_6609,N_6466,N_6331);
and U6610 (N_6610,N_6100,N_6334);
nor U6611 (N_6611,N_6494,N_6364);
nor U6612 (N_6612,N_6325,N_6149);
nor U6613 (N_6613,N_6477,N_6305);
or U6614 (N_6614,N_6006,N_6177);
or U6615 (N_6615,N_6459,N_6273);
or U6616 (N_6616,N_6008,N_6240);
and U6617 (N_6617,N_6157,N_6126);
and U6618 (N_6618,N_6341,N_6333);
xnor U6619 (N_6619,N_6155,N_6327);
nor U6620 (N_6620,N_6431,N_6162);
nand U6621 (N_6621,N_6235,N_6489);
nor U6622 (N_6622,N_6398,N_6419);
and U6623 (N_6623,N_6024,N_6355);
nor U6624 (N_6624,N_6178,N_6302);
or U6625 (N_6625,N_6483,N_6381);
nor U6626 (N_6626,N_6059,N_6255);
and U6627 (N_6627,N_6241,N_6400);
and U6628 (N_6628,N_6499,N_6108);
xor U6629 (N_6629,N_6430,N_6396);
xor U6630 (N_6630,N_6456,N_6441);
xnor U6631 (N_6631,N_6125,N_6420);
nor U6632 (N_6632,N_6225,N_6007);
and U6633 (N_6633,N_6200,N_6406);
xnor U6634 (N_6634,N_6145,N_6245);
nand U6635 (N_6635,N_6362,N_6003);
or U6636 (N_6636,N_6234,N_6174);
nand U6637 (N_6637,N_6087,N_6069);
xnor U6638 (N_6638,N_6306,N_6248);
nor U6639 (N_6639,N_6107,N_6160);
and U6640 (N_6640,N_6493,N_6342);
nand U6641 (N_6641,N_6182,N_6010);
nor U6642 (N_6642,N_6307,N_6437);
and U6643 (N_6643,N_6202,N_6005);
nand U6644 (N_6644,N_6236,N_6301);
and U6645 (N_6645,N_6313,N_6184);
and U6646 (N_6646,N_6290,N_6075);
xnor U6647 (N_6647,N_6021,N_6279);
xor U6648 (N_6648,N_6088,N_6216);
nor U6649 (N_6649,N_6242,N_6068);
nand U6650 (N_6650,N_6451,N_6074);
nor U6651 (N_6651,N_6417,N_6030);
nor U6652 (N_6652,N_6188,N_6222);
and U6653 (N_6653,N_6332,N_6190);
nand U6654 (N_6654,N_6223,N_6233);
nand U6655 (N_6655,N_6300,N_6104);
xnor U6656 (N_6656,N_6056,N_6448);
or U6657 (N_6657,N_6259,N_6105);
nand U6658 (N_6658,N_6311,N_6375);
or U6659 (N_6659,N_6414,N_6218);
xor U6660 (N_6660,N_6292,N_6025);
xnor U6661 (N_6661,N_6367,N_6052);
nor U6662 (N_6662,N_6022,N_6421);
xor U6663 (N_6663,N_6215,N_6495);
nor U6664 (N_6664,N_6395,N_6081);
nor U6665 (N_6665,N_6091,N_6344);
and U6666 (N_6666,N_6131,N_6144);
xnor U6667 (N_6667,N_6193,N_6137);
nor U6668 (N_6668,N_6031,N_6049);
xor U6669 (N_6669,N_6001,N_6205);
nand U6670 (N_6670,N_6454,N_6491);
xnor U6671 (N_6671,N_6023,N_6166);
xor U6672 (N_6672,N_6361,N_6278);
xor U6673 (N_6673,N_6409,N_6132);
and U6674 (N_6674,N_6309,N_6067);
nand U6675 (N_6675,N_6452,N_6498);
nor U6676 (N_6676,N_6080,N_6009);
nor U6677 (N_6677,N_6310,N_6229);
xor U6678 (N_6678,N_6261,N_6207);
and U6679 (N_6679,N_6004,N_6013);
nor U6680 (N_6680,N_6247,N_6073);
nand U6681 (N_6681,N_6422,N_6323);
xnor U6682 (N_6682,N_6260,N_6321);
and U6683 (N_6683,N_6429,N_6257);
or U6684 (N_6684,N_6382,N_6083);
or U6685 (N_6685,N_6206,N_6418);
or U6686 (N_6686,N_6349,N_6468);
and U6687 (N_6687,N_6358,N_6037);
xor U6688 (N_6688,N_6312,N_6265);
xnor U6689 (N_6689,N_6096,N_6461);
xnor U6690 (N_6690,N_6357,N_6191);
xor U6691 (N_6691,N_6072,N_6179);
nor U6692 (N_6692,N_6365,N_6221);
and U6693 (N_6693,N_6425,N_6258);
xnor U6694 (N_6694,N_6407,N_6356);
or U6695 (N_6695,N_6293,N_6442);
nor U6696 (N_6696,N_6319,N_6326);
or U6697 (N_6697,N_6181,N_6438);
xor U6698 (N_6698,N_6117,N_6199);
and U6699 (N_6699,N_6402,N_6450);
and U6700 (N_6700,N_6385,N_6038);
nor U6701 (N_6701,N_6164,N_6147);
or U6702 (N_6702,N_6416,N_6053);
or U6703 (N_6703,N_6211,N_6043);
nor U6704 (N_6704,N_6343,N_6379);
nor U6705 (N_6705,N_6176,N_6252);
nor U6706 (N_6706,N_6018,N_6308);
nand U6707 (N_6707,N_6254,N_6220);
nor U6708 (N_6708,N_6449,N_6287);
and U6709 (N_6709,N_6106,N_6217);
xor U6710 (N_6710,N_6486,N_6180);
nand U6711 (N_6711,N_6154,N_6134);
and U6712 (N_6712,N_6138,N_6373);
nand U6713 (N_6713,N_6127,N_6175);
or U6714 (N_6714,N_6384,N_6213);
or U6715 (N_6715,N_6201,N_6353);
nor U6716 (N_6716,N_6141,N_6393);
and U6717 (N_6717,N_6473,N_6463);
and U6718 (N_6718,N_6159,N_6065);
and U6719 (N_6719,N_6487,N_6277);
nor U6720 (N_6720,N_6262,N_6122);
nand U6721 (N_6721,N_6251,N_6046);
and U6722 (N_6722,N_6465,N_6113);
nor U6723 (N_6723,N_6172,N_6054);
nand U6724 (N_6724,N_6082,N_6228);
nor U6725 (N_6725,N_6443,N_6270);
nor U6726 (N_6726,N_6064,N_6231);
nand U6727 (N_6727,N_6351,N_6114);
xnor U6728 (N_6728,N_6210,N_6453);
nand U6729 (N_6729,N_6136,N_6426);
and U6730 (N_6730,N_6224,N_6042);
and U6731 (N_6731,N_6482,N_6434);
nor U6732 (N_6732,N_6044,N_6047);
nand U6733 (N_6733,N_6322,N_6020);
or U6734 (N_6734,N_6467,N_6412);
and U6735 (N_6735,N_6034,N_6066);
nor U6736 (N_6736,N_6272,N_6089);
nand U6737 (N_6737,N_6060,N_6153);
xnor U6738 (N_6738,N_6411,N_6244);
xnor U6739 (N_6739,N_6253,N_6246);
nand U6740 (N_6740,N_6280,N_6485);
or U6741 (N_6741,N_6150,N_6471);
xor U6742 (N_6742,N_6462,N_6378);
and U6743 (N_6743,N_6156,N_6360);
xnor U6744 (N_6744,N_6055,N_6399);
and U6745 (N_6745,N_6158,N_6460);
nand U6746 (N_6746,N_6488,N_6394);
nor U6747 (N_6747,N_6484,N_6028);
or U6748 (N_6748,N_6432,N_6120);
and U6749 (N_6749,N_6372,N_6276);
nor U6750 (N_6750,N_6434,N_6025);
nand U6751 (N_6751,N_6133,N_6091);
nand U6752 (N_6752,N_6134,N_6464);
nand U6753 (N_6753,N_6095,N_6166);
nor U6754 (N_6754,N_6161,N_6081);
nand U6755 (N_6755,N_6232,N_6059);
and U6756 (N_6756,N_6036,N_6333);
nor U6757 (N_6757,N_6312,N_6007);
xor U6758 (N_6758,N_6035,N_6477);
xnor U6759 (N_6759,N_6323,N_6246);
nor U6760 (N_6760,N_6415,N_6187);
or U6761 (N_6761,N_6387,N_6329);
and U6762 (N_6762,N_6301,N_6219);
nand U6763 (N_6763,N_6266,N_6487);
nor U6764 (N_6764,N_6043,N_6210);
xnor U6765 (N_6765,N_6416,N_6092);
nand U6766 (N_6766,N_6254,N_6454);
xnor U6767 (N_6767,N_6225,N_6336);
nor U6768 (N_6768,N_6434,N_6236);
nor U6769 (N_6769,N_6260,N_6117);
or U6770 (N_6770,N_6133,N_6184);
xnor U6771 (N_6771,N_6223,N_6130);
and U6772 (N_6772,N_6445,N_6292);
and U6773 (N_6773,N_6109,N_6335);
nor U6774 (N_6774,N_6438,N_6123);
xor U6775 (N_6775,N_6291,N_6268);
nor U6776 (N_6776,N_6216,N_6390);
nand U6777 (N_6777,N_6441,N_6110);
and U6778 (N_6778,N_6128,N_6349);
nor U6779 (N_6779,N_6092,N_6366);
or U6780 (N_6780,N_6097,N_6475);
nor U6781 (N_6781,N_6028,N_6091);
or U6782 (N_6782,N_6205,N_6026);
nand U6783 (N_6783,N_6350,N_6193);
nand U6784 (N_6784,N_6260,N_6267);
and U6785 (N_6785,N_6401,N_6275);
nor U6786 (N_6786,N_6214,N_6243);
nand U6787 (N_6787,N_6249,N_6436);
nand U6788 (N_6788,N_6416,N_6370);
xor U6789 (N_6789,N_6492,N_6440);
nand U6790 (N_6790,N_6152,N_6326);
and U6791 (N_6791,N_6221,N_6250);
xor U6792 (N_6792,N_6030,N_6490);
nand U6793 (N_6793,N_6280,N_6494);
or U6794 (N_6794,N_6387,N_6458);
nor U6795 (N_6795,N_6216,N_6187);
or U6796 (N_6796,N_6031,N_6272);
nand U6797 (N_6797,N_6234,N_6072);
and U6798 (N_6798,N_6203,N_6473);
xnor U6799 (N_6799,N_6340,N_6326);
xor U6800 (N_6800,N_6167,N_6464);
xor U6801 (N_6801,N_6394,N_6375);
or U6802 (N_6802,N_6051,N_6076);
nand U6803 (N_6803,N_6476,N_6219);
nor U6804 (N_6804,N_6383,N_6488);
or U6805 (N_6805,N_6264,N_6348);
and U6806 (N_6806,N_6051,N_6350);
xor U6807 (N_6807,N_6002,N_6234);
nor U6808 (N_6808,N_6431,N_6072);
or U6809 (N_6809,N_6165,N_6070);
or U6810 (N_6810,N_6467,N_6111);
nand U6811 (N_6811,N_6261,N_6493);
or U6812 (N_6812,N_6074,N_6180);
and U6813 (N_6813,N_6226,N_6006);
and U6814 (N_6814,N_6361,N_6080);
and U6815 (N_6815,N_6045,N_6498);
nor U6816 (N_6816,N_6016,N_6267);
nand U6817 (N_6817,N_6222,N_6421);
and U6818 (N_6818,N_6290,N_6345);
nand U6819 (N_6819,N_6028,N_6227);
or U6820 (N_6820,N_6134,N_6275);
and U6821 (N_6821,N_6249,N_6054);
or U6822 (N_6822,N_6318,N_6193);
nor U6823 (N_6823,N_6286,N_6145);
xnor U6824 (N_6824,N_6343,N_6193);
nor U6825 (N_6825,N_6445,N_6108);
or U6826 (N_6826,N_6318,N_6441);
nand U6827 (N_6827,N_6032,N_6002);
and U6828 (N_6828,N_6253,N_6146);
and U6829 (N_6829,N_6390,N_6439);
or U6830 (N_6830,N_6059,N_6486);
and U6831 (N_6831,N_6001,N_6452);
and U6832 (N_6832,N_6187,N_6371);
nor U6833 (N_6833,N_6220,N_6228);
nor U6834 (N_6834,N_6049,N_6198);
nor U6835 (N_6835,N_6252,N_6480);
nor U6836 (N_6836,N_6373,N_6150);
nand U6837 (N_6837,N_6440,N_6247);
xnor U6838 (N_6838,N_6132,N_6272);
xnor U6839 (N_6839,N_6226,N_6104);
xor U6840 (N_6840,N_6370,N_6336);
xor U6841 (N_6841,N_6025,N_6401);
nand U6842 (N_6842,N_6192,N_6252);
nand U6843 (N_6843,N_6485,N_6490);
and U6844 (N_6844,N_6202,N_6010);
and U6845 (N_6845,N_6202,N_6141);
or U6846 (N_6846,N_6190,N_6324);
or U6847 (N_6847,N_6261,N_6209);
nor U6848 (N_6848,N_6350,N_6008);
or U6849 (N_6849,N_6417,N_6431);
nor U6850 (N_6850,N_6241,N_6384);
nor U6851 (N_6851,N_6403,N_6106);
xnor U6852 (N_6852,N_6083,N_6002);
nor U6853 (N_6853,N_6496,N_6289);
nand U6854 (N_6854,N_6046,N_6118);
or U6855 (N_6855,N_6370,N_6169);
xor U6856 (N_6856,N_6249,N_6175);
or U6857 (N_6857,N_6357,N_6203);
or U6858 (N_6858,N_6147,N_6096);
or U6859 (N_6859,N_6028,N_6189);
nand U6860 (N_6860,N_6337,N_6367);
nand U6861 (N_6861,N_6220,N_6326);
or U6862 (N_6862,N_6232,N_6075);
and U6863 (N_6863,N_6000,N_6002);
or U6864 (N_6864,N_6326,N_6297);
xnor U6865 (N_6865,N_6179,N_6158);
or U6866 (N_6866,N_6337,N_6051);
or U6867 (N_6867,N_6033,N_6244);
xor U6868 (N_6868,N_6115,N_6261);
nand U6869 (N_6869,N_6080,N_6105);
nand U6870 (N_6870,N_6288,N_6073);
or U6871 (N_6871,N_6325,N_6197);
nor U6872 (N_6872,N_6088,N_6445);
and U6873 (N_6873,N_6211,N_6162);
nor U6874 (N_6874,N_6477,N_6163);
nor U6875 (N_6875,N_6496,N_6008);
xor U6876 (N_6876,N_6174,N_6032);
nand U6877 (N_6877,N_6186,N_6178);
or U6878 (N_6878,N_6446,N_6127);
and U6879 (N_6879,N_6022,N_6213);
nor U6880 (N_6880,N_6019,N_6260);
xor U6881 (N_6881,N_6002,N_6280);
xnor U6882 (N_6882,N_6381,N_6238);
nand U6883 (N_6883,N_6240,N_6040);
nor U6884 (N_6884,N_6124,N_6007);
and U6885 (N_6885,N_6480,N_6133);
and U6886 (N_6886,N_6411,N_6403);
or U6887 (N_6887,N_6109,N_6330);
and U6888 (N_6888,N_6271,N_6325);
nor U6889 (N_6889,N_6445,N_6281);
and U6890 (N_6890,N_6213,N_6401);
nor U6891 (N_6891,N_6081,N_6178);
and U6892 (N_6892,N_6280,N_6149);
nand U6893 (N_6893,N_6146,N_6286);
nand U6894 (N_6894,N_6133,N_6067);
or U6895 (N_6895,N_6091,N_6358);
nor U6896 (N_6896,N_6384,N_6048);
nor U6897 (N_6897,N_6470,N_6294);
or U6898 (N_6898,N_6475,N_6240);
xnor U6899 (N_6899,N_6357,N_6313);
or U6900 (N_6900,N_6149,N_6181);
and U6901 (N_6901,N_6041,N_6093);
or U6902 (N_6902,N_6130,N_6001);
and U6903 (N_6903,N_6158,N_6472);
nor U6904 (N_6904,N_6470,N_6251);
and U6905 (N_6905,N_6338,N_6170);
nor U6906 (N_6906,N_6104,N_6485);
and U6907 (N_6907,N_6025,N_6079);
and U6908 (N_6908,N_6061,N_6334);
or U6909 (N_6909,N_6052,N_6021);
xnor U6910 (N_6910,N_6221,N_6260);
and U6911 (N_6911,N_6078,N_6040);
or U6912 (N_6912,N_6227,N_6159);
xor U6913 (N_6913,N_6365,N_6002);
or U6914 (N_6914,N_6366,N_6479);
nor U6915 (N_6915,N_6068,N_6104);
xnor U6916 (N_6916,N_6305,N_6392);
nor U6917 (N_6917,N_6298,N_6009);
or U6918 (N_6918,N_6262,N_6346);
or U6919 (N_6919,N_6148,N_6115);
nand U6920 (N_6920,N_6016,N_6185);
xor U6921 (N_6921,N_6424,N_6108);
nand U6922 (N_6922,N_6073,N_6451);
xnor U6923 (N_6923,N_6175,N_6389);
nor U6924 (N_6924,N_6133,N_6463);
and U6925 (N_6925,N_6284,N_6344);
or U6926 (N_6926,N_6327,N_6346);
and U6927 (N_6927,N_6020,N_6119);
or U6928 (N_6928,N_6464,N_6286);
or U6929 (N_6929,N_6194,N_6431);
and U6930 (N_6930,N_6125,N_6489);
nor U6931 (N_6931,N_6016,N_6342);
xor U6932 (N_6932,N_6193,N_6091);
or U6933 (N_6933,N_6008,N_6128);
and U6934 (N_6934,N_6293,N_6336);
xor U6935 (N_6935,N_6202,N_6029);
xnor U6936 (N_6936,N_6172,N_6000);
and U6937 (N_6937,N_6126,N_6290);
and U6938 (N_6938,N_6443,N_6137);
or U6939 (N_6939,N_6263,N_6217);
nand U6940 (N_6940,N_6268,N_6352);
and U6941 (N_6941,N_6379,N_6186);
and U6942 (N_6942,N_6317,N_6252);
and U6943 (N_6943,N_6298,N_6472);
xor U6944 (N_6944,N_6218,N_6211);
and U6945 (N_6945,N_6333,N_6408);
and U6946 (N_6946,N_6201,N_6428);
and U6947 (N_6947,N_6291,N_6089);
xor U6948 (N_6948,N_6366,N_6059);
or U6949 (N_6949,N_6083,N_6173);
nand U6950 (N_6950,N_6183,N_6032);
or U6951 (N_6951,N_6430,N_6029);
or U6952 (N_6952,N_6345,N_6158);
nor U6953 (N_6953,N_6036,N_6201);
xor U6954 (N_6954,N_6020,N_6225);
nand U6955 (N_6955,N_6185,N_6497);
xor U6956 (N_6956,N_6495,N_6316);
xor U6957 (N_6957,N_6484,N_6431);
and U6958 (N_6958,N_6142,N_6384);
nor U6959 (N_6959,N_6354,N_6498);
or U6960 (N_6960,N_6081,N_6492);
nor U6961 (N_6961,N_6165,N_6139);
xnor U6962 (N_6962,N_6116,N_6423);
and U6963 (N_6963,N_6297,N_6367);
nand U6964 (N_6964,N_6482,N_6117);
nor U6965 (N_6965,N_6211,N_6390);
nor U6966 (N_6966,N_6128,N_6119);
and U6967 (N_6967,N_6207,N_6345);
nand U6968 (N_6968,N_6033,N_6439);
xor U6969 (N_6969,N_6334,N_6206);
or U6970 (N_6970,N_6215,N_6086);
nor U6971 (N_6971,N_6067,N_6448);
xor U6972 (N_6972,N_6385,N_6358);
or U6973 (N_6973,N_6037,N_6310);
or U6974 (N_6974,N_6147,N_6301);
or U6975 (N_6975,N_6279,N_6206);
xnor U6976 (N_6976,N_6179,N_6447);
nand U6977 (N_6977,N_6353,N_6144);
nand U6978 (N_6978,N_6453,N_6013);
and U6979 (N_6979,N_6271,N_6235);
nor U6980 (N_6980,N_6034,N_6146);
or U6981 (N_6981,N_6201,N_6250);
nor U6982 (N_6982,N_6137,N_6165);
or U6983 (N_6983,N_6176,N_6057);
nor U6984 (N_6984,N_6433,N_6155);
nand U6985 (N_6985,N_6429,N_6333);
nor U6986 (N_6986,N_6221,N_6012);
nor U6987 (N_6987,N_6081,N_6495);
nand U6988 (N_6988,N_6052,N_6070);
nand U6989 (N_6989,N_6281,N_6270);
and U6990 (N_6990,N_6349,N_6097);
xnor U6991 (N_6991,N_6474,N_6343);
nand U6992 (N_6992,N_6256,N_6396);
or U6993 (N_6993,N_6238,N_6069);
and U6994 (N_6994,N_6159,N_6169);
and U6995 (N_6995,N_6199,N_6428);
nand U6996 (N_6996,N_6379,N_6306);
and U6997 (N_6997,N_6270,N_6199);
and U6998 (N_6998,N_6308,N_6108);
xor U6999 (N_6999,N_6357,N_6105);
or U7000 (N_7000,N_6747,N_6505);
xor U7001 (N_7001,N_6774,N_6500);
or U7002 (N_7002,N_6905,N_6887);
xor U7003 (N_7003,N_6904,N_6892);
nor U7004 (N_7004,N_6609,N_6736);
nor U7005 (N_7005,N_6829,N_6949);
nand U7006 (N_7006,N_6832,N_6742);
or U7007 (N_7007,N_6955,N_6557);
nor U7008 (N_7008,N_6817,N_6737);
or U7009 (N_7009,N_6794,N_6782);
nand U7010 (N_7010,N_6992,N_6978);
xnor U7011 (N_7011,N_6997,N_6944);
nand U7012 (N_7012,N_6532,N_6523);
or U7013 (N_7013,N_6787,N_6819);
or U7014 (N_7014,N_6545,N_6508);
xor U7015 (N_7015,N_6743,N_6839);
nand U7016 (N_7016,N_6648,N_6823);
or U7017 (N_7017,N_6756,N_6726);
and U7018 (N_7018,N_6600,N_6682);
nor U7019 (N_7019,N_6546,N_6598);
nor U7020 (N_7020,N_6588,N_6512);
nand U7021 (N_7021,N_6681,N_6964);
nor U7022 (N_7022,N_6719,N_6547);
nand U7023 (N_7023,N_6601,N_6750);
or U7024 (N_7024,N_6927,N_6740);
or U7025 (N_7025,N_6801,N_6699);
or U7026 (N_7026,N_6816,N_6886);
xnor U7027 (N_7027,N_6834,N_6570);
or U7028 (N_7028,N_6773,N_6748);
or U7029 (N_7029,N_6576,N_6830);
xnor U7030 (N_7030,N_6614,N_6530);
and U7031 (N_7031,N_6898,N_6919);
and U7032 (N_7032,N_6804,N_6565);
and U7033 (N_7033,N_6651,N_6504);
nor U7034 (N_7034,N_6718,N_6684);
or U7035 (N_7035,N_6999,N_6710);
or U7036 (N_7036,N_6515,N_6907);
nor U7037 (N_7037,N_6826,N_6783);
nor U7038 (N_7038,N_6555,N_6874);
xor U7039 (N_7039,N_6779,N_6825);
and U7040 (N_7040,N_6702,N_6940);
xor U7041 (N_7041,N_6861,N_6608);
nand U7042 (N_7042,N_6833,N_6688);
or U7043 (N_7043,N_6679,N_6948);
nand U7044 (N_7044,N_6900,N_6667);
or U7045 (N_7045,N_6752,N_6594);
xor U7046 (N_7046,N_6820,N_6522);
nor U7047 (N_7047,N_6633,N_6622);
and U7048 (N_7048,N_6569,N_6507);
or U7049 (N_7049,N_6597,N_6984);
nand U7050 (N_7050,N_6706,N_6968);
and U7051 (N_7051,N_6627,N_6923);
xnor U7052 (N_7052,N_6800,N_6666);
and U7053 (N_7053,N_6631,N_6730);
nor U7054 (N_7054,N_6806,N_6851);
nor U7055 (N_7055,N_6521,N_6761);
or U7056 (N_7056,N_6632,N_6925);
nor U7057 (N_7057,N_6722,N_6689);
nor U7058 (N_7058,N_6864,N_6640);
nor U7059 (N_7059,N_6603,N_6813);
or U7060 (N_7060,N_6916,N_6815);
nand U7061 (N_7061,N_6653,N_6906);
nor U7062 (N_7062,N_6553,N_6974);
nand U7063 (N_7063,N_6858,N_6767);
or U7064 (N_7064,N_6996,N_6528);
xnor U7065 (N_7065,N_6837,N_6797);
nand U7066 (N_7066,N_6639,N_6953);
or U7067 (N_7067,N_6717,N_6994);
nand U7068 (N_7068,N_6912,N_6729);
nor U7069 (N_7069,N_6960,N_6971);
xor U7070 (N_7070,N_6791,N_6929);
and U7071 (N_7071,N_6693,N_6979);
nand U7072 (N_7072,N_6764,N_6728);
xnor U7073 (N_7073,N_6866,N_6962);
xnor U7074 (N_7074,N_6928,N_6604);
nand U7075 (N_7075,N_6692,N_6672);
xnor U7076 (N_7076,N_6655,N_6535);
or U7077 (N_7077,N_6758,N_6674);
xnor U7078 (N_7078,N_6937,N_6678);
nand U7079 (N_7079,N_6664,N_6592);
and U7080 (N_7080,N_6540,N_6510);
or U7081 (N_7081,N_6513,N_6757);
xor U7082 (N_7082,N_6981,N_6503);
nand U7083 (N_7083,N_6646,N_6642);
nand U7084 (N_7084,N_6776,N_6768);
nor U7085 (N_7085,N_6873,N_6760);
nand U7086 (N_7086,N_6876,N_6753);
nand U7087 (N_7087,N_6720,N_6769);
and U7088 (N_7088,N_6824,N_6903);
nand U7089 (N_7089,N_6685,N_6607);
nand U7090 (N_7090,N_6613,N_6550);
or U7091 (N_7091,N_6660,N_6657);
nand U7092 (N_7092,N_6599,N_6775);
xor U7093 (N_7093,N_6854,N_6872);
or U7094 (N_7094,N_6561,N_6635);
or U7095 (N_7095,N_6654,N_6509);
xor U7096 (N_7096,N_6727,N_6590);
or U7097 (N_7097,N_6698,N_6884);
xor U7098 (N_7098,N_6969,N_6715);
and U7099 (N_7099,N_6784,N_6985);
xor U7100 (N_7100,N_6630,N_6763);
nor U7101 (N_7101,N_6786,N_6889);
nor U7102 (N_7102,N_6993,N_6890);
nor U7103 (N_7103,N_6694,N_6792);
and U7104 (N_7104,N_6951,N_6871);
nor U7105 (N_7105,N_6788,N_6911);
xor U7106 (N_7106,N_6983,N_6947);
nor U7107 (N_7107,N_6785,N_6998);
or U7108 (N_7108,N_6957,N_6665);
xnor U7109 (N_7109,N_6582,N_6567);
xnor U7110 (N_7110,N_6879,N_6914);
or U7111 (N_7111,N_6564,N_6683);
nor U7112 (N_7112,N_6842,N_6661);
or U7113 (N_7113,N_6812,N_6650);
nand U7114 (N_7114,N_6897,N_6853);
nand U7115 (N_7115,N_6860,N_6502);
nand U7116 (N_7116,N_6739,N_6668);
xor U7117 (N_7117,N_6881,N_6705);
and U7118 (N_7118,N_6732,N_6566);
xnor U7119 (N_7119,N_6605,N_6647);
nand U7120 (N_7120,N_6893,N_6697);
xnor U7121 (N_7121,N_6525,N_6716);
nor U7122 (N_7122,N_6931,N_6803);
xor U7123 (N_7123,N_6615,N_6933);
nor U7124 (N_7124,N_6882,N_6932);
nand U7125 (N_7125,N_6934,N_6585);
or U7126 (N_7126,N_6634,N_6506);
or U7127 (N_7127,N_6659,N_6680);
and U7128 (N_7128,N_6913,N_6552);
and U7129 (N_7129,N_6943,N_6524);
xnor U7130 (N_7130,N_6908,N_6875);
nor U7131 (N_7131,N_6840,N_6749);
xnor U7132 (N_7132,N_6616,N_6618);
xnor U7133 (N_7133,N_6821,N_6623);
or U7134 (N_7134,N_6894,N_6789);
and U7135 (N_7135,N_6568,N_6930);
or U7136 (N_7136,N_6878,N_6731);
nand U7137 (N_7137,N_6844,N_6514);
and U7138 (N_7138,N_6636,N_6865);
nand U7139 (N_7139,N_6518,N_6563);
nor U7140 (N_7140,N_6670,N_6755);
nor U7141 (N_7141,N_6556,N_6920);
and U7142 (N_7142,N_6793,N_6909);
xor U7143 (N_7143,N_6695,N_6602);
nor U7144 (N_7144,N_6558,N_6808);
nor U7145 (N_7145,N_6662,N_6754);
nand U7146 (N_7146,N_6579,N_6707);
or U7147 (N_7147,N_6675,N_6644);
nor U7148 (N_7148,N_6572,N_6533);
xnor U7149 (N_7149,N_6629,N_6536);
or U7150 (N_7150,N_6977,N_6501);
xor U7151 (N_7151,N_6852,N_6584);
nor U7152 (N_7152,N_6899,N_6966);
and U7153 (N_7153,N_6586,N_6845);
and U7154 (N_7154,N_6721,N_6959);
and U7155 (N_7155,N_6888,N_6798);
xor U7156 (N_7156,N_6885,N_6970);
or U7157 (N_7157,N_6935,N_6686);
xnor U7158 (N_7158,N_6945,N_6902);
nor U7159 (N_7159,N_6676,N_6963);
nand U7160 (N_7160,N_6723,N_6895);
nor U7161 (N_7161,N_6863,N_6796);
nor U7162 (N_7162,N_6538,N_6652);
nand U7163 (N_7163,N_6551,N_6939);
and U7164 (N_7164,N_6520,N_6734);
and U7165 (N_7165,N_6746,N_6841);
and U7166 (N_7166,N_6526,N_6738);
nand U7167 (N_7167,N_6573,N_6814);
and U7168 (N_7168,N_6663,N_6641);
nor U7169 (N_7169,N_6703,N_6915);
xnor U7170 (N_7170,N_6700,N_6967);
or U7171 (N_7171,N_6539,N_6965);
nand U7172 (N_7172,N_6809,N_6917);
nor U7173 (N_7173,N_6958,N_6612);
nand U7174 (N_7174,N_6952,N_6790);
or U7175 (N_7175,N_6918,N_6571);
xnor U7176 (N_7176,N_6701,N_6938);
nor U7177 (N_7177,N_6687,N_6862);
or U7178 (N_7178,N_6973,N_6946);
and U7179 (N_7179,N_6542,N_6744);
or U7180 (N_7180,N_6531,N_6577);
and U7181 (N_7181,N_6516,N_6870);
or U7182 (N_7182,N_6926,N_6762);
or U7183 (N_7183,N_6989,N_6777);
nand U7184 (N_7184,N_6578,N_6975);
or U7185 (N_7185,N_6541,N_6991);
nor U7186 (N_7186,N_6581,N_6529);
nor U7187 (N_7187,N_6606,N_6910);
or U7188 (N_7188,N_6982,N_6580);
or U7189 (N_7189,N_6610,N_6591);
or U7190 (N_7190,N_6691,N_6519);
nand U7191 (N_7191,N_6950,N_6990);
nand U7192 (N_7192,N_6517,N_6741);
and U7193 (N_7193,N_6619,N_6795);
and U7194 (N_7194,N_6677,N_6867);
or U7195 (N_7195,N_6596,N_6690);
or U7196 (N_7196,N_6843,N_6869);
nand U7197 (N_7197,N_6624,N_6712);
or U7198 (N_7198,N_6877,N_6544);
xnor U7199 (N_7199,N_6835,N_6818);
nand U7200 (N_7200,N_6656,N_6759);
nor U7201 (N_7201,N_6827,N_6976);
or U7202 (N_7202,N_6626,N_6559);
and U7203 (N_7203,N_6637,N_6987);
or U7204 (N_7204,N_6658,N_6611);
or U7205 (N_7205,N_6537,N_6534);
xor U7206 (N_7206,N_6595,N_6988);
or U7207 (N_7207,N_6822,N_6617);
nand U7208 (N_7208,N_6671,N_6621);
nor U7209 (N_7209,N_6714,N_6956);
nor U7210 (N_7210,N_6961,N_6805);
nor U7211 (N_7211,N_6780,N_6924);
nand U7212 (N_7212,N_6511,N_6896);
or U7213 (N_7213,N_6857,N_6980);
or U7214 (N_7214,N_6936,N_6649);
nor U7215 (N_7215,N_6709,N_6807);
nand U7216 (N_7216,N_6575,N_6847);
nor U7217 (N_7217,N_6733,N_6745);
and U7218 (N_7218,N_6673,N_6799);
nand U7219 (N_7219,N_6589,N_6724);
nand U7220 (N_7220,N_6554,N_6891);
xnor U7221 (N_7221,N_6811,N_6725);
xnor U7222 (N_7222,N_6562,N_6669);
or U7223 (N_7223,N_6828,N_6766);
xor U7224 (N_7224,N_6778,N_6765);
or U7225 (N_7225,N_6901,N_6883);
nand U7226 (N_7226,N_6527,N_6859);
or U7227 (N_7227,N_6849,N_6735);
or U7228 (N_7228,N_6770,N_6838);
nand U7229 (N_7229,N_6549,N_6868);
and U7230 (N_7230,N_6856,N_6711);
xnor U7231 (N_7231,N_6850,N_6941);
nand U7232 (N_7232,N_6696,N_6995);
or U7233 (N_7233,N_6954,N_6628);
xnor U7234 (N_7234,N_6548,N_6781);
or U7235 (N_7235,N_6848,N_6643);
nand U7236 (N_7236,N_6583,N_6543);
nand U7237 (N_7237,N_6810,N_6638);
nand U7238 (N_7238,N_6574,N_6880);
nand U7239 (N_7239,N_6625,N_6771);
nand U7240 (N_7240,N_6986,N_6836);
xnor U7241 (N_7241,N_6772,N_6855);
or U7242 (N_7242,N_6831,N_6620);
and U7243 (N_7243,N_6645,N_6593);
nand U7244 (N_7244,N_6587,N_6704);
xor U7245 (N_7245,N_6846,N_6708);
nor U7246 (N_7246,N_6921,N_6802);
or U7247 (N_7247,N_6942,N_6713);
nor U7248 (N_7248,N_6560,N_6922);
nand U7249 (N_7249,N_6972,N_6751);
nor U7250 (N_7250,N_6921,N_6947);
nand U7251 (N_7251,N_6799,N_6560);
xor U7252 (N_7252,N_6809,N_6538);
nand U7253 (N_7253,N_6902,N_6761);
nor U7254 (N_7254,N_6577,N_6981);
or U7255 (N_7255,N_6983,N_6674);
or U7256 (N_7256,N_6939,N_6590);
nor U7257 (N_7257,N_6865,N_6649);
and U7258 (N_7258,N_6751,N_6670);
nor U7259 (N_7259,N_6850,N_6663);
xor U7260 (N_7260,N_6775,N_6813);
or U7261 (N_7261,N_6547,N_6714);
nand U7262 (N_7262,N_6555,N_6600);
xnor U7263 (N_7263,N_6736,N_6902);
nor U7264 (N_7264,N_6708,N_6762);
and U7265 (N_7265,N_6696,N_6566);
or U7266 (N_7266,N_6664,N_6841);
nand U7267 (N_7267,N_6724,N_6633);
nand U7268 (N_7268,N_6580,N_6911);
or U7269 (N_7269,N_6650,N_6915);
xnor U7270 (N_7270,N_6536,N_6610);
xor U7271 (N_7271,N_6542,N_6896);
or U7272 (N_7272,N_6592,N_6937);
nor U7273 (N_7273,N_6767,N_6688);
or U7274 (N_7274,N_6543,N_6747);
nor U7275 (N_7275,N_6535,N_6987);
xnor U7276 (N_7276,N_6789,N_6931);
or U7277 (N_7277,N_6796,N_6762);
or U7278 (N_7278,N_6564,N_6795);
nor U7279 (N_7279,N_6636,N_6875);
nor U7280 (N_7280,N_6615,N_6513);
and U7281 (N_7281,N_6558,N_6758);
or U7282 (N_7282,N_6895,N_6992);
xor U7283 (N_7283,N_6689,N_6870);
and U7284 (N_7284,N_6727,N_6532);
nor U7285 (N_7285,N_6559,N_6877);
nand U7286 (N_7286,N_6635,N_6535);
nand U7287 (N_7287,N_6721,N_6837);
or U7288 (N_7288,N_6956,N_6639);
or U7289 (N_7289,N_6975,N_6949);
nand U7290 (N_7290,N_6993,N_6749);
nand U7291 (N_7291,N_6668,N_6750);
xnor U7292 (N_7292,N_6802,N_6929);
nor U7293 (N_7293,N_6836,N_6525);
nand U7294 (N_7294,N_6507,N_6954);
xnor U7295 (N_7295,N_6770,N_6991);
and U7296 (N_7296,N_6794,N_6509);
nor U7297 (N_7297,N_6624,N_6830);
nand U7298 (N_7298,N_6828,N_6991);
or U7299 (N_7299,N_6918,N_6788);
or U7300 (N_7300,N_6758,N_6950);
and U7301 (N_7301,N_6672,N_6972);
or U7302 (N_7302,N_6685,N_6932);
nand U7303 (N_7303,N_6527,N_6913);
xor U7304 (N_7304,N_6623,N_6690);
xor U7305 (N_7305,N_6726,N_6695);
nand U7306 (N_7306,N_6861,N_6650);
xor U7307 (N_7307,N_6983,N_6707);
xor U7308 (N_7308,N_6918,N_6710);
xor U7309 (N_7309,N_6569,N_6886);
xnor U7310 (N_7310,N_6636,N_6515);
nor U7311 (N_7311,N_6734,N_6874);
nand U7312 (N_7312,N_6508,N_6671);
nor U7313 (N_7313,N_6961,N_6958);
nor U7314 (N_7314,N_6773,N_6871);
xnor U7315 (N_7315,N_6640,N_6760);
xnor U7316 (N_7316,N_6539,N_6611);
nor U7317 (N_7317,N_6874,N_6564);
xnor U7318 (N_7318,N_6784,N_6553);
or U7319 (N_7319,N_6613,N_6600);
nand U7320 (N_7320,N_6505,N_6920);
or U7321 (N_7321,N_6645,N_6866);
nand U7322 (N_7322,N_6982,N_6653);
xor U7323 (N_7323,N_6937,N_6824);
and U7324 (N_7324,N_6890,N_6846);
nand U7325 (N_7325,N_6652,N_6958);
or U7326 (N_7326,N_6850,N_6882);
and U7327 (N_7327,N_6568,N_6813);
nor U7328 (N_7328,N_6696,N_6919);
xor U7329 (N_7329,N_6605,N_6902);
and U7330 (N_7330,N_6701,N_6559);
nor U7331 (N_7331,N_6615,N_6596);
and U7332 (N_7332,N_6739,N_6908);
and U7333 (N_7333,N_6507,N_6641);
nor U7334 (N_7334,N_6772,N_6660);
or U7335 (N_7335,N_6736,N_6930);
and U7336 (N_7336,N_6560,N_6949);
and U7337 (N_7337,N_6764,N_6845);
xor U7338 (N_7338,N_6677,N_6900);
xor U7339 (N_7339,N_6840,N_6933);
nand U7340 (N_7340,N_6977,N_6730);
nand U7341 (N_7341,N_6648,N_6585);
xor U7342 (N_7342,N_6527,N_6808);
xnor U7343 (N_7343,N_6689,N_6604);
nor U7344 (N_7344,N_6895,N_6637);
or U7345 (N_7345,N_6953,N_6759);
nor U7346 (N_7346,N_6975,N_6913);
and U7347 (N_7347,N_6977,N_6651);
or U7348 (N_7348,N_6784,N_6825);
nor U7349 (N_7349,N_6670,N_6972);
or U7350 (N_7350,N_6753,N_6663);
nor U7351 (N_7351,N_6720,N_6515);
nand U7352 (N_7352,N_6513,N_6625);
nand U7353 (N_7353,N_6966,N_6667);
nand U7354 (N_7354,N_6903,N_6882);
nand U7355 (N_7355,N_6735,N_6689);
nand U7356 (N_7356,N_6714,N_6632);
or U7357 (N_7357,N_6655,N_6946);
nand U7358 (N_7358,N_6782,N_6881);
and U7359 (N_7359,N_6921,N_6948);
xor U7360 (N_7360,N_6904,N_6867);
nor U7361 (N_7361,N_6512,N_6582);
nand U7362 (N_7362,N_6852,N_6731);
nor U7363 (N_7363,N_6598,N_6506);
xor U7364 (N_7364,N_6798,N_6927);
nand U7365 (N_7365,N_6775,N_6719);
nand U7366 (N_7366,N_6703,N_6621);
or U7367 (N_7367,N_6797,N_6665);
nor U7368 (N_7368,N_6920,N_6543);
xnor U7369 (N_7369,N_6509,N_6893);
or U7370 (N_7370,N_6606,N_6974);
or U7371 (N_7371,N_6951,N_6674);
nor U7372 (N_7372,N_6574,N_6840);
and U7373 (N_7373,N_6716,N_6778);
xnor U7374 (N_7374,N_6846,N_6849);
or U7375 (N_7375,N_6716,N_6564);
nand U7376 (N_7376,N_6865,N_6666);
xor U7377 (N_7377,N_6541,N_6812);
or U7378 (N_7378,N_6693,N_6908);
xor U7379 (N_7379,N_6985,N_6514);
nand U7380 (N_7380,N_6694,N_6668);
nor U7381 (N_7381,N_6896,N_6675);
and U7382 (N_7382,N_6678,N_6651);
or U7383 (N_7383,N_6772,N_6853);
nor U7384 (N_7384,N_6746,N_6905);
nand U7385 (N_7385,N_6770,N_6643);
nand U7386 (N_7386,N_6751,N_6910);
or U7387 (N_7387,N_6547,N_6684);
xor U7388 (N_7388,N_6860,N_6707);
or U7389 (N_7389,N_6913,N_6634);
nand U7390 (N_7390,N_6656,N_6732);
xor U7391 (N_7391,N_6562,N_6871);
nand U7392 (N_7392,N_6648,N_6668);
nor U7393 (N_7393,N_6643,N_6750);
and U7394 (N_7394,N_6976,N_6993);
xor U7395 (N_7395,N_6616,N_6823);
or U7396 (N_7396,N_6687,N_6762);
xnor U7397 (N_7397,N_6547,N_6723);
nor U7398 (N_7398,N_6788,N_6754);
nand U7399 (N_7399,N_6984,N_6739);
nor U7400 (N_7400,N_6626,N_6709);
nor U7401 (N_7401,N_6885,N_6660);
or U7402 (N_7402,N_6952,N_6727);
xor U7403 (N_7403,N_6982,N_6913);
and U7404 (N_7404,N_6523,N_6775);
or U7405 (N_7405,N_6693,N_6607);
or U7406 (N_7406,N_6810,N_6911);
or U7407 (N_7407,N_6911,N_6922);
nor U7408 (N_7408,N_6677,N_6516);
and U7409 (N_7409,N_6585,N_6584);
and U7410 (N_7410,N_6657,N_6724);
and U7411 (N_7411,N_6658,N_6754);
xnor U7412 (N_7412,N_6837,N_6809);
nor U7413 (N_7413,N_6616,N_6607);
nand U7414 (N_7414,N_6667,N_6641);
nor U7415 (N_7415,N_6649,N_6709);
or U7416 (N_7416,N_6716,N_6827);
nor U7417 (N_7417,N_6848,N_6974);
nor U7418 (N_7418,N_6875,N_6715);
nor U7419 (N_7419,N_6661,N_6799);
nand U7420 (N_7420,N_6852,N_6683);
xor U7421 (N_7421,N_6892,N_6638);
or U7422 (N_7422,N_6977,N_6598);
nand U7423 (N_7423,N_6863,N_6598);
xnor U7424 (N_7424,N_6594,N_6514);
or U7425 (N_7425,N_6556,N_6568);
or U7426 (N_7426,N_6882,N_6560);
or U7427 (N_7427,N_6716,N_6622);
nand U7428 (N_7428,N_6591,N_6600);
and U7429 (N_7429,N_6576,N_6618);
and U7430 (N_7430,N_6937,N_6915);
xnor U7431 (N_7431,N_6850,N_6586);
and U7432 (N_7432,N_6534,N_6824);
xor U7433 (N_7433,N_6501,N_6770);
xnor U7434 (N_7434,N_6909,N_6512);
or U7435 (N_7435,N_6913,N_6795);
and U7436 (N_7436,N_6675,N_6965);
or U7437 (N_7437,N_6970,N_6851);
nand U7438 (N_7438,N_6951,N_6913);
nor U7439 (N_7439,N_6816,N_6658);
and U7440 (N_7440,N_6889,N_6823);
nor U7441 (N_7441,N_6910,N_6760);
xor U7442 (N_7442,N_6519,N_6958);
and U7443 (N_7443,N_6544,N_6601);
nor U7444 (N_7444,N_6991,N_6901);
xor U7445 (N_7445,N_6876,N_6543);
nand U7446 (N_7446,N_6880,N_6983);
or U7447 (N_7447,N_6682,N_6565);
or U7448 (N_7448,N_6655,N_6697);
or U7449 (N_7449,N_6682,N_6716);
xor U7450 (N_7450,N_6974,N_6617);
xnor U7451 (N_7451,N_6507,N_6854);
or U7452 (N_7452,N_6617,N_6611);
or U7453 (N_7453,N_6979,N_6852);
nor U7454 (N_7454,N_6879,N_6997);
xor U7455 (N_7455,N_6527,N_6738);
and U7456 (N_7456,N_6922,N_6598);
or U7457 (N_7457,N_6596,N_6849);
and U7458 (N_7458,N_6712,N_6538);
nor U7459 (N_7459,N_6933,N_6730);
and U7460 (N_7460,N_6911,N_6736);
or U7461 (N_7461,N_6918,N_6668);
nor U7462 (N_7462,N_6694,N_6717);
nand U7463 (N_7463,N_6588,N_6968);
xnor U7464 (N_7464,N_6985,N_6892);
nand U7465 (N_7465,N_6645,N_6898);
and U7466 (N_7466,N_6589,N_6736);
nor U7467 (N_7467,N_6774,N_6976);
or U7468 (N_7468,N_6634,N_6567);
xor U7469 (N_7469,N_6561,N_6968);
or U7470 (N_7470,N_6760,N_6604);
nor U7471 (N_7471,N_6587,N_6950);
or U7472 (N_7472,N_6674,N_6639);
or U7473 (N_7473,N_6899,N_6504);
or U7474 (N_7474,N_6823,N_6555);
nor U7475 (N_7475,N_6899,N_6821);
and U7476 (N_7476,N_6684,N_6567);
xor U7477 (N_7477,N_6591,N_6731);
and U7478 (N_7478,N_6747,N_6545);
and U7479 (N_7479,N_6799,N_6603);
xor U7480 (N_7480,N_6781,N_6530);
and U7481 (N_7481,N_6769,N_6848);
and U7482 (N_7482,N_6967,N_6669);
or U7483 (N_7483,N_6645,N_6622);
or U7484 (N_7484,N_6973,N_6725);
or U7485 (N_7485,N_6857,N_6960);
nor U7486 (N_7486,N_6806,N_6706);
xor U7487 (N_7487,N_6978,N_6857);
nor U7488 (N_7488,N_6521,N_6986);
or U7489 (N_7489,N_6543,N_6717);
xnor U7490 (N_7490,N_6836,N_6682);
xnor U7491 (N_7491,N_6793,N_6589);
nand U7492 (N_7492,N_6588,N_6858);
and U7493 (N_7493,N_6964,N_6680);
and U7494 (N_7494,N_6803,N_6955);
and U7495 (N_7495,N_6670,N_6760);
xor U7496 (N_7496,N_6953,N_6851);
nand U7497 (N_7497,N_6795,N_6657);
and U7498 (N_7498,N_6980,N_6569);
xor U7499 (N_7499,N_6703,N_6549);
nand U7500 (N_7500,N_7210,N_7022);
and U7501 (N_7501,N_7331,N_7252);
xor U7502 (N_7502,N_7434,N_7037);
and U7503 (N_7503,N_7380,N_7046);
xnor U7504 (N_7504,N_7276,N_7197);
nor U7505 (N_7505,N_7065,N_7288);
nand U7506 (N_7506,N_7034,N_7374);
nor U7507 (N_7507,N_7042,N_7077);
nand U7508 (N_7508,N_7397,N_7257);
xor U7509 (N_7509,N_7471,N_7137);
xnor U7510 (N_7510,N_7268,N_7202);
nor U7511 (N_7511,N_7057,N_7153);
and U7512 (N_7512,N_7053,N_7302);
and U7513 (N_7513,N_7320,N_7349);
or U7514 (N_7514,N_7182,N_7185);
xnor U7515 (N_7515,N_7047,N_7396);
and U7516 (N_7516,N_7300,N_7145);
nand U7517 (N_7517,N_7492,N_7128);
and U7518 (N_7518,N_7371,N_7081);
and U7519 (N_7519,N_7166,N_7376);
nor U7520 (N_7520,N_7438,N_7466);
nand U7521 (N_7521,N_7060,N_7458);
xor U7522 (N_7522,N_7385,N_7002);
and U7523 (N_7523,N_7196,N_7323);
or U7524 (N_7524,N_7248,N_7461);
and U7525 (N_7525,N_7398,N_7410);
nand U7526 (N_7526,N_7058,N_7220);
xnor U7527 (N_7527,N_7284,N_7488);
or U7528 (N_7528,N_7425,N_7119);
or U7529 (N_7529,N_7099,N_7489);
and U7530 (N_7530,N_7150,N_7225);
nand U7531 (N_7531,N_7351,N_7219);
xor U7532 (N_7532,N_7105,N_7129);
nand U7533 (N_7533,N_7122,N_7319);
and U7534 (N_7534,N_7352,N_7080);
nand U7535 (N_7535,N_7148,N_7406);
xnor U7536 (N_7536,N_7072,N_7340);
xnor U7537 (N_7537,N_7298,N_7023);
xor U7538 (N_7538,N_7010,N_7250);
nand U7539 (N_7539,N_7030,N_7031);
nand U7540 (N_7540,N_7305,N_7071);
and U7541 (N_7541,N_7278,N_7116);
nor U7542 (N_7542,N_7096,N_7452);
or U7543 (N_7543,N_7008,N_7270);
nor U7544 (N_7544,N_7063,N_7440);
or U7545 (N_7545,N_7241,N_7067);
nor U7546 (N_7546,N_7416,N_7100);
nand U7547 (N_7547,N_7372,N_7159);
nand U7548 (N_7548,N_7490,N_7136);
xor U7549 (N_7549,N_7226,N_7249);
or U7550 (N_7550,N_7429,N_7297);
and U7551 (N_7551,N_7135,N_7019);
or U7552 (N_7552,N_7259,N_7369);
and U7553 (N_7553,N_7269,N_7328);
xor U7554 (N_7554,N_7024,N_7256);
or U7555 (N_7555,N_7321,N_7164);
nor U7556 (N_7556,N_7357,N_7098);
nand U7557 (N_7557,N_7353,N_7485);
or U7558 (N_7558,N_7059,N_7222);
or U7559 (N_7559,N_7375,N_7232);
nor U7560 (N_7560,N_7127,N_7432);
nand U7561 (N_7561,N_7332,N_7187);
or U7562 (N_7562,N_7192,N_7223);
and U7563 (N_7563,N_7016,N_7462);
and U7564 (N_7564,N_7258,N_7117);
nand U7565 (N_7565,N_7061,N_7191);
nand U7566 (N_7566,N_7475,N_7444);
or U7567 (N_7567,N_7313,N_7048);
xor U7568 (N_7568,N_7303,N_7068);
or U7569 (N_7569,N_7402,N_7000);
nor U7570 (N_7570,N_7110,N_7275);
or U7571 (N_7571,N_7206,N_7230);
or U7572 (N_7572,N_7106,N_7170);
nor U7573 (N_7573,N_7162,N_7107);
xor U7574 (N_7574,N_7463,N_7428);
nor U7575 (N_7575,N_7295,N_7012);
and U7576 (N_7576,N_7384,N_7496);
nor U7577 (N_7577,N_7090,N_7464);
nor U7578 (N_7578,N_7198,N_7215);
nand U7579 (N_7579,N_7358,N_7377);
xor U7580 (N_7580,N_7188,N_7142);
and U7581 (N_7581,N_7325,N_7073);
nor U7582 (N_7582,N_7498,N_7004);
and U7583 (N_7583,N_7155,N_7407);
xor U7584 (N_7584,N_7238,N_7265);
nor U7585 (N_7585,N_7160,N_7460);
or U7586 (N_7586,N_7224,N_7163);
nor U7587 (N_7587,N_7382,N_7003);
xor U7588 (N_7588,N_7386,N_7263);
nand U7589 (N_7589,N_7472,N_7345);
nor U7590 (N_7590,N_7271,N_7218);
nand U7591 (N_7591,N_7495,N_7074);
nand U7592 (N_7592,N_7304,N_7337);
nand U7593 (N_7593,N_7028,N_7038);
nor U7594 (N_7594,N_7333,N_7070);
or U7595 (N_7595,N_7497,N_7367);
nor U7596 (N_7596,N_7242,N_7350);
nand U7597 (N_7597,N_7158,N_7040);
xor U7598 (N_7598,N_7180,N_7095);
and U7599 (N_7599,N_7126,N_7045);
xor U7600 (N_7600,N_7032,N_7368);
nand U7601 (N_7601,N_7113,N_7005);
or U7602 (N_7602,N_7186,N_7214);
xnor U7603 (N_7603,N_7262,N_7112);
or U7604 (N_7604,N_7413,N_7207);
nor U7605 (N_7605,N_7189,N_7433);
xnor U7606 (N_7606,N_7245,N_7317);
xnor U7607 (N_7607,N_7293,N_7181);
nor U7608 (N_7608,N_7283,N_7143);
xor U7609 (N_7609,N_7289,N_7013);
nor U7610 (N_7610,N_7007,N_7479);
xor U7611 (N_7611,N_7442,N_7450);
nand U7612 (N_7612,N_7322,N_7235);
or U7613 (N_7613,N_7287,N_7405);
nor U7614 (N_7614,N_7473,N_7393);
nor U7615 (N_7615,N_7394,N_7221);
nand U7616 (N_7616,N_7335,N_7430);
xor U7617 (N_7617,N_7216,N_7121);
xor U7618 (N_7618,N_7292,N_7446);
and U7619 (N_7619,N_7373,N_7193);
nand U7620 (N_7620,N_7360,N_7036);
or U7621 (N_7621,N_7194,N_7114);
or U7622 (N_7622,N_7228,N_7343);
nor U7623 (N_7623,N_7487,N_7029);
or U7624 (N_7624,N_7329,N_7138);
and U7625 (N_7625,N_7423,N_7139);
or U7626 (N_7626,N_7001,N_7173);
nand U7627 (N_7627,N_7195,N_7285);
xnor U7628 (N_7628,N_7379,N_7062);
nand U7629 (N_7629,N_7491,N_7154);
and U7630 (N_7630,N_7169,N_7212);
xor U7631 (N_7631,N_7172,N_7174);
or U7632 (N_7632,N_7441,N_7391);
or U7633 (N_7633,N_7456,N_7254);
nor U7634 (N_7634,N_7326,N_7033);
nand U7635 (N_7635,N_7403,N_7315);
and U7636 (N_7636,N_7086,N_7286);
nand U7637 (N_7637,N_7251,N_7338);
xnor U7638 (N_7638,N_7474,N_7296);
nor U7639 (N_7639,N_7205,N_7334);
and U7640 (N_7640,N_7015,N_7017);
nand U7641 (N_7641,N_7344,N_7267);
and U7642 (N_7642,N_7294,N_7299);
and U7643 (N_7643,N_7243,N_7209);
and U7644 (N_7644,N_7356,N_7097);
or U7645 (N_7645,N_7435,N_7177);
and U7646 (N_7646,N_7078,N_7408);
and U7647 (N_7647,N_7364,N_7347);
nor U7648 (N_7648,N_7484,N_7457);
nand U7649 (N_7649,N_7400,N_7124);
or U7650 (N_7650,N_7076,N_7167);
xnor U7651 (N_7651,N_7021,N_7176);
or U7652 (N_7652,N_7211,N_7156);
nor U7653 (N_7653,N_7476,N_7208);
nand U7654 (N_7654,N_7041,N_7079);
nand U7655 (N_7655,N_7141,N_7094);
xor U7656 (N_7656,N_7161,N_7201);
xor U7657 (N_7657,N_7436,N_7018);
and U7658 (N_7658,N_7200,N_7418);
or U7659 (N_7659,N_7327,N_7020);
or U7660 (N_7660,N_7417,N_7227);
and U7661 (N_7661,N_7363,N_7051);
nor U7662 (N_7662,N_7237,N_7101);
nor U7663 (N_7663,N_7125,N_7307);
nand U7664 (N_7664,N_7109,N_7027);
xor U7665 (N_7665,N_7451,N_7318);
nand U7666 (N_7666,N_7420,N_7240);
xnor U7667 (N_7667,N_7108,N_7316);
xor U7668 (N_7668,N_7151,N_7395);
nand U7669 (N_7669,N_7039,N_7431);
or U7670 (N_7670,N_7118,N_7467);
nor U7671 (N_7671,N_7272,N_7104);
and U7672 (N_7672,N_7115,N_7229);
nor U7673 (N_7673,N_7359,N_7389);
xor U7674 (N_7674,N_7260,N_7203);
xnor U7675 (N_7675,N_7341,N_7006);
nor U7676 (N_7676,N_7082,N_7244);
xor U7677 (N_7677,N_7330,N_7348);
nor U7678 (N_7678,N_7044,N_7165);
and U7679 (N_7679,N_7459,N_7277);
or U7680 (N_7680,N_7468,N_7054);
or U7681 (N_7681,N_7247,N_7049);
or U7682 (N_7682,N_7231,N_7093);
or U7683 (N_7683,N_7469,N_7362);
xor U7684 (N_7684,N_7217,N_7131);
xnor U7685 (N_7685,N_7253,N_7144);
xor U7686 (N_7686,N_7483,N_7411);
nand U7687 (N_7687,N_7306,N_7361);
or U7688 (N_7688,N_7422,N_7091);
nand U7689 (N_7689,N_7401,N_7453);
or U7690 (N_7690,N_7064,N_7087);
nand U7691 (N_7691,N_7449,N_7152);
or U7692 (N_7692,N_7239,N_7443);
nor U7693 (N_7693,N_7234,N_7454);
or U7694 (N_7694,N_7419,N_7482);
nor U7695 (N_7695,N_7404,N_7204);
xnor U7696 (N_7696,N_7480,N_7084);
nor U7697 (N_7697,N_7415,N_7183);
nand U7698 (N_7698,N_7346,N_7092);
xor U7699 (N_7699,N_7336,N_7056);
or U7700 (N_7700,N_7414,N_7448);
or U7701 (N_7701,N_7370,N_7310);
xnor U7702 (N_7702,N_7179,N_7261);
xnor U7703 (N_7703,N_7421,N_7133);
or U7704 (N_7704,N_7388,N_7255);
xnor U7705 (N_7705,N_7424,N_7168);
or U7706 (N_7706,N_7014,N_7111);
nor U7707 (N_7707,N_7069,N_7123);
xnor U7708 (N_7708,N_7387,N_7342);
nand U7709 (N_7709,N_7291,N_7146);
nand U7710 (N_7710,N_7383,N_7178);
and U7711 (N_7711,N_7282,N_7439);
nor U7712 (N_7712,N_7009,N_7365);
nand U7713 (N_7713,N_7290,N_7083);
nor U7714 (N_7714,N_7478,N_7399);
or U7715 (N_7715,N_7011,N_7309);
xnor U7716 (N_7716,N_7381,N_7266);
or U7717 (N_7717,N_7494,N_7426);
nand U7718 (N_7718,N_7311,N_7075);
or U7719 (N_7719,N_7190,N_7171);
and U7720 (N_7720,N_7412,N_7354);
or U7721 (N_7721,N_7455,N_7324);
xor U7722 (N_7722,N_7366,N_7312);
or U7723 (N_7723,N_7233,N_7066);
nand U7724 (N_7724,N_7273,N_7378);
xor U7725 (N_7725,N_7085,N_7103);
and U7726 (N_7726,N_7157,N_7493);
or U7727 (N_7727,N_7052,N_7055);
or U7728 (N_7728,N_7025,N_7314);
nor U7729 (N_7729,N_7140,N_7130);
and U7730 (N_7730,N_7089,N_7447);
nand U7731 (N_7731,N_7390,N_7409);
xor U7732 (N_7732,N_7213,N_7392);
nor U7733 (N_7733,N_7355,N_7050);
nor U7734 (N_7734,N_7246,N_7134);
nor U7735 (N_7735,N_7465,N_7026);
nor U7736 (N_7736,N_7486,N_7199);
nor U7737 (N_7737,N_7035,N_7427);
or U7738 (N_7738,N_7445,N_7102);
nor U7739 (N_7739,N_7280,N_7339);
or U7740 (N_7740,N_7437,N_7236);
and U7741 (N_7741,N_7149,N_7088);
xnor U7742 (N_7742,N_7132,N_7147);
nor U7743 (N_7743,N_7281,N_7120);
nand U7744 (N_7744,N_7477,N_7184);
nor U7745 (N_7745,N_7279,N_7308);
nor U7746 (N_7746,N_7274,N_7470);
nor U7747 (N_7747,N_7499,N_7481);
nand U7748 (N_7748,N_7264,N_7301);
xor U7749 (N_7749,N_7175,N_7043);
and U7750 (N_7750,N_7272,N_7473);
nand U7751 (N_7751,N_7014,N_7319);
nor U7752 (N_7752,N_7246,N_7042);
or U7753 (N_7753,N_7144,N_7210);
or U7754 (N_7754,N_7163,N_7477);
or U7755 (N_7755,N_7014,N_7210);
or U7756 (N_7756,N_7394,N_7488);
or U7757 (N_7757,N_7306,N_7054);
nor U7758 (N_7758,N_7473,N_7162);
or U7759 (N_7759,N_7104,N_7296);
nand U7760 (N_7760,N_7187,N_7009);
nor U7761 (N_7761,N_7352,N_7221);
nand U7762 (N_7762,N_7154,N_7339);
and U7763 (N_7763,N_7496,N_7032);
xnor U7764 (N_7764,N_7187,N_7434);
and U7765 (N_7765,N_7361,N_7458);
or U7766 (N_7766,N_7190,N_7428);
or U7767 (N_7767,N_7282,N_7228);
xnor U7768 (N_7768,N_7259,N_7426);
nor U7769 (N_7769,N_7239,N_7302);
nor U7770 (N_7770,N_7210,N_7046);
nand U7771 (N_7771,N_7439,N_7091);
and U7772 (N_7772,N_7058,N_7405);
and U7773 (N_7773,N_7419,N_7003);
and U7774 (N_7774,N_7473,N_7492);
or U7775 (N_7775,N_7066,N_7301);
xor U7776 (N_7776,N_7469,N_7489);
or U7777 (N_7777,N_7464,N_7365);
nand U7778 (N_7778,N_7017,N_7330);
xor U7779 (N_7779,N_7472,N_7004);
or U7780 (N_7780,N_7137,N_7377);
nand U7781 (N_7781,N_7277,N_7411);
and U7782 (N_7782,N_7353,N_7379);
and U7783 (N_7783,N_7142,N_7197);
and U7784 (N_7784,N_7393,N_7172);
xor U7785 (N_7785,N_7057,N_7159);
and U7786 (N_7786,N_7092,N_7043);
or U7787 (N_7787,N_7094,N_7308);
and U7788 (N_7788,N_7008,N_7467);
or U7789 (N_7789,N_7116,N_7215);
nor U7790 (N_7790,N_7195,N_7133);
xor U7791 (N_7791,N_7314,N_7499);
and U7792 (N_7792,N_7470,N_7171);
nand U7793 (N_7793,N_7026,N_7283);
nand U7794 (N_7794,N_7354,N_7228);
or U7795 (N_7795,N_7176,N_7402);
nor U7796 (N_7796,N_7333,N_7392);
xor U7797 (N_7797,N_7393,N_7222);
nor U7798 (N_7798,N_7340,N_7286);
nand U7799 (N_7799,N_7361,N_7003);
nor U7800 (N_7800,N_7111,N_7138);
xnor U7801 (N_7801,N_7242,N_7052);
xnor U7802 (N_7802,N_7478,N_7028);
xor U7803 (N_7803,N_7388,N_7386);
xnor U7804 (N_7804,N_7411,N_7145);
or U7805 (N_7805,N_7304,N_7119);
nand U7806 (N_7806,N_7072,N_7239);
nor U7807 (N_7807,N_7003,N_7466);
xor U7808 (N_7808,N_7344,N_7345);
nor U7809 (N_7809,N_7359,N_7204);
nand U7810 (N_7810,N_7420,N_7353);
nand U7811 (N_7811,N_7063,N_7047);
and U7812 (N_7812,N_7335,N_7447);
or U7813 (N_7813,N_7108,N_7219);
xor U7814 (N_7814,N_7226,N_7386);
xnor U7815 (N_7815,N_7138,N_7411);
and U7816 (N_7816,N_7132,N_7118);
and U7817 (N_7817,N_7338,N_7455);
or U7818 (N_7818,N_7082,N_7296);
and U7819 (N_7819,N_7421,N_7461);
and U7820 (N_7820,N_7187,N_7239);
nand U7821 (N_7821,N_7257,N_7199);
or U7822 (N_7822,N_7019,N_7119);
and U7823 (N_7823,N_7371,N_7451);
or U7824 (N_7824,N_7215,N_7253);
nor U7825 (N_7825,N_7214,N_7410);
xor U7826 (N_7826,N_7340,N_7276);
nand U7827 (N_7827,N_7135,N_7496);
nor U7828 (N_7828,N_7344,N_7178);
nor U7829 (N_7829,N_7189,N_7256);
nor U7830 (N_7830,N_7346,N_7449);
nor U7831 (N_7831,N_7147,N_7061);
xnor U7832 (N_7832,N_7047,N_7190);
and U7833 (N_7833,N_7073,N_7013);
nor U7834 (N_7834,N_7182,N_7359);
and U7835 (N_7835,N_7443,N_7238);
nand U7836 (N_7836,N_7095,N_7387);
xor U7837 (N_7837,N_7075,N_7037);
xnor U7838 (N_7838,N_7028,N_7330);
xor U7839 (N_7839,N_7367,N_7334);
nor U7840 (N_7840,N_7303,N_7079);
and U7841 (N_7841,N_7356,N_7412);
nor U7842 (N_7842,N_7427,N_7009);
and U7843 (N_7843,N_7064,N_7436);
nand U7844 (N_7844,N_7077,N_7332);
and U7845 (N_7845,N_7091,N_7133);
nor U7846 (N_7846,N_7410,N_7258);
and U7847 (N_7847,N_7340,N_7386);
and U7848 (N_7848,N_7283,N_7185);
or U7849 (N_7849,N_7120,N_7354);
and U7850 (N_7850,N_7110,N_7109);
xnor U7851 (N_7851,N_7308,N_7046);
and U7852 (N_7852,N_7213,N_7075);
and U7853 (N_7853,N_7468,N_7147);
nand U7854 (N_7854,N_7160,N_7216);
nor U7855 (N_7855,N_7346,N_7438);
or U7856 (N_7856,N_7417,N_7060);
nand U7857 (N_7857,N_7010,N_7153);
or U7858 (N_7858,N_7277,N_7339);
xor U7859 (N_7859,N_7168,N_7196);
xor U7860 (N_7860,N_7477,N_7128);
xor U7861 (N_7861,N_7292,N_7189);
or U7862 (N_7862,N_7004,N_7478);
xor U7863 (N_7863,N_7408,N_7276);
nor U7864 (N_7864,N_7035,N_7026);
and U7865 (N_7865,N_7059,N_7094);
and U7866 (N_7866,N_7058,N_7226);
xor U7867 (N_7867,N_7297,N_7085);
nand U7868 (N_7868,N_7194,N_7059);
nor U7869 (N_7869,N_7133,N_7422);
and U7870 (N_7870,N_7340,N_7052);
and U7871 (N_7871,N_7340,N_7217);
and U7872 (N_7872,N_7244,N_7422);
nor U7873 (N_7873,N_7132,N_7104);
and U7874 (N_7874,N_7402,N_7034);
or U7875 (N_7875,N_7229,N_7027);
xor U7876 (N_7876,N_7200,N_7455);
nand U7877 (N_7877,N_7225,N_7097);
xor U7878 (N_7878,N_7168,N_7023);
or U7879 (N_7879,N_7115,N_7143);
and U7880 (N_7880,N_7456,N_7063);
nand U7881 (N_7881,N_7357,N_7492);
and U7882 (N_7882,N_7439,N_7131);
and U7883 (N_7883,N_7066,N_7123);
and U7884 (N_7884,N_7163,N_7152);
nor U7885 (N_7885,N_7368,N_7120);
or U7886 (N_7886,N_7390,N_7074);
or U7887 (N_7887,N_7202,N_7366);
nand U7888 (N_7888,N_7483,N_7326);
and U7889 (N_7889,N_7050,N_7201);
and U7890 (N_7890,N_7167,N_7202);
xor U7891 (N_7891,N_7257,N_7297);
nor U7892 (N_7892,N_7329,N_7334);
nor U7893 (N_7893,N_7367,N_7382);
nand U7894 (N_7894,N_7379,N_7329);
nand U7895 (N_7895,N_7053,N_7108);
or U7896 (N_7896,N_7172,N_7186);
xor U7897 (N_7897,N_7437,N_7483);
nand U7898 (N_7898,N_7407,N_7018);
and U7899 (N_7899,N_7138,N_7110);
xnor U7900 (N_7900,N_7332,N_7248);
nor U7901 (N_7901,N_7396,N_7191);
nand U7902 (N_7902,N_7318,N_7400);
xor U7903 (N_7903,N_7072,N_7379);
and U7904 (N_7904,N_7482,N_7209);
xnor U7905 (N_7905,N_7332,N_7345);
and U7906 (N_7906,N_7275,N_7238);
or U7907 (N_7907,N_7493,N_7005);
nand U7908 (N_7908,N_7137,N_7023);
nand U7909 (N_7909,N_7104,N_7437);
or U7910 (N_7910,N_7201,N_7213);
nor U7911 (N_7911,N_7172,N_7198);
or U7912 (N_7912,N_7128,N_7265);
nor U7913 (N_7913,N_7475,N_7235);
nor U7914 (N_7914,N_7421,N_7485);
nor U7915 (N_7915,N_7086,N_7109);
or U7916 (N_7916,N_7064,N_7491);
nor U7917 (N_7917,N_7460,N_7161);
nand U7918 (N_7918,N_7233,N_7477);
and U7919 (N_7919,N_7419,N_7332);
xnor U7920 (N_7920,N_7467,N_7212);
or U7921 (N_7921,N_7194,N_7489);
nor U7922 (N_7922,N_7218,N_7208);
or U7923 (N_7923,N_7395,N_7193);
nand U7924 (N_7924,N_7484,N_7489);
nor U7925 (N_7925,N_7399,N_7425);
and U7926 (N_7926,N_7417,N_7189);
nor U7927 (N_7927,N_7263,N_7027);
xnor U7928 (N_7928,N_7364,N_7172);
xor U7929 (N_7929,N_7258,N_7103);
xor U7930 (N_7930,N_7235,N_7082);
nor U7931 (N_7931,N_7163,N_7354);
or U7932 (N_7932,N_7104,N_7110);
nand U7933 (N_7933,N_7156,N_7185);
xor U7934 (N_7934,N_7452,N_7040);
nand U7935 (N_7935,N_7420,N_7215);
and U7936 (N_7936,N_7174,N_7187);
nor U7937 (N_7937,N_7270,N_7101);
nor U7938 (N_7938,N_7103,N_7267);
or U7939 (N_7939,N_7369,N_7456);
nand U7940 (N_7940,N_7388,N_7028);
or U7941 (N_7941,N_7192,N_7224);
xnor U7942 (N_7942,N_7498,N_7207);
and U7943 (N_7943,N_7483,N_7098);
or U7944 (N_7944,N_7081,N_7312);
xor U7945 (N_7945,N_7420,N_7308);
or U7946 (N_7946,N_7066,N_7444);
xor U7947 (N_7947,N_7378,N_7287);
xnor U7948 (N_7948,N_7326,N_7476);
nor U7949 (N_7949,N_7334,N_7121);
nand U7950 (N_7950,N_7363,N_7402);
xnor U7951 (N_7951,N_7444,N_7495);
xnor U7952 (N_7952,N_7369,N_7134);
or U7953 (N_7953,N_7213,N_7450);
or U7954 (N_7954,N_7205,N_7231);
nor U7955 (N_7955,N_7037,N_7017);
nor U7956 (N_7956,N_7151,N_7074);
nor U7957 (N_7957,N_7480,N_7066);
or U7958 (N_7958,N_7165,N_7086);
and U7959 (N_7959,N_7207,N_7217);
nand U7960 (N_7960,N_7239,N_7154);
and U7961 (N_7961,N_7130,N_7237);
and U7962 (N_7962,N_7174,N_7254);
xnor U7963 (N_7963,N_7366,N_7399);
and U7964 (N_7964,N_7040,N_7134);
or U7965 (N_7965,N_7306,N_7087);
or U7966 (N_7966,N_7197,N_7023);
nand U7967 (N_7967,N_7151,N_7202);
and U7968 (N_7968,N_7340,N_7371);
nor U7969 (N_7969,N_7239,N_7406);
or U7970 (N_7970,N_7413,N_7286);
nand U7971 (N_7971,N_7288,N_7003);
nand U7972 (N_7972,N_7464,N_7070);
and U7973 (N_7973,N_7097,N_7042);
nor U7974 (N_7974,N_7028,N_7440);
nand U7975 (N_7975,N_7262,N_7186);
and U7976 (N_7976,N_7284,N_7085);
nor U7977 (N_7977,N_7229,N_7452);
or U7978 (N_7978,N_7428,N_7182);
and U7979 (N_7979,N_7190,N_7013);
and U7980 (N_7980,N_7312,N_7076);
xor U7981 (N_7981,N_7136,N_7183);
or U7982 (N_7982,N_7269,N_7031);
nand U7983 (N_7983,N_7095,N_7328);
nand U7984 (N_7984,N_7495,N_7442);
xor U7985 (N_7985,N_7126,N_7453);
xor U7986 (N_7986,N_7371,N_7452);
or U7987 (N_7987,N_7119,N_7105);
nor U7988 (N_7988,N_7017,N_7217);
and U7989 (N_7989,N_7399,N_7450);
and U7990 (N_7990,N_7397,N_7410);
nor U7991 (N_7991,N_7196,N_7473);
or U7992 (N_7992,N_7430,N_7214);
nand U7993 (N_7993,N_7285,N_7283);
nand U7994 (N_7994,N_7282,N_7163);
nand U7995 (N_7995,N_7331,N_7061);
or U7996 (N_7996,N_7296,N_7425);
nor U7997 (N_7997,N_7374,N_7047);
xor U7998 (N_7998,N_7387,N_7186);
nand U7999 (N_7999,N_7161,N_7065);
xnor U8000 (N_8000,N_7530,N_7656);
or U8001 (N_8001,N_7519,N_7978);
xnor U8002 (N_8002,N_7990,N_7674);
nand U8003 (N_8003,N_7755,N_7665);
xor U8004 (N_8004,N_7794,N_7948);
nand U8005 (N_8005,N_7911,N_7883);
or U8006 (N_8006,N_7657,N_7541);
nand U8007 (N_8007,N_7787,N_7810);
xor U8008 (N_8008,N_7969,N_7870);
or U8009 (N_8009,N_7539,N_7570);
nand U8010 (N_8010,N_7563,N_7798);
and U8011 (N_8011,N_7716,N_7630);
nand U8012 (N_8012,N_7724,N_7583);
or U8013 (N_8013,N_7981,N_7825);
nor U8014 (N_8014,N_7706,N_7954);
nor U8015 (N_8015,N_7604,N_7664);
nand U8016 (N_8016,N_7722,N_7717);
and U8017 (N_8017,N_7641,N_7997);
nor U8018 (N_8018,N_7579,N_7844);
or U8019 (N_8019,N_7565,N_7955);
or U8020 (N_8020,N_7538,N_7669);
nand U8021 (N_8021,N_7741,N_7915);
and U8022 (N_8022,N_7984,N_7584);
nand U8023 (N_8023,N_7805,N_7887);
nand U8024 (N_8024,N_7617,N_7876);
or U8025 (N_8025,N_7660,N_7698);
and U8026 (N_8026,N_7725,N_7838);
or U8027 (N_8027,N_7742,N_7675);
nor U8028 (N_8028,N_7754,N_7983);
nor U8029 (N_8029,N_7547,N_7644);
or U8030 (N_8030,N_7551,N_7543);
and U8031 (N_8031,N_7513,N_7816);
or U8032 (N_8032,N_7790,N_7917);
xnor U8033 (N_8033,N_7612,N_7671);
xnor U8034 (N_8034,N_7756,N_7763);
nor U8035 (N_8035,N_7855,N_7828);
and U8036 (N_8036,N_7836,N_7931);
or U8037 (N_8037,N_7616,N_7945);
nor U8038 (N_8038,N_7542,N_7628);
and U8039 (N_8039,N_7764,N_7893);
nand U8040 (N_8040,N_7729,N_7767);
or U8041 (N_8041,N_7700,N_7517);
nand U8042 (N_8042,N_7928,N_7834);
nand U8043 (N_8043,N_7822,N_7553);
nor U8044 (N_8044,N_7548,N_7976);
or U8045 (N_8045,N_7869,N_7625);
nor U8046 (N_8046,N_7898,N_7765);
and U8047 (N_8047,N_7562,N_7919);
nand U8048 (N_8048,N_7676,N_7649);
and U8049 (N_8049,N_7932,N_7780);
xor U8050 (N_8050,N_7685,N_7505);
and U8051 (N_8051,N_7621,N_7620);
nor U8052 (N_8052,N_7958,N_7723);
nor U8053 (N_8053,N_7515,N_7732);
nor U8054 (N_8054,N_7710,N_7652);
xor U8055 (N_8055,N_7874,N_7827);
nor U8056 (N_8056,N_7709,N_7786);
nand U8057 (N_8057,N_7529,N_7525);
xor U8058 (N_8058,N_7602,N_7615);
and U8059 (N_8059,N_7566,N_7956);
xnor U8060 (N_8060,N_7728,N_7559);
nor U8061 (N_8061,N_7689,N_7719);
and U8062 (N_8062,N_7618,N_7885);
or U8063 (N_8063,N_7904,N_7776);
nor U8064 (N_8064,N_7532,N_7992);
or U8065 (N_8065,N_7801,N_7534);
or U8066 (N_8066,N_7711,N_7817);
xor U8067 (N_8067,N_7878,N_7820);
or U8068 (N_8068,N_7629,N_7961);
nor U8069 (N_8069,N_7858,N_7989);
nor U8070 (N_8070,N_7731,N_7987);
or U8071 (N_8071,N_7707,N_7662);
and U8072 (N_8072,N_7651,N_7939);
or U8073 (N_8073,N_7909,N_7753);
nor U8074 (N_8074,N_7688,N_7906);
nor U8075 (N_8075,N_7704,N_7854);
xnor U8076 (N_8076,N_7596,N_7933);
xor U8077 (N_8077,N_7937,N_7952);
nand U8078 (N_8078,N_7872,N_7973);
xnor U8079 (N_8079,N_7891,N_7775);
and U8080 (N_8080,N_7504,N_7666);
nor U8081 (N_8081,N_7789,N_7899);
nand U8082 (N_8082,N_7727,N_7781);
xnor U8083 (N_8083,N_7924,N_7636);
nor U8084 (N_8084,N_7808,N_7800);
nor U8085 (N_8085,N_7545,N_7622);
nand U8086 (N_8086,N_7582,N_7569);
nor U8087 (N_8087,N_7748,N_7733);
or U8088 (N_8088,N_7726,N_7892);
or U8089 (N_8089,N_7735,N_7634);
nor U8090 (N_8090,N_7848,N_7577);
and U8091 (N_8091,N_7925,N_7920);
and U8092 (N_8092,N_7561,N_7743);
nand U8093 (N_8093,N_7701,N_7610);
nor U8094 (N_8094,N_7777,N_7687);
nand U8095 (N_8095,N_7575,N_7979);
nand U8096 (N_8096,N_7739,N_7645);
nor U8097 (N_8097,N_7960,N_7560);
nor U8098 (N_8098,N_7703,N_7771);
and U8099 (N_8099,N_7690,N_7884);
nor U8100 (N_8100,N_7788,N_7850);
and U8101 (N_8101,N_7684,N_7982);
and U8102 (N_8102,N_7528,N_7957);
nand U8103 (N_8103,N_7994,N_7962);
xor U8104 (N_8104,N_7877,N_7988);
and U8105 (N_8105,N_7804,N_7890);
and U8106 (N_8106,N_7867,N_7943);
nor U8107 (N_8107,N_7557,N_7766);
or U8108 (N_8108,N_7695,N_7968);
or U8109 (N_8109,N_7759,N_7832);
nand U8110 (N_8110,N_7736,N_7809);
xnor U8111 (N_8111,N_7694,N_7847);
or U8112 (N_8112,N_7587,N_7871);
and U8113 (N_8113,N_7679,N_7910);
nor U8114 (N_8114,N_7738,N_7894);
and U8115 (N_8115,N_7993,N_7552);
nor U8116 (N_8116,N_7995,N_7571);
or U8117 (N_8117,N_7998,N_7807);
or U8118 (N_8118,N_7830,N_7673);
or U8119 (N_8119,N_7901,N_7715);
nand U8120 (N_8120,N_7923,N_7974);
or U8121 (N_8121,N_7692,N_7813);
or U8122 (N_8122,N_7837,N_7599);
nand U8123 (N_8123,N_7677,N_7845);
nor U8124 (N_8124,N_7773,N_7611);
xnor U8125 (N_8125,N_7510,N_7812);
nor U8126 (N_8126,N_7918,N_7768);
nand U8127 (N_8127,N_7799,N_7903);
xnor U8128 (N_8128,N_7966,N_7908);
nand U8129 (N_8129,N_7506,N_7900);
nor U8130 (N_8130,N_7654,N_7934);
xnor U8131 (N_8131,N_7600,N_7856);
xnor U8132 (N_8132,N_7581,N_7550);
nand U8133 (N_8133,N_7949,N_7970);
or U8134 (N_8134,N_7627,N_7824);
xor U8135 (N_8135,N_7971,N_7686);
and U8136 (N_8136,N_7697,N_7886);
nor U8137 (N_8137,N_7866,N_7792);
and U8138 (N_8138,N_7947,N_7926);
nor U8139 (N_8139,N_7522,N_7638);
nor U8140 (N_8140,N_7626,N_7624);
and U8141 (N_8141,N_7940,N_7589);
nor U8142 (N_8142,N_7914,N_7784);
and U8143 (N_8143,N_7929,N_7942);
or U8144 (N_8144,N_7986,N_7556);
nand U8145 (N_8145,N_7647,N_7520);
nand U8146 (N_8146,N_7500,N_7721);
nand U8147 (N_8147,N_7774,N_7831);
nand U8148 (N_8148,N_7533,N_7803);
nand U8149 (N_8149,N_7922,N_7779);
and U8150 (N_8150,N_7950,N_7859);
or U8151 (N_8151,N_7758,N_7916);
nor U8152 (N_8152,N_7796,N_7718);
and U8153 (N_8153,N_7623,N_7594);
and U8154 (N_8154,N_7588,N_7591);
xnor U8155 (N_8155,N_7509,N_7637);
nand U8156 (N_8156,N_7632,N_7605);
and U8157 (N_8157,N_7964,N_7935);
nor U8158 (N_8158,N_7558,N_7860);
and U8159 (N_8159,N_7702,N_7699);
and U8160 (N_8160,N_7875,N_7593);
nand U8161 (N_8161,N_7567,N_7770);
and U8162 (N_8162,N_7667,N_7842);
xnor U8163 (N_8163,N_7586,N_7905);
or U8164 (N_8164,N_7524,N_7639);
or U8165 (N_8165,N_7888,N_7846);
nand U8166 (N_8166,N_7833,N_7633);
or U8167 (N_8167,N_7503,N_7572);
and U8168 (N_8168,N_7857,N_7554);
and U8169 (N_8169,N_7841,N_7744);
nand U8170 (N_8170,N_7714,N_7585);
nand U8171 (N_8171,N_7720,N_7868);
xor U8172 (N_8172,N_7745,N_7913);
or U8173 (N_8173,N_7889,N_7646);
nor U8174 (N_8174,N_7555,N_7653);
or U8175 (N_8175,N_7549,N_7705);
xor U8176 (N_8176,N_7516,N_7682);
xnor U8177 (N_8177,N_7752,N_7546);
and U8178 (N_8178,N_7712,N_7791);
xnor U8179 (N_8179,N_7861,N_7873);
or U8180 (N_8180,N_7769,N_7648);
or U8181 (N_8181,N_7762,N_7749);
and U8182 (N_8182,N_7501,N_7897);
nor U8183 (N_8183,N_7521,N_7595);
xor U8184 (N_8184,N_7696,N_7607);
and U8185 (N_8185,N_7921,N_7863);
or U8186 (N_8186,N_7975,N_7977);
nor U8187 (N_8187,N_7938,N_7750);
and U8188 (N_8188,N_7761,N_7614);
or U8189 (N_8189,N_7640,N_7881);
nand U8190 (N_8190,N_7663,N_7751);
nor U8191 (N_8191,N_7912,N_7965);
nand U8192 (N_8192,N_7806,N_7793);
nor U8193 (N_8193,N_7659,N_7760);
and U8194 (N_8194,N_7502,N_7598);
xnor U8195 (N_8195,N_7568,N_7693);
xnor U8196 (N_8196,N_7544,N_7980);
and U8197 (N_8197,N_7609,N_7590);
or U8198 (N_8198,N_7658,N_7747);
and U8199 (N_8199,N_7523,N_7597);
nor U8200 (N_8200,N_7999,N_7811);
nand U8201 (N_8201,N_7592,N_7650);
nor U8202 (N_8202,N_7681,N_7996);
and U8203 (N_8203,N_7951,N_7536);
nor U8204 (N_8204,N_7511,N_7852);
or U8205 (N_8205,N_7691,N_7815);
nand U8206 (N_8206,N_7907,N_7531);
nand U8207 (N_8207,N_7672,N_7851);
nand U8208 (N_8208,N_7527,N_7655);
and U8209 (N_8209,N_7514,N_7613);
or U8210 (N_8210,N_7835,N_7826);
nor U8211 (N_8211,N_7829,N_7576);
nor U8212 (N_8212,N_7606,N_7713);
xnor U8213 (N_8213,N_7865,N_7927);
and U8214 (N_8214,N_7631,N_7839);
and U8215 (N_8215,N_7708,N_7535);
xnor U8216 (N_8216,N_7730,N_7772);
xor U8217 (N_8217,N_7507,N_7608);
nor U8218 (N_8218,N_7896,N_7963);
xnor U8219 (N_8219,N_7864,N_7953);
xor U8220 (N_8220,N_7619,N_7814);
xor U8221 (N_8221,N_7819,N_7526);
xnor U8222 (N_8222,N_7740,N_7785);
nand U8223 (N_8223,N_7853,N_7985);
nor U8224 (N_8224,N_7840,N_7518);
nand U8225 (N_8225,N_7642,N_7967);
and U8226 (N_8226,N_7823,N_7678);
nor U8227 (N_8227,N_7930,N_7778);
xor U8228 (N_8228,N_7578,N_7797);
nand U8229 (N_8229,N_7540,N_7783);
and U8230 (N_8230,N_7802,N_7895);
or U8231 (N_8231,N_7734,N_7941);
or U8232 (N_8232,N_7564,N_7821);
nor U8233 (N_8233,N_7879,N_7580);
xor U8234 (N_8234,N_7661,N_7959);
and U8235 (N_8235,N_7603,N_7635);
or U8236 (N_8236,N_7880,N_7573);
nand U8237 (N_8237,N_7795,N_7670);
or U8238 (N_8238,N_7601,N_7643);
or U8239 (N_8239,N_7944,N_7680);
xor U8240 (N_8240,N_7757,N_7849);
and U8241 (N_8241,N_7668,N_7936);
or U8242 (N_8242,N_7737,N_7972);
xnor U8243 (N_8243,N_7782,N_7902);
xor U8244 (N_8244,N_7882,N_7508);
xnor U8245 (N_8245,N_7862,N_7683);
nand U8246 (N_8246,N_7574,N_7818);
nand U8247 (N_8247,N_7512,N_7843);
nor U8248 (N_8248,N_7946,N_7746);
nand U8249 (N_8249,N_7537,N_7991);
xor U8250 (N_8250,N_7631,N_7504);
xor U8251 (N_8251,N_7848,N_7777);
nor U8252 (N_8252,N_7771,N_7592);
nor U8253 (N_8253,N_7981,N_7840);
and U8254 (N_8254,N_7689,N_7771);
and U8255 (N_8255,N_7528,N_7856);
xor U8256 (N_8256,N_7785,N_7828);
nor U8257 (N_8257,N_7503,N_7702);
or U8258 (N_8258,N_7584,N_7770);
and U8259 (N_8259,N_7713,N_7907);
and U8260 (N_8260,N_7891,N_7573);
and U8261 (N_8261,N_7996,N_7800);
nor U8262 (N_8262,N_7819,N_7624);
and U8263 (N_8263,N_7671,N_7866);
or U8264 (N_8264,N_7592,N_7781);
nor U8265 (N_8265,N_7877,N_7868);
nor U8266 (N_8266,N_7998,N_7726);
and U8267 (N_8267,N_7723,N_7500);
xnor U8268 (N_8268,N_7641,N_7998);
or U8269 (N_8269,N_7632,N_7976);
or U8270 (N_8270,N_7934,N_7793);
nand U8271 (N_8271,N_7597,N_7792);
xor U8272 (N_8272,N_7916,N_7859);
or U8273 (N_8273,N_7700,N_7705);
or U8274 (N_8274,N_7916,N_7938);
xor U8275 (N_8275,N_7610,N_7532);
xnor U8276 (N_8276,N_7642,N_7658);
nor U8277 (N_8277,N_7894,N_7817);
nand U8278 (N_8278,N_7795,N_7885);
nand U8279 (N_8279,N_7842,N_7711);
xnor U8280 (N_8280,N_7741,N_7547);
and U8281 (N_8281,N_7838,N_7877);
xnor U8282 (N_8282,N_7789,N_7748);
nand U8283 (N_8283,N_7835,N_7611);
and U8284 (N_8284,N_7772,N_7852);
nor U8285 (N_8285,N_7972,N_7967);
and U8286 (N_8286,N_7908,N_7729);
nand U8287 (N_8287,N_7744,N_7896);
or U8288 (N_8288,N_7772,N_7879);
nand U8289 (N_8289,N_7508,N_7884);
nand U8290 (N_8290,N_7519,N_7571);
nor U8291 (N_8291,N_7868,N_7693);
nor U8292 (N_8292,N_7633,N_7664);
nand U8293 (N_8293,N_7819,N_7885);
nor U8294 (N_8294,N_7864,N_7704);
or U8295 (N_8295,N_7782,N_7628);
xnor U8296 (N_8296,N_7591,N_7989);
or U8297 (N_8297,N_7767,N_7726);
nor U8298 (N_8298,N_7552,N_7955);
nor U8299 (N_8299,N_7827,N_7694);
or U8300 (N_8300,N_7825,N_7702);
nor U8301 (N_8301,N_7711,N_7862);
and U8302 (N_8302,N_7595,N_7571);
and U8303 (N_8303,N_7706,N_7633);
nor U8304 (N_8304,N_7858,N_7818);
and U8305 (N_8305,N_7670,N_7514);
xor U8306 (N_8306,N_7574,N_7715);
or U8307 (N_8307,N_7963,N_7664);
and U8308 (N_8308,N_7780,N_7568);
nand U8309 (N_8309,N_7929,N_7638);
and U8310 (N_8310,N_7935,N_7773);
xor U8311 (N_8311,N_7756,N_7710);
or U8312 (N_8312,N_7540,N_7775);
and U8313 (N_8313,N_7852,N_7700);
xor U8314 (N_8314,N_7768,N_7831);
nand U8315 (N_8315,N_7714,N_7875);
and U8316 (N_8316,N_7932,N_7740);
and U8317 (N_8317,N_7873,N_7927);
or U8318 (N_8318,N_7519,N_7530);
nor U8319 (N_8319,N_7681,N_7677);
or U8320 (N_8320,N_7923,N_7798);
nor U8321 (N_8321,N_7877,N_7735);
or U8322 (N_8322,N_7528,N_7803);
xnor U8323 (N_8323,N_7735,N_7934);
or U8324 (N_8324,N_7535,N_7761);
xor U8325 (N_8325,N_7814,N_7579);
xor U8326 (N_8326,N_7785,N_7651);
or U8327 (N_8327,N_7888,N_7620);
or U8328 (N_8328,N_7997,N_7789);
nor U8329 (N_8329,N_7721,N_7905);
nand U8330 (N_8330,N_7624,N_7695);
xor U8331 (N_8331,N_7683,N_7988);
or U8332 (N_8332,N_7707,N_7766);
and U8333 (N_8333,N_7920,N_7793);
or U8334 (N_8334,N_7594,N_7929);
and U8335 (N_8335,N_7605,N_7749);
nor U8336 (N_8336,N_7513,N_7700);
nand U8337 (N_8337,N_7556,N_7697);
or U8338 (N_8338,N_7710,N_7709);
nor U8339 (N_8339,N_7858,N_7824);
xor U8340 (N_8340,N_7671,N_7510);
or U8341 (N_8341,N_7524,N_7858);
and U8342 (N_8342,N_7828,N_7833);
nor U8343 (N_8343,N_7975,N_7981);
and U8344 (N_8344,N_7892,N_7687);
and U8345 (N_8345,N_7725,N_7689);
and U8346 (N_8346,N_7966,N_7764);
or U8347 (N_8347,N_7915,N_7729);
and U8348 (N_8348,N_7984,N_7759);
nor U8349 (N_8349,N_7877,N_7777);
xnor U8350 (N_8350,N_7957,N_7745);
nand U8351 (N_8351,N_7613,N_7765);
nor U8352 (N_8352,N_7502,N_7657);
and U8353 (N_8353,N_7816,N_7736);
nand U8354 (N_8354,N_7888,N_7770);
or U8355 (N_8355,N_7806,N_7984);
nor U8356 (N_8356,N_7514,N_7729);
nand U8357 (N_8357,N_7954,N_7520);
nand U8358 (N_8358,N_7932,N_7553);
xnor U8359 (N_8359,N_7995,N_7703);
or U8360 (N_8360,N_7596,N_7739);
and U8361 (N_8361,N_7861,N_7564);
or U8362 (N_8362,N_7765,N_7970);
or U8363 (N_8363,N_7905,N_7785);
or U8364 (N_8364,N_7531,N_7769);
or U8365 (N_8365,N_7668,N_7964);
and U8366 (N_8366,N_7938,N_7841);
nor U8367 (N_8367,N_7932,N_7986);
and U8368 (N_8368,N_7976,N_7554);
or U8369 (N_8369,N_7975,N_7618);
or U8370 (N_8370,N_7561,N_7918);
xor U8371 (N_8371,N_7676,N_7944);
or U8372 (N_8372,N_7947,N_7916);
or U8373 (N_8373,N_7949,N_7652);
xor U8374 (N_8374,N_7698,N_7526);
nor U8375 (N_8375,N_7572,N_7758);
nand U8376 (N_8376,N_7799,N_7653);
nor U8377 (N_8377,N_7568,N_7781);
or U8378 (N_8378,N_7543,N_7698);
and U8379 (N_8379,N_7594,N_7856);
nor U8380 (N_8380,N_7669,N_7926);
xnor U8381 (N_8381,N_7809,N_7764);
xnor U8382 (N_8382,N_7840,N_7987);
or U8383 (N_8383,N_7954,N_7808);
and U8384 (N_8384,N_7852,N_7719);
or U8385 (N_8385,N_7954,N_7732);
xnor U8386 (N_8386,N_7945,N_7826);
xor U8387 (N_8387,N_7738,N_7653);
nor U8388 (N_8388,N_7967,N_7896);
or U8389 (N_8389,N_7566,N_7787);
or U8390 (N_8390,N_7918,N_7603);
or U8391 (N_8391,N_7815,N_7763);
nor U8392 (N_8392,N_7618,N_7940);
nor U8393 (N_8393,N_7899,N_7620);
or U8394 (N_8394,N_7796,N_7568);
nand U8395 (N_8395,N_7964,N_7517);
nand U8396 (N_8396,N_7685,N_7942);
xor U8397 (N_8397,N_7842,N_7656);
nand U8398 (N_8398,N_7646,N_7581);
nor U8399 (N_8399,N_7775,N_7503);
nand U8400 (N_8400,N_7646,N_7807);
or U8401 (N_8401,N_7835,N_7596);
nand U8402 (N_8402,N_7978,N_7965);
or U8403 (N_8403,N_7555,N_7717);
nand U8404 (N_8404,N_7554,N_7968);
and U8405 (N_8405,N_7890,N_7907);
nand U8406 (N_8406,N_7839,N_7979);
nand U8407 (N_8407,N_7508,N_7776);
nand U8408 (N_8408,N_7632,N_7763);
or U8409 (N_8409,N_7819,N_7545);
xnor U8410 (N_8410,N_7890,N_7883);
nand U8411 (N_8411,N_7968,N_7655);
nor U8412 (N_8412,N_7746,N_7691);
and U8413 (N_8413,N_7903,N_7864);
xor U8414 (N_8414,N_7777,N_7699);
and U8415 (N_8415,N_7814,N_7611);
and U8416 (N_8416,N_7767,N_7733);
nor U8417 (N_8417,N_7698,N_7511);
and U8418 (N_8418,N_7936,N_7708);
and U8419 (N_8419,N_7914,N_7947);
and U8420 (N_8420,N_7590,N_7732);
and U8421 (N_8421,N_7611,N_7669);
xor U8422 (N_8422,N_7814,N_7923);
and U8423 (N_8423,N_7581,N_7949);
nand U8424 (N_8424,N_7519,N_7696);
nor U8425 (N_8425,N_7744,N_7968);
nand U8426 (N_8426,N_7966,N_7819);
or U8427 (N_8427,N_7906,N_7989);
nor U8428 (N_8428,N_7614,N_7626);
xnor U8429 (N_8429,N_7896,N_7779);
xor U8430 (N_8430,N_7557,N_7783);
or U8431 (N_8431,N_7970,N_7777);
nand U8432 (N_8432,N_7825,N_7819);
nor U8433 (N_8433,N_7595,N_7919);
or U8434 (N_8434,N_7706,N_7704);
nand U8435 (N_8435,N_7613,N_7795);
nor U8436 (N_8436,N_7991,N_7781);
or U8437 (N_8437,N_7866,N_7503);
and U8438 (N_8438,N_7640,N_7871);
xnor U8439 (N_8439,N_7827,N_7979);
xor U8440 (N_8440,N_7560,N_7607);
or U8441 (N_8441,N_7601,N_7529);
and U8442 (N_8442,N_7992,N_7518);
or U8443 (N_8443,N_7819,N_7724);
nand U8444 (N_8444,N_7982,N_7965);
nand U8445 (N_8445,N_7579,N_7831);
and U8446 (N_8446,N_7520,N_7544);
nor U8447 (N_8447,N_7958,N_7957);
or U8448 (N_8448,N_7504,N_7915);
nand U8449 (N_8449,N_7786,N_7621);
nand U8450 (N_8450,N_7843,N_7825);
xor U8451 (N_8451,N_7778,N_7626);
or U8452 (N_8452,N_7705,N_7875);
or U8453 (N_8453,N_7516,N_7962);
and U8454 (N_8454,N_7855,N_7773);
and U8455 (N_8455,N_7878,N_7941);
nor U8456 (N_8456,N_7612,N_7787);
or U8457 (N_8457,N_7919,N_7807);
nand U8458 (N_8458,N_7608,N_7830);
and U8459 (N_8459,N_7922,N_7520);
and U8460 (N_8460,N_7602,N_7516);
xnor U8461 (N_8461,N_7888,N_7946);
nor U8462 (N_8462,N_7673,N_7889);
and U8463 (N_8463,N_7504,N_7880);
or U8464 (N_8464,N_7527,N_7590);
and U8465 (N_8465,N_7577,N_7789);
nor U8466 (N_8466,N_7869,N_7800);
nand U8467 (N_8467,N_7671,N_7716);
xor U8468 (N_8468,N_7917,N_7731);
nor U8469 (N_8469,N_7821,N_7511);
or U8470 (N_8470,N_7502,N_7631);
xor U8471 (N_8471,N_7941,N_7852);
or U8472 (N_8472,N_7852,N_7856);
nor U8473 (N_8473,N_7861,N_7765);
nand U8474 (N_8474,N_7711,N_7763);
and U8475 (N_8475,N_7570,N_7606);
nand U8476 (N_8476,N_7620,N_7961);
or U8477 (N_8477,N_7792,N_7957);
nand U8478 (N_8478,N_7543,N_7508);
nor U8479 (N_8479,N_7832,N_7997);
nor U8480 (N_8480,N_7673,N_7790);
and U8481 (N_8481,N_7642,N_7764);
nand U8482 (N_8482,N_7869,N_7932);
nand U8483 (N_8483,N_7695,N_7512);
nor U8484 (N_8484,N_7618,N_7586);
xor U8485 (N_8485,N_7882,N_7903);
nor U8486 (N_8486,N_7596,N_7569);
or U8487 (N_8487,N_7993,N_7963);
xnor U8488 (N_8488,N_7738,N_7841);
xnor U8489 (N_8489,N_7907,N_7994);
or U8490 (N_8490,N_7840,N_7538);
and U8491 (N_8491,N_7799,N_7710);
nand U8492 (N_8492,N_7661,N_7872);
nand U8493 (N_8493,N_7820,N_7881);
nand U8494 (N_8494,N_7710,N_7959);
and U8495 (N_8495,N_7849,N_7719);
nand U8496 (N_8496,N_7713,N_7655);
nand U8497 (N_8497,N_7935,N_7594);
xor U8498 (N_8498,N_7567,N_7704);
nand U8499 (N_8499,N_7509,N_7898);
nor U8500 (N_8500,N_8001,N_8185);
or U8501 (N_8501,N_8342,N_8041);
nand U8502 (N_8502,N_8307,N_8121);
or U8503 (N_8503,N_8306,N_8471);
and U8504 (N_8504,N_8440,N_8132);
and U8505 (N_8505,N_8479,N_8034);
and U8506 (N_8506,N_8272,N_8357);
nand U8507 (N_8507,N_8350,N_8370);
nor U8508 (N_8508,N_8255,N_8300);
xor U8509 (N_8509,N_8367,N_8207);
nand U8510 (N_8510,N_8012,N_8196);
nand U8511 (N_8511,N_8403,N_8019);
nor U8512 (N_8512,N_8401,N_8213);
and U8513 (N_8513,N_8105,N_8150);
xnor U8514 (N_8514,N_8188,N_8358);
or U8515 (N_8515,N_8483,N_8275);
xnor U8516 (N_8516,N_8436,N_8478);
and U8517 (N_8517,N_8294,N_8347);
nand U8518 (N_8518,N_8052,N_8181);
xor U8519 (N_8519,N_8262,N_8464);
xor U8520 (N_8520,N_8455,N_8140);
xor U8521 (N_8521,N_8382,N_8108);
or U8522 (N_8522,N_8462,N_8032);
and U8523 (N_8523,N_8095,N_8092);
nand U8524 (N_8524,N_8399,N_8428);
nor U8525 (N_8525,N_8119,N_8496);
and U8526 (N_8526,N_8433,N_8003);
xor U8527 (N_8527,N_8424,N_8045);
or U8528 (N_8528,N_8091,N_8419);
or U8529 (N_8529,N_8125,N_8058);
xor U8530 (N_8530,N_8426,N_8258);
nand U8531 (N_8531,N_8490,N_8302);
nor U8532 (N_8532,N_8099,N_8212);
and U8533 (N_8533,N_8271,N_8182);
nand U8534 (N_8534,N_8210,N_8482);
xnor U8535 (N_8535,N_8187,N_8222);
and U8536 (N_8536,N_8248,N_8197);
or U8537 (N_8537,N_8253,N_8221);
xnor U8538 (N_8538,N_8036,N_8466);
or U8539 (N_8539,N_8240,N_8093);
or U8540 (N_8540,N_8329,N_8154);
and U8541 (N_8541,N_8035,N_8468);
nand U8542 (N_8542,N_8441,N_8249);
and U8543 (N_8543,N_8220,N_8410);
nor U8544 (N_8544,N_8322,N_8214);
nand U8545 (N_8545,N_8086,N_8340);
xnor U8546 (N_8546,N_8224,N_8163);
nor U8547 (N_8547,N_8394,N_8420);
and U8548 (N_8548,N_8051,N_8028);
nand U8549 (N_8549,N_8276,N_8391);
or U8550 (N_8550,N_8386,N_8193);
or U8551 (N_8551,N_8067,N_8319);
nand U8552 (N_8552,N_8373,N_8065);
nand U8553 (N_8553,N_8075,N_8388);
or U8554 (N_8554,N_8260,N_8409);
or U8555 (N_8555,N_8149,N_8209);
xor U8556 (N_8556,N_8082,N_8002);
and U8557 (N_8557,N_8195,N_8328);
nand U8558 (N_8558,N_8161,N_8492);
and U8559 (N_8559,N_8009,N_8166);
or U8560 (N_8560,N_8162,N_8283);
nand U8561 (N_8561,N_8005,N_8458);
nor U8562 (N_8562,N_8407,N_8024);
or U8563 (N_8563,N_8070,N_8349);
nor U8564 (N_8564,N_8006,N_8025);
and U8565 (N_8565,N_8172,N_8241);
xnor U8566 (N_8566,N_8296,N_8178);
nand U8567 (N_8567,N_8146,N_8079);
or U8568 (N_8568,N_8174,N_8189);
nor U8569 (N_8569,N_8153,N_8447);
nand U8570 (N_8570,N_8397,N_8497);
and U8571 (N_8571,N_8372,N_8413);
xnor U8572 (N_8572,N_8218,N_8083);
or U8573 (N_8573,N_8327,N_8049);
nor U8574 (N_8574,N_8033,N_8074);
xnor U8575 (N_8575,N_8402,N_8011);
xor U8576 (N_8576,N_8008,N_8280);
xor U8577 (N_8577,N_8434,N_8359);
nand U8578 (N_8578,N_8289,N_8109);
xnor U8579 (N_8579,N_8158,N_8183);
nand U8580 (N_8580,N_8425,N_8336);
xor U8581 (N_8581,N_8156,N_8416);
nor U8582 (N_8582,N_8341,N_8363);
nand U8583 (N_8583,N_8287,N_8481);
nor U8584 (N_8584,N_8208,N_8216);
nand U8585 (N_8585,N_8064,N_8127);
nor U8586 (N_8586,N_8485,N_8236);
xnor U8587 (N_8587,N_8384,N_8202);
xor U8588 (N_8588,N_8459,N_8152);
nor U8589 (N_8589,N_8335,N_8239);
xor U8590 (N_8590,N_8446,N_8332);
and U8591 (N_8591,N_8203,N_8164);
xor U8592 (N_8592,N_8057,N_8250);
or U8593 (N_8593,N_8257,N_8321);
or U8594 (N_8594,N_8219,N_8405);
nor U8595 (N_8595,N_8389,N_8415);
or U8596 (N_8596,N_8398,N_8039);
nor U8597 (N_8597,N_8072,N_8017);
nand U8598 (N_8598,N_8225,N_8138);
nor U8599 (N_8599,N_8487,N_8282);
nand U8600 (N_8600,N_8310,N_8047);
and U8601 (N_8601,N_8186,N_8097);
or U8602 (N_8602,N_8068,N_8110);
nand U8603 (N_8603,N_8043,N_8114);
and U8604 (N_8604,N_8026,N_8376);
and U8605 (N_8605,N_8274,N_8015);
and U8606 (N_8606,N_8361,N_8444);
nand U8607 (N_8607,N_8493,N_8211);
and U8608 (N_8608,N_8309,N_8046);
and U8609 (N_8609,N_8264,N_8023);
nor U8610 (N_8610,N_8044,N_8390);
nor U8611 (N_8611,N_8170,N_8355);
nor U8612 (N_8612,N_8456,N_8432);
nand U8613 (N_8613,N_8270,N_8293);
or U8614 (N_8614,N_8457,N_8465);
nand U8615 (N_8615,N_8469,N_8404);
or U8616 (N_8616,N_8206,N_8438);
and U8617 (N_8617,N_8038,N_8247);
nand U8618 (N_8618,N_8325,N_8489);
nand U8619 (N_8619,N_8215,N_8256);
xnor U8620 (N_8620,N_8037,N_8266);
xor U8621 (N_8621,N_8194,N_8245);
nor U8622 (N_8622,N_8124,N_8176);
nor U8623 (N_8623,N_8159,N_8131);
and U8624 (N_8624,N_8050,N_8055);
and U8625 (N_8625,N_8141,N_8071);
and U8626 (N_8626,N_8130,N_8380);
nand U8627 (N_8627,N_8004,N_8175);
nor U8628 (N_8628,N_8360,N_8246);
nor U8629 (N_8629,N_8148,N_8334);
nor U8630 (N_8630,N_8313,N_8348);
or U8631 (N_8631,N_8470,N_8123);
xnor U8632 (N_8632,N_8463,N_8229);
nor U8633 (N_8633,N_8308,N_8018);
nand U8634 (N_8634,N_8155,N_8273);
and U8635 (N_8635,N_8443,N_8031);
nor U8636 (N_8636,N_8473,N_8377);
or U8637 (N_8637,N_8339,N_8021);
nand U8638 (N_8638,N_8192,N_8198);
xor U8639 (N_8639,N_8134,N_8251);
nor U8640 (N_8640,N_8383,N_8118);
nor U8641 (N_8641,N_8412,N_8160);
xnor U8642 (N_8642,N_8318,N_8151);
or U8643 (N_8643,N_8199,N_8356);
xor U8644 (N_8644,N_8261,N_8385);
xnor U8645 (N_8645,N_8450,N_8263);
and U8646 (N_8646,N_8452,N_8277);
xnor U8647 (N_8647,N_8379,N_8323);
xnor U8648 (N_8648,N_8467,N_8486);
nor U8649 (N_8649,N_8352,N_8088);
nor U8650 (N_8650,N_8429,N_8291);
xor U8651 (N_8651,N_8406,N_8040);
xor U8652 (N_8652,N_8242,N_8312);
and U8653 (N_8653,N_8364,N_8314);
nand U8654 (N_8654,N_8366,N_8101);
or U8655 (N_8655,N_8080,N_8030);
nor U8656 (N_8656,N_8104,N_8371);
or U8657 (N_8657,N_8085,N_8103);
or U8658 (N_8658,N_8311,N_8157);
xor U8659 (N_8659,N_8354,N_8115);
nor U8660 (N_8660,N_8237,N_8096);
nand U8661 (N_8661,N_8442,N_8090);
and U8662 (N_8662,N_8252,N_8167);
nor U8663 (N_8663,N_8353,N_8298);
or U8664 (N_8664,N_8474,N_8062);
and U8665 (N_8665,N_8351,N_8396);
or U8666 (N_8666,N_8027,N_8393);
and U8667 (N_8667,N_8437,N_8439);
nand U8668 (N_8668,N_8331,N_8147);
and U8669 (N_8669,N_8244,N_8061);
xnor U8670 (N_8670,N_8000,N_8400);
and U8671 (N_8671,N_8133,N_8461);
and U8672 (N_8672,N_8292,N_8265);
nand U8673 (N_8673,N_8137,N_8381);
xnor U8674 (N_8674,N_8077,N_8191);
xnor U8675 (N_8675,N_8087,N_8168);
and U8676 (N_8676,N_8020,N_8453);
nor U8677 (N_8677,N_8117,N_8078);
nand U8678 (N_8678,N_8480,N_8427);
xnor U8679 (N_8679,N_8238,N_8171);
or U8680 (N_8680,N_8144,N_8414);
and U8681 (N_8681,N_8243,N_8076);
nand U8682 (N_8682,N_8418,N_8116);
nor U8683 (N_8683,N_8284,N_8343);
or U8684 (N_8684,N_8136,N_8476);
nand U8685 (N_8685,N_8295,N_8337);
or U8686 (N_8686,N_8042,N_8226);
and U8687 (N_8687,N_8281,N_8217);
and U8688 (N_8688,N_8190,N_8315);
or U8689 (N_8689,N_8177,N_8059);
xnor U8690 (N_8690,N_8056,N_8233);
nand U8691 (N_8691,N_8454,N_8165);
xor U8692 (N_8692,N_8200,N_8112);
xor U8693 (N_8693,N_8128,N_8324);
nand U8694 (N_8694,N_8430,N_8326);
nand U8695 (N_8695,N_8344,N_8053);
nor U8696 (N_8696,N_8346,N_8107);
xor U8697 (N_8697,N_8232,N_8016);
nand U8698 (N_8698,N_8301,N_8378);
xnor U8699 (N_8699,N_8169,N_8231);
nor U8700 (N_8700,N_8368,N_8054);
or U8701 (N_8701,N_8084,N_8320);
and U8702 (N_8702,N_8369,N_8048);
nand U8703 (N_8703,N_8254,N_8305);
nor U8704 (N_8704,N_8488,N_8421);
and U8705 (N_8705,N_8408,N_8477);
nand U8706 (N_8706,N_8451,N_8268);
or U8707 (N_8707,N_8139,N_8374);
xor U8708 (N_8708,N_8495,N_8010);
and U8709 (N_8709,N_8297,N_8435);
nand U8710 (N_8710,N_8205,N_8106);
xnor U8711 (N_8711,N_8345,N_8460);
nor U8712 (N_8712,N_8286,N_8223);
nor U8713 (N_8713,N_8235,N_8303);
xor U8714 (N_8714,N_8100,N_8316);
or U8715 (N_8715,N_8029,N_8288);
nor U8716 (N_8716,N_8431,N_8069);
xnor U8717 (N_8717,N_8299,N_8362);
nor U8718 (N_8718,N_8259,N_8073);
nor U8719 (N_8719,N_8081,N_8113);
and U8720 (N_8720,N_8475,N_8122);
and U8721 (N_8721,N_8304,N_8066);
or U8722 (N_8722,N_8089,N_8126);
nand U8723 (N_8723,N_8472,N_8094);
nand U8724 (N_8724,N_8423,N_8120);
or U8725 (N_8725,N_8448,N_8142);
xnor U8726 (N_8726,N_8230,N_8278);
nand U8727 (N_8727,N_8173,N_8375);
or U8728 (N_8728,N_8102,N_8111);
nor U8729 (N_8729,N_8365,N_8484);
nor U8730 (N_8730,N_8180,N_8228);
or U8731 (N_8731,N_8494,N_8063);
or U8732 (N_8732,N_8060,N_8267);
xor U8733 (N_8733,N_8234,N_8129);
nand U8734 (N_8734,N_8179,N_8499);
and U8735 (N_8735,N_8269,N_8022);
and U8736 (N_8736,N_8279,N_8498);
and U8737 (N_8737,N_8411,N_8145);
nor U8738 (N_8738,N_8143,N_8392);
or U8739 (N_8739,N_8014,N_8338);
and U8740 (N_8740,N_8387,N_8317);
xor U8741 (N_8741,N_8098,N_8395);
and U8742 (N_8742,N_8201,N_8290);
xnor U8743 (N_8743,N_8417,N_8491);
xor U8744 (N_8744,N_8330,N_8007);
xor U8745 (N_8745,N_8333,N_8445);
or U8746 (N_8746,N_8204,N_8013);
xor U8747 (N_8747,N_8227,N_8184);
and U8748 (N_8748,N_8422,N_8449);
and U8749 (N_8749,N_8285,N_8135);
xor U8750 (N_8750,N_8076,N_8026);
nand U8751 (N_8751,N_8486,N_8281);
xnor U8752 (N_8752,N_8413,N_8460);
nor U8753 (N_8753,N_8021,N_8229);
or U8754 (N_8754,N_8286,N_8344);
nor U8755 (N_8755,N_8406,N_8325);
nand U8756 (N_8756,N_8488,N_8124);
nor U8757 (N_8757,N_8057,N_8458);
or U8758 (N_8758,N_8117,N_8109);
xnor U8759 (N_8759,N_8363,N_8362);
xor U8760 (N_8760,N_8206,N_8048);
and U8761 (N_8761,N_8194,N_8446);
nor U8762 (N_8762,N_8427,N_8417);
and U8763 (N_8763,N_8001,N_8417);
xnor U8764 (N_8764,N_8084,N_8408);
nor U8765 (N_8765,N_8463,N_8434);
or U8766 (N_8766,N_8065,N_8208);
or U8767 (N_8767,N_8328,N_8260);
and U8768 (N_8768,N_8245,N_8116);
and U8769 (N_8769,N_8266,N_8352);
xnor U8770 (N_8770,N_8353,N_8236);
xnor U8771 (N_8771,N_8138,N_8393);
xor U8772 (N_8772,N_8200,N_8289);
nor U8773 (N_8773,N_8098,N_8248);
or U8774 (N_8774,N_8329,N_8213);
or U8775 (N_8775,N_8113,N_8362);
xnor U8776 (N_8776,N_8327,N_8371);
and U8777 (N_8777,N_8119,N_8446);
nand U8778 (N_8778,N_8056,N_8080);
and U8779 (N_8779,N_8207,N_8055);
nand U8780 (N_8780,N_8049,N_8372);
and U8781 (N_8781,N_8310,N_8171);
nor U8782 (N_8782,N_8286,N_8200);
or U8783 (N_8783,N_8367,N_8231);
and U8784 (N_8784,N_8077,N_8333);
and U8785 (N_8785,N_8216,N_8171);
xor U8786 (N_8786,N_8215,N_8008);
nor U8787 (N_8787,N_8366,N_8164);
xnor U8788 (N_8788,N_8292,N_8390);
nor U8789 (N_8789,N_8249,N_8360);
or U8790 (N_8790,N_8189,N_8348);
xor U8791 (N_8791,N_8203,N_8393);
or U8792 (N_8792,N_8027,N_8193);
nor U8793 (N_8793,N_8363,N_8280);
nor U8794 (N_8794,N_8118,N_8310);
xnor U8795 (N_8795,N_8222,N_8151);
nor U8796 (N_8796,N_8438,N_8431);
or U8797 (N_8797,N_8037,N_8305);
nor U8798 (N_8798,N_8270,N_8382);
nor U8799 (N_8799,N_8201,N_8194);
nand U8800 (N_8800,N_8292,N_8212);
or U8801 (N_8801,N_8001,N_8114);
nand U8802 (N_8802,N_8332,N_8485);
xnor U8803 (N_8803,N_8175,N_8324);
xor U8804 (N_8804,N_8019,N_8461);
nand U8805 (N_8805,N_8390,N_8431);
nor U8806 (N_8806,N_8310,N_8332);
xnor U8807 (N_8807,N_8130,N_8424);
nor U8808 (N_8808,N_8379,N_8246);
or U8809 (N_8809,N_8357,N_8486);
nor U8810 (N_8810,N_8173,N_8493);
nand U8811 (N_8811,N_8468,N_8294);
xor U8812 (N_8812,N_8491,N_8420);
nor U8813 (N_8813,N_8255,N_8023);
nand U8814 (N_8814,N_8034,N_8445);
and U8815 (N_8815,N_8410,N_8010);
nor U8816 (N_8816,N_8034,N_8058);
nor U8817 (N_8817,N_8160,N_8183);
nand U8818 (N_8818,N_8122,N_8093);
nor U8819 (N_8819,N_8331,N_8014);
or U8820 (N_8820,N_8486,N_8448);
and U8821 (N_8821,N_8100,N_8488);
nand U8822 (N_8822,N_8486,N_8222);
nor U8823 (N_8823,N_8340,N_8397);
or U8824 (N_8824,N_8016,N_8449);
or U8825 (N_8825,N_8089,N_8062);
nand U8826 (N_8826,N_8289,N_8046);
xnor U8827 (N_8827,N_8467,N_8200);
nand U8828 (N_8828,N_8152,N_8170);
xor U8829 (N_8829,N_8084,N_8344);
nand U8830 (N_8830,N_8343,N_8112);
xnor U8831 (N_8831,N_8322,N_8347);
and U8832 (N_8832,N_8176,N_8282);
or U8833 (N_8833,N_8422,N_8012);
nor U8834 (N_8834,N_8099,N_8378);
nor U8835 (N_8835,N_8293,N_8281);
nand U8836 (N_8836,N_8403,N_8329);
xnor U8837 (N_8837,N_8341,N_8079);
xnor U8838 (N_8838,N_8250,N_8034);
nand U8839 (N_8839,N_8211,N_8338);
nor U8840 (N_8840,N_8197,N_8350);
or U8841 (N_8841,N_8282,N_8455);
and U8842 (N_8842,N_8139,N_8337);
nand U8843 (N_8843,N_8296,N_8329);
and U8844 (N_8844,N_8314,N_8355);
and U8845 (N_8845,N_8306,N_8053);
or U8846 (N_8846,N_8323,N_8369);
xnor U8847 (N_8847,N_8315,N_8343);
nor U8848 (N_8848,N_8282,N_8322);
nor U8849 (N_8849,N_8372,N_8325);
and U8850 (N_8850,N_8173,N_8456);
nand U8851 (N_8851,N_8057,N_8483);
and U8852 (N_8852,N_8096,N_8321);
and U8853 (N_8853,N_8044,N_8491);
nor U8854 (N_8854,N_8497,N_8448);
xnor U8855 (N_8855,N_8136,N_8009);
xnor U8856 (N_8856,N_8240,N_8438);
or U8857 (N_8857,N_8007,N_8001);
xor U8858 (N_8858,N_8200,N_8426);
xnor U8859 (N_8859,N_8340,N_8047);
nand U8860 (N_8860,N_8134,N_8025);
nand U8861 (N_8861,N_8417,N_8228);
and U8862 (N_8862,N_8101,N_8414);
nor U8863 (N_8863,N_8271,N_8274);
nand U8864 (N_8864,N_8335,N_8340);
or U8865 (N_8865,N_8224,N_8127);
and U8866 (N_8866,N_8238,N_8335);
nand U8867 (N_8867,N_8141,N_8334);
nor U8868 (N_8868,N_8158,N_8116);
xor U8869 (N_8869,N_8373,N_8049);
xnor U8870 (N_8870,N_8400,N_8356);
nand U8871 (N_8871,N_8279,N_8412);
or U8872 (N_8872,N_8143,N_8163);
xor U8873 (N_8873,N_8287,N_8153);
or U8874 (N_8874,N_8069,N_8450);
and U8875 (N_8875,N_8459,N_8216);
or U8876 (N_8876,N_8032,N_8068);
nand U8877 (N_8877,N_8188,N_8384);
and U8878 (N_8878,N_8481,N_8438);
or U8879 (N_8879,N_8267,N_8153);
xnor U8880 (N_8880,N_8300,N_8291);
nand U8881 (N_8881,N_8201,N_8212);
and U8882 (N_8882,N_8474,N_8142);
nand U8883 (N_8883,N_8348,N_8466);
nand U8884 (N_8884,N_8195,N_8283);
nor U8885 (N_8885,N_8232,N_8209);
xor U8886 (N_8886,N_8233,N_8457);
xor U8887 (N_8887,N_8331,N_8309);
xnor U8888 (N_8888,N_8427,N_8351);
xor U8889 (N_8889,N_8293,N_8327);
nand U8890 (N_8890,N_8011,N_8079);
xor U8891 (N_8891,N_8039,N_8148);
or U8892 (N_8892,N_8034,N_8242);
nor U8893 (N_8893,N_8229,N_8471);
xor U8894 (N_8894,N_8232,N_8098);
nand U8895 (N_8895,N_8267,N_8340);
nand U8896 (N_8896,N_8201,N_8090);
and U8897 (N_8897,N_8008,N_8343);
and U8898 (N_8898,N_8141,N_8177);
and U8899 (N_8899,N_8225,N_8328);
xnor U8900 (N_8900,N_8228,N_8316);
xor U8901 (N_8901,N_8328,N_8274);
xor U8902 (N_8902,N_8160,N_8212);
and U8903 (N_8903,N_8115,N_8111);
nor U8904 (N_8904,N_8466,N_8067);
xnor U8905 (N_8905,N_8088,N_8021);
xnor U8906 (N_8906,N_8342,N_8214);
and U8907 (N_8907,N_8276,N_8345);
nand U8908 (N_8908,N_8089,N_8190);
or U8909 (N_8909,N_8031,N_8012);
nor U8910 (N_8910,N_8045,N_8089);
or U8911 (N_8911,N_8489,N_8465);
and U8912 (N_8912,N_8350,N_8114);
xnor U8913 (N_8913,N_8487,N_8405);
xnor U8914 (N_8914,N_8044,N_8454);
xor U8915 (N_8915,N_8169,N_8256);
and U8916 (N_8916,N_8370,N_8377);
nand U8917 (N_8917,N_8257,N_8107);
xor U8918 (N_8918,N_8015,N_8427);
or U8919 (N_8919,N_8412,N_8436);
nand U8920 (N_8920,N_8020,N_8080);
or U8921 (N_8921,N_8205,N_8423);
xnor U8922 (N_8922,N_8477,N_8014);
and U8923 (N_8923,N_8467,N_8298);
xor U8924 (N_8924,N_8218,N_8324);
nor U8925 (N_8925,N_8363,N_8382);
xnor U8926 (N_8926,N_8010,N_8433);
or U8927 (N_8927,N_8161,N_8352);
xnor U8928 (N_8928,N_8254,N_8371);
or U8929 (N_8929,N_8063,N_8209);
nor U8930 (N_8930,N_8161,N_8041);
xor U8931 (N_8931,N_8124,N_8013);
nor U8932 (N_8932,N_8484,N_8050);
nand U8933 (N_8933,N_8492,N_8493);
nand U8934 (N_8934,N_8230,N_8383);
and U8935 (N_8935,N_8326,N_8212);
nor U8936 (N_8936,N_8426,N_8444);
nor U8937 (N_8937,N_8145,N_8470);
and U8938 (N_8938,N_8001,N_8378);
nor U8939 (N_8939,N_8455,N_8029);
and U8940 (N_8940,N_8145,N_8200);
nor U8941 (N_8941,N_8084,N_8303);
and U8942 (N_8942,N_8390,N_8163);
nor U8943 (N_8943,N_8289,N_8280);
xor U8944 (N_8944,N_8381,N_8477);
and U8945 (N_8945,N_8392,N_8481);
or U8946 (N_8946,N_8375,N_8148);
xor U8947 (N_8947,N_8096,N_8304);
or U8948 (N_8948,N_8301,N_8262);
or U8949 (N_8949,N_8017,N_8311);
and U8950 (N_8950,N_8289,N_8369);
nand U8951 (N_8951,N_8441,N_8143);
nand U8952 (N_8952,N_8307,N_8178);
nor U8953 (N_8953,N_8170,N_8428);
xor U8954 (N_8954,N_8322,N_8424);
and U8955 (N_8955,N_8257,N_8323);
and U8956 (N_8956,N_8494,N_8048);
nand U8957 (N_8957,N_8425,N_8390);
nand U8958 (N_8958,N_8080,N_8258);
or U8959 (N_8959,N_8464,N_8042);
xor U8960 (N_8960,N_8291,N_8014);
and U8961 (N_8961,N_8018,N_8226);
nor U8962 (N_8962,N_8381,N_8347);
nand U8963 (N_8963,N_8394,N_8462);
and U8964 (N_8964,N_8351,N_8241);
nand U8965 (N_8965,N_8290,N_8321);
or U8966 (N_8966,N_8099,N_8443);
xor U8967 (N_8967,N_8350,N_8383);
nand U8968 (N_8968,N_8213,N_8232);
xor U8969 (N_8969,N_8322,N_8488);
and U8970 (N_8970,N_8035,N_8321);
and U8971 (N_8971,N_8130,N_8096);
and U8972 (N_8972,N_8366,N_8166);
xor U8973 (N_8973,N_8267,N_8033);
and U8974 (N_8974,N_8349,N_8416);
and U8975 (N_8975,N_8307,N_8496);
nand U8976 (N_8976,N_8153,N_8460);
and U8977 (N_8977,N_8205,N_8130);
nor U8978 (N_8978,N_8000,N_8103);
or U8979 (N_8979,N_8146,N_8190);
nand U8980 (N_8980,N_8463,N_8219);
nor U8981 (N_8981,N_8273,N_8430);
and U8982 (N_8982,N_8493,N_8068);
xor U8983 (N_8983,N_8386,N_8465);
xnor U8984 (N_8984,N_8292,N_8056);
and U8985 (N_8985,N_8489,N_8142);
nor U8986 (N_8986,N_8197,N_8397);
or U8987 (N_8987,N_8093,N_8034);
nand U8988 (N_8988,N_8387,N_8180);
or U8989 (N_8989,N_8287,N_8415);
nor U8990 (N_8990,N_8488,N_8461);
and U8991 (N_8991,N_8104,N_8248);
nor U8992 (N_8992,N_8230,N_8184);
nor U8993 (N_8993,N_8327,N_8237);
nand U8994 (N_8994,N_8220,N_8096);
nor U8995 (N_8995,N_8264,N_8054);
nand U8996 (N_8996,N_8177,N_8314);
or U8997 (N_8997,N_8235,N_8414);
xnor U8998 (N_8998,N_8495,N_8066);
nand U8999 (N_8999,N_8278,N_8053);
nor U9000 (N_9000,N_8642,N_8629);
or U9001 (N_9001,N_8754,N_8821);
and U9002 (N_9002,N_8625,N_8747);
or U9003 (N_9003,N_8717,N_8977);
nand U9004 (N_9004,N_8501,N_8579);
nor U9005 (N_9005,N_8780,N_8775);
and U9006 (N_9006,N_8656,N_8819);
nand U9007 (N_9007,N_8841,N_8830);
and U9008 (N_9008,N_8544,N_8556);
nand U9009 (N_9009,N_8768,N_8619);
nor U9010 (N_9010,N_8985,N_8992);
and U9011 (N_9011,N_8870,N_8912);
nor U9012 (N_9012,N_8998,N_8837);
or U9013 (N_9013,N_8962,N_8741);
or U9014 (N_9014,N_8878,N_8887);
xnor U9015 (N_9015,N_8602,N_8618);
nor U9016 (N_9016,N_8785,N_8990);
nor U9017 (N_9017,N_8971,N_8514);
and U9018 (N_9018,N_8527,N_8667);
and U9019 (N_9019,N_8925,N_8574);
xnor U9020 (N_9020,N_8773,N_8926);
xor U9021 (N_9021,N_8682,N_8562);
and U9022 (N_9022,N_8970,N_8729);
nor U9023 (N_9023,N_8645,N_8955);
nor U9024 (N_9024,N_8897,N_8695);
or U9025 (N_9025,N_8718,N_8877);
and U9026 (N_9026,N_8883,N_8793);
xor U9027 (N_9027,N_8829,N_8942);
and U9028 (N_9028,N_8908,N_8731);
nand U9029 (N_9029,N_8694,N_8523);
or U9030 (N_9030,N_8563,N_8834);
nor U9031 (N_9031,N_8928,N_8687);
or U9032 (N_9032,N_8999,N_8838);
nor U9033 (N_9033,N_8650,N_8605);
or U9034 (N_9034,N_8533,N_8993);
or U9035 (N_9035,N_8854,N_8587);
nor U9036 (N_9036,N_8689,N_8658);
and U9037 (N_9037,N_8572,N_8916);
or U9038 (N_9038,N_8759,N_8657);
or U9039 (N_9039,N_8545,N_8714);
and U9040 (N_9040,N_8525,N_8716);
nand U9041 (N_9041,N_8739,N_8839);
nor U9042 (N_9042,N_8835,N_8910);
and U9043 (N_9043,N_8935,N_8715);
and U9044 (N_9044,N_8982,N_8799);
or U9045 (N_9045,N_8530,N_8790);
and U9046 (N_9046,N_8844,N_8875);
nand U9047 (N_9047,N_8507,N_8610);
and U9048 (N_9048,N_8711,N_8763);
nor U9049 (N_9049,N_8526,N_8691);
xnor U9050 (N_9050,N_8896,N_8934);
nand U9051 (N_9051,N_8669,N_8807);
nand U9052 (N_9052,N_8590,N_8538);
and U9053 (N_9053,N_8709,N_8930);
or U9054 (N_9054,N_8980,N_8564);
nor U9055 (N_9055,N_8802,N_8913);
or U9056 (N_9056,N_8660,N_8893);
xor U9057 (N_9057,N_8614,N_8789);
and U9058 (N_9058,N_8510,N_8520);
and U9059 (N_9059,N_8621,N_8920);
or U9060 (N_9060,N_8596,N_8818);
xnor U9061 (N_9061,N_8787,N_8532);
nand U9062 (N_9062,N_8863,N_8640);
nand U9063 (N_9063,N_8606,N_8932);
nand U9064 (N_9064,N_8652,N_8987);
or U9065 (N_9065,N_8542,N_8655);
xor U9066 (N_9066,N_8812,N_8937);
and U9067 (N_9067,N_8984,N_8794);
or U9068 (N_9068,N_8943,N_8751);
and U9069 (N_9069,N_8728,N_8866);
nand U9070 (N_9070,N_8949,N_8541);
xor U9071 (N_9071,N_8557,N_8677);
xor U9072 (N_9072,N_8588,N_8852);
xor U9073 (N_9073,N_8504,N_8659);
xor U9074 (N_9074,N_8769,N_8534);
nor U9075 (N_9075,N_8784,N_8688);
or U9076 (N_9076,N_8743,N_8700);
nand U9077 (N_9077,N_8989,N_8933);
nand U9078 (N_9078,N_8749,N_8840);
and U9079 (N_9079,N_8918,N_8549);
and U9080 (N_9080,N_8696,N_8617);
or U9081 (N_9081,N_8948,N_8740);
nor U9082 (N_9082,N_8733,N_8959);
and U9083 (N_9083,N_8853,N_8960);
nor U9084 (N_9084,N_8742,N_8552);
xnor U9085 (N_9085,N_8566,N_8692);
and U9086 (N_9086,N_8901,N_8737);
nor U9087 (N_9087,N_8974,N_8967);
nor U9088 (N_9088,N_8503,N_8808);
nand U9089 (N_9089,N_8979,N_8651);
nor U9090 (N_9090,N_8881,N_8641);
nor U9091 (N_9091,N_8771,N_8836);
and U9092 (N_9092,N_8864,N_8941);
and U9093 (N_9093,N_8813,N_8531);
xnor U9094 (N_9094,N_8903,N_8976);
nor U9095 (N_9095,N_8663,N_8585);
and U9096 (N_9096,N_8828,N_8764);
and U9097 (N_9097,N_8738,N_8861);
or U9098 (N_9098,N_8888,N_8608);
or U9099 (N_9099,N_8953,N_8902);
nor U9100 (N_9100,N_8680,N_8859);
xor U9101 (N_9101,N_8584,N_8851);
or U9102 (N_9102,N_8911,N_8515);
nor U9103 (N_9103,N_8800,N_8643);
xor U9104 (N_9104,N_8620,N_8710);
nand U9105 (N_9105,N_8712,N_8543);
xnor U9106 (N_9106,N_8699,N_8683);
or U9107 (N_9107,N_8755,N_8644);
xnor U9108 (N_9108,N_8779,N_8513);
xor U9109 (N_9109,N_8831,N_8529);
and U9110 (N_9110,N_8867,N_8871);
or U9111 (N_9111,N_8704,N_8891);
nand U9112 (N_9112,N_8786,N_8589);
nor U9113 (N_9113,N_8547,N_8665);
xnor U9114 (N_9114,N_8637,N_8686);
xnor U9115 (N_9115,N_8791,N_8517);
or U9116 (N_9116,N_8539,N_8627);
or U9117 (N_9117,N_8805,N_8772);
and U9118 (N_9118,N_8612,N_8862);
or U9119 (N_9119,N_8890,N_8796);
nor U9120 (N_9120,N_8849,N_8598);
or U9121 (N_9121,N_8915,N_8604);
xnor U9122 (N_9122,N_8927,N_8846);
and U9123 (N_9123,N_8622,N_8647);
or U9124 (N_9124,N_8899,N_8646);
or U9125 (N_9125,N_8944,N_8703);
and U9126 (N_9126,N_8810,N_8636);
nor U9127 (N_9127,N_8550,N_8994);
nor U9128 (N_9128,N_8511,N_8963);
or U9129 (N_9129,N_8827,N_8991);
nand U9130 (N_9130,N_8792,N_8988);
nand U9131 (N_9131,N_8500,N_8983);
nand U9132 (N_9132,N_8653,N_8869);
or U9133 (N_9133,N_8968,N_8560);
xnor U9134 (N_9134,N_8630,N_8874);
or U9135 (N_9135,N_8900,N_8732);
nand U9136 (N_9136,N_8722,N_8516);
or U9137 (N_9137,N_8776,N_8756);
and U9138 (N_9138,N_8996,N_8767);
nand U9139 (N_9139,N_8624,N_8761);
nor U9140 (N_9140,N_8894,N_8597);
and U9141 (N_9141,N_8826,N_8553);
nor U9142 (N_9142,N_8748,N_8832);
xnor U9143 (N_9143,N_8924,N_8952);
nor U9144 (N_9144,N_8676,N_8664);
and U9145 (N_9145,N_8847,N_8518);
and U9146 (N_9146,N_8957,N_8734);
nor U9147 (N_9147,N_8939,N_8986);
xnor U9148 (N_9148,N_8966,N_8762);
xnor U9149 (N_9149,N_8524,N_8678);
nand U9150 (N_9150,N_8746,N_8634);
xor U9151 (N_9151,N_8577,N_8855);
and U9152 (N_9152,N_8843,N_8744);
or U9153 (N_9153,N_8626,N_8884);
nand U9154 (N_9154,N_8633,N_8546);
or U9155 (N_9155,N_8995,N_8567);
and U9156 (N_9156,N_8551,N_8945);
or U9157 (N_9157,N_8758,N_8907);
or U9158 (N_9158,N_8508,N_8820);
or U9159 (N_9159,N_8565,N_8795);
and U9160 (N_9160,N_8599,N_8661);
nand U9161 (N_9161,N_8909,N_8725);
nand U9162 (N_9162,N_8917,N_8554);
nand U9163 (N_9163,N_8639,N_8860);
xnor U9164 (N_9164,N_8815,N_8735);
and U9165 (N_9165,N_8865,N_8705);
or U9166 (N_9166,N_8940,N_8506);
nand U9167 (N_9167,N_8671,N_8628);
and U9168 (N_9168,N_8736,N_8923);
or U9169 (N_9169,N_8842,N_8593);
xnor U9170 (N_9170,N_8981,N_8580);
and U9171 (N_9171,N_8889,N_8919);
and U9172 (N_9172,N_8607,N_8753);
or U9173 (N_9173,N_8929,N_8898);
or U9174 (N_9174,N_8635,N_8964);
and U9175 (N_9175,N_8649,N_8783);
nor U9176 (N_9176,N_8814,N_8594);
and U9177 (N_9177,N_8956,N_8951);
xnor U9178 (N_9178,N_8719,N_8879);
nor U9179 (N_9179,N_8528,N_8936);
or U9180 (N_9180,N_8723,N_8782);
or U9181 (N_9181,N_8535,N_8882);
xor U9182 (N_9182,N_8601,N_8648);
or U9183 (N_9183,N_8578,N_8858);
xnor U9184 (N_9184,N_8904,N_8781);
xnor U9185 (N_9185,N_8555,N_8672);
and U9186 (N_9186,N_8536,N_8857);
nor U9187 (N_9187,N_8707,N_8674);
and U9188 (N_9188,N_8788,N_8752);
nor U9189 (N_9189,N_8922,N_8745);
nand U9190 (N_9190,N_8825,N_8569);
nor U9191 (N_9191,N_8872,N_8950);
xnor U9192 (N_9192,N_8679,N_8631);
or U9193 (N_9193,N_8681,N_8575);
or U9194 (N_9194,N_8573,N_8623);
nand U9195 (N_9195,N_8519,N_8522);
or U9196 (N_9196,N_8568,N_8978);
nand U9197 (N_9197,N_8662,N_8559);
nor U9198 (N_9198,N_8811,N_8921);
nor U9199 (N_9199,N_8880,N_8586);
nor U9200 (N_9200,N_8931,N_8774);
nor U9201 (N_9201,N_8505,N_8850);
and U9202 (N_9202,N_8581,N_8613);
xor U9203 (N_9203,N_8886,N_8797);
nand U9204 (N_9204,N_8592,N_8778);
or U9205 (N_9205,N_8502,N_8892);
nand U9206 (N_9206,N_8697,N_8973);
or U9207 (N_9207,N_8673,N_8666);
and U9208 (N_9208,N_8609,N_8750);
and U9209 (N_9209,N_8969,N_8954);
nand U9210 (N_9210,N_8856,N_8720);
nor U9211 (N_9211,N_8512,N_8509);
nand U9212 (N_9212,N_8684,N_8914);
and U9213 (N_9213,N_8706,N_8845);
nand U9214 (N_9214,N_8961,N_8876);
nand U9215 (N_9215,N_8997,N_8611);
xnor U9216 (N_9216,N_8702,N_8972);
and U9217 (N_9217,N_8873,N_8801);
nand U9218 (N_9218,N_8561,N_8708);
or U9219 (N_9219,N_8693,N_8537);
xor U9220 (N_9220,N_8721,N_8570);
and U9221 (N_9221,N_8591,N_8803);
xor U9222 (N_9222,N_8603,N_8975);
nor U9223 (N_9223,N_8654,N_8548);
or U9224 (N_9224,N_8816,N_8824);
xor U9225 (N_9225,N_8946,N_8765);
and U9226 (N_9226,N_8848,N_8895);
nor U9227 (N_9227,N_8600,N_8868);
or U9228 (N_9228,N_8632,N_8713);
nor U9229 (N_9229,N_8906,N_8576);
nor U9230 (N_9230,N_8615,N_8583);
nor U9231 (N_9231,N_8595,N_8806);
xnor U9232 (N_9232,N_8726,N_8670);
nor U9233 (N_9233,N_8798,N_8730);
nand U9234 (N_9234,N_8905,N_8558);
or U9235 (N_9235,N_8766,N_8965);
xnor U9236 (N_9236,N_8770,N_8701);
and U9237 (N_9237,N_8690,N_8833);
or U9238 (N_9238,N_8885,N_8777);
xor U9239 (N_9239,N_8804,N_8698);
nand U9240 (N_9240,N_8958,N_8582);
xor U9241 (N_9241,N_8521,N_8817);
and U9242 (N_9242,N_8685,N_8757);
nor U9243 (N_9243,N_8638,N_8540);
or U9244 (N_9244,N_8668,N_8822);
nor U9245 (N_9245,N_8938,N_8760);
and U9246 (N_9246,N_8675,N_8947);
and U9247 (N_9247,N_8823,N_8809);
nand U9248 (N_9248,N_8724,N_8616);
and U9249 (N_9249,N_8571,N_8727);
xnor U9250 (N_9250,N_8973,N_8914);
and U9251 (N_9251,N_8574,N_8991);
nor U9252 (N_9252,N_8558,N_8798);
nand U9253 (N_9253,N_8945,N_8951);
xor U9254 (N_9254,N_8806,N_8582);
and U9255 (N_9255,N_8832,N_8584);
or U9256 (N_9256,N_8626,N_8835);
nand U9257 (N_9257,N_8964,N_8600);
xor U9258 (N_9258,N_8932,N_8753);
and U9259 (N_9259,N_8675,N_8636);
or U9260 (N_9260,N_8827,N_8935);
nor U9261 (N_9261,N_8641,N_8593);
and U9262 (N_9262,N_8978,N_8684);
nor U9263 (N_9263,N_8718,N_8967);
nand U9264 (N_9264,N_8633,N_8817);
nand U9265 (N_9265,N_8524,N_8560);
and U9266 (N_9266,N_8884,N_8638);
xnor U9267 (N_9267,N_8940,N_8616);
nor U9268 (N_9268,N_8880,N_8760);
xnor U9269 (N_9269,N_8799,N_8678);
nand U9270 (N_9270,N_8545,N_8889);
xor U9271 (N_9271,N_8857,N_8952);
and U9272 (N_9272,N_8566,N_8713);
xor U9273 (N_9273,N_8649,N_8549);
nand U9274 (N_9274,N_8941,N_8847);
or U9275 (N_9275,N_8827,N_8777);
xor U9276 (N_9276,N_8829,N_8902);
nand U9277 (N_9277,N_8999,N_8509);
and U9278 (N_9278,N_8558,N_8788);
nand U9279 (N_9279,N_8715,N_8820);
and U9280 (N_9280,N_8955,N_8963);
and U9281 (N_9281,N_8969,N_8641);
nand U9282 (N_9282,N_8861,N_8676);
xnor U9283 (N_9283,N_8559,N_8513);
or U9284 (N_9284,N_8995,N_8890);
and U9285 (N_9285,N_8876,N_8614);
or U9286 (N_9286,N_8820,N_8568);
nand U9287 (N_9287,N_8931,N_8554);
nor U9288 (N_9288,N_8678,N_8956);
and U9289 (N_9289,N_8917,N_8726);
and U9290 (N_9290,N_8508,N_8804);
nand U9291 (N_9291,N_8944,N_8555);
nand U9292 (N_9292,N_8720,N_8679);
xor U9293 (N_9293,N_8512,N_8620);
nand U9294 (N_9294,N_8842,N_8973);
or U9295 (N_9295,N_8999,N_8532);
xnor U9296 (N_9296,N_8706,N_8939);
or U9297 (N_9297,N_8610,N_8745);
nand U9298 (N_9298,N_8995,N_8751);
and U9299 (N_9299,N_8740,N_8602);
and U9300 (N_9300,N_8516,N_8880);
or U9301 (N_9301,N_8806,N_8897);
or U9302 (N_9302,N_8743,N_8814);
xnor U9303 (N_9303,N_8736,N_8552);
nand U9304 (N_9304,N_8504,N_8543);
xnor U9305 (N_9305,N_8580,N_8972);
and U9306 (N_9306,N_8537,N_8622);
xnor U9307 (N_9307,N_8781,N_8636);
and U9308 (N_9308,N_8808,N_8532);
nand U9309 (N_9309,N_8793,N_8966);
nand U9310 (N_9310,N_8558,N_8859);
nor U9311 (N_9311,N_8555,N_8786);
nand U9312 (N_9312,N_8760,N_8915);
nand U9313 (N_9313,N_8500,N_8503);
nand U9314 (N_9314,N_8540,N_8676);
nor U9315 (N_9315,N_8990,N_8652);
or U9316 (N_9316,N_8531,N_8988);
nand U9317 (N_9317,N_8562,N_8870);
nand U9318 (N_9318,N_8513,N_8632);
and U9319 (N_9319,N_8549,N_8874);
or U9320 (N_9320,N_8832,N_8573);
nand U9321 (N_9321,N_8812,N_8509);
nand U9322 (N_9322,N_8977,N_8575);
or U9323 (N_9323,N_8550,N_8507);
and U9324 (N_9324,N_8778,N_8881);
or U9325 (N_9325,N_8875,N_8511);
or U9326 (N_9326,N_8898,N_8861);
and U9327 (N_9327,N_8868,N_8542);
or U9328 (N_9328,N_8805,N_8950);
nand U9329 (N_9329,N_8926,N_8986);
or U9330 (N_9330,N_8942,N_8775);
xor U9331 (N_9331,N_8579,N_8742);
and U9332 (N_9332,N_8753,N_8751);
nor U9333 (N_9333,N_8813,N_8536);
or U9334 (N_9334,N_8610,N_8539);
xor U9335 (N_9335,N_8867,N_8528);
xnor U9336 (N_9336,N_8730,N_8979);
nand U9337 (N_9337,N_8965,N_8856);
xnor U9338 (N_9338,N_8906,N_8992);
xor U9339 (N_9339,N_8607,N_8903);
nor U9340 (N_9340,N_8583,N_8983);
xnor U9341 (N_9341,N_8536,N_8918);
or U9342 (N_9342,N_8818,N_8553);
nand U9343 (N_9343,N_8673,N_8933);
nand U9344 (N_9344,N_8577,N_8696);
or U9345 (N_9345,N_8824,N_8955);
or U9346 (N_9346,N_8526,N_8629);
or U9347 (N_9347,N_8900,N_8743);
nand U9348 (N_9348,N_8632,N_8878);
nor U9349 (N_9349,N_8880,N_8841);
and U9350 (N_9350,N_8638,N_8652);
and U9351 (N_9351,N_8810,N_8827);
nor U9352 (N_9352,N_8982,N_8565);
nor U9353 (N_9353,N_8914,N_8927);
xnor U9354 (N_9354,N_8605,N_8897);
nor U9355 (N_9355,N_8674,N_8615);
or U9356 (N_9356,N_8779,N_8577);
nand U9357 (N_9357,N_8831,N_8739);
nor U9358 (N_9358,N_8740,N_8919);
xnor U9359 (N_9359,N_8762,N_8607);
nor U9360 (N_9360,N_8738,N_8826);
nand U9361 (N_9361,N_8973,N_8846);
and U9362 (N_9362,N_8999,N_8964);
nor U9363 (N_9363,N_8624,N_8641);
nand U9364 (N_9364,N_8685,N_8663);
xor U9365 (N_9365,N_8862,N_8684);
or U9366 (N_9366,N_8518,N_8761);
xnor U9367 (N_9367,N_8525,N_8631);
xor U9368 (N_9368,N_8957,N_8607);
or U9369 (N_9369,N_8581,N_8680);
nand U9370 (N_9370,N_8646,N_8740);
xor U9371 (N_9371,N_8656,N_8578);
or U9372 (N_9372,N_8799,N_8757);
nor U9373 (N_9373,N_8850,N_8720);
xor U9374 (N_9374,N_8933,N_8777);
xor U9375 (N_9375,N_8526,N_8639);
xor U9376 (N_9376,N_8561,N_8988);
and U9377 (N_9377,N_8825,N_8867);
nor U9378 (N_9378,N_8996,N_8571);
and U9379 (N_9379,N_8997,N_8850);
nor U9380 (N_9380,N_8930,N_8902);
nor U9381 (N_9381,N_8865,N_8761);
nand U9382 (N_9382,N_8915,N_8831);
and U9383 (N_9383,N_8936,N_8651);
nor U9384 (N_9384,N_8859,N_8935);
xor U9385 (N_9385,N_8930,N_8745);
and U9386 (N_9386,N_8863,N_8989);
nand U9387 (N_9387,N_8787,N_8864);
xnor U9388 (N_9388,N_8892,N_8750);
and U9389 (N_9389,N_8906,N_8825);
nor U9390 (N_9390,N_8600,N_8639);
nand U9391 (N_9391,N_8852,N_8841);
nand U9392 (N_9392,N_8561,N_8717);
nor U9393 (N_9393,N_8639,N_8819);
nor U9394 (N_9394,N_8501,N_8840);
or U9395 (N_9395,N_8723,N_8955);
and U9396 (N_9396,N_8600,N_8566);
xor U9397 (N_9397,N_8841,N_8807);
or U9398 (N_9398,N_8773,N_8586);
and U9399 (N_9399,N_8817,N_8801);
or U9400 (N_9400,N_8981,N_8548);
and U9401 (N_9401,N_8735,N_8989);
and U9402 (N_9402,N_8515,N_8555);
xnor U9403 (N_9403,N_8980,N_8814);
nand U9404 (N_9404,N_8995,N_8673);
xnor U9405 (N_9405,N_8592,N_8700);
xnor U9406 (N_9406,N_8974,N_8543);
nand U9407 (N_9407,N_8911,N_8733);
or U9408 (N_9408,N_8639,N_8723);
or U9409 (N_9409,N_8586,N_8689);
and U9410 (N_9410,N_8843,N_8802);
xnor U9411 (N_9411,N_8545,N_8928);
nand U9412 (N_9412,N_8713,N_8753);
and U9413 (N_9413,N_8994,N_8854);
or U9414 (N_9414,N_8725,N_8960);
or U9415 (N_9415,N_8559,N_8527);
nor U9416 (N_9416,N_8893,N_8631);
xnor U9417 (N_9417,N_8923,N_8554);
nand U9418 (N_9418,N_8541,N_8561);
xnor U9419 (N_9419,N_8794,N_8625);
nor U9420 (N_9420,N_8516,N_8768);
or U9421 (N_9421,N_8846,N_8605);
and U9422 (N_9422,N_8827,N_8867);
and U9423 (N_9423,N_8605,N_8767);
and U9424 (N_9424,N_8733,N_8624);
and U9425 (N_9425,N_8954,N_8699);
nor U9426 (N_9426,N_8931,N_8720);
xor U9427 (N_9427,N_8516,N_8863);
and U9428 (N_9428,N_8987,N_8548);
xnor U9429 (N_9429,N_8770,N_8618);
and U9430 (N_9430,N_8887,N_8526);
xnor U9431 (N_9431,N_8949,N_8925);
or U9432 (N_9432,N_8771,N_8745);
and U9433 (N_9433,N_8927,N_8820);
xor U9434 (N_9434,N_8622,N_8970);
or U9435 (N_9435,N_8546,N_8928);
and U9436 (N_9436,N_8644,N_8614);
nand U9437 (N_9437,N_8749,N_8649);
xnor U9438 (N_9438,N_8858,N_8693);
xnor U9439 (N_9439,N_8650,N_8612);
nand U9440 (N_9440,N_8922,N_8919);
and U9441 (N_9441,N_8569,N_8667);
or U9442 (N_9442,N_8518,N_8683);
xnor U9443 (N_9443,N_8668,N_8965);
nand U9444 (N_9444,N_8912,N_8670);
nand U9445 (N_9445,N_8850,N_8729);
or U9446 (N_9446,N_8675,N_8522);
and U9447 (N_9447,N_8695,N_8987);
and U9448 (N_9448,N_8928,N_8818);
and U9449 (N_9449,N_8574,N_8652);
nor U9450 (N_9450,N_8803,N_8895);
xnor U9451 (N_9451,N_8925,N_8645);
or U9452 (N_9452,N_8533,N_8566);
or U9453 (N_9453,N_8912,N_8937);
or U9454 (N_9454,N_8621,N_8738);
xor U9455 (N_9455,N_8919,N_8965);
nand U9456 (N_9456,N_8614,N_8747);
nand U9457 (N_9457,N_8621,N_8732);
nor U9458 (N_9458,N_8984,N_8885);
or U9459 (N_9459,N_8537,N_8788);
and U9460 (N_9460,N_8630,N_8542);
nand U9461 (N_9461,N_8964,N_8943);
nand U9462 (N_9462,N_8781,N_8736);
and U9463 (N_9463,N_8595,N_8767);
nand U9464 (N_9464,N_8962,N_8620);
nand U9465 (N_9465,N_8670,N_8984);
nor U9466 (N_9466,N_8897,N_8999);
xnor U9467 (N_9467,N_8668,N_8776);
nor U9468 (N_9468,N_8759,N_8770);
nand U9469 (N_9469,N_8609,N_8672);
or U9470 (N_9470,N_8543,N_8732);
nor U9471 (N_9471,N_8837,N_8559);
or U9472 (N_9472,N_8758,N_8577);
nand U9473 (N_9473,N_8845,N_8993);
nand U9474 (N_9474,N_8533,N_8900);
and U9475 (N_9475,N_8543,N_8921);
or U9476 (N_9476,N_8882,N_8780);
nor U9477 (N_9477,N_8768,N_8582);
nand U9478 (N_9478,N_8638,N_8576);
nor U9479 (N_9479,N_8559,N_8698);
nand U9480 (N_9480,N_8837,N_8788);
nor U9481 (N_9481,N_8514,N_8561);
nor U9482 (N_9482,N_8543,N_8682);
nand U9483 (N_9483,N_8587,N_8685);
and U9484 (N_9484,N_8763,N_8897);
xor U9485 (N_9485,N_8652,N_8928);
and U9486 (N_9486,N_8687,N_8959);
or U9487 (N_9487,N_8909,N_8619);
or U9488 (N_9488,N_8880,N_8631);
xnor U9489 (N_9489,N_8576,N_8733);
nor U9490 (N_9490,N_8655,N_8851);
xor U9491 (N_9491,N_8628,N_8773);
or U9492 (N_9492,N_8953,N_8839);
or U9493 (N_9493,N_8892,N_8673);
nand U9494 (N_9494,N_8850,N_8681);
or U9495 (N_9495,N_8819,N_8893);
xor U9496 (N_9496,N_8802,N_8687);
nand U9497 (N_9497,N_8782,N_8745);
xnor U9498 (N_9498,N_8738,N_8579);
and U9499 (N_9499,N_8984,N_8655);
xnor U9500 (N_9500,N_9111,N_9402);
nand U9501 (N_9501,N_9366,N_9206);
nand U9502 (N_9502,N_9310,N_9261);
xor U9503 (N_9503,N_9121,N_9247);
nand U9504 (N_9504,N_9046,N_9107);
and U9505 (N_9505,N_9217,N_9409);
nand U9506 (N_9506,N_9249,N_9243);
nor U9507 (N_9507,N_9327,N_9049);
xnor U9508 (N_9508,N_9382,N_9087);
and U9509 (N_9509,N_9151,N_9275);
nand U9510 (N_9510,N_9127,N_9112);
xnor U9511 (N_9511,N_9152,N_9140);
nand U9512 (N_9512,N_9285,N_9317);
and U9513 (N_9513,N_9101,N_9043);
nor U9514 (N_9514,N_9018,N_9166);
xor U9515 (N_9515,N_9067,N_9244);
or U9516 (N_9516,N_9021,N_9191);
nor U9517 (N_9517,N_9408,N_9135);
nand U9518 (N_9518,N_9209,N_9444);
or U9519 (N_9519,N_9313,N_9024);
nor U9520 (N_9520,N_9042,N_9485);
xor U9521 (N_9521,N_9189,N_9429);
xnor U9522 (N_9522,N_9009,N_9404);
nand U9523 (N_9523,N_9267,N_9386);
xnor U9524 (N_9524,N_9268,N_9475);
nand U9525 (N_9525,N_9202,N_9023);
xnor U9526 (N_9526,N_9416,N_9484);
xor U9527 (N_9527,N_9194,N_9048);
and U9528 (N_9528,N_9224,N_9302);
xor U9529 (N_9529,N_9421,N_9155);
nand U9530 (N_9530,N_9073,N_9103);
nand U9531 (N_9531,N_9392,N_9447);
and U9532 (N_9532,N_9056,N_9315);
nor U9533 (N_9533,N_9329,N_9074);
nand U9534 (N_9534,N_9358,N_9040);
or U9535 (N_9535,N_9175,N_9367);
and U9536 (N_9536,N_9230,N_9430);
nand U9537 (N_9537,N_9352,N_9168);
or U9538 (N_9538,N_9470,N_9420);
xor U9539 (N_9539,N_9171,N_9034);
nand U9540 (N_9540,N_9381,N_9290);
nor U9541 (N_9541,N_9214,N_9344);
nand U9542 (N_9542,N_9493,N_9143);
xnor U9543 (N_9543,N_9241,N_9498);
xnor U9544 (N_9544,N_9343,N_9406);
nand U9545 (N_9545,N_9384,N_9086);
nor U9546 (N_9546,N_9089,N_9085);
xor U9547 (N_9547,N_9099,N_9237);
or U9548 (N_9548,N_9288,N_9026);
nand U9549 (N_9549,N_9170,N_9012);
nor U9550 (N_9550,N_9326,N_9466);
xor U9551 (N_9551,N_9298,N_9115);
nand U9552 (N_9552,N_9178,N_9004);
and U9553 (N_9553,N_9393,N_9277);
and U9554 (N_9554,N_9254,N_9307);
nor U9555 (N_9555,N_9279,N_9452);
or U9556 (N_9556,N_9010,N_9163);
xnor U9557 (N_9557,N_9453,N_9105);
xnor U9558 (N_9558,N_9177,N_9415);
xnor U9559 (N_9559,N_9192,N_9119);
nand U9560 (N_9560,N_9469,N_9499);
nor U9561 (N_9561,N_9422,N_9319);
and U9562 (N_9562,N_9014,N_9320);
nand U9563 (N_9563,N_9379,N_9066);
or U9564 (N_9564,N_9487,N_9193);
nor U9565 (N_9565,N_9272,N_9286);
nand U9566 (N_9566,N_9456,N_9443);
and U9567 (N_9567,N_9227,N_9492);
or U9568 (N_9568,N_9291,N_9325);
nor U9569 (N_9569,N_9308,N_9176);
xor U9570 (N_9570,N_9390,N_9208);
or U9571 (N_9571,N_9183,N_9281);
xnor U9572 (N_9572,N_9036,N_9207);
nand U9573 (N_9573,N_9410,N_9116);
nor U9574 (N_9574,N_9395,N_9013);
nor U9575 (N_9575,N_9118,N_9011);
xor U9576 (N_9576,N_9129,N_9084);
nand U9577 (N_9577,N_9486,N_9432);
nor U9578 (N_9578,N_9374,N_9083);
xor U9579 (N_9579,N_9231,N_9264);
and U9580 (N_9580,N_9394,N_9082);
and U9581 (N_9581,N_9333,N_9215);
nand U9582 (N_9582,N_9289,N_9365);
nor U9583 (N_9583,N_9239,N_9106);
nor U9584 (N_9584,N_9283,N_9134);
or U9585 (N_9585,N_9482,N_9445);
nor U9586 (N_9586,N_9007,N_9360);
or U9587 (N_9587,N_9180,N_9167);
nand U9588 (N_9588,N_9423,N_9258);
xnor U9589 (N_9589,N_9050,N_9158);
nor U9590 (N_9590,N_9147,N_9266);
nor U9591 (N_9591,N_9160,N_9433);
nand U9592 (N_9592,N_9462,N_9037);
or U9593 (N_9593,N_9001,N_9335);
nand U9594 (N_9594,N_9076,N_9132);
nand U9595 (N_9595,N_9095,N_9378);
xor U9596 (N_9596,N_9376,N_9490);
nor U9597 (N_9597,N_9297,N_9117);
or U9598 (N_9598,N_9156,N_9269);
and U9599 (N_9599,N_9454,N_9077);
xor U9600 (N_9600,N_9448,N_9164);
and U9601 (N_9601,N_9091,N_9015);
nor U9602 (N_9602,N_9041,N_9293);
nor U9603 (N_9603,N_9418,N_9185);
xor U9604 (N_9604,N_9491,N_9441);
and U9605 (N_9605,N_9316,N_9424);
and U9606 (N_9606,N_9232,N_9383);
nor U9607 (N_9607,N_9407,N_9350);
xnor U9608 (N_9608,N_9022,N_9030);
nor U9609 (N_9609,N_9380,N_9070);
nor U9610 (N_9610,N_9186,N_9341);
nand U9611 (N_9611,N_9033,N_9114);
xor U9612 (N_9612,N_9346,N_9262);
or U9613 (N_9613,N_9439,N_9304);
or U9614 (N_9614,N_9172,N_9467);
or U9615 (N_9615,N_9057,N_9081);
nand U9616 (N_9616,N_9233,N_9228);
and U9617 (N_9617,N_9354,N_9045);
nor U9618 (N_9618,N_9110,N_9252);
xnor U9619 (N_9619,N_9436,N_9154);
and U9620 (N_9620,N_9385,N_9100);
nor U9621 (N_9621,N_9488,N_9413);
or U9622 (N_9622,N_9223,N_9179);
nand U9623 (N_9623,N_9200,N_9016);
or U9624 (N_9624,N_9460,N_9464);
nand U9625 (N_9625,N_9075,N_9032);
nand U9626 (N_9626,N_9028,N_9002);
nand U9627 (N_9627,N_9065,N_9256);
nor U9628 (N_9628,N_9027,N_9356);
xor U9629 (N_9629,N_9145,N_9113);
nor U9630 (N_9630,N_9280,N_9238);
nand U9631 (N_9631,N_9161,N_9006);
nor U9632 (N_9632,N_9124,N_9338);
nand U9633 (N_9633,N_9332,N_9093);
nor U9634 (N_9634,N_9182,N_9403);
and U9635 (N_9635,N_9199,N_9253);
nand U9636 (N_9636,N_9351,N_9483);
xor U9637 (N_9637,N_9039,N_9471);
xor U9638 (N_9638,N_9094,N_9072);
nand U9639 (N_9639,N_9062,N_9029);
or U9640 (N_9640,N_9157,N_9468);
xnor U9641 (N_9641,N_9052,N_9263);
nand U9642 (N_9642,N_9148,N_9440);
nand U9643 (N_9643,N_9031,N_9340);
nor U9644 (N_9644,N_9273,N_9146);
nor U9645 (N_9645,N_9188,N_9400);
xnor U9646 (N_9646,N_9497,N_9229);
nor U9647 (N_9647,N_9349,N_9477);
and U9648 (N_9648,N_9345,N_9035);
nor U9649 (N_9649,N_9153,N_9270);
nor U9650 (N_9650,N_9248,N_9125);
xor U9651 (N_9651,N_9219,N_9292);
xor U9652 (N_9652,N_9080,N_9213);
or U9653 (N_9653,N_9435,N_9417);
nand U9654 (N_9654,N_9060,N_9159);
xnor U9655 (N_9655,N_9481,N_9071);
nor U9656 (N_9656,N_9278,N_9328);
nor U9657 (N_9657,N_9398,N_9479);
nand U9658 (N_9658,N_9449,N_9212);
xor U9659 (N_9659,N_9437,N_9296);
nand U9660 (N_9660,N_9412,N_9226);
nand U9661 (N_9661,N_9257,N_9184);
or U9662 (N_9662,N_9434,N_9122);
nand U9663 (N_9663,N_9210,N_9342);
and U9664 (N_9664,N_9299,N_9123);
and U9665 (N_9665,N_9051,N_9388);
and U9666 (N_9666,N_9368,N_9088);
and U9667 (N_9667,N_9419,N_9369);
xnor U9668 (N_9668,N_9245,N_9323);
and U9669 (N_9669,N_9274,N_9405);
or U9670 (N_9670,N_9090,N_9427);
and U9671 (N_9671,N_9098,N_9187);
nor U9672 (N_9672,N_9054,N_9181);
and U9673 (N_9673,N_9139,N_9204);
or U9674 (N_9674,N_9203,N_9355);
nand U9675 (N_9675,N_9225,N_9331);
nor U9676 (N_9676,N_9472,N_9311);
nand U9677 (N_9677,N_9463,N_9334);
xnor U9678 (N_9678,N_9426,N_9008);
or U9679 (N_9679,N_9138,N_9330);
and U9680 (N_9680,N_9240,N_9205);
or U9681 (N_9681,N_9120,N_9372);
xnor U9682 (N_9682,N_9260,N_9347);
nor U9683 (N_9683,N_9431,N_9371);
xnor U9684 (N_9684,N_9038,N_9130);
xor U9685 (N_9685,N_9251,N_9461);
and U9686 (N_9686,N_9465,N_9321);
xor U9687 (N_9687,N_9312,N_9020);
nand U9688 (N_9688,N_9473,N_9142);
xnor U9689 (N_9689,N_9457,N_9190);
and U9690 (N_9690,N_9496,N_9357);
and U9691 (N_9691,N_9019,N_9414);
and U9692 (N_9692,N_9364,N_9373);
xnor U9693 (N_9693,N_9389,N_9494);
xnor U9694 (N_9694,N_9391,N_9131);
nor U9695 (N_9695,N_9450,N_9149);
or U9696 (N_9696,N_9362,N_9102);
nor U9697 (N_9697,N_9195,N_9211);
xor U9698 (N_9698,N_9476,N_9198);
xor U9699 (N_9699,N_9336,N_9282);
nand U9700 (N_9700,N_9144,N_9220);
nand U9701 (N_9701,N_9458,N_9363);
nand U9702 (N_9702,N_9162,N_9305);
nand U9703 (N_9703,N_9339,N_9459);
nor U9704 (N_9704,N_9061,N_9397);
nand U9705 (N_9705,N_9000,N_9265);
or U9706 (N_9706,N_9411,N_9318);
nor U9707 (N_9707,N_9303,N_9174);
or U9708 (N_9708,N_9235,N_9387);
nand U9709 (N_9709,N_9401,N_9255);
or U9710 (N_9710,N_9300,N_9455);
nand U9711 (N_9711,N_9322,N_9474);
or U9712 (N_9712,N_9495,N_9047);
and U9713 (N_9713,N_9221,N_9246);
nor U9714 (N_9714,N_9294,N_9348);
nand U9715 (N_9715,N_9069,N_9337);
and U9716 (N_9716,N_9306,N_9063);
nand U9717 (N_9717,N_9137,N_9092);
nand U9718 (N_9718,N_9324,N_9058);
nor U9719 (N_9719,N_9242,N_9222);
xor U9720 (N_9720,N_9096,N_9287);
and U9721 (N_9721,N_9314,N_9309);
or U9722 (N_9722,N_9250,N_9399);
or U9723 (N_9723,N_9271,N_9442);
nand U9724 (N_9724,N_9059,N_9017);
xor U9725 (N_9725,N_9428,N_9108);
xnor U9726 (N_9726,N_9377,N_9375);
and U9727 (N_9727,N_9295,N_9259);
xnor U9728 (N_9728,N_9197,N_9451);
xnor U9729 (N_9729,N_9201,N_9003);
and U9730 (N_9730,N_9425,N_9109);
or U9731 (N_9731,N_9128,N_9480);
xor U9732 (N_9732,N_9079,N_9173);
nor U9733 (N_9733,N_9136,N_9361);
or U9734 (N_9734,N_9353,N_9104);
and U9735 (N_9735,N_9005,N_9044);
nor U9736 (N_9736,N_9216,N_9025);
nor U9737 (N_9737,N_9165,N_9370);
nor U9738 (N_9738,N_9218,N_9301);
nor U9739 (N_9739,N_9097,N_9359);
nor U9740 (N_9740,N_9126,N_9169);
nand U9741 (N_9741,N_9055,N_9068);
nor U9742 (N_9742,N_9234,N_9438);
and U9743 (N_9743,N_9284,N_9053);
nand U9744 (N_9744,N_9064,N_9141);
or U9745 (N_9745,N_9078,N_9236);
or U9746 (N_9746,N_9396,N_9150);
and U9747 (N_9747,N_9133,N_9276);
nor U9748 (N_9748,N_9446,N_9196);
xnor U9749 (N_9749,N_9489,N_9478);
nor U9750 (N_9750,N_9147,N_9380);
xnor U9751 (N_9751,N_9452,N_9074);
or U9752 (N_9752,N_9316,N_9379);
nor U9753 (N_9753,N_9469,N_9069);
xnor U9754 (N_9754,N_9139,N_9294);
nor U9755 (N_9755,N_9020,N_9220);
nand U9756 (N_9756,N_9363,N_9302);
xnor U9757 (N_9757,N_9271,N_9391);
or U9758 (N_9758,N_9191,N_9324);
xor U9759 (N_9759,N_9255,N_9459);
or U9760 (N_9760,N_9447,N_9229);
xor U9761 (N_9761,N_9498,N_9289);
nand U9762 (N_9762,N_9382,N_9021);
and U9763 (N_9763,N_9276,N_9177);
and U9764 (N_9764,N_9437,N_9464);
nand U9765 (N_9765,N_9094,N_9481);
xor U9766 (N_9766,N_9191,N_9468);
nand U9767 (N_9767,N_9423,N_9436);
nor U9768 (N_9768,N_9233,N_9094);
or U9769 (N_9769,N_9390,N_9392);
nor U9770 (N_9770,N_9350,N_9199);
nor U9771 (N_9771,N_9304,N_9362);
and U9772 (N_9772,N_9122,N_9050);
nor U9773 (N_9773,N_9466,N_9176);
or U9774 (N_9774,N_9168,N_9140);
or U9775 (N_9775,N_9104,N_9043);
or U9776 (N_9776,N_9445,N_9439);
nor U9777 (N_9777,N_9223,N_9260);
nor U9778 (N_9778,N_9297,N_9361);
or U9779 (N_9779,N_9062,N_9192);
xor U9780 (N_9780,N_9201,N_9269);
nand U9781 (N_9781,N_9266,N_9141);
nand U9782 (N_9782,N_9211,N_9021);
xor U9783 (N_9783,N_9310,N_9112);
nand U9784 (N_9784,N_9474,N_9498);
or U9785 (N_9785,N_9040,N_9282);
nor U9786 (N_9786,N_9334,N_9356);
nand U9787 (N_9787,N_9036,N_9396);
xnor U9788 (N_9788,N_9118,N_9404);
and U9789 (N_9789,N_9370,N_9353);
xnor U9790 (N_9790,N_9373,N_9332);
or U9791 (N_9791,N_9456,N_9479);
nand U9792 (N_9792,N_9185,N_9048);
xor U9793 (N_9793,N_9211,N_9152);
or U9794 (N_9794,N_9415,N_9372);
and U9795 (N_9795,N_9375,N_9086);
nor U9796 (N_9796,N_9186,N_9412);
nor U9797 (N_9797,N_9214,N_9112);
nor U9798 (N_9798,N_9370,N_9115);
or U9799 (N_9799,N_9112,N_9223);
and U9800 (N_9800,N_9222,N_9357);
or U9801 (N_9801,N_9340,N_9221);
and U9802 (N_9802,N_9381,N_9115);
xnor U9803 (N_9803,N_9470,N_9165);
nand U9804 (N_9804,N_9182,N_9056);
xnor U9805 (N_9805,N_9415,N_9462);
nor U9806 (N_9806,N_9083,N_9329);
nand U9807 (N_9807,N_9244,N_9206);
and U9808 (N_9808,N_9422,N_9344);
nand U9809 (N_9809,N_9476,N_9039);
nor U9810 (N_9810,N_9273,N_9058);
xor U9811 (N_9811,N_9226,N_9450);
nor U9812 (N_9812,N_9080,N_9327);
or U9813 (N_9813,N_9075,N_9411);
xor U9814 (N_9814,N_9348,N_9423);
and U9815 (N_9815,N_9448,N_9481);
and U9816 (N_9816,N_9388,N_9219);
nand U9817 (N_9817,N_9393,N_9174);
nand U9818 (N_9818,N_9034,N_9264);
or U9819 (N_9819,N_9182,N_9319);
or U9820 (N_9820,N_9386,N_9487);
xor U9821 (N_9821,N_9220,N_9367);
and U9822 (N_9822,N_9305,N_9195);
xnor U9823 (N_9823,N_9015,N_9328);
xnor U9824 (N_9824,N_9092,N_9255);
nand U9825 (N_9825,N_9387,N_9037);
and U9826 (N_9826,N_9368,N_9373);
nand U9827 (N_9827,N_9260,N_9410);
or U9828 (N_9828,N_9238,N_9330);
xor U9829 (N_9829,N_9074,N_9243);
nand U9830 (N_9830,N_9331,N_9472);
xnor U9831 (N_9831,N_9407,N_9361);
or U9832 (N_9832,N_9361,N_9193);
nand U9833 (N_9833,N_9210,N_9377);
xnor U9834 (N_9834,N_9031,N_9188);
or U9835 (N_9835,N_9496,N_9020);
nand U9836 (N_9836,N_9343,N_9283);
and U9837 (N_9837,N_9459,N_9433);
nand U9838 (N_9838,N_9280,N_9166);
or U9839 (N_9839,N_9347,N_9221);
xnor U9840 (N_9840,N_9218,N_9224);
nand U9841 (N_9841,N_9001,N_9205);
nor U9842 (N_9842,N_9028,N_9164);
and U9843 (N_9843,N_9466,N_9152);
or U9844 (N_9844,N_9214,N_9237);
nor U9845 (N_9845,N_9302,N_9486);
or U9846 (N_9846,N_9377,N_9001);
and U9847 (N_9847,N_9088,N_9236);
nor U9848 (N_9848,N_9382,N_9254);
or U9849 (N_9849,N_9115,N_9197);
and U9850 (N_9850,N_9085,N_9078);
xor U9851 (N_9851,N_9467,N_9176);
nand U9852 (N_9852,N_9089,N_9422);
xor U9853 (N_9853,N_9101,N_9206);
nor U9854 (N_9854,N_9469,N_9240);
nor U9855 (N_9855,N_9499,N_9289);
nand U9856 (N_9856,N_9125,N_9153);
or U9857 (N_9857,N_9093,N_9234);
or U9858 (N_9858,N_9337,N_9149);
or U9859 (N_9859,N_9396,N_9261);
nand U9860 (N_9860,N_9469,N_9277);
and U9861 (N_9861,N_9377,N_9084);
or U9862 (N_9862,N_9290,N_9415);
and U9863 (N_9863,N_9350,N_9414);
xnor U9864 (N_9864,N_9419,N_9348);
nand U9865 (N_9865,N_9011,N_9141);
xor U9866 (N_9866,N_9267,N_9054);
nand U9867 (N_9867,N_9305,N_9360);
xnor U9868 (N_9868,N_9183,N_9279);
nand U9869 (N_9869,N_9063,N_9272);
nand U9870 (N_9870,N_9063,N_9200);
and U9871 (N_9871,N_9188,N_9192);
or U9872 (N_9872,N_9397,N_9281);
nor U9873 (N_9873,N_9106,N_9063);
or U9874 (N_9874,N_9324,N_9031);
nor U9875 (N_9875,N_9260,N_9083);
nor U9876 (N_9876,N_9113,N_9048);
and U9877 (N_9877,N_9350,N_9013);
and U9878 (N_9878,N_9296,N_9421);
and U9879 (N_9879,N_9112,N_9097);
nor U9880 (N_9880,N_9243,N_9347);
nor U9881 (N_9881,N_9145,N_9237);
nand U9882 (N_9882,N_9105,N_9266);
and U9883 (N_9883,N_9262,N_9111);
nor U9884 (N_9884,N_9340,N_9430);
or U9885 (N_9885,N_9333,N_9038);
or U9886 (N_9886,N_9269,N_9028);
nor U9887 (N_9887,N_9373,N_9470);
and U9888 (N_9888,N_9079,N_9180);
and U9889 (N_9889,N_9426,N_9424);
nor U9890 (N_9890,N_9488,N_9096);
nand U9891 (N_9891,N_9345,N_9264);
or U9892 (N_9892,N_9432,N_9062);
nor U9893 (N_9893,N_9141,N_9441);
nand U9894 (N_9894,N_9209,N_9168);
or U9895 (N_9895,N_9496,N_9281);
xor U9896 (N_9896,N_9230,N_9131);
and U9897 (N_9897,N_9176,N_9324);
xnor U9898 (N_9898,N_9017,N_9044);
and U9899 (N_9899,N_9426,N_9483);
xor U9900 (N_9900,N_9116,N_9261);
xor U9901 (N_9901,N_9458,N_9419);
or U9902 (N_9902,N_9209,N_9115);
nand U9903 (N_9903,N_9301,N_9304);
and U9904 (N_9904,N_9228,N_9144);
or U9905 (N_9905,N_9228,N_9254);
or U9906 (N_9906,N_9310,N_9276);
nand U9907 (N_9907,N_9332,N_9446);
xnor U9908 (N_9908,N_9470,N_9310);
xnor U9909 (N_9909,N_9252,N_9423);
nor U9910 (N_9910,N_9011,N_9468);
and U9911 (N_9911,N_9196,N_9105);
and U9912 (N_9912,N_9373,N_9158);
nand U9913 (N_9913,N_9101,N_9178);
nand U9914 (N_9914,N_9143,N_9288);
or U9915 (N_9915,N_9088,N_9126);
xnor U9916 (N_9916,N_9132,N_9271);
xor U9917 (N_9917,N_9451,N_9024);
and U9918 (N_9918,N_9292,N_9267);
or U9919 (N_9919,N_9215,N_9422);
nand U9920 (N_9920,N_9487,N_9076);
and U9921 (N_9921,N_9410,N_9191);
nor U9922 (N_9922,N_9365,N_9235);
and U9923 (N_9923,N_9397,N_9220);
nand U9924 (N_9924,N_9160,N_9245);
or U9925 (N_9925,N_9242,N_9368);
nor U9926 (N_9926,N_9369,N_9370);
or U9927 (N_9927,N_9477,N_9326);
xor U9928 (N_9928,N_9074,N_9204);
xnor U9929 (N_9929,N_9365,N_9045);
and U9930 (N_9930,N_9099,N_9009);
nor U9931 (N_9931,N_9177,N_9365);
nand U9932 (N_9932,N_9387,N_9293);
or U9933 (N_9933,N_9263,N_9214);
nor U9934 (N_9934,N_9057,N_9255);
xnor U9935 (N_9935,N_9062,N_9108);
nand U9936 (N_9936,N_9318,N_9426);
or U9937 (N_9937,N_9310,N_9018);
nand U9938 (N_9938,N_9308,N_9272);
nand U9939 (N_9939,N_9215,N_9219);
xor U9940 (N_9940,N_9104,N_9468);
xor U9941 (N_9941,N_9499,N_9449);
nand U9942 (N_9942,N_9312,N_9117);
or U9943 (N_9943,N_9499,N_9165);
or U9944 (N_9944,N_9215,N_9161);
and U9945 (N_9945,N_9265,N_9124);
or U9946 (N_9946,N_9075,N_9178);
and U9947 (N_9947,N_9105,N_9112);
nor U9948 (N_9948,N_9263,N_9159);
or U9949 (N_9949,N_9196,N_9134);
xnor U9950 (N_9950,N_9492,N_9109);
nand U9951 (N_9951,N_9134,N_9142);
nand U9952 (N_9952,N_9255,N_9346);
nand U9953 (N_9953,N_9106,N_9290);
xor U9954 (N_9954,N_9098,N_9185);
and U9955 (N_9955,N_9083,N_9095);
nand U9956 (N_9956,N_9091,N_9151);
nand U9957 (N_9957,N_9453,N_9096);
nor U9958 (N_9958,N_9000,N_9220);
and U9959 (N_9959,N_9348,N_9436);
xnor U9960 (N_9960,N_9193,N_9044);
nand U9961 (N_9961,N_9491,N_9074);
nand U9962 (N_9962,N_9336,N_9374);
xor U9963 (N_9963,N_9035,N_9028);
nand U9964 (N_9964,N_9379,N_9065);
nor U9965 (N_9965,N_9466,N_9458);
and U9966 (N_9966,N_9179,N_9052);
nand U9967 (N_9967,N_9122,N_9164);
nor U9968 (N_9968,N_9446,N_9389);
xor U9969 (N_9969,N_9097,N_9091);
xnor U9970 (N_9970,N_9085,N_9253);
or U9971 (N_9971,N_9328,N_9414);
xnor U9972 (N_9972,N_9072,N_9194);
and U9973 (N_9973,N_9150,N_9402);
xnor U9974 (N_9974,N_9467,N_9026);
nand U9975 (N_9975,N_9323,N_9365);
xnor U9976 (N_9976,N_9235,N_9306);
nor U9977 (N_9977,N_9123,N_9317);
nand U9978 (N_9978,N_9074,N_9429);
nand U9979 (N_9979,N_9243,N_9435);
nor U9980 (N_9980,N_9049,N_9012);
and U9981 (N_9981,N_9497,N_9159);
xnor U9982 (N_9982,N_9246,N_9461);
nor U9983 (N_9983,N_9008,N_9198);
nor U9984 (N_9984,N_9487,N_9148);
nor U9985 (N_9985,N_9275,N_9326);
xnor U9986 (N_9986,N_9326,N_9370);
nand U9987 (N_9987,N_9125,N_9387);
nand U9988 (N_9988,N_9000,N_9305);
nor U9989 (N_9989,N_9024,N_9180);
and U9990 (N_9990,N_9208,N_9133);
nand U9991 (N_9991,N_9352,N_9006);
and U9992 (N_9992,N_9145,N_9361);
xor U9993 (N_9993,N_9346,N_9138);
or U9994 (N_9994,N_9230,N_9395);
and U9995 (N_9995,N_9212,N_9115);
nand U9996 (N_9996,N_9181,N_9410);
nor U9997 (N_9997,N_9362,N_9124);
nand U9998 (N_9998,N_9365,N_9256);
nand U9999 (N_9999,N_9278,N_9211);
nand U10000 (N_10000,N_9884,N_9726);
nand U10001 (N_10001,N_9710,N_9854);
or U10002 (N_10002,N_9679,N_9993);
or U10003 (N_10003,N_9719,N_9590);
and U10004 (N_10004,N_9800,N_9995);
nor U10005 (N_10005,N_9727,N_9621);
nand U10006 (N_10006,N_9616,N_9777);
nor U10007 (N_10007,N_9694,N_9661);
nand U10008 (N_10008,N_9671,N_9909);
nand U10009 (N_10009,N_9957,N_9749);
xor U10010 (N_10010,N_9662,N_9807);
and U10011 (N_10011,N_9925,N_9723);
xor U10012 (N_10012,N_9740,N_9778);
nand U10013 (N_10013,N_9941,N_9891);
and U10014 (N_10014,N_9715,N_9663);
xor U10015 (N_10015,N_9923,N_9522);
nand U10016 (N_10016,N_9573,N_9689);
or U10017 (N_10017,N_9893,N_9823);
xnor U10018 (N_10018,N_9566,N_9978);
nor U10019 (N_10019,N_9652,N_9531);
nand U10020 (N_10020,N_9561,N_9655);
and U10021 (N_10021,N_9805,N_9820);
and U10022 (N_10022,N_9707,N_9812);
xor U10023 (N_10023,N_9587,N_9589);
xnor U10024 (N_10024,N_9792,N_9739);
or U10025 (N_10025,N_9708,N_9511);
nand U10026 (N_10026,N_9861,N_9610);
and U10027 (N_10027,N_9628,N_9956);
or U10028 (N_10028,N_9517,N_9967);
nor U10029 (N_10029,N_9542,N_9701);
and U10030 (N_10030,N_9819,N_9575);
xnor U10031 (N_10031,N_9580,N_9979);
nand U10032 (N_10032,N_9693,N_9874);
or U10033 (N_10033,N_9848,N_9545);
and U10034 (N_10034,N_9975,N_9653);
or U10035 (N_10035,N_9981,N_9798);
xor U10036 (N_10036,N_9834,N_9936);
and U10037 (N_10037,N_9548,N_9670);
nor U10038 (N_10038,N_9885,N_9878);
nand U10039 (N_10039,N_9674,N_9875);
and U10040 (N_10040,N_9571,N_9592);
nor U10041 (N_10041,N_9900,N_9976);
nand U10042 (N_10042,N_9583,N_9562);
or U10043 (N_10043,N_9998,N_9731);
nor U10044 (N_10044,N_9618,N_9504);
nand U10045 (N_10045,N_9572,N_9604);
nor U10046 (N_10046,N_9609,N_9700);
or U10047 (N_10047,N_9595,N_9619);
nor U10048 (N_10048,N_9530,N_9507);
nand U10049 (N_10049,N_9950,N_9990);
xor U10050 (N_10050,N_9747,N_9643);
nand U10051 (N_10051,N_9680,N_9744);
and U10052 (N_10052,N_9963,N_9793);
xor U10053 (N_10053,N_9540,N_9758);
xnor U10054 (N_10054,N_9804,N_9977);
and U10055 (N_10055,N_9980,N_9772);
or U10056 (N_10056,N_9912,N_9883);
and U10057 (N_10057,N_9702,N_9742);
xnor U10058 (N_10058,N_9968,N_9853);
nand U10059 (N_10059,N_9826,N_9965);
nand U10060 (N_10060,N_9879,N_9811);
nand U10061 (N_10061,N_9942,N_9829);
xnor U10062 (N_10062,N_9771,N_9533);
and U10063 (N_10063,N_9622,N_9565);
and U10064 (N_10064,N_9645,N_9905);
and U10065 (N_10065,N_9703,N_9728);
nand U10066 (N_10066,N_9928,N_9974);
or U10067 (N_10067,N_9781,N_9896);
xor U10068 (N_10068,N_9560,N_9871);
xor U10069 (N_10069,N_9596,N_9602);
xor U10070 (N_10070,N_9746,N_9847);
xnor U10071 (N_10071,N_9509,N_9922);
and U10072 (N_10072,N_9631,N_9765);
nand U10073 (N_10073,N_9852,N_9649);
and U10074 (N_10074,N_9784,N_9620);
and U10075 (N_10075,N_9924,N_9763);
nor U10076 (N_10076,N_9897,N_9822);
and U10077 (N_10077,N_9837,N_9770);
and U10078 (N_10078,N_9817,N_9872);
and U10079 (N_10079,N_9699,N_9555);
or U10080 (N_10080,N_9659,N_9697);
nor U10081 (N_10081,N_9717,N_9796);
and U10082 (N_10082,N_9557,N_9678);
and U10083 (N_10083,N_9667,N_9984);
xor U10084 (N_10084,N_9564,N_9598);
xor U10085 (N_10085,N_9868,N_9886);
nor U10086 (N_10086,N_9828,N_9532);
xnor U10087 (N_10087,N_9787,N_9791);
and U10088 (N_10088,N_9552,N_9790);
xnor U10089 (N_10089,N_9973,N_9913);
xnor U10090 (N_10090,N_9730,N_9529);
xor U10091 (N_10091,N_9937,N_9716);
xor U10092 (N_10092,N_9690,N_9558);
nor U10093 (N_10093,N_9762,N_9961);
xnor U10094 (N_10094,N_9753,N_9698);
nor U10095 (N_10095,N_9806,N_9623);
or U10096 (N_10096,N_9676,N_9944);
or U10097 (N_10097,N_9513,N_9563);
xnor U10098 (N_10098,N_9991,N_9989);
nor U10099 (N_10099,N_9982,N_9721);
and U10100 (N_10100,N_9514,N_9919);
xor U10101 (N_10101,N_9759,N_9752);
nor U10102 (N_10102,N_9684,N_9915);
and U10103 (N_10103,N_9794,N_9890);
nor U10104 (N_10104,N_9866,N_9613);
nand U10105 (N_10105,N_9988,N_9803);
nand U10106 (N_10106,N_9881,N_9786);
nor U10107 (N_10107,N_9855,N_9953);
nor U10108 (N_10108,N_9931,N_9783);
or U10109 (N_10109,N_9764,N_9551);
and U10110 (N_10110,N_9947,N_9642);
and U10111 (N_10111,N_9591,N_9748);
nand U10112 (N_10112,N_9999,N_9627);
nand U10113 (N_10113,N_9519,N_9683);
nor U10114 (N_10114,N_9775,N_9608);
nand U10115 (N_10115,N_9646,N_9756);
xnor U10116 (N_10116,N_9711,N_9525);
or U10117 (N_10117,N_9894,N_9789);
or U10118 (N_10118,N_9629,N_9994);
nor U10119 (N_10119,N_9932,N_9839);
nor U10120 (N_10120,N_9503,N_9594);
and U10121 (N_10121,N_9945,N_9538);
and U10122 (N_10122,N_9992,N_9766);
nand U10123 (N_10123,N_9718,N_9722);
nand U10124 (N_10124,N_9779,N_9506);
or U10125 (N_10125,N_9732,N_9996);
xnor U10126 (N_10126,N_9987,N_9750);
xnor U10127 (N_10127,N_9734,N_9810);
xor U10128 (N_10128,N_9933,N_9813);
xor U10129 (N_10129,N_9962,N_9949);
nor U10130 (N_10130,N_9851,N_9665);
nor U10131 (N_10131,N_9735,N_9971);
xor U10132 (N_10132,N_9910,N_9876);
nor U10133 (N_10133,N_9599,N_9640);
nand U10134 (N_10134,N_9677,N_9626);
nor U10135 (N_10135,N_9911,N_9773);
or U10136 (N_10136,N_9802,N_9939);
xor U10137 (N_10137,N_9835,N_9914);
xnor U10138 (N_10138,N_9669,N_9641);
or U10139 (N_10139,N_9743,N_9510);
xnor U10140 (N_10140,N_9808,N_9624);
nor U10141 (N_10141,N_9706,N_9559);
xnor U10142 (N_10142,N_9570,N_9658);
or U10143 (N_10143,N_9831,N_9569);
nand U10144 (N_10144,N_9768,N_9825);
or U10145 (N_10145,N_9859,N_9651);
or U10146 (N_10146,N_9568,N_9929);
nand U10147 (N_10147,N_9958,N_9755);
xnor U10148 (N_10148,N_9918,N_9880);
and U10149 (N_10149,N_9581,N_9774);
nand U10150 (N_10150,N_9654,N_9597);
xnor U10151 (N_10151,N_9741,N_9636);
xnor U10152 (N_10152,N_9867,N_9983);
or U10153 (N_10153,N_9537,N_9827);
nor U10154 (N_10154,N_9738,N_9712);
and U10155 (N_10155,N_9672,N_9769);
nand U10156 (N_10156,N_9902,N_9841);
xor U10157 (N_10157,N_9611,N_9660);
nor U10158 (N_10158,N_9901,N_9898);
or U10159 (N_10159,N_9857,N_9903);
nor U10160 (N_10160,N_9948,N_9632);
and U10161 (N_10161,N_9917,N_9985);
and U10162 (N_10162,N_9964,N_9795);
xnor U10163 (N_10163,N_9927,N_9724);
xnor U10164 (N_10164,N_9547,N_9585);
nand U10165 (N_10165,N_9668,N_9904);
nand U10166 (N_10166,N_9930,N_9567);
nand U10167 (N_10167,N_9960,N_9780);
and U10168 (N_10168,N_9926,N_9887);
or U10169 (N_10169,N_9695,N_9696);
or U10170 (N_10170,N_9846,N_9681);
or U10171 (N_10171,N_9554,N_9600);
and U10172 (N_10172,N_9954,N_9637);
nor U10173 (N_10173,N_9615,N_9970);
or U10174 (N_10174,N_9934,N_9785);
nand U10175 (N_10175,N_9832,N_9850);
nand U10176 (N_10176,N_9634,N_9729);
xor U10177 (N_10177,N_9951,N_9907);
nor U10178 (N_10178,N_9736,N_9704);
nor U10179 (N_10179,N_9997,N_9656);
nor U10180 (N_10180,N_9843,N_9916);
and U10181 (N_10181,N_9691,N_9809);
and U10182 (N_10182,N_9788,N_9675);
nor U10183 (N_10183,N_9844,N_9920);
or U10184 (N_10184,N_9577,N_9799);
xor U10185 (N_10185,N_9528,N_9574);
xnor U10186 (N_10186,N_9754,N_9539);
xor U10187 (N_10187,N_9638,N_9607);
or U10188 (N_10188,N_9849,N_9955);
or U10189 (N_10189,N_9972,N_9836);
nor U10190 (N_10190,N_9863,N_9524);
nand U10191 (N_10191,N_9761,N_9969);
and U10192 (N_10192,N_9523,N_9612);
nor U10193 (N_10193,N_9737,N_9639);
or U10194 (N_10194,N_9906,N_9521);
nand U10195 (N_10195,N_9685,N_9818);
xor U10196 (N_10196,N_9614,N_9873);
nand U10197 (N_10197,N_9688,N_9546);
nand U10198 (N_10198,N_9536,N_9544);
or U10199 (N_10199,N_9648,N_9518);
xnor U10200 (N_10200,N_9856,N_9865);
nor U10201 (N_10201,N_9888,N_9588);
and U10202 (N_10202,N_9657,N_9757);
xor U10203 (N_10203,N_9720,N_9801);
or U10204 (N_10204,N_9650,N_9733);
and U10205 (N_10205,N_9858,N_9860);
xor U10206 (N_10206,N_9635,N_9601);
xnor U10207 (N_10207,N_9705,N_9578);
and U10208 (N_10208,N_9593,N_9966);
or U10209 (N_10209,N_9633,N_9814);
nand U10210 (N_10210,N_9797,N_9842);
or U10211 (N_10211,N_9556,N_9606);
or U10212 (N_10212,N_9745,N_9776);
or U10213 (N_10213,N_9647,N_9520);
nor U10214 (N_10214,N_9840,N_9673);
or U10215 (N_10215,N_9869,N_9664);
or U10216 (N_10216,N_9549,N_9833);
or U10217 (N_10217,N_9725,N_9935);
xor U10218 (N_10218,N_9692,N_9899);
nand U10219 (N_10219,N_9502,N_9877);
and U10220 (N_10220,N_9644,N_9959);
nand U10221 (N_10221,N_9870,N_9625);
or U10222 (N_10222,N_9682,N_9543);
or U10223 (N_10223,N_9576,N_9892);
nand U10224 (N_10224,N_9527,N_9882);
nor U10225 (N_10225,N_9824,N_9952);
or U10226 (N_10226,N_9782,N_9862);
or U10227 (N_10227,N_9686,N_9889);
nor U10228 (N_10228,N_9586,N_9751);
xor U10229 (N_10229,N_9541,N_9550);
nor U10230 (N_10230,N_9943,N_9534);
xor U10231 (N_10231,N_9845,N_9500);
and U10232 (N_10232,N_9526,N_9864);
nand U10233 (N_10233,N_9986,N_9821);
nor U10234 (N_10234,N_9535,N_9713);
or U10235 (N_10235,N_9895,N_9630);
nor U10236 (N_10236,N_9605,N_9709);
nand U10237 (N_10237,N_9908,N_9830);
and U10238 (N_10238,N_9501,N_9767);
xor U10239 (N_10239,N_9946,N_9816);
nand U10240 (N_10240,N_9940,N_9579);
and U10241 (N_10241,N_9687,N_9505);
xor U10242 (N_10242,N_9516,N_9921);
nand U10243 (N_10243,N_9515,N_9508);
xnor U10244 (N_10244,N_9815,N_9582);
nand U10245 (N_10245,N_9714,N_9666);
xor U10246 (N_10246,N_9512,N_9617);
xnor U10247 (N_10247,N_9838,N_9603);
or U10248 (N_10248,N_9584,N_9938);
nand U10249 (N_10249,N_9760,N_9553);
xor U10250 (N_10250,N_9801,N_9779);
and U10251 (N_10251,N_9522,N_9847);
xnor U10252 (N_10252,N_9753,N_9906);
nand U10253 (N_10253,N_9609,N_9585);
xnor U10254 (N_10254,N_9584,N_9791);
and U10255 (N_10255,N_9815,N_9852);
nand U10256 (N_10256,N_9599,N_9712);
nor U10257 (N_10257,N_9685,N_9696);
and U10258 (N_10258,N_9716,N_9598);
xnor U10259 (N_10259,N_9511,N_9769);
or U10260 (N_10260,N_9743,N_9583);
and U10261 (N_10261,N_9856,N_9656);
xnor U10262 (N_10262,N_9549,N_9966);
or U10263 (N_10263,N_9959,N_9802);
nand U10264 (N_10264,N_9882,N_9666);
nor U10265 (N_10265,N_9522,N_9920);
and U10266 (N_10266,N_9714,N_9845);
xor U10267 (N_10267,N_9852,N_9950);
or U10268 (N_10268,N_9936,N_9627);
or U10269 (N_10269,N_9611,N_9995);
nand U10270 (N_10270,N_9716,N_9597);
and U10271 (N_10271,N_9706,N_9914);
or U10272 (N_10272,N_9590,N_9804);
xnor U10273 (N_10273,N_9659,N_9732);
xnor U10274 (N_10274,N_9903,N_9945);
xnor U10275 (N_10275,N_9749,N_9559);
or U10276 (N_10276,N_9711,N_9644);
and U10277 (N_10277,N_9533,N_9600);
nand U10278 (N_10278,N_9714,N_9902);
nand U10279 (N_10279,N_9509,N_9760);
nor U10280 (N_10280,N_9665,N_9554);
or U10281 (N_10281,N_9878,N_9622);
and U10282 (N_10282,N_9598,N_9643);
nor U10283 (N_10283,N_9642,N_9752);
xor U10284 (N_10284,N_9815,N_9627);
or U10285 (N_10285,N_9541,N_9778);
xnor U10286 (N_10286,N_9815,N_9565);
and U10287 (N_10287,N_9764,N_9654);
or U10288 (N_10288,N_9934,N_9919);
xnor U10289 (N_10289,N_9681,N_9586);
nor U10290 (N_10290,N_9668,N_9724);
nor U10291 (N_10291,N_9538,N_9786);
and U10292 (N_10292,N_9665,N_9708);
or U10293 (N_10293,N_9590,N_9725);
or U10294 (N_10294,N_9959,N_9625);
or U10295 (N_10295,N_9645,N_9614);
nand U10296 (N_10296,N_9871,N_9878);
and U10297 (N_10297,N_9954,N_9651);
nand U10298 (N_10298,N_9663,N_9928);
xor U10299 (N_10299,N_9509,N_9766);
nor U10300 (N_10300,N_9912,N_9556);
nand U10301 (N_10301,N_9582,N_9849);
nand U10302 (N_10302,N_9787,N_9835);
or U10303 (N_10303,N_9910,N_9516);
xor U10304 (N_10304,N_9507,N_9721);
and U10305 (N_10305,N_9808,N_9526);
or U10306 (N_10306,N_9749,N_9730);
nand U10307 (N_10307,N_9884,N_9731);
nor U10308 (N_10308,N_9610,N_9800);
xnor U10309 (N_10309,N_9834,N_9587);
nor U10310 (N_10310,N_9593,N_9713);
or U10311 (N_10311,N_9527,N_9753);
xor U10312 (N_10312,N_9621,N_9915);
or U10313 (N_10313,N_9980,N_9770);
xor U10314 (N_10314,N_9507,N_9786);
xor U10315 (N_10315,N_9693,N_9669);
nor U10316 (N_10316,N_9849,N_9753);
or U10317 (N_10317,N_9574,N_9712);
nor U10318 (N_10318,N_9846,N_9878);
or U10319 (N_10319,N_9574,N_9585);
or U10320 (N_10320,N_9680,N_9847);
or U10321 (N_10321,N_9863,N_9725);
nand U10322 (N_10322,N_9525,N_9519);
or U10323 (N_10323,N_9915,N_9919);
nor U10324 (N_10324,N_9524,N_9708);
xnor U10325 (N_10325,N_9897,N_9986);
nor U10326 (N_10326,N_9652,N_9877);
or U10327 (N_10327,N_9958,N_9938);
nor U10328 (N_10328,N_9919,N_9898);
xnor U10329 (N_10329,N_9864,N_9758);
nor U10330 (N_10330,N_9950,N_9528);
nand U10331 (N_10331,N_9527,N_9725);
and U10332 (N_10332,N_9810,N_9602);
and U10333 (N_10333,N_9907,N_9965);
nand U10334 (N_10334,N_9683,N_9736);
or U10335 (N_10335,N_9605,N_9522);
nand U10336 (N_10336,N_9573,N_9727);
xnor U10337 (N_10337,N_9985,N_9797);
nand U10338 (N_10338,N_9720,N_9692);
nand U10339 (N_10339,N_9784,N_9809);
and U10340 (N_10340,N_9725,N_9938);
nand U10341 (N_10341,N_9542,N_9767);
and U10342 (N_10342,N_9804,N_9999);
nand U10343 (N_10343,N_9832,N_9600);
or U10344 (N_10344,N_9566,N_9774);
xnor U10345 (N_10345,N_9694,N_9667);
or U10346 (N_10346,N_9986,N_9530);
nor U10347 (N_10347,N_9812,N_9579);
nor U10348 (N_10348,N_9862,N_9605);
nor U10349 (N_10349,N_9938,N_9548);
xor U10350 (N_10350,N_9992,N_9616);
nand U10351 (N_10351,N_9894,N_9890);
nand U10352 (N_10352,N_9767,N_9557);
or U10353 (N_10353,N_9648,N_9543);
nand U10354 (N_10354,N_9810,N_9877);
or U10355 (N_10355,N_9901,N_9678);
nand U10356 (N_10356,N_9743,N_9806);
nand U10357 (N_10357,N_9820,N_9976);
xnor U10358 (N_10358,N_9898,N_9985);
or U10359 (N_10359,N_9915,N_9985);
nor U10360 (N_10360,N_9986,N_9885);
and U10361 (N_10361,N_9591,N_9611);
and U10362 (N_10362,N_9712,N_9726);
nor U10363 (N_10363,N_9636,N_9814);
or U10364 (N_10364,N_9851,N_9572);
and U10365 (N_10365,N_9869,N_9552);
nor U10366 (N_10366,N_9595,N_9699);
and U10367 (N_10367,N_9521,N_9834);
nand U10368 (N_10368,N_9528,N_9707);
xor U10369 (N_10369,N_9926,N_9949);
or U10370 (N_10370,N_9803,N_9750);
and U10371 (N_10371,N_9883,N_9819);
nand U10372 (N_10372,N_9839,N_9692);
nor U10373 (N_10373,N_9836,N_9890);
xor U10374 (N_10374,N_9860,N_9920);
nor U10375 (N_10375,N_9720,N_9901);
and U10376 (N_10376,N_9803,N_9741);
xnor U10377 (N_10377,N_9874,N_9709);
nor U10378 (N_10378,N_9866,N_9586);
nand U10379 (N_10379,N_9905,N_9884);
nand U10380 (N_10380,N_9588,N_9732);
and U10381 (N_10381,N_9755,N_9561);
xnor U10382 (N_10382,N_9822,N_9797);
nor U10383 (N_10383,N_9846,N_9736);
nand U10384 (N_10384,N_9712,N_9958);
xor U10385 (N_10385,N_9618,N_9748);
and U10386 (N_10386,N_9659,N_9757);
nand U10387 (N_10387,N_9661,N_9942);
xnor U10388 (N_10388,N_9628,N_9953);
nand U10389 (N_10389,N_9932,N_9923);
and U10390 (N_10390,N_9787,N_9544);
nand U10391 (N_10391,N_9861,N_9766);
nand U10392 (N_10392,N_9659,N_9536);
nand U10393 (N_10393,N_9512,N_9938);
nand U10394 (N_10394,N_9997,N_9501);
or U10395 (N_10395,N_9712,N_9906);
xor U10396 (N_10396,N_9857,N_9741);
and U10397 (N_10397,N_9547,N_9581);
nor U10398 (N_10398,N_9678,N_9951);
and U10399 (N_10399,N_9824,N_9886);
xnor U10400 (N_10400,N_9937,N_9571);
and U10401 (N_10401,N_9737,N_9815);
nor U10402 (N_10402,N_9872,N_9735);
or U10403 (N_10403,N_9698,N_9604);
xnor U10404 (N_10404,N_9636,N_9608);
and U10405 (N_10405,N_9815,N_9671);
or U10406 (N_10406,N_9803,N_9936);
nand U10407 (N_10407,N_9620,N_9670);
or U10408 (N_10408,N_9584,N_9781);
and U10409 (N_10409,N_9636,N_9816);
or U10410 (N_10410,N_9972,N_9897);
nand U10411 (N_10411,N_9742,N_9515);
xnor U10412 (N_10412,N_9824,N_9825);
xnor U10413 (N_10413,N_9592,N_9736);
nand U10414 (N_10414,N_9686,N_9565);
nand U10415 (N_10415,N_9882,N_9809);
and U10416 (N_10416,N_9570,N_9591);
xor U10417 (N_10417,N_9753,N_9608);
and U10418 (N_10418,N_9743,N_9717);
and U10419 (N_10419,N_9600,N_9559);
or U10420 (N_10420,N_9725,N_9866);
nor U10421 (N_10421,N_9761,N_9541);
xor U10422 (N_10422,N_9957,N_9763);
nand U10423 (N_10423,N_9637,N_9768);
nand U10424 (N_10424,N_9670,N_9892);
nor U10425 (N_10425,N_9950,N_9520);
xor U10426 (N_10426,N_9850,N_9745);
nor U10427 (N_10427,N_9684,N_9742);
nor U10428 (N_10428,N_9718,N_9671);
or U10429 (N_10429,N_9708,N_9623);
nand U10430 (N_10430,N_9556,N_9722);
xor U10431 (N_10431,N_9902,N_9944);
nand U10432 (N_10432,N_9977,N_9627);
nor U10433 (N_10433,N_9927,N_9744);
and U10434 (N_10434,N_9545,N_9966);
nand U10435 (N_10435,N_9826,N_9542);
nand U10436 (N_10436,N_9645,N_9944);
xnor U10437 (N_10437,N_9783,N_9612);
or U10438 (N_10438,N_9603,N_9544);
and U10439 (N_10439,N_9937,N_9630);
nor U10440 (N_10440,N_9806,N_9653);
nand U10441 (N_10441,N_9990,N_9558);
or U10442 (N_10442,N_9541,N_9645);
or U10443 (N_10443,N_9731,N_9750);
or U10444 (N_10444,N_9716,N_9689);
or U10445 (N_10445,N_9672,N_9512);
nor U10446 (N_10446,N_9859,N_9551);
xnor U10447 (N_10447,N_9600,N_9858);
and U10448 (N_10448,N_9809,N_9859);
nand U10449 (N_10449,N_9926,N_9671);
and U10450 (N_10450,N_9561,N_9894);
nor U10451 (N_10451,N_9926,N_9773);
and U10452 (N_10452,N_9983,N_9794);
or U10453 (N_10453,N_9913,N_9652);
and U10454 (N_10454,N_9909,N_9534);
xnor U10455 (N_10455,N_9953,N_9863);
and U10456 (N_10456,N_9541,N_9809);
and U10457 (N_10457,N_9510,N_9628);
and U10458 (N_10458,N_9974,N_9914);
nor U10459 (N_10459,N_9576,N_9595);
nand U10460 (N_10460,N_9786,N_9888);
nor U10461 (N_10461,N_9626,N_9976);
nor U10462 (N_10462,N_9974,N_9899);
or U10463 (N_10463,N_9962,N_9895);
or U10464 (N_10464,N_9766,N_9638);
nand U10465 (N_10465,N_9778,N_9802);
nor U10466 (N_10466,N_9793,N_9524);
nand U10467 (N_10467,N_9537,N_9744);
nand U10468 (N_10468,N_9639,N_9960);
nand U10469 (N_10469,N_9991,N_9955);
or U10470 (N_10470,N_9985,N_9771);
nor U10471 (N_10471,N_9696,N_9580);
or U10472 (N_10472,N_9815,N_9629);
xnor U10473 (N_10473,N_9821,N_9792);
xnor U10474 (N_10474,N_9512,N_9636);
nor U10475 (N_10475,N_9628,N_9840);
and U10476 (N_10476,N_9633,N_9954);
or U10477 (N_10477,N_9951,N_9860);
nor U10478 (N_10478,N_9736,N_9676);
nand U10479 (N_10479,N_9534,N_9697);
nor U10480 (N_10480,N_9688,N_9835);
and U10481 (N_10481,N_9860,N_9595);
or U10482 (N_10482,N_9604,N_9563);
nand U10483 (N_10483,N_9776,N_9545);
nor U10484 (N_10484,N_9714,N_9779);
and U10485 (N_10485,N_9824,N_9941);
nand U10486 (N_10486,N_9873,N_9513);
and U10487 (N_10487,N_9598,N_9608);
xor U10488 (N_10488,N_9641,N_9549);
and U10489 (N_10489,N_9601,N_9571);
nand U10490 (N_10490,N_9626,N_9943);
nor U10491 (N_10491,N_9780,N_9903);
or U10492 (N_10492,N_9532,N_9735);
nor U10493 (N_10493,N_9559,N_9516);
and U10494 (N_10494,N_9614,N_9707);
and U10495 (N_10495,N_9701,N_9741);
or U10496 (N_10496,N_9902,N_9865);
or U10497 (N_10497,N_9722,N_9986);
nor U10498 (N_10498,N_9619,N_9994);
and U10499 (N_10499,N_9821,N_9553);
nor U10500 (N_10500,N_10042,N_10406);
and U10501 (N_10501,N_10118,N_10228);
or U10502 (N_10502,N_10262,N_10235);
or U10503 (N_10503,N_10227,N_10185);
nor U10504 (N_10504,N_10096,N_10080);
xnor U10505 (N_10505,N_10303,N_10046);
xnor U10506 (N_10506,N_10022,N_10157);
xor U10507 (N_10507,N_10246,N_10033);
nand U10508 (N_10508,N_10137,N_10336);
nand U10509 (N_10509,N_10317,N_10029);
or U10510 (N_10510,N_10256,N_10363);
nor U10511 (N_10511,N_10209,N_10208);
and U10512 (N_10512,N_10155,N_10180);
or U10513 (N_10513,N_10011,N_10001);
and U10514 (N_10514,N_10100,N_10438);
nand U10515 (N_10515,N_10364,N_10481);
xor U10516 (N_10516,N_10172,N_10062);
or U10517 (N_10517,N_10082,N_10486);
xnor U10518 (N_10518,N_10237,N_10400);
nor U10519 (N_10519,N_10485,N_10123);
nand U10520 (N_10520,N_10439,N_10404);
nor U10521 (N_10521,N_10091,N_10177);
nor U10522 (N_10522,N_10450,N_10179);
or U10523 (N_10523,N_10099,N_10036);
nand U10524 (N_10524,N_10419,N_10347);
and U10525 (N_10525,N_10075,N_10412);
nor U10526 (N_10526,N_10018,N_10337);
or U10527 (N_10527,N_10340,N_10395);
xnor U10528 (N_10528,N_10349,N_10092);
nor U10529 (N_10529,N_10003,N_10013);
or U10530 (N_10530,N_10221,N_10020);
and U10531 (N_10531,N_10121,N_10356);
nand U10532 (N_10532,N_10264,N_10304);
nor U10533 (N_10533,N_10078,N_10050);
nand U10534 (N_10534,N_10371,N_10352);
or U10535 (N_10535,N_10226,N_10272);
and U10536 (N_10536,N_10282,N_10066);
nor U10537 (N_10537,N_10051,N_10278);
xor U10538 (N_10538,N_10341,N_10276);
or U10539 (N_10539,N_10016,N_10335);
nor U10540 (N_10540,N_10087,N_10027);
and U10541 (N_10541,N_10086,N_10232);
xnor U10542 (N_10542,N_10354,N_10108);
nor U10543 (N_10543,N_10383,N_10071);
nor U10544 (N_10544,N_10409,N_10328);
or U10545 (N_10545,N_10152,N_10048);
xnor U10546 (N_10546,N_10343,N_10401);
nand U10547 (N_10547,N_10240,N_10259);
xor U10548 (N_10548,N_10195,N_10134);
and U10549 (N_10549,N_10479,N_10132);
nor U10550 (N_10550,N_10370,N_10368);
nand U10551 (N_10551,N_10088,N_10425);
or U10552 (N_10552,N_10037,N_10420);
xnor U10553 (N_10553,N_10427,N_10355);
xor U10554 (N_10554,N_10012,N_10116);
nor U10555 (N_10555,N_10248,N_10320);
and U10556 (N_10556,N_10098,N_10417);
and U10557 (N_10557,N_10442,N_10010);
nor U10558 (N_10558,N_10330,N_10498);
nor U10559 (N_10559,N_10149,N_10476);
or U10560 (N_10560,N_10094,N_10223);
nand U10561 (N_10561,N_10423,N_10459);
xnor U10562 (N_10562,N_10113,N_10421);
and U10563 (N_10563,N_10426,N_10418);
or U10564 (N_10564,N_10194,N_10253);
nand U10565 (N_10565,N_10252,N_10153);
and U10566 (N_10566,N_10057,N_10230);
and U10567 (N_10567,N_10119,N_10374);
nor U10568 (N_10568,N_10321,N_10162);
xnor U10569 (N_10569,N_10133,N_10008);
or U10570 (N_10570,N_10458,N_10261);
nand U10571 (N_10571,N_10385,N_10025);
nor U10572 (N_10572,N_10480,N_10126);
or U10573 (N_10573,N_10039,N_10318);
xnor U10574 (N_10574,N_10166,N_10073);
or U10575 (N_10575,N_10410,N_10451);
nor U10576 (N_10576,N_10396,N_10483);
or U10577 (N_10577,N_10461,N_10372);
and U10578 (N_10578,N_10081,N_10064);
xnor U10579 (N_10579,N_10314,N_10366);
nand U10580 (N_10580,N_10296,N_10411);
nor U10581 (N_10581,N_10300,N_10173);
or U10582 (N_10582,N_10467,N_10229);
nand U10583 (N_10583,N_10138,N_10097);
and U10584 (N_10584,N_10084,N_10324);
or U10585 (N_10585,N_10146,N_10357);
or U10586 (N_10586,N_10487,N_10198);
nand U10587 (N_10587,N_10147,N_10076);
or U10588 (N_10588,N_10367,N_10224);
or U10589 (N_10589,N_10074,N_10361);
or U10590 (N_10590,N_10435,N_10142);
xnor U10591 (N_10591,N_10388,N_10284);
nor U10592 (N_10592,N_10181,N_10322);
and U10593 (N_10593,N_10305,N_10291);
and U10594 (N_10594,N_10275,N_10164);
xor U10595 (N_10595,N_10218,N_10333);
nor U10596 (N_10596,N_10308,N_10058);
and U10597 (N_10597,N_10006,N_10053);
nor U10598 (N_10598,N_10306,N_10413);
and U10599 (N_10599,N_10429,N_10403);
and U10600 (N_10600,N_10007,N_10151);
or U10601 (N_10601,N_10307,N_10462);
and U10602 (N_10602,N_10184,N_10054);
or U10603 (N_10603,N_10129,N_10312);
nand U10604 (N_10604,N_10326,N_10494);
nor U10605 (N_10605,N_10024,N_10477);
or U10606 (N_10606,N_10251,N_10216);
or U10607 (N_10607,N_10424,N_10289);
or U10608 (N_10608,N_10070,N_10431);
xnor U10609 (N_10609,N_10441,N_10068);
or U10610 (N_10610,N_10298,N_10271);
nor U10611 (N_10611,N_10452,N_10052);
nand U10612 (N_10612,N_10169,N_10122);
nor U10613 (N_10613,N_10249,N_10473);
or U10614 (N_10614,N_10145,N_10117);
nand U10615 (N_10615,N_10263,N_10041);
or U10616 (N_10616,N_10375,N_10200);
nand U10617 (N_10617,N_10201,N_10474);
xnor U10618 (N_10618,N_10447,N_10014);
xor U10619 (N_10619,N_10197,N_10238);
xor U10620 (N_10620,N_10277,N_10475);
or U10621 (N_10621,N_10236,N_10205);
xnor U10622 (N_10622,N_10241,N_10378);
nand U10623 (N_10623,N_10286,N_10090);
nand U10624 (N_10624,N_10199,N_10215);
and U10625 (N_10625,N_10156,N_10083);
or U10626 (N_10626,N_10433,N_10471);
nor U10627 (N_10627,N_10416,N_10055);
and U10628 (N_10628,N_10407,N_10136);
or U10629 (N_10629,N_10004,N_10430);
nor U10630 (N_10630,N_10239,N_10247);
xnor U10631 (N_10631,N_10186,N_10065);
xor U10632 (N_10632,N_10482,N_10288);
xor U10633 (N_10633,N_10369,N_10168);
or U10634 (N_10634,N_10207,N_10379);
xor U10635 (N_10635,N_10044,N_10023);
nand U10636 (N_10636,N_10171,N_10351);
or U10637 (N_10637,N_10219,N_10102);
nand U10638 (N_10638,N_10456,N_10444);
xnor U10639 (N_10639,N_10030,N_10455);
nand U10640 (N_10640,N_10414,N_10028);
nand U10641 (N_10641,N_10124,N_10213);
xnor U10642 (N_10642,N_10301,N_10472);
and U10643 (N_10643,N_10127,N_10188);
or U10644 (N_10644,N_10394,N_10329);
nand U10645 (N_10645,N_10267,N_10047);
or U10646 (N_10646,N_10376,N_10273);
nand U10647 (N_10647,N_10035,N_10254);
nand U10648 (N_10648,N_10101,N_10270);
nor U10649 (N_10649,N_10085,N_10290);
nand U10650 (N_10650,N_10021,N_10178);
nor U10651 (N_10651,N_10191,N_10210);
xor U10652 (N_10652,N_10144,N_10107);
xor U10653 (N_10653,N_10049,N_10359);
nor U10654 (N_10654,N_10389,N_10139);
nor U10655 (N_10655,N_10358,N_10390);
nor U10656 (N_10656,N_10295,N_10225);
and U10657 (N_10657,N_10422,N_10231);
and U10658 (N_10658,N_10280,N_10141);
and U10659 (N_10659,N_10294,N_10060);
and U10660 (N_10660,N_10387,N_10381);
nand U10661 (N_10661,N_10000,N_10077);
nor U10662 (N_10662,N_10265,N_10495);
xor U10663 (N_10663,N_10464,N_10182);
nand U10664 (N_10664,N_10135,N_10061);
or U10665 (N_10665,N_10040,N_10334);
and U10666 (N_10666,N_10203,N_10316);
and U10667 (N_10667,N_10384,N_10457);
or U10668 (N_10668,N_10323,N_10345);
and U10669 (N_10669,N_10446,N_10373);
and U10670 (N_10670,N_10143,N_10104);
xnor U10671 (N_10671,N_10017,N_10103);
or U10672 (N_10672,N_10031,N_10437);
xor U10673 (N_10673,N_10258,N_10204);
nand U10674 (N_10674,N_10015,N_10443);
nand U10675 (N_10675,N_10362,N_10163);
nand U10676 (N_10676,N_10377,N_10148);
xor U10677 (N_10677,N_10034,N_10242);
nand U10678 (N_10678,N_10285,N_10342);
or U10679 (N_10679,N_10468,N_10257);
nand U10680 (N_10680,N_10283,N_10313);
and U10681 (N_10681,N_10069,N_10130);
nor U10682 (N_10682,N_10339,N_10274);
or U10683 (N_10683,N_10331,N_10344);
nand U10684 (N_10684,N_10287,N_10310);
and U10685 (N_10685,N_10009,N_10160);
nor U10686 (N_10686,N_10038,N_10279);
xor U10687 (N_10687,N_10222,N_10250);
and U10688 (N_10688,N_10319,N_10445);
or U10689 (N_10689,N_10002,N_10165);
nor U10690 (N_10690,N_10365,N_10187);
or U10691 (N_10691,N_10478,N_10175);
xor U10692 (N_10692,N_10183,N_10491);
nand U10693 (N_10693,N_10089,N_10393);
nor U10694 (N_10694,N_10346,N_10269);
or U10695 (N_10695,N_10161,N_10245);
xor U10696 (N_10696,N_10402,N_10492);
and U10697 (N_10697,N_10399,N_10244);
nor U10698 (N_10698,N_10105,N_10415);
nand U10699 (N_10699,N_10348,N_10111);
nor U10700 (N_10700,N_10154,N_10120);
or U10701 (N_10701,N_10350,N_10260);
nor U10702 (N_10702,N_10234,N_10428);
xnor U10703 (N_10703,N_10436,N_10174);
xor U10704 (N_10704,N_10360,N_10128);
and U10705 (N_10705,N_10332,N_10448);
xnor U10706 (N_10706,N_10176,N_10211);
nand U10707 (N_10707,N_10386,N_10170);
nor U10708 (N_10708,N_10408,N_10380);
or U10709 (N_10709,N_10093,N_10026);
or U10710 (N_10710,N_10391,N_10214);
xor U10711 (N_10711,N_10397,N_10140);
nand U10712 (N_10712,N_10095,N_10114);
and U10713 (N_10713,N_10338,N_10382);
nor U10714 (N_10714,N_10353,N_10243);
or U10715 (N_10715,N_10398,N_10465);
or U10716 (N_10716,N_10192,N_10206);
or U10717 (N_10717,N_10109,N_10189);
nor U10718 (N_10718,N_10150,N_10067);
or U10719 (N_10719,N_10266,N_10217);
nor U10720 (N_10720,N_10292,N_10496);
nand U10721 (N_10721,N_10045,N_10255);
nand U10722 (N_10722,N_10466,N_10112);
nor U10723 (N_10723,N_10005,N_10315);
xnor U10724 (N_10724,N_10159,N_10470);
xor U10725 (N_10725,N_10131,N_10490);
nor U10726 (N_10726,N_10453,N_10299);
xor U10727 (N_10727,N_10059,N_10405);
or U10728 (N_10728,N_10434,N_10110);
or U10729 (N_10729,N_10079,N_10449);
and U10730 (N_10730,N_10106,N_10489);
nor U10731 (N_10731,N_10484,N_10019);
xor U10732 (N_10732,N_10220,N_10460);
and U10733 (N_10733,N_10325,N_10497);
and U10734 (N_10734,N_10115,N_10469);
nor U10735 (N_10735,N_10463,N_10125);
and U10736 (N_10736,N_10440,N_10499);
xnor U10737 (N_10737,N_10309,N_10268);
or U10738 (N_10738,N_10190,N_10493);
and U10739 (N_10739,N_10281,N_10072);
and U10740 (N_10740,N_10297,N_10032);
or U10741 (N_10741,N_10454,N_10043);
and U10742 (N_10742,N_10302,N_10158);
nor U10743 (N_10743,N_10167,N_10196);
or U10744 (N_10744,N_10311,N_10392);
xor U10745 (N_10745,N_10202,N_10327);
or U10746 (N_10746,N_10193,N_10233);
nand U10747 (N_10747,N_10056,N_10432);
xor U10748 (N_10748,N_10488,N_10212);
nor U10749 (N_10749,N_10293,N_10063);
xnor U10750 (N_10750,N_10252,N_10464);
and U10751 (N_10751,N_10355,N_10409);
nor U10752 (N_10752,N_10369,N_10425);
or U10753 (N_10753,N_10427,N_10482);
nand U10754 (N_10754,N_10050,N_10206);
nor U10755 (N_10755,N_10499,N_10068);
xor U10756 (N_10756,N_10341,N_10390);
nor U10757 (N_10757,N_10275,N_10264);
xnor U10758 (N_10758,N_10464,N_10128);
xor U10759 (N_10759,N_10473,N_10375);
or U10760 (N_10760,N_10130,N_10201);
or U10761 (N_10761,N_10340,N_10367);
or U10762 (N_10762,N_10156,N_10111);
xnor U10763 (N_10763,N_10068,N_10335);
xnor U10764 (N_10764,N_10189,N_10485);
nor U10765 (N_10765,N_10281,N_10306);
and U10766 (N_10766,N_10030,N_10357);
nor U10767 (N_10767,N_10114,N_10207);
xor U10768 (N_10768,N_10195,N_10420);
nor U10769 (N_10769,N_10365,N_10078);
and U10770 (N_10770,N_10094,N_10115);
and U10771 (N_10771,N_10299,N_10280);
nand U10772 (N_10772,N_10118,N_10200);
xor U10773 (N_10773,N_10275,N_10095);
and U10774 (N_10774,N_10355,N_10207);
nor U10775 (N_10775,N_10177,N_10293);
nor U10776 (N_10776,N_10061,N_10101);
and U10777 (N_10777,N_10432,N_10151);
nor U10778 (N_10778,N_10188,N_10176);
xor U10779 (N_10779,N_10456,N_10166);
nor U10780 (N_10780,N_10055,N_10063);
xor U10781 (N_10781,N_10146,N_10422);
xor U10782 (N_10782,N_10497,N_10486);
nor U10783 (N_10783,N_10308,N_10344);
and U10784 (N_10784,N_10046,N_10055);
nor U10785 (N_10785,N_10430,N_10202);
nor U10786 (N_10786,N_10007,N_10427);
and U10787 (N_10787,N_10341,N_10435);
and U10788 (N_10788,N_10121,N_10290);
nand U10789 (N_10789,N_10227,N_10261);
nand U10790 (N_10790,N_10404,N_10387);
and U10791 (N_10791,N_10116,N_10158);
and U10792 (N_10792,N_10066,N_10169);
xor U10793 (N_10793,N_10255,N_10401);
or U10794 (N_10794,N_10467,N_10302);
xor U10795 (N_10795,N_10482,N_10107);
xnor U10796 (N_10796,N_10362,N_10049);
nor U10797 (N_10797,N_10114,N_10269);
nand U10798 (N_10798,N_10315,N_10139);
and U10799 (N_10799,N_10246,N_10138);
nand U10800 (N_10800,N_10270,N_10435);
or U10801 (N_10801,N_10212,N_10433);
nand U10802 (N_10802,N_10207,N_10039);
or U10803 (N_10803,N_10315,N_10105);
nor U10804 (N_10804,N_10465,N_10307);
nor U10805 (N_10805,N_10325,N_10358);
nor U10806 (N_10806,N_10223,N_10077);
xnor U10807 (N_10807,N_10001,N_10369);
nand U10808 (N_10808,N_10007,N_10402);
nand U10809 (N_10809,N_10208,N_10197);
or U10810 (N_10810,N_10337,N_10117);
and U10811 (N_10811,N_10111,N_10272);
and U10812 (N_10812,N_10488,N_10180);
xnor U10813 (N_10813,N_10080,N_10219);
xor U10814 (N_10814,N_10099,N_10148);
or U10815 (N_10815,N_10203,N_10378);
or U10816 (N_10816,N_10497,N_10093);
and U10817 (N_10817,N_10404,N_10422);
nor U10818 (N_10818,N_10358,N_10459);
or U10819 (N_10819,N_10302,N_10414);
and U10820 (N_10820,N_10442,N_10319);
nand U10821 (N_10821,N_10201,N_10437);
xnor U10822 (N_10822,N_10011,N_10360);
or U10823 (N_10823,N_10318,N_10077);
nor U10824 (N_10824,N_10252,N_10362);
or U10825 (N_10825,N_10115,N_10018);
xor U10826 (N_10826,N_10234,N_10432);
and U10827 (N_10827,N_10045,N_10418);
and U10828 (N_10828,N_10351,N_10127);
nand U10829 (N_10829,N_10009,N_10006);
or U10830 (N_10830,N_10483,N_10229);
or U10831 (N_10831,N_10009,N_10127);
and U10832 (N_10832,N_10317,N_10147);
or U10833 (N_10833,N_10065,N_10001);
or U10834 (N_10834,N_10312,N_10017);
and U10835 (N_10835,N_10258,N_10102);
and U10836 (N_10836,N_10293,N_10366);
nor U10837 (N_10837,N_10213,N_10269);
nand U10838 (N_10838,N_10072,N_10135);
and U10839 (N_10839,N_10199,N_10155);
nand U10840 (N_10840,N_10005,N_10237);
or U10841 (N_10841,N_10051,N_10276);
xnor U10842 (N_10842,N_10377,N_10241);
nor U10843 (N_10843,N_10156,N_10040);
nand U10844 (N_10844,N_10139,N_10206);
nand U10845 (N_10845,N_10280,N_10292);
nand U10846 (N_10846,N_10015,N_10021);
or U10847 (N_10847,N_10232,N_10135);
and U10848 (N_10848,N_10382,N_10209);
xor U10849 (N_10849,N_10415,N_10059);
nor U10850 (N_10850,N_10082,N_10006);
and U10851 (N_10851,N_10055,N_10317);
xor U10852 (N_10852,N_10224,N_10431);
and U10853 (N_10853,N_10031,N_10298);
nand U10854 (N_10854,N_10324,N_10358);
nand U10855 (N_10855,N_10108,N_10011);
xor U10856 (N_10856,N_10412,N_10113);
nor U10857 (N_10857,N_10121,N_10314);
xnor U10858 (N_10858,N_10134,N_10203);
xor U10859 (N_10859,N_10355,N_10038);
nor U10860 (N_10860,N_10150,N_10406);
xor U10861 (N_10861,N_10034,N_10426);
or U10862 (N_10862,N_10310,N_10059);
nor U10863 (N_10863,N_10276,N_10499);
and U10864 (N_10864,N_10184,N_10102);
xnor U10865 (N_10865,N_10402,N_10381);
and U10866 (N_10866,N_10080,N_10396);
nand U10867 (N_10867,N_10474,N_10340);
and U10868 (N_10868,N_10095,N_10391);
xor U10869 (N_10869,N_10402,N_10191);
nand U10870 (N_10870,N_10118,N_10099);
nor U10871 (N_10871,N_10162,N_10427);
or U10872 (N_10872,N_10427,N_10159);
nor U10873 (N_10873,N_10178,N_10418);
nor U10874 (N_10874,N_10400,N_10406);
or U10875 (N_10875,N_10231,N_10360);
or U10876 (N_10876,N_10308,N_10375);
or U10877 (N_10877,N_10346,N_10477);
or U10878 (N_10878,N_10053,N_10102);
or U10879 (N_10879,N_10285,N_10089);
xor U10880 (N_10880,N_10431,N_10177);
and U10881 (N_10881,N_10480,N_10287);
xor U10882 (N_10882,N_10283,N_10335);
nor U10883 (N_10883,N_10406,N_10431);
nand U10884 (N_10884,N_10493,N_10268);
or U10885 (N_10885,N_10140,N_10176);
xor U10886 (N_10886,N_10170,N_10145);
xnor U10887 (N_10887,N_10146,N_10457);
nor U10888 (N_10888,N_10112,N_10294);
xnor U10889 (N_10889,N_10130,N_10251);
or U10890 (N_10890,N_10120,N_10428);
nor U10891 (N_10891,N_10170,N_10025);
or U10892 (N_10892,N_10449,N_10454);
xor U10893 (N_10893,N_10160,N_10320);
or U10894 (N_10894,N_10315,N_10115);
nor U10895 (N_10895,N_10479,N_10120);
nand U10896 (N_10896,N_10146,N_10351);
nand U10897 (N_10897,N_10268,N_10015);
nand U10898 (N_10898,N_10022,N_10442);
nand U10899 (N_10899,N_10152,N_10299);
and U10900 (N_10900,N_10060,N_10469);
and U10901 (N_10901,N_10418,N_10458);
nand U10902 (N_10902,N_10349,N_10195);
nand U10903 (N_10903,N_10389,N_10496);
nand U10904 (N_10904,N_10254,N_10151);
and U10905 (N_10905,N_10025,N_10178);
nor U10906 (N_10906,N_10439,N_10379);
nor U10907 (N_10907,N_10124,N_10499);
nor U10908 (N_10908,N_10337,N_10320);
nand U10909 (N_10909,N_10182,N_10055);
or U10910 (N_10910,N_10146,N_10380);
nor U10911 (N_10911,N_10234,N_10032);
or U10912 (N_10912,N_10050,N_10294);
nor U10913 (N_10913,N_10290,N_10149);
nor U10914 (N_10914,N_10211,N_10494);
and U10915 (N_10915,N_10352,N_10115);
xor U10916 (N_10916,N_10062,N_10051);
or U10917 (N_10917,N_10053,N_10247);
xnor U10918 (N_10918,N_10176,N_10040);
nand U10919 (N_10919,N_10358,N_10170);
or U10920 (N_10920,N_10259,N_10478);
and U10921 (N_10921,N_10187,N_10253);
nand U10922 (N_10922,N_10028,N_10144);
or U10923 (N_10923,N_10156,N_10327);
and U10924 (N_10924,N_10469,N_10347);
nor U10925 (N_10925,N_10403,N_10441);
and U10926 (N_10926,N_10396,N_10448);
nor U10927 (N_10927,N_10284,N_10353);
and U10928 (N_10928,N_10395,N_10379);
or U10929 (N_10929,N_10176,N_10332);
nand U10930 (N_10930,N_10332,N_10368);
and U10931 (N_10931,N_10330,N_10445);
or U10932 (N_10932,N_10281,N_10058);
xnor U10933 (N_10933,N_10001,N_10096);
xnor U10934 (N_10934,N_10004,N_10333);
xnor U10935 (N_10935,N_10310,N_10241);
nor U10936 (N_10936,N_10025,N_10378);
nand U10937 (N_10937,N_10067,N_10439);
and U10938 (N_10938,N_10019,N_10420);
nor U10939 (N_10939,N_10482,N_10253);
and U10940 (N_10940,N_10186,N_10208);
xor U10941 (N_10941,N_10282,N_10170);
xnor U10942 (N_10942,N_10429,N_10336);
xor U10943 (N_10943,N_10269,N_10319);
xor U10944 (N_10944,N_10218,N_10179);
xnor U10945 (N_10945,N_10106,N_10493);
and U10946 (N_10946,N_10119,N_10476);
and U10947 (N_10947,N_10218,N_10276);
nand U10948 (N_10948,N_10010,N_10276);
and U10949 (N_10949,N_10498,N_10050);
and U10950 (N_10950,N_10077,N_10487);
nand U10951 (N_10951,N_10263,N_10092);
nor U10952 (N_10952,N_10135,N_10297);
nand U10953 (N_10953,N_10055,N_10246);
xnor U10954 (N_10954,N_10046,N_10313);
nor U10955 (N_10955,N_10183,N_10088);
or U10956 (N_10956,N_10393,N_10415);
xnor U10957 (N_10957,N_10159,N_10314);
and U10958 (N_10958,N_10396,N_10001);
and U10959 (N_10959,N_10204,N_10092);
xor U10960 (N_10960,N_10327,N_10453);
and U10961 (N_10961,N_10065,N_10166);
nand U10962 (N_10962,N_10219,N_10170);
or U10963 (N_10963,N_10234,N_10436);
xnor U10964 (N_10964,N_10410,N_10087);
or U10965 (N_10965,N_10276,N_10128);
and U10966 (N_10966,N_10425,N_10134);
or U10967 (N_10967,N_10441,N_10012);
nor U10968 (N_10968,N_10054,N_10186);
nor U10969 (N_10969,N_10491,N_10078);
nor U10970 (N_10970,N_10039,N_10259);
or U10971 (N_10971,N_10239,N_10084);
nor U10972 (N_10972,N_10406,N_10477);
nand U10973 (N_10973,N_10480,N_10035);
nand U10974 (N_10974,N_10367,N_10356);
or U10975 (N_10975,N_10372,N_10181);
xnor U10976 (N_10976,N_10404,N_10372);
and U10977 (N_10977,N_10045,N_10350);
and U10978 (N_10978,N_10033,N_10249);
or U10979 (N_10979,N_10206,N_10143);
and U10980 (N_10980,N_10199,N_10498);
and U10981 (N_10981,N_10276,N_10285);
or U10982 (N_10982,N_10271,N_10032);
xor U10983 (N_10983,N_10037,N_10032);
nand U10984 (N_10984,N_10212,N_10078);
or U10985 (N_10985,N_10225,N_10421);
or U10986 (N_10986,N_10395,N_10015);
nor U10987 (N_10987,N_10355,N_10024);
xor U10988 (N_10988,N_10400,N_10019);
or U10989 (N_10989,N_10195,N_10065);
and U10990 (N_10990,N_10134,N_10182);
nor U10991 (N_10991,N_10089,N_10169);
xor U10992 (N_10992,N_10039,N_10129);
or U10993 (N_10993,N_10454,N_10498);
nand U10994 (N_10994,N_10432,N_10476);
and U10995 (N_10995,N_10450,N_10394);
xor U10996 (N_10996,N_10181,N_10216);
and U10997 (N_10997,N_10292,N_10365);
or U10998 (N_10998,N_10050,N_10313);
nor U10999 (N_10999,N_10276,N_10177);
or U11000 (N_11000,N_10877,N_10568);
xnor U11001 (N_11001,N_10904,N_10572);
and U11002 (N_11002,N_10977,N_10872);
or U11003 (N_11003,N_10703,N_10503);
or U11004 (N_11004,N_10693,N_10878);
and U11005 (N_11005,N_10643,N_10774);
and U11006 (N_11006,N_10667,N_10853);
and U11007 (N_11007,N_10580,N_10788);
nor U11008 (N_11008,N_10954,N_10661);
and U11009 (N_11009,N_10502,N_10755);
and U11010 (N_11010,N_10586,N_10929);
or U11011 (N_11011,N_10922,N_10850);
and U11012 (N_11012,N_10711,N_10972);
nor U11013 (N_11013,N_10543,N_10974);
xnor U11014 (N_11014,N_10575,N_10544);
and U11015 (N_11015,N_10961,N_10671);
nand U11016 (N_11016,N_10776,N_10807);
xnor U11017 (N_11017,N_10861,N_10556);
xor U11018 (N_11018,N_10604,N_10690);
nor U11019 (N_11019,N_10800,N_10862);
or U11020 (N_11020,N_10958,N_10557);
nand U11021 (N_11021,N_10946,N_10910);
and U11022 (N_11022,N_10682,N_10723);
or U11023 (N_11023,N_10719,N_10883);
and U11024 (N_11024,N_10510,N_10907);
and U11025 (N_11025,N_10651,N_10798);
xor U11026 (N_11026,N_10647,N_10678);
xor U11027 (N_11027,N_10691,N_10621);
nand U11028 (N_11028,N_10845,N_10710);
and U11029 (N_11029,N_10911,N_10595);
nand U11030 (N_11030,N_10786,N_10822);
nor U11031 (N_11031,N_10813,N_10593);
nand U11032 (N_11032,N_10629,N_10736);
or U11033 (N_11033,N_10914,N_10857);
nor U11034 (N_11034,N_10842,N_10831);
or U11035 (N_11035,N_10576,N_10803);
and U11036 (N_11036,N_10535,N_10749);
or U11037 (N_11037,N_10863,N_10740);
or U11038 (N_11038,N_10625,N_10865);
nand U11039 (N_11039,N_10789,N_10584);
nand U11040 (N_11040,N_10591,N_10882);
nor U11041 (N_11041,N_10553,N_10517);
xor U11042 (N_11042,N_10832,N_10988);
xor U11043 (N_11043,N_10953,N_10607);
xor U11044 (N_11044,N_10712,N_10927);
nor U11045 (N_11045,N_10708,N_10631);
or U11046 (N_11046,N_10658,N_10968);
nor U11047 (N_11047,N_10934,N_10936);
and U11048 (N_11048,N_10947,N_10819);
and U11049 (N_11049,N_10602,N_10512);
nand U11050 (N_11050,N_10537,N_10999);
nand U11051 (N_11051,N_10672,N_10742);
nand U11052 (N_11052,N_10841,N_10756);
xor U11053 (N_11053,N_10814,N_10697);
or U11054 (N_11054,N_10777,N_10992);
nand U11055 (N_11055,N_10815,N_10871);
and U11056 (N_11056,N_10555,N_10799);
or U11057 (N_11057,N_10599,N_10967);
xor U11058 (N_11058,N_10897,N_10791);
nor U11059 (N_11059,N_10852,N_10830);
or U11060 (N_11060,N_10998,N_10955);
and U11061 (N_11061,N_10731,N_10884);
xnor U11062 (N_11062,N_10713,N_10728);
xor U11063 (N_11063,N_10895,N_10560);
nand U11064 (N_11064,N_10804,N_10894);
nand U11065 (N_11065,N_10592,N_10991);
or U11066 (N_11066,N_10551,N_10913);
nand U11067 (N_11067,N_10596,N_10696);
nand U11068 (N_11068,N_10754,N_10617);
nand U11069 (N_11069,N_10552,N_10650);
nand U11070 (N_11070,N_10851,N_10585);
nor U11071 (N_11071,N_10680,N_10635);
and U11072 (N_11072,N_10717,N_10790);
nand U11073 (N_11073,N_10674,N_10699);
xnor U11074 (N_11074,N_10539,N_10589);
xnor U11075 (N_11075,N_10834,N_10866);
nor U11076 (N_11076,N_10981,N_10745);
nor U11077 (N_11077,N_10610,N_10869);
and U11078 (N_11078,N_10627,N_10513);
nand U11079 (N_11079,N_10638,N_10917);
nand U11080 (N_11080,N_10566,N_10924);
and U11081 (N_11081,N_10630,N_10701);
nand U11082 (N_11082,N_10901,N_10893);
nor U11083 (N_11083,N_10536,N_10854);
or U11084 (N_11084,N_10752,N_10709);
nor U11085 (N_11085,N_10562,N_10781);
nand U11086 (N_11086,N_10944,N_10778);
or U11087 (N_11087,N_10903,N_10888);
and U11088 (N_11088,N_10826,N_10677);
and U11089 (N_11089,N_10545,N_10547);
nand U11090 (N_11090,N_10770,N_10590);
nand U11091 (N_11091,N_10806,N_10577);
xnor U11092 (N_11092,N_10567,N_10724);
xnor U11093 (N_11093,N_10849,N_10608);
xnor U11094 (N_11094,N_10726,N_10676);
nand U11095 (N_11095,N_10687,N_10941);
and U11096 (N_11096,N_10619,N_10960);
or U11097 (N_11097,N_10730,N_10835);
nand U11098 (N_11098,N_10615,N_10642);
and U11099 (N_11099,N_10645,N_10675);
nor U11100 (N_11100,N_10542,N_10594);
or U11101 (N_11101,N_10732,N_10876);
xor U11102 (N_11102,N_10973,N_10660);
and U11103 (N_11103,N_10980,N_10810);
nand U11104 (N_11104,N_10932,N_10987);
xnor U11105 (N_11105,N_10505,N_10964);
xnor U11106 (N_11106,N_10860,N_10959);
nand U11107 (N_11107,N_10758,N_10735);
and U11108 (N_11108,N_10796,N_10765);
xnor U11109 (N_11109,N_10507,N_10880);
nor U11110 (N_11110,N_10905,N_10684);
nand U11111 (N_11111,N_10673,N_10978);
or U11112 (N_11112,N_10773,N_10870);
nor U11113 (N_11113,N_10686,N_10771);
nand U11114 (N_11114,N_10744,N_10506);
nor U11115 (N_11115,N_10700,N_10784);
and U11116 (N_11116,N_10706,N_10679);
nor U11117 (N_11117,N_10548,N_10581);
nand U11118 (N_11118,N_10601,N_10989);
and U11119 (N_11119,N_10632,N_10899);
xor U11120 (N_11120,N_10836,N_10926);
xnor U11121 (N_11121,N_10587,N_10793);
and U11122 (N_11122,N_10855,N_10856);
and U11123 (N_11123,N_10875,N_10763);
or U11124 (N_11124,N_10702,N_10962);
or U11125 (N_11125,N_10616,N_10994);
nand U11126 (N_11126,N_10530,N_10569);
and U11127 (N_11127,N_10746,N_10683);
and U11128 (N_11128,N_10761,N_10727);
nor U11129 (N_11129,N_10531,N_10816);
or U11130 (N_11130,N_10943,N_10634);
and U11131 (N_11131,N_10896,N_10885);
nand U11132 (N_11132,N_10670,N_10747);
nor U11133 (N_11133,N_10707,N_10718);
xor U11134 (N_11134,N_10753,N_10809);
or U11135 (N_11135,N_10688,N_10808);
and U11136 (N_11136,N_10858,N_10821);
xnor U11137 (N_11137,N_10983,N_10504);
xnor U11138 (N_11138,N_10757,N_10890);
or U11139 (N_11139,N_10963,N_10583);
xnor U11140 (N_11140,N_10802,N_10633);
xnor U11141 (N_11141,N_10952,N_10668);
xnor U11142 (N_11142,N_10823,N_10501);
nand U11143 (N_11143,N_10532,N_10550);
and U11144 (N_11144,N_10611,N_10571);
nand U11145 (N_11145,N_10541,N_10665);
xor U11146 (N_11146,N_10887,N_10521);
nor U11147 (N_11147,N_10805,N_10868);
nor U11148 (N_11148,N_10751,N_10825);
or U11149 (N_11149,N_10563,N_10511);
xnor U11150 (N_11150,N_10840,N_10915);
nor U11151 (N_11151,N_10957,N_10985);
nor U11152 (N_11152,N_10829,N_10935);
xor U11153 (N_11153,N_10626,N_10846);
and U11154 (N_11154,N_10729,N_10818);
and U11155 (N_11155,N_10613,N_10623);
nor U11156 (N_11156,N_10663,N_10659);
or U11157 (N_11157,N_10522,N_10928);
nand U11158 (N_11158,N_10787,N_10656);
xor U11159 (N_11159,N_10867,N_10889);
nand U11160 (N_11160,N_10750,N_10618);
nand U11161 (N_11161,N_10741,N_10641);
or U11162 (N_11162,N_10892,N_10780);
xor U11163 (N_11163,N_10909,N_10533);
and U11164 (N_11164,N_10655,N_10767);
or U11165 (N_11165,N_10933,N_10538);
nand U11166 (N_11166,N_10820,N_10508);
xnor U11167 (N_11167,N_10579,N_10636);
nor U11168 (N_11168,N_10738,N_10785);
and U11169 (N_11169,N_10605,N_10879);
nor U11170 (N_11170,N_10603,N_10639);
nor U11171 (N_11171,N_10681,N_10812);
nor U11172 (N_11172,N_10597,N_10839);
nor U11173 (N_11173,N_10720,N_10649);
or U11174 (N_11174,N_10902,N_10722);
xor U11175 (N_11175,N_10827,N_10881);
and U11176 (N_11176,N_10725,N_10509);
or U11177 (N_11177,N_10956,N_10769);
or U11178 (N_11178,N_10705,N_10516);
and U11179 (N_11179,N_10921,N_10794);
xor U11180 (N_11180,N_10931,N_10966);
and U11181 (N_11181,N_10971,N_10937);
and U11182 (N_11182,N_10939,N_10715);
nand U11183 (N_11183,N_10652,N_10716);
xor U11184 (N_11184,N_10559,N_10524);
nand U11185 (N_11185,N_10768,N_10982);
or U11186 (N_11186,N_10734,N_10523);
nor U11187 (N_11187,N_10996,N_10546);
and U11188 (N_11188,N_10993,N_10515);
nor U11189 (N_11189,N_10886,N_10527);
and U11190 (N_11190,N_10653,N_10704);
xnor U11191 (N_11191,N_10795,N_10561);
or U11192 (N_11192,N_10644,N_10549);
xnor U11193 (N_11193,N_10669,N_10824);
nor U11194 (N_11194,N_10938,N_10970);
nor U11195 (N_11195,N_10588,N_10775);
xor U11196 (N_11196,N_10578,N_10646);
nor U11197 (N_11197,N_10570,N_10759);
nand U11198 (N_11198,N_10748,N_10828);
and U11199 (N_11199,N_10692,N_10843);
nor U11200 (N_11200,N_10792,N_10648);
xnor U11201 (N_11201,N_10975,N_10997);
nor U11202 (N_11202,N_10772,N_10518);
and U11203 (N_11203,N_10666,N_10891);
xnor U11204 (N_11204,N_10540,N_10609);
and U11205 (N_11205,N_10898,N_10624);
nand U11206 (N_11206,N_10766,N_10500);
nor U11207 (N_11207,N_10664,N_10783);
and U11208 (N_11208,N_10918,N_10698);
xor U11209 (N_11209,N_10612,N_10519);
or U11210 (N_11210,N_10940,N_10598);
xnor U11211 (N_11211,N_10733,N_10514);
or U11212 (N_11212,N_10995,N_10912);
and U11213 (N_11213,N_10779,N_10574);
nand U11214 (N_11214,N_10526,N_10714);
and U11215 (N_11215,N_10948,N_10573);
xnor U11216 (N_11216,N_10529,N_10762);
xor U11217 (N_11217,N_10990,N_10906);
xnor U11218 (N_11218,N_10534,N_10695);
and U11219 (N_11219,N_10737,N_10950);
and U11220 (N_11220,N_10622,N_10844);
nor U11221 (N_11221,N_10847,N_10965);
nand U11222 (N_11222,N_10916,N_10760);
and U11223 (N_11223,N_10657,N_10919);
or U11224 (N_11224,N_10859,N_10640);
and U11225 (N_11225,N_10743,N_10801);
and U11226 (N_11226,N_10662,N_10925);
and U11227 (N_11227,N_10864,N_10848);
nor U11228 (N_11228,N_10620,N_10951);
nor U11229 (N_11229,N_10837,N_10565);
nor U11230 (N_11230,N_10817,N_10979);
and U11231 (N_11231,N_10600,N_10942);
and U11232 (N_11232,N_10811,N_10654);
or U11233 (N_11233,N_10685,N_10628);
xnor U11234 (N_11234,N_10873,N_10614);
xor U11235 (N_11235,N_10908,N_10900);
nand U11236 (N_11236,N_10969,N_10554);
or U11237 (N_11237,N_10838,N_10945);
or U11238 (N_11238,N_10582,N_10833);
nand U11239 (N_11239,N_10874,N_10564);
nand U11240 (N_11240,N_10520,N_10984);
nand U11241 (N_11241,N_10976,N_10797);
nor U11242 (N_11242,N_10606,N_10764);
nand U11243 (N_11243,N_10694,N_10558);
xor U11244 (N_11244,N_10525,N_10920);
nand U11245 (N_11245,N_10739,N_10986);
nor U11246 (N_11246,N_10782,N_10923);
nor U11247 (N_11247,N_10689,N_10528);
or U11248 (N_11248,N_10949,N_10721);
xor U11249 (N_11249,N_10637,N_10930);
and U11250 (N_11250,N_10962,N_10841);
and U11251 (N_11251,N_10700,N_10890);
and U11252 (N_11252,N_10668,N_10957);
xnor U11253 (N_11253,N_10550,N_10988);
nand U11254 (N_11254,N_10894,N_10547);
and U11255 (N_11255,N_10724,N_10963);
xor U11256 (N_11256,N_10784,N_10643);
or U11257 (N_11257,N_10593,N_10773);
nor U11258 (N_11258,N_10780,N_10595);
and U11259 (N_11259,N_10800,N_10622);
nor U11260 (N_11260,N_10815,N_10555);
nor U11261 (N_11261,N_10629,N_10983);
xnor U11262 (N_11262,N_10595,N_10893);
or U11263 (N_11263,N_10778,N_10947);
nand U11264 (N_11264,N_10769,N_10702);
nor U11265 (N_11265,N_10823,N_10692);
nor U11266 (N_11266,N_10534,N_10954);
and U11267 (N_11267,N_10544,N_10647);
nor U11268 (N_11268,N_10773,N_10938);
and U11269 (N_11269,N_10593,N_10538);
xor U11270 (N_11270,N_10521,N_10945);
and U11271 (N_11271,N_10594,N_10739);
nor U11272 (N_11272,N_10932,N_10670);
xnor U11273 (N_11273,N_10725,N_10919);
nor U11274 (N_11274,N_10765,N_10740);
nor U11275 (N_11275,N_10550,N_10674);
xnor U11276 (N_11276,N_10599,N_10802);
xnor U11277 (N_11277,N_10783,N_10868);
nand U11278 (N_11278,N_10564,N_10504);
or U11279 (N_11279,N_10988,N_10957);
xnor U11280 (N_11280,N_10909,N_10785);
and U11281 (N_11281,N_10801,N_10915);
or U11282 (N_11282,N_10953,N_10546);
and U11283 (N_11283,N_10648,N_10751);
or U11284 (N_11284,N_10890,N_10535);
nor U11285 (N_11285,N_10690,N_10978);
nand U11286 (N_11286,N_10963,N_10524);
and U11287 (N_11287,N_10814,N_10851);
nor U11288 (N_11288,N_10613,N_10694);
xor U11289 (N_11289,N_10698,N_10919);
nand U11290 (N_11290,N_10595,N_10648);
or U11291 (N_11291,N_10788,N_10988);
xor U11292 (N_11292,N_10568,N_10939);
or U11293 (N_11293,N_10783,N_10977);
and U11294 (N_11294,N_10804,N_10842);
xnor U11295 (N_11295,N_10840,N_10808);
nor U11296 (N_11296,N_10664,N_10654);
nor U11297 (N_11297,N_10797,N_10871);
nor U11298 (N_11298,N_10686,N_10850);
xor U11299 (N_11299,N_10972,N_10801);
xor U11300 (N_11300,N_10667,N_10644);
nand U11301 (N_11301,N_10521,N_10830);
nor U11302 (N_11302,N_10713,N_10847);
or U11303 (N_11303,N_10511,N_10941);
nor U11304 (N_11304,N_10532,N_10655);
nor U11305 (N_11305,N_10998,N_10889);
nand U11306 (N_11306,N_10836,N_10862);
nor U11307 (N_11307,N_10851,N_10599);
and U11308 (N_11308,N_10549,N_10931);
nand U11309 (N_11309,N_10580,N_10576);
xor U11310 (N_11310,N_10785,N_10564);
nand U11311 (N_11311,N_10952,N_10954);
nor U11312 (N_11312,N_10517,N_10502);
nand U11313 (N_11313,N_10950,N_10580);
xnor U11314 (N_11314,N_10948,N_10923);
nand U11315 (N_11315,N_10563,N_10708);
xor U11316 (N_11316,N_10905,N_10548);
and U11317 (N_11317,N_10524,N_10772);
xor U11318 (N_11318,N_10537,N_10775);
or U11319 (N_11319,N_10516,N_10550);
nor U11320 (N_11320,N_10568,N_10791);
nor U11321 (N_11321,N_10719,N_10657);
or U11322 (N_11322,N_10649,N_10623);
nand U11323 (N_11323,N_10575,N_10966);
or U11324 (N_11324,N_10906,N_10576);
nor U11325 (N_11325,N_10733,N_10695);
nand U11326 (N_11326,N_10934,N_10622);
xnor U11327 (N_11327,N_10821,N_10744);
nand U11328 (N_11328,N_10905,N_10645);
nor U11329 (N_11329,N_10680,N_10790);
nand U11330 (N_11330,N_10503,N_10616);
nand U11331 (N_11331,N_10702,N_10688);
and U11332 (N_11332,N_10963,N_10837);
and U11333 (N_11333,N_10887,N_10745);
or U11334 (N_11334,N_10583,N_10614);
nor U11335 (N_11335,N_10917,N_10935);
and U11336 (N_11336,N_10956,N_10837);
xnor U11337 (N_11337,N_10828,N_10879);
nand U11338 (N_11338,N_10852,N_10621);
nand U11339 (N_11339,N_10645,N_10850);
nor U11340 (N_11340,N_10814,N_10844);
nor U11341 (N_11341,N_10946,N_10816);
and U11342 (N_11342,N_10913,N_10841);
nor U11343 (N_11343,N_10761,N_10868);
nor U11344 (N_11344,N_10686,N_10658);
nor U11345 (N_11345,N_10670,N_10551);
xor U11346 (N_11346,N_10685,N_10942);
or U11347 (N_11347,N_10606,N_10530);
xor U11348 (N_11348,N_10899,N_10690);
nand U11349 (N_11349,N_10945,N_10611);
and U11350 (N_11350,N_10548,N_10627);
or U11351 (N_11351,N_10773,N_10989);
and U11352 (N_11352,N_10565,N_10626);
xor U11353 (N_11353,N_10659,N_10979);
xor U11354 (N_11354,N_10975,N_10844);
or U11355 (N_11355,N_10597,N_10729);
nand U11356 (N_11356,N_10535,N_10949);
and U11357 (N_11357,N_10987,N_10676);
nand U11358 (N_11358,N_10680,N_10839);
nor U11359 (N_11359,N_10971,N_10605);
and U11360 (N_11360,N_10608,N_10600);
and U11361 (N_11361,N_10664,N_10978);
xnor U11362 (N_11362,N_10890,N_10951);
and U11363 (N_11363,N_10783,N_10696);
or U11364 (N_11364,N_10894,N_10506);
or U11365 (N_11365,N_10612,N_10604);
nor U11366 (N_11366,N_10970,N_10633);
or U11367 (N_11367,N_10503,N_10548);
nor U11368 (N_11368,N_10649,N_10725);
and U11369 (N_11369,N_10618,N_10706);
nand U11370 (N_11370,N_10997,N_10810);
xnor U11371 (N_11371,N_10944,N_10844);
nand U11372 (N_11372,N_10550,N_10812);
nor U11373 (N_11373,N_10578,N_10841);
and U11374 (N_11374,N_10671,N_10845);
nand U11375 (N_11375,N_10517,N_10608);
or U11376 (N_11376,N_10933,N_10573);
and U11377 (N_11377,N_10639,N_10923);
xor U11378 (N_11378,N_10990,N_10776);
xor U11379 (N_11379,N_10793,N_10934);
nor U11380 (N_11380,N_10958,N_10593);
and U11381 (N_11381,N_10791,N_10582);
nor U11382 (N_11382,N_10809,N_10730);
nor U11383 (N_11383,N_10959,N_10523);
xnor U11384 (N_11384,N_10548,N_10552);
or U11385 (N_11385,N_10627,N_10874);
xnor U11386 (N_11386,N_10923,N_10760);
and U11387 (N_11387,N_10986,N_10920);
or U11388 (N_11388,N_10812,N_10830);
nand U11389 (N_11389,N_10672,N_10782);
and U11390 (N_11390,N_10536,N_10610);
and U11391 (N_11391,N_10593,N_10569);
nand U11392 (N_11392,N_10923,N_10723);
nand U11393 (N_11393,N_10976,N_10596);
and U11394 (N_11394,N_10653,N_10545);
nor U11395 (N_11395,N_10506,N_10619);
nor U11396 (N_11396,N_10853,N_10517);
and U11397 (N_11397,N_10935,N_10796);
xor U11398 (N_11398,N_10985,N_10964);
xnor U11399 (N_11399,N_10613,N_10609);
nand U11400 (N_11400,N_10605,N_10751);
nand U11401 (N_11401,N_10516,N_10537);
and U11402 (N_11402,N_10930,N_10843);
nand U11403 (N_11403,N_10802,N_10969);
and U11404 (N_11404,N_10595,N_10637);
nor U11405 (N_11405,N_10618,N_10796);
nand U11406 (N_11406,N_10974,N_10604);
and U11407 (N_11407,N_10763,N_10682);
or U11408 (N_11408,N_10696,N_10738);
nor U11409 (N_11409,N_10968,N_10589);
nand U11410 (N_11410,N_10696,N_10817);
nand U11411 (N_11411,N_10873,N_10787);
xnor U11412 (N_11412,N_10761,N_10524);
or U11413 (N_11413,N_10542,N_10633);
xor U11414 (N_11414,N_10947,N_10934);
nand U11415 (N_11415,N_10836,N_10811);
nand U11416 (N_11416,N_10815,N_10514);
and U11417 (N_11417,N_10701,N_10835);
or U11418 (N_11418,N_10594,N_10703);
nand U11419 (N_11419,N_10675,N_10611);
nand U11420 (N_11420,N_10677,N_10580);
xnor U11421 (N_11421,N_10508,N_10990);
or U11422 (N_11422,N_10794,N_10552);
or U11423 (N_11423,N_10692,N_10879);
and U11424 (N_11424,N_10588,N_10702);
nor U11425 (N_11425,N_10897,N_10718);
nand U11426 (N_11426,N_10637,N_10915);
and U11427 (N_11427,N_10797,N_10582);
xnor U11428 (N_11428,N_10601,N_10842);
and U11429 (N_11429,N_10502,N_10757);
xor U11430 (N_11430,N_10845,N_10750);
nor U11431 (N_11431,N_10752,N_10657);
nor U11432 (N_11432,N_10608,N_10986);
nor U11433 (N_11433,N_10607,N_10716);
nand U11434 (N_11434,N_10996,N_10920);
nand U11435 (N_11435,N_10602,N_10898);
nor U11436 (N_11436,N_10624,N_10712);
or U11437 (N_11437,N_10951,N_10985);
nand U11438 (N_11438,N_10699,N_10721);
nand U11439 (N_11439,N_10527,N_10915);
xor U11440 (N_11440,N_10935,N_10556);
or U11441 (N_11441,N_10707,N_10642);
and U11442 (N_11442,N_10936,N_10877);
and U11443 (N_11443,N_10950,N_10798);
nor U11444 (N_11444,N_10868,N_10664);
xor U11445 (N_11445,N_10894,N_10670);
and U11446 (N_11446,N_10700,N_10661);
or U11447 (N_11447,N_10612,N_10864);
xnor U11448 (N_11448,N_10816,N_10981);
xor U11449 (N_11449,N_10970,N_10704);
nand U11450 (N_11450,N_10973,N_10590);
or U11451 (N_11451,N_10928,N_10992);
and U11452 (N_11452,N_10934,N_10984);
nor U11453 (N_11453,N_10715,N_10875);
and U11454 (N_11454,N_10534,N_10911);
and U11455 (N_11455,N_10986,N_10661);
xor U11456 (N_11456,N_10631,N_10882);
and U11457 (N_11457,N_10621,N_10717);
xnor U11458 (N_11458,N_10905,N_10903);
nand U11459 (N_11459,N_10755,N_10999);
nand U11460 (N_11460,N_10524,N_10598);
nand U11461 (N_11461,N_10864,N_10717);
xnor U11462 (N_11462,N_10792,N_10734);
and U11463 (N_11463,N_10660,N_10947);
nor U11464 (N_11464,N_10738,N_10778);
and U11465 (N_11465,N_10861,N_10619);
or U11466 (N_11466,N_10889,N_10788);
xor U11467 (N_11467,N_10509,N_10954);
nor U11468 (N_11468,N_10861,N_10677);
xnor U11469 (N_11469,N_10854,N_10695);
and U11470 (N_11470,N_10846,N_10575);
xor U11471 (N_11471,N_10619,N_10533);
xnor U11472 (N_11472,N_10965,N_10530);
nand U11473 (N_11473,N_10517,N_10787);
nand U11474 (N_11474,N_10705,N_10742);
nand U11475 (N_11475,N_10639,N_10906);
nand U11476 (N_11476,N_10591,N_10844);
nor U11477 (N_11477,N_10629,N_10687);
nor U11478 (N_11478,N_10859,N_10794);
and U11479 (N_11479,N_10835,N_10610);
and U11480 (N_11480,N_10834,N_10746);
xor U11481 (N_11481,N_10947,N_10961);
nor U11482 (N_11482,N_10648,N_10905);
nand U11483 (N_11483,N_10681,N_10804);
or U11484 (N_11484,N_10831,N_10850);
xor U11485 (N_11485,N_10815,N_10761);
xor U11486 (N_11486,N_10567,N_10542);
or U11487 (N_11487,N_10802,N_10872);
or U11488 (N_11488,N_10727,N_10754);
or U11489 (N_11489,N_10740,N_10972);
nor U11490 (N_11490,N_10849,N_10594);
nand U11491 (N_11491,N_10656,N_10923);
and U11492 (N_11492,N_10550,N_10871);
and U11493 (N_11493,N_10534,N_10853);
nand U11494 (N_11494,N_10725,N_10909);
xor U11495 (N_11495,N_10750,N_10651);
and U11496 (N_11496,N_10697,N_10597);
xnor U11497 (N_11497,N_10704,N_10951);
and U11498 (N_11498,N_10611,N_10707);
xor U11499 (N_11499,N_10590,N_10593);
nor U11500 (N_11500,N_11051,N_11364);
nand U11501 (N_11501,N_11137,N_11159);
nand U11502 (N_11502,N_11122,N_11308);
nand U11503 (N_11503,N_11081,N_11176);
or U11504 (N_11504,N_11464,N_11312);
nand U11505 (N_11505,N_11160,N_11438);
or U11506 (N_11506,N_11385,N_11384);
or U11507 (N_11507,N_11274,N_11409);
and U11508 (N_11508,N_11413,N_11365);
nor U11509 (N_11509,N_11469,N_11231);
xnor U11510 (N_11510,N_11104,N_11338);
and U11511 (N_11511,N_11287,N_11116);
nor U11512 (N_11512,N_11099,N_11052);
or U11513 (N_11513,N_11107,N_11360);
nand U11514 (N_11514,N_11218,N_11079);
xnor U11515 (N_11515,N_11016,N_11309);
nor U11516 (N_11516,N_11432,N_11246);
xnor U11517 (N_11517,N_11336,N_11013);
xnor U11518 (N_11518,N_11084,N_11205);
nand U11519 (N_11519,N_11319,N_11020);
and U11520 (N_11520,N_11070,N_11283);
or U11521 (N_11521,N_11425,N_11109);
nand U11522 (N_11522,N_11374,N_11294);
nand U11523 (N_11523,N_11194,N_11396);
xnor U11524 (N_11524,N_11221,N_11430);
and U11525 (N_11525,N_11474,N_11427);
nor U11526 (N_11526,N_11045,N_11375);
nor U11527 (N_11527,N_11290,N_11224);
xnor U11528 (N_11528,N_11034,N_11225);
nor U11529 (N_11529,N_11350,N_11382);
nor U11530 (N_11530,N_11050,N_11462);
nand U11531 (N_11531,N_11297,N_11219);
nor U11532 (N_11532,N_11289,N_11090);
xor U11533 (N_11533,N_11471,N_11491);
xor U11534 (N_11534,N_11422,N_11124);
xnor U11535 (N_11535,N_11402,N_11239);
nor U11536 (N_11536,N_11447,N_11486);
or U11537 (N_11537,N_11242,N_11273);
nand U11538 (N_11538,N_11435,N_11479);
or U11539 (N_11539,N_11354,N_11378);
or U11540 (N_11540,N_11390,N_11161);
nor U11541 (N_11541,N_11493,N_11015);
xnor U11542 (N_11542,N_11085,N_11183);
or U11543 (N_11543,N_11062,N_11391);
nor U11544 (N_11544,N_11482,N_11128);
or U11545 (N_11545,N_11293,N_11281);
xnor U11546 (N_11546,N_11089,N_11178);
or U11547 (N_11547,N_11200,N_11111);
nand U11548 (N_11548,N_11358,N_11035);
and U11549 (N_11549,N_11172,N_11499);
nor U11550 (N_11550,N_11496,N_11315);
xnor U11551 (N_11551,N_11278,N_11222);
and U11552 (N_11552,N_11484,N_11343);
xnor U11553 (N_11553,N_11068,N_11276);
nand U11554 (N_11554,N_11423,N_11450);
xnor U11555 (N_11555,N_11215,N_11249);
xnor U11556 (N_11556,N_11304,N_11127);
or U11557 (N_11557,N_11216,N_11414);
nand U11558 (N_11558,N_11237,N_11025);
nor U11559 (N_11559,N_11386,N_11371);
and U11560 (N_11560,N_11042,N_11400);
xnor U11561 (N_11561,N_11142,N_11320);
nor U11562 (N_11562,N_11195,N_11286);
or U11563 (N_11563,N_11057,N_11188);
or U11564 (N_11564,N_11133,N_11008);
and U11565 (N_11565,N_11258,N_11058);
xnor U11566 (N_11566,N_11348,N_11497);
nand U11567 (N_11567,N_11055,N_11149);
xor U11568 (N_11568,N_11038,N_11442);
nand U11569 (N_11569,N_11202,N_11119);
xor U11570 (N_11570,N_11210,N_11046);
and U11571 (N_11571,N_11363,N_11305);
xor U11572 (N_11572,N_11233,N_11303);
and U11573 (N_11573,N_11306,N_11096);
or U11574 (N_11574,N_11129,N_11033);
nand U11575 (N_11575,N_11039,N_11190);
and U11576 (N_11576,N_11477,N_11492);
or U11577 (N_11577,N_11389,N_11284);
or U11578 (N_11578,N_11475,N_11362);
nand U11579 (N_11579,N_11141,N_11466);
and U11580 (N_11580,N_11175,N_11316);
or U11581 (N_11581,N_11048,N_11162);
or U11582 (N_11582,N_11135,N_11376);
nor U11583 (N_11583,N_11226,N_11014);
and U11584 (N_11584,N_11490,N_11445);
xnor U11585 (N_11585,N_11214,N_11080);
nor U11586 (N_11586,N_11408,N_11227);
xnor U11587 (N_11587,N_11005,N_11076);
nor U11588 (N_11588,N_11317,N_11481);
xnor U11589 (N_11589,N_11032,N_11411);
and U11590 (N_11590,N_11023,N_11480);
nand U11591 (N_11591,N_11110,N_11465);
nand U11592 (N_11592,N_11105,N_11017);
xnor U11593 (N_11593,N_11407,N_11060);
nand U11594 (N_11594,N_11072,N_11456);
or U11595 (N_11595,N_11311,N_11054);
nand U11596 (N_11596,N_11207,N_11313);
xnor U11597 (N_11597,N_11457,N_11361);
or U11598 (N_11598,N_11332,N_11208);
nand U11599 (N_11599,N_11347,N_11426);
nand U11600 (N_11600,N_11260,N_11399);
nand U11601 (N_11601,N_11185,N_11428);
xnor U11602 (N_11602,N_11117,N_11342);
xor U11603 (N_11603,N_11270,N_11229);
nand U11604 (N_11604,N_11279,N_11130);
nor U11605 (N_11605,N_11146,N_11071);
nor U11606 (N_11606,N_11394,N_11377);
and U11607 (N_11607,N_11082,N_11108);
xnor U11608 (N_11608,N_11275,N_11417);
nor U11609 (N_11609,N_11243,N_11369);
and U11610 (N_11610,N_11395,N_11381);
and U11611 (N_11611,N_11180,N_11257);
and U11612 (N_11612,N_11168,N_11251);
nand U11613 (N_11613,N_11167,N_11198);
nor U11614 (N_11614,N_11467,N_11223);
nand U11615 (N_11615,N_11461,N_11255);
nor U11616 (N_11616,N_11291,N_11310);
nand U11617 (N_11617,N_11346,N_11123);
or U11618 (N_11618,N_11006,N_11157);
or U11619 (N_11619,N_11134,N_11148);
nor U11620 (N_11620,N_11418,N_11019);
nand U11621 (N_11621,N_11101,N_11166);
and U11622 (N_11622,N_11196,N_11182);
or U11623 (N_11623,N_11087,N_11069);
or U11624 (N_11624,N_11329,N_11476);
xor U11625 (N_11625,N_11106,N_11063);
and U11626 (N_11626,N_11184,N_11126);
and U11627 (N_11627,N_11001,N_11029);
nor U11628 (N_11628,N_11355,N_11259);
and U11629 (N_11629,N_11352,N_11212);
nor U11630 (N_11630,N_11236,N_11372);
and U11631 (N_11631,N_11366,N_11356);
nor U11632 (N_11632,N_11125,N_11324);
xnor U11633 (N_11633,N_11451,N_11150);
or U11634 (N_11634,N_11170,N_11353);
or U11635 (N_11635,N_11049,N_11272);
nand U11636 (N_11636,N_11383,N_11392);
and U11637 (N_11637,N_11269,N_11268);
xnor U11638 (N_11638,N_11488,N_11398);
xnor U11639 (N_11639,N_11410,N_11191);
and U11640 (N_11640,N_11163,N_11250);
nand U11641 (N_11641,N_11120,N_11244);
nand U11642 (N_11642,N_11021,N_11439);
and U11643 (N_11643,N_11373,N_11186);
nand U11644 (N_11644,N_11240,N_11264);
nor U11645 (N_11645,N_11300,N_11351);
xnor U11646 (N_11646,N_11066,N_11091);
nor U11647 (N_11647,N_11199,N_11112);
nand U11648 (N_11648,N_11098,N_11282);
xnor U11649 (N_11649,N_11139,N_11368);
nand U11650 (N_11650,N_11179,N_11280);
nand U11651 (N_11651,N_11132,N_11165);
or U11652 (N_11652,N_11012,N_11040);
or U11653 (N_11653,N_11024,N_11073);
and U11654 (N_11654,N_11036,N_11174);
or U11655 (N_11655,N_11173,N_11230);
nand U11656 (N_11656,N_11065,N_11086);
nand U11657 (N_11657,N_11341,N_11113);
xnor U11658 (N_11658,N_11404,N_11143);
or U11659 (N_11659,N_11463,N_11302);
or U11660 (N_11660,N_11131,N_11437);
nand U11661 (N_11661,N_11261,N_11328);
and U11662 (N_11662,N_11429,N_11235);
and U11663 (N_11663,N_11446,N_11228);
nand U11664 (N_11664,N_11443,N_11421);
nand U11665 (N_11665,N_11292,N_11318);
or U11666 (N_11666,N_11405,N_11441);
nand U11667 (N_11667,N_11415,N_11043);
nand U11668 (N_11668,N_11193,N_11431);
xnor U11669 (N_11669,N_11201,N_11151);
nand U11670 (N_11670,N_11053,N_11000);
nor U11671 (N_11671,N_11002,N_11004);
nand U11672 (N_11672,N_11047,N_11209);
or U11673 (N_11673,N_11296,N_11092);
or U11674 (N_11674,N_11144,N_11453);
xnor U11675 (N_11675,N_11097,N_11169);
or U11676 (N_11676,N_11262,N_11075);
and U11677 (N_11677,N_11380,N_11436);
and U11678 (N_11678,N_11056,N_11121);
nand U11679 (N_11679,N_11103,N_11397);
nor U11680 (N_11680,N_11030,N_11321);
nand U11681 (N_11681,N_11064,N_11189);
nor U11682 (N_11682,N_11478,N_11078);
xnor U11683 (N_11683,N_11011,N_11147);
or U11684 (N_11684,N_11095,N_11455);
nor U11685 (N_11685,N_11155,N_11158);
nor U11686 (N_11686,N_11138,N_11181);
and U11687 (N_11687,N_11118,N_11494);
or U11688 (N_11688,N_11234,N_11263);
or U11689 (N_11689,N_11154,N_11026);
nor U11690 (N_11690,N_11449,N_11213);
xor U11691 (N_11691,N_11485,N_11256);
and U11692 (N_11692,N_11211,N_11031);
and U11693 (N_11693,N_11440,N_11285);
xor U11694 (N_11694,N_11460,N_11330);
nor U11695 (N_11695,N_11061,N_11498);
nand U11696 (N_11696,N_11314,N_11406);
xnor U11697 (N_11697,N_11177,N_11018);
nand U11698 (N_11698,N_11206,N_11367);
nor U11699 (N_11699,N_11295,N_11335);
nand U11700 (N_11700,N_11254,N_11483);
nand U11701 (N_11701,N_11037,N_11331);
nor U11702 (N_11702,N_11349,N_11114);
nand U11703 (N_11703,N_11388,N_11452);
and U11704 (N_11704,N_11299,N_11322);
or U11705 (N_11705,N_11059,N_11434);
xor U11706 (N_11706,N_11252,N_11379);
nand U11707 (N_11707,N_11473,N_11267);
nor U11708 (N_11708,N_11145,N_11327);
nand U11709 (N_11709,N_11102,N_11495);
or U11710 (N_11710,N_11156,N_11403);
and U11711 (N_11711,N_11326,N_11044);
or U11712 (N_11712,N_11164,N_11359);
and U11713 (N_11713,N_11153,N_11253);
or U11714 (N_11714,N_11470,N_11266);
or U11715 (N_11715,N_11074,N_11340);
nor U11716 (N_11716,N_11344,N_11136);
nor U11717 (N_11717,N_11100,N_11247);
or U11718 (N_11718,N_11472,N_11241);
nor U11719 (N_11719,N_11245,N_11009);
nor U11720 (N_11720,N_11307,N_11115);
nor U11721 (N_11721,N_11203,N_11444);
nand U11722 (N_11722,N_11337,N_11277);
nor U11723 (N_11723,N_11459,N_11468);
and U11724 (N_11724,N_11007,N_11152);
xnor U11725 (N_11725,N_11093,N_11041);
nor U11726 (N_11726,N_11077,N_11370);
nand U11727 (N_11727,N_11454,N_11140);
nand U11728 (N_11728,N_11192,N_11028);
and U11729 (N_11729,N_11298,N_11323);
nor U11730 (N_11730,N_11416,N_11204);
and U11731 (N_11731,N_11010,N_11265);
xor U11732 (N_11732,N_11067,N_11420);
xor U11733 (N_11733,N_11238,N_11448);
and U11734 (N_11734,N_11027,N_11220);
xor U11735 (N_11735,N_11232,N_11171);
xor U11736 (N_11736,N_11022,N_11088);
nand U11737 (N_11737,N_11489,N_11419);
xnor U11738 (N_11738,N_11339,N_11325);
or U11739 (N_11739,N_11458,N_11393);
and U11740 (N_11740,N_11094,N_11433);
xnor U11741 (N_11741,N_11357,N_11217);
nand U11742 (N_11742,N_11345,N_11424);
or U11743 (N_11743,N_11301,N_11187);
nor U11744 (N_11744,N_11288,N_11003);
and U11745 (N_11745,N_11083,N_11412);
and U11746 (N_11746,N_11401,N_11387);
xnor U11747 (N_11747,N_11487,N_11334);
nor U11748 (N_11748,N_11248,N_11333);
or U11749 (N_11749,N_11197,N_11271);
nor U11750 (N_11750,N_11243,N_11220);
nand U11751 (N_11751,N_11243,N_11164);
or U11752 (N_11752,N_11141,N_11084);
xnor U11753 (N_11753,N_11361,N_11335);
nand U11754 (N_11754,N_11278,N_11361);
nor U11755 (N_11755,N_11092,N_11468);
or U11756 (N_11756,N_11114,N_11402);
nor U11757 (N_11757,N_11425,N_11463);
nand U11758 (N_11758,N_11039,N_11440);
nor U11759 (N_11759,N_11381,N_11378);
or U11760 (N_11760,N_11409,N_11338);
or U11761 (N_11761,N_11051,N_11208);
nor U11762 (N_11762,N_11089,N_11374);
nor U11763 (N_11763,N_11119,N_11427);
or U11764 (N_11764,N_11141,N_11032);
xor U11765 (N_11765,N_11487,N_11055);
and U11766 (N_11766,N_11271,N_11455);
nor U11767 (N_11767,N_11253,N_11297);
nand U11768 (N_11768,N_11119,N_11452);
xnor U11769 (N_11769,N_11351,N_11293);
nor U11770 (N_11770,N_11149,N_11126);
and U11771 (N_11771,N_11188,N_11380);
and U11772 (N_11772,N_11430,N_11272);
or U11773 (N_11773,N_11082,N_11171);
xor U11774 (N_11774,N_11352,N_11229);
and U11775 (N_11775,N_11459,N_11051);
xnor U11776 (N_11776,N_11415,N_11072);
and U11777 (N_11777,N_11114,N_11391);
or U11778 (N_11778,N_11229,N_11334);
and U11779 (N_11779,N_11090,N_11013);
and U11780 (N_11780,N_11256,N_11332);
or U11781 (N_11781,N_11451,N_11180);
or U11782 (N_11782,N_11357,N_11285);
xor U11783 (N_11783,N_11248,N_11027);
or U11784 (N_11784,N_11463,N_11234);
or U11785 (N_11785,N_11329,N_11409);
nor U11786 (N_11786,N_11261,N_11267);
xor U11787 (N_11787,N_11009,N_11139);
nand U11788 (N_11788,N_11429,N_11422);
nand U11789 (N_11789,N_11027,N_11463);
or U11790 (N_11790,N_11473,N_11180);
nor U11791 (N_11791,N_11445,N_11235);
nand U11792 (N_11792,N_11219,N_11064);
nand U11793 (N_11793,N_11227,N_11233);
nor U11794 (N_11794,N_11403,N_11236);
nor U11795 (N_11795,N_11198,N_11489);
nand U11796 (N_11796,N_11053,N_11282);
xor U11797 (N_11797,N_11081,N_11059);
xor U11798 (N_11798,N_11216,N_11499);
or U11799 (N_11799,N_11361,N_11301);
nand U11800 (N_11800,N_11399,N_11482);
xor U11801 (N_11801,N_11201,N_11474);
or U11802 (N_11802,N_11285,N_11115);
xnor U11803 (N_11803,N_11264,N_11321);
and U11804 (N_11804,N_11452,N_11194);
nand U11805 (N_11805,N_11377,N_11277);
nor U11806 (N_11806,N_11415,N_11350);
nand U11807 (N_11807,N_11483,N_11213);
nand U11808 (N_11808,N_11107,N_11203);
xor U11809 (N_11809,N_11389,N_11344);
nand U11810 (N_11810,N_11133,N_11354);
and U11811 (N_11811,N_11181,N_11275);
or U11812 (N_11812,N_11191,N_11424);
xnor U11813 (N_11813,N_11130,N_11495);
and U11814 (N_11814,N_11261,N_11252);
nor U11815 (N_11815,N_11270,N_11412);
and U11816 (N_11816,N_11353,N_11307);
or U11817 (N_11817,N_11429,N_11049);
and U11818 (N_11818,N_11386,N_11050);
and U11819 (N_11819,N_11136,N_11086);
nor U11820 (N_11820,N_11068,N_11290);
nor U11821 (N_11821,N_11237,N_11026);
or U11822 (N_11822,N_11424,N_11404);
nor U11823 (N_11823,N_11103,N_11101);
xor U11824 (N_11824,N_11082,N_11295);
or U11825 (N_11825,N_11217,N_11458);
nor U11826 (N_11826,N_11192,N_11492);
xnor U11827 (N_11827,N_11478,N_11442);
or U11828 (N_11828,N_11443,N_11049);
xnor U11829 (N_11829,N_11457,N_11423);
nor U11830 (N_11830,N_11173,N_11220);
nand U11831 (N_11831,N_11110,N_11372);
and U11832 (N_11832,N_11249,N_11378);
xnor U11833 (N_11833,N_11330,N_11411);
xor U11834 (N_11834,N_11300,N_11393);
xnor U11835 (N_11835,N_11304,N_11448);
nor U11836 (N_11836,N_11268,N_11164);
and U11837 (N_11837,N_11103,N_11339);
or U11838 (N_11838,N_11128,N_11135);
nor U11839 (N_11839,N_11350,N_11375);
or U11840 (N_11840,N_11295,N_11127);
or U11841 (N_11841,N_11364,N_11176);
nor U11842 (N_11842,N_11215,N_11362);
nor U11843 (N_11843,N_11323,N_11204);
and U11844 (N_11844,N_11365,N_11074);
and U11845 (N_11845,N_11430,N_11015);
or U11846 (N_11846,N_11118,N_11284);
nor U11847 (N_11847,N_11236,N_11228);
or U11848 (N_11848,N_11203,N_11038);
xor U11849 (N_11849,N_11186,N_11277);
nor U11850 (N_11850,N_11167,N_11200);
xnor U11851 (N_11851,N_11007,N_11017);
and U11852 (N_11852,N_11228,N_11268);
nor U11853 (N_11853,N_11140,N_11356);
nor U11854 (N_11854,N_11325,N_11193);
or U11855 (N_11855,N_11086,N_11473);
xor U11856 (N_11856,N_11382,N_11286);
and U11857 (N_11857,N_11390,N_11473);
and U11858 (N_11858,N_11092,N_11118);
nand U11859 (N_11859,N_11017,N_11375);
and U11860 (N_11860,N_11345,N_11070);
and U11861 (N_11861,N_11299,N_11000);
nor U11862 (N_11862,N_11168,N_11486);
xnor U11863 (N_11863,N_11231,N_11131);
xnor U11864 (N_11864,N_11442,N_11284);
and U11865 (N_11865,N_11491,N_11442);
nor U11866 (N_11866,N_11426,N_11367);
or U11867 (N_11867,N_11308,N_11147);
and U11868 (N_11868,N_11323,N_11056);
and U11869 (N_11869,N_11046,N_11280);
nand U11870 (N_11870,N_11122,N_11288);
and U11871 (N_11871,N_11189,N_11289);
and U11872 (N_11872,N_11182,N_11294);
nand U11873 (N_11873,N_11211,N_11071);
nand U11874 (N_11874,N_11330,N_11435);
nor U11875 (N_11875,N_11259,N_11275);
nand U11876 (N_11876,N_11111,N_11220);
nand U11877 (N_11877,N_11488,N_11360);
and U11878 (N_11878,N_11259,N_11100);
nand U11879 (N_11879,N_11168,N_11165);
nor U11880 (N_11880,N_11210,N_11446);
nor U11881 (N_11881,N_11287,N_11437);
or U11882 (N_11882,N_11030,N_11420);
and U11883 (N_11883,N_11415,N_11352);
and U11884 (N_11884,N_11022,N_11205);
nand U11885 (N_11885,N_11012,N_11375);
xnor U11886 (N_11886,N_11219,N_11225);
and U11887 (N_11887,N_11255,N_11094);
and U11888 (N_11888,N_11000,N_11016);
nand U11889 (N_11889,N_11414,N_11410);
nand U11890 (N_11890,N_11402,N_11381);
nor U11891 (N_11891,N_11284,N_11316);
xnor U11892 (N_11892,N_11147,N_11478);
nor U11893 (N_11893,N_11344,N_11248);
nand U11894 (N_11894,N_11169,N_11086);
xor U11895 (N_11895,N_11257,N_11112);
and U11896 (N_11896,N_11373,N_11030);
xor U11897 (N_11897,N_11182,N_11006);
nand U11898 (N_11898,N_11050,N_11455);
nor U11899 (N_11899,N_11006,N_11446);
and U11900 (N_11900,N_11202,N_11280);
xor U11901 (N_11901,N_11365,N_11247);
or U11902 (N_11902,N_11023,N_11462);
nand U11903 (N_11903,N_11427,N_11000);
nand U11904 (N_11904,N_11186,N_11495);
nor U11905 (N_11905,N_11041,N_11434);
nor U11906 (N_11906,N_11296,N_11433);
or U11907 (N_11907,N_11394,N_11038);
and U11908 (N_11908,N_11445,N_11373);
nor U11909 (N_11909,N_11298,N_11304);
or U11910 (N_11910,N_11161,N_11058);
nand U11911 (N_11911,N_11237,N_11084);
or U11912 (N_11912,N_11294,N_11429);
nand U11913 (N_11913,N_11096,N_11182);
xnor U11914 (N_11914,N_11322,N_11265);
or U11915 (N_11915,N_11425,N_11401);
nor U11916 (N_11916,N_11203,N_11300);
and U11917 (N_11917,N_11239,N_11032);
nor U11918 (N_11918,N_11175,N_11177);
xor U11919 (N_11919,N_11488,N_11040);
or U11920 (N_11920,N_11008,N_11092);
and U11921 (N_11921,N_11307,N_11232);
nand U11922 (N_11922,N_11059,N_11469);
xnor U11923 (N_11923,N_11439,N_11201);
nand U11924 (N_11924,N_11098,N_11005);
and U11925 (N_11925,N_11445,N_11081);
and U11926 (N_11926,N_11139,N_11126);
xor U11927 (N_11927,N_11333,N_11169);
nand U11928 (N_11928,N_11247,N_11126);
nand U11929 (N_11929,N_11382,N_11495);
or U11930 (N_11930,N_11005,N_11299);
xor U11931 (N_11931,N_11164,N_11112);
and U11932 (N_11932,N_11428,N_11456);
nand U11933 (N_11933,N_11297,N_11380);
xor U11934 (N_11934,N_11381,N_11400);
and U11935 (N_11935,N_11091,N_11155);
nand U11936 (N_11936,N_11020,N_11118);
xor U11937 (N_11937,N_11224,N_11464);
or U11938 (N_11938,N_11337,N_11055);
and U11939 (N_11939,N_11369,N_11165);
nor U11940 (N_11940,N_11488,N_11099);
and U11941 (N_11941,N_11044,N_11320);
nand U11942 (N_11942,N_11253,N_11047);
nand U11943 (N_11943,N_11186,N_11247);
nand U11944 (N_11944,N_11052,N_11457);
xnor U11945 (N_11945,N_11148,N_11495);
nor U11946 (N_11946,N_11055,N_11128);
or U11947 (N_11947,N_11429,N_11455);
xnor U11948 (N_11948,N_11422,N_11475);
or U11949 (N_11949,N_11082,N_11076);
xor U11950 (N_11950,N_11488,N_11306);
nor U11951 (N_11951,N_11257,N_11318);
and U11952 (N_11952,N_11117,N_11367);
nor U11953 (N_11953,N_11033,N_11278);
nand U11954 (N_11954,N_11272,N_11442);
nand U11955 (N_11955,N_11248,N_11144);
nor U11956 (N_11956,N_11008,N_11228);
or U11957 (N_11957,N_11160,N_11422);
nand U11958 (N_11958,N_11012,N_11007);
xnor U11959 (N_11959,N_11107,N_11220);
xnor U11960 (N_11960,N_11296,N_11254);
and U11961 (N_11961,N_11035,N_11437);
nor U11962 (N_11962,N_11433,N_11319);
xnor U11963 (N_11963,N_11376,N_11412);
xor U11964 (N_11964,N_11030,N_11354);
xor U11965 (N_11965,N_11089,N_11018);
xnor U11966 (N_11966,N_11436,N_11083);
nor U11967 (N_11967,N_11238,N_11207);
or U11968 (N_11968,N_11365,N_11163);
or U11969 (N_11969,N_11241,N_11415);
or U11970 (N_11970,N_11440,N_11091);
nor U11971 (N_11971,N_11335,N_11203);
or U11972 (N_11972,N_11057,N_11331);
nand U11973 (N_11973,N_11161,N_11467);
and U11974 (N_11974,N_11005,N_11226);
and U11975 (N_11975,N_11307,N_11395);
or U11976 (N_11976,N_11079,N_11073);
and U11977 (N_11977,N_11306,N_11149);
nand U11978 (N_11978,N_11047,N_11004);
and U11979 (N_11979,N_11325,N_11047);
nor U11980 (N_11980,N_11412,N_11447);
and U11981 (N_11981,N_11068,N_11220);
or U11982 (N_11982,N_11246,N_11495);
xor U11983 (N_11983,N_11180,N_11373);
nand U11984 (N_11984,N_11070,N_11491);
nand U11985 (N_11985,N_11422,N_11198);
nor U11986 (N_11986,N_11271,N_11105);
or U11987 (N_11987,N_11444,N_11231);
nand U11988 (N_11988,N_11491,N_11215);
nand U11989 (N_11989,N_11421,N_11307);
xnor U11990 (N_11990,N_11374,N_11402);
nor U11991 (N_11991,N_11487,N_11112);
and U11992 (N_11992,N_11344,N_11392);
and U11993 (N_11993,N_11346,N_11301);
nand U11994 (N_11994,N_11066,N_11423);
and U11995 (N_11995,N_11217,N_11312);
xor U11996 (N_11996,N_11044,N_11416);
nand U11997 (N_11997,N_11403,N_11266);
and U11998 (N_11998,N_11214,N_11060);
nand U11999 (N_11999,N_11115,N_11068);
and U12000 (N_12000,N_11801,N_11796);
or U12001 (N_12001,N_11651,N_11533);
xor U12002 (N_12002,N_11863,N_11840);
or U12003 (N_12003,N_11734,N_11810);
nand U12004 (N_12004,N_11973,N_11527);
or U12005 (N_12005,N_11701,N_11592);
nor U12006 (N_12006,N_11587,N_11511);
nor U12007 (N_12007,N_11871,N_11659);
nor U12008 (N_12008,N_11784,N_11621);
and U12009 (N_12009,N_11697,N_11931);
nand U12010 (N_12010,N_11635,N_11661);
nor U12011 (N_12011,N_11685,N_11773);
nand U12012 (N_12012,N_11769,N_11662);
nand U12013 (N_12013,N_11905,N_11792);
and U12014 (N_12014,N_11517,N_11892);
xor U12015 (N_12015,N_11770,N_11934);
xnor U12016 (N_12016,N_11790,N_11837);
and U12017 (N_12017,N_11620,N_11829);
nand U12018 (N_12018,N_11704,N_11855);
nor U12019 (N_12019,N_11739,N_11648);
nor U12020 (N_12020,N_11509,N_11588);
or U12021 (N_12021,N_11961,N_11619);
nand U12022 (N_12022,N_11921,N_11660);
nor U12023 (N_12023,N_11839,N_11761);
and U12024 (N_12024,N_11713,N_11766);
nand U12025 (N_12025,N_11938,N_11847);
xnor U12026 (N_12026,N_11678,N_11927);
nand U12027 (N_12027,N_11512,N_11744);
or U12028 (N_12028,N_11644,N_11836);
xor U12029 (N_12029,N_11671,N_11747);
nand U12030 (N_12030,N_11756,N_11989);
and U12031 (N_12031,N_11788,N_11578);
and U12032 (N_12032,N_11876,N_11960);
nand U12033 (N_12033,N_11835,N_11944);
or U12034 (N_12034,N_11866,N_11502);
nand U12035 (N_12035,N_11958,N_11872);
and U12036 (N_12036,N_11825,N_11986);
nor U12037 (N_12037,N_11993,N_11643);
xor U12038 (N_12038,N_11645,N_11904);
or U12039 (N_12039,N_11504,N_11545);
xor U12040 (N_12040,N_11560,N_11575);
nor U12041 (N_12041,N_11748,N_11615);
or U12042 (N_12042,N_11966,N_11984);
or U12043 (N_12043,N_11548,N_11689);
xor U12044 (N_12044,N_11817,N_11983);
nor U12045 (N_12045,N_11994,N_11918);
and U12046 (N_12046,N_11637,N_11561);
and U12047 (N_12047,N_11922,N_11742);
and U12048 (N_12048,N_11719,N_11636);
xor U12049 (N_12049,N_11864,N_11534);
xor U12050 (N_12050,N_11939,N_11752);
or U12051 (N_12051,N_11813,N_11577);
or U12052 (N_12052,N_11584,N_11711);
and U12053 (N_12053,N_11672,N_11781);
nand U12054 (N_12054,N_11702,N_11946);
and U12055 (N_12055,N_11755,N_11674);
nor U12056 (N_12056,N_11928,N_11873);
or U12057 (N_12057,N_11599,N_11915);
nand U12058 (N_12058,N_11795,N_11731);
nand U12059 (N_12059,N_11604,N_11688);
or U12060 (N_12060,N_11594,N_11874);
nand U12061 (N_12061,N_11799,N_11505);
and U12062 (N_12062,N_11543,N_11700);
nand U12063 (N_12063,N_11771,N_11694);
nor U12064 (N_12064,N_11733,N_11858);
nand U12065 (N_12065,N_11913,N_11664);
nor U12066 (N_12066,N_11881,N_11880);
nand U12067 (N_12067,N_11978,N_11554);
and U12068 (N_12068,N_11628,N_11914);
nor U12069 (N_12069,N_11806,N_11573);
and U12070 (N_12070,N_11682,N_11895);
nand U12071 (N_12071,N_11617,N_11725);
or U12072 (N_12072,N_11624,N_11550);
nor U12073 (N_12073,N_11528,N_11998);
and U12074 (N_12074,N_11859,N_11764);
nand U12075 (N_12075,N_11917,N_11687);
xor U12076 (N_12076,N_11544,N_11708);
and U12077 (N_12077,N_11970,N_11805);
and U12078 (N_12078,N_11997,N_11727);
and U12079 (N_12079,N_11540,N_11558);
nor U12080 (N_12080,N_11783,N_11654);
and U12081 (N_12081,N_11794,N_11536);
nor U12082 (N_12082,N_11812,N_11878);
and U12083 (N_12083,N_11759,N_11572);
and U12084 (N_12084,N_11570,N_11912);
nand U12085 (N_12085,N_11598,N_11862);
and U12086 (N_12086,N_11525,N_11516);
nor U12087 (N_12087,N_11832,N_11552);
and U12088 (N_12088,N_11924,N_11556);
xnor U12089 (N_12089,N_11894,N_11684);
xnor U12090 (N_12090,N_11768,N_11630);
and U12091 (N_12091,N_11853,N_11987);
nor U12092 (N_12092,N_11699,N_11633);
or U12093 (N_12093,N_11816,N_11721);
xnor U12094 (N_12094,N_11948,N_11562);
nor U12095 (N_12095,N_11585,N_11597);
nor U12096 (N_12096,N_11860,N_11897);
or U12097 (N_12097,N_11683,N_11532);
xnor U12098 (N_12098,N_11740,N_11510);
xnor U12099 (N_12099,N_11717,N_11798);
nand U12100 (N_12100,N_11963,N_11696);
or U12101 (N_12101,N_11977,N_11808);
or U12102 (N_12102,N_11907,N_11567);
or U12103 (N_12103,N_11888,N_11580);
nor U12104 (N_12104,N_11618,N_11555);
nor U12105 (N_12105,N_11677,N_11531);
and U12106 (N_12106,N_11841,N_11911);
nor U12107 (N_12107,N_11551,N_11830);
and U12108 (N_12108,N_11842,N_11953);
xor U12109 (N_12109,N_11564,N_11667);
nor U12110 (N_12110,N_11823,N_11956);
and U12111 (N_12111,N_11899,N_11736);
nor U12112 (N_12112,N_11519,N_11668);
and U12113 (N_12113,N_11666,N_11879);
nand U12114 (N_12114,N_11906,N_11967);
and U12115 (N_12115,N_11760,N_11965);
nor U12116 (N_12116,N_11869,N_11609);
or U12117 (N_12117,N_11949,N_11820);
nor U12118 (N_12118,N_11779,N_11821);
nand U12119 (N_12119,N_11925,N_11882);
xor U12120 (N_12120,N_11542,N_11732);
and U12121 (N_12121,N_11896,N_11787);
nor U12122 (N_12122,N_11908,N_11652);
or U12123 (N_12123,N_11990,N_11501);
xor U12124 (N_12124,N_11523,N_11707);
nand U12125 (N_12125,N_11613,N_11591);
xor U12126 (N_12126,N_11933,N_11951);
and U12127 (N_12127,N_11901,N_11774);
nand U12128 (N_12128,N_11526,N_11935);
nor U12129 (N_12129,N_11930,N_11690);
or U12130 (N_12130,N_11507,N_11607);
and U12131 (N_12131,N_11920,N_11681);
and U12132 (N_12132,N_11581,N_11718);
and U12133 (N_12133,N_11898,N_11947);
xnor U12134 (N_12134,N_11834,N_11815);
nor U12135 (N_12135,N_11601,N_11658);
and U12136 (N_12136,N_11614,N_11706);
nor U12137 (N_12137,N_11826,N_11665);
xor U12138 (N_12138,N_11969,N_11565);
or U12139 (N_12139,N_11656,N_11720);
nor U12140 (N_12140,N_11846,N_11524);
or U12141 (N_12141,N_11877,N_11539);
nor U12142 (N_12142,N_11715,N_11566);
nand U12143 (N_12143,N_11843,N_11680);
and U12144 (N_12144,N_11714,N_11802);
nand U12145 (N_12145,N_11549,N_11576);
nor U12146 (N_12146,N_11596,N_11698);
nor U12147 (N_12147,N_11608,N_11778);
xor U12148 (N_12148,N_11603,N_11776);
nor U12149 (N_12149,N_11522,N_11849);
or U12150 (N_12150,N_11735,N_11968);
and U12151 (N_12151,N_11809,N_11940);
and U12152 (N_12152,N_11828,N_11950);
xor U12153 (N_12153,N_11926,N_11954);
and U12154 (N_12154,N_11765,N_11515);
and U12155 (N_12155,N_11503,N_11602);
and U12156 (N_12156,N_11647,N_11582);
or U12157 (N_12157,N_11612,N_11606);
and U12158 (N_12158,N_11883,N_11945);
nand U12159 (N_12159,N_11807,N_11762);
and U12160 (N_12160,N_11500,N_11589);
and U12161 (N_12161,N_11791,N_11722);
or U12162 (N_12162,N_11590,N_11514);
or U12163 (N_12163,N_11726,N_11831);
or U12164 (N_12164,N_11982,N_11646);
nor U12165 (N_12165,N_11738,N_11886);
and U12166 (N_12166,N_11691,N_11639);
xnor U12167 (N_12167,N_11610,N_11669);
or U12168 (N_12168,N_11593,N_11657);
and U12169 (N_12169,N_11673,N_11981);
nand U12170 (N_12170,N_11936,N_11793);
or U12171 (N_12171,N_11955,N_11723);
nand U12172 (N_12172,N_11885,N_11749);
or U12173 (N_12173,N_11976,N_11838);
nand U12174 (N_12174,N_11586,N_11649);
and U12175 (N_12175,N_11746,N_11557);
and U12176 (N_12176,N_11579,N_11979);
nand U12177 (N_12177,N_11985,N_11916);
xor U12178 (N_12178,N_11852,N_11663);
or U12179 (N_12179,N_11757,N_11943);
xnor U12180 (N_12180,N_11937,N_11992);
and U12181 (N_12181,N_11754,N_11942);
nand U12182 (N_12182,N_11632,N_11775);
xor U12183 (N_12183,N_11919,N_11634);
and U12184 (N_12184,N_11971,N_11996);
or U12185 (N_12185,N_11767,N_11571);
xor U12186 (N_12186,N_11785,N_11959);
and U12187 (N_12187,N_11583,N_11642);
and U12188 (N_12188,N_11595,N_11811);
nand U12189 (N_12189,N_11988,N_11854);
nor U12190 (N_12190,N_11626,N_11995);
and U12191 (N_12191,N_11695,N_11513);
or U12192 (N_12192,N_11909,N_11903);
and U12193 (N_12193,N_11709,N_11716);
and U12194 (N_12194,N_11743,N_11758);
or U12195 (N_12195,N_11848,N_11991);
or U12196 (N_12196,N_11975,N_11563);
and U12197 (N_12197,N_11675,N_11999);
nand U12198 (N_12198,N_11900,N_11623);
nor U12199 (N_12199,N_11941,N_11627);
nand U12200 (N_12200,N_11867,N_11751);
nand U12201 (N_12201,N_11692,N_11957);
and U12202 (N_12202,N_11889,N_11833);
xnor U12203 (N_12203,N_11962,N_11710);
or U12204 (N_12204,N_11875,N_11803);
or U12205 (N_12205,N_11737,N_11753);
nand U12206 (N_12206,N_11827,N_11508);
or U12207 (N_12207,N_11529,N_11800);
or U12208 (N_12208,N_11891,N_11728);
or U12209 (N_12209,N_11605,N_11670);
nor U12210 (N_12210,N_11521,N_11676);
and U12211 (N_12211,N_11535,N_11686);
nor U12212 (N_12212,N_11655,N_11818);
or U12213 (N_12213,N_11705,N_11520);
and U12214 (N_12214,N_11845,N_11822);
nand U12215 (N_12215,N_11629,N_11729);
nor U12216 (N_12216,N_11538,N_11641);
or U12217 (N_12217,N_11972,N_11763);
or U12218 (N_12218,N_11750,N_11547);
and U12219 (N_12219,N_11964,N_11703);
and U12220 (N_12220,N_11797,N_11541);
xor U12221 (N_12221,N_11884,N_11786);
and U12222 (N_12222,N_11518,N_11851);
nor U12223 (N_12223,N_11625,N_11653);
nand U12224 (N_12224,N_11923,N_11824);
nand U12225 (N_12225,N_11569,N_11910);
or U12226 (N_12226,N_11616,N_11780);
and U12227 (N_12227,N_11568,N_11857);
nand U12228 (N_12228,N_11574,N_11902);
nor U12229 (N_12229,N_11952,N_11782);
nor U12230 (N_12230,N_11600,N_11819);
nand U12231 (N_12231,N_11932,N_11804);
xor U12232 (N_12232,N_11865,N_11506);
or U12233 (N_12233,N_11559,N_11929);
nand U12234 (N_12234,N_11814,N_11530);
and U12235 (N_12235,N_11638,N_11844);
or U12236 (N_12236,N_11890,N_11745);
xor U12237 (N_12237,N_11650,N_11611);
and U12238 (N_12238,N_11679,N_11546);
nand U12239 (N_12239,N_11789,N_11870);
nand U12240 (N_12240,N_11631,N_11693);
or U12241 (N_12241,N_11537,N_11893);
xnor U12242 (N_12242,N_11980,N_11868);
nand U12243 (N_12243,N_11640,N_11712);
nor U12244 (N_12244,N_11730,N_11741);
nor U12245 (N_12245,N_11887,N_11622);
or U12246 (N_12246,N_11861,N_11974);
nor U12247 (N_12247,N_11856,N_11850);
nor U12248 (N_12248,N_11724,N_11553);
xor U12249 (N_12249,N_11772,N_11777);
or U12250 (N_12250,N_11737,N_11865);
xnor U12251 (N_12251,N_11897,N_11793);
nor U12252 (N_12252,N_11520,N_11693);
or U12253 (N_12253,N_11655,N_11887);
nand U12254 (N_12254,N_11932,N_11887);
and U12255 (N_12255,N_11617,N_11515);
or U12256 (N_12256,N_11680,N_11799);
or U12257 (N_12257,N_11868,N_11832);
and U12258 (N_12258,N_11999,N_11613);
xor U12259 (N_12259,N_11728,N_11745);
xor U12260 (N_12260,N_11851,N_11598);
or U12261 (N_12261,N_11831,N_11657);
nand U12262 (N_12262,N_11574,N_11706);
nor U12263 (N_12263,N_11506,N_11690);
xor U12264 (N_12264,N_11539,N_11956);
or U12265 (N_12265,N_11634,N_11898);
or U12266 (N_12266,N_11583,N_11633);
nor U12267 (N_12267,N_11874,N_11717);
xor U12268 (N_12268,N_11584,N_11960);
nor U12269 (N_12269,N_11659,N_11865);
nand U12270 (N_12270,N_11721,N_11588);
xnor U12271 (N_12271,N_11993,N_11615);
xor U12272 (N_12272,N_11699,N_11862);
and U12273 (N_12273,N_11947,N_11844);
or U12274 (N_12274,N_11853,N_11916);
xor U12275 (N_12275,N_11743,N_11765);
or U12276 (N_12276,N_11717,N_11556);
xor U12277 (N_12277,N_11788,N_11773);
nand U12278 (N_12278,N_11533,N_11657);
nand U12279 (N_12279,N_11628,N_11500);
and U12280 (N_12280,N_11920,N_11864);
or U12281 (N_12281,N_11872,N_11639);
and U12282 (N_12282,N_11613,N_11635);
nand U12283 (N_12283,N_11869,N_11649);
nor U12284 (N_12284,N_11542,N_11814);
nand U12285 (N_12285,N_11801,N_11967);
nand U12286 (N_12286,N_11657,N_11806);
xnor U12287 (N_12287,N_11701,N_11652);
xor U12288 (N_12288,N_11639,N_11503);
nor U12289 (N_12289,N_11568,N_11528);
nor U12290 (N_12290,N_11734,N_11630);
and U12291 (N_12291,N_11729,N_11717);
xor U12292 (N_12292,N_11503,N_11598);
xor U12293 (N_12293,N_11515,N_11545);
nor U12294 (N_12294,N_11731,N_11580);
nor U12295 (N_12295,N_11766,N_11530);
or U12296 (N_12296,N_11591,N_11717);
nor U12297 (N_12297,N_11571,N_11720);
xor U12298 (N_12298,N_11572,N_11702);
or U12299 (N_12299,N_11674,N_11739);
and U12300 (N_12300,N_11689,N_11960);
and U12301 (N_12301,N_11832,N_11654);
or U12302 (N_12302,N_11643,N_11674);
or U12303 (N_12303,N_11898,N_11817);
or U12304 (N_12304,N_11976,N_11874);
xor U12305 (N_12305,N_11664,N_11511);
and U12306 (N_12306,N_11720,N_11744);
or U12307 (N_12307,N_11633,N_11952);
or U12308 (N_12308,N_11745,N_11945);
nand U12309 (N_12309,N_11619,N_11527);
and U12310 (N_12310,N_11651,N_11550);
xnor U12311 (N_12311,N_11979,N_11877);
and U12312 (N_12312,N_11939,N_11839);
or U12313 (N_12313,N_11903,N_11623);
nor U12314 (N_12314,N_11904,N_11712);
nor U12315 (N_12315,N_11568,N_11804);
xor U12316 (N_12316,N_11658,N_11798);
nor U12317 (N_12317,N_11762,N_11684);
nand U12318 (N_12318,N_11605,N_11689);
or U12319 (N_12319,N_11502,N_11653);
or U12320 (N_12320,N_11731,N_11707);
nand U12321 (N_12321,N_11765,N_11694);
nand U12322 (N_12322,N_11793,N_11611);
or U12323 (N_12323,N_11570,N_11833);
or U12324 (N_12324,N_11928,N_11661);
or U12325 (N_12325,N_11525,N_11707);
and U12326 (N_12326,N_11830,N_11619);
xor U12327 (N_12327,N_11510,N_11798);
nand U12328 (N_12328,N_11644,N_11556);
nand U12329 (N_12329,N_11710,N_11977);
and U12330 (N_12330,N_11958,N_11579);
and U12331 (N_12331,N_11640,N_11636);
or U12332 (N_12332,N_11697,N_11520);
nand U12333 (N_12333,N_11598,N_11601);
and U12334 (N_12334,N_11621,N_11945);
nor U12335 (N_12335,N_11624,N_11836);
or U12336 (N_12336,N_11635,N_11504);
or U12337 (N_12337,N_11751,N_11585);
or U12338 (N_12338,N_11796,N_11531);
xnor U12339 (N_12339,N_11533,N_11807);
xor U12340 (N_12340,N_11590,N_11745);
or U12341 (N_12341,N_11646,N_11915);
nand U12342 (N_12342,N_11823,N_11765);
nor U12343 (N_12343,N_11950,N_11599);
or U12344 (N_12344,N_11878,N_11918);
or U12345 (N_12345,N_11937,N_11576);
xnor U12346 (N_12346,N_11534,N_11772);
and U12347 (N_12347,N_11805,N_11995);
nor U12348 (N_12348,N_11996,N_11796);
nand U12349 (N_12349,N_11567,N_11816);
and U12350 (N_12350,N_11987,N_11678);
nor U12351 (N_12351,N_11872,N_11819);
or U12352 (N_12352,N_11831,N_11834);
nand U12353 (N_12353,N_11707,N_11955);
xnor U12354 (N_12354,N_11987,N_11605);
xnor U12355 (N_12355,N_11767,N_11901);
xnor U12356 (N_12356,N_11945,N_11781);
nand U12357 (N_12357,N_11826,N_11556);
nor U12358 (N_12358,N_11510,N_11795);
nor U12359 (N_12359,N_11568,N_11961);
nor U12360 (N_12360,N_11795,N_11547);
nor U12361 (N_12361,N_11714,N_11583);
nand U12362 (N_12362,N_11801,N_11662);
xnor U12363 (N_12363,N_11653,N_11772);
nand U12364 (N_12364,N_11687,N_11708);
or U12365 (N_12365,N_11923,N_11992);
or U12366 (N_12366,N_11624,N_11757);
or U12367 (N_12367,N_11973,N_11989);
nor U12368 (N_12368,N_11933,N_11961);
nand U12369 (N_12369,N_11862,N_11962);
or U12370 (N_12370,N_11641,N_11837);
and U12371 (N_12371,N_11644,N_11883);
nor U12372 (N_12372,N_11626,N_11828);
and U12373 (N_12373,N_11788,N_11569);
and U12374 (N_12374,N_11953,N_11617);
xnor U12375 (N_12375,N_11584,N_11988);
and U12376 (N_12376,N_11939,N_11623);
nor U12377 (N_12377,N_11617,N_11934);
nand U12378 (N_12378,N_11848,N_11644);
xor U12379 (N_12379,N_11836,N_11956);
nand U12380 (N_12380,N_11673,N_11535);
nor U12381 (N_12381,N_11705,N_11771);
or U12382 (N_12382,N_11933,N_11545);
nor U12383 (N_12383,N_11710,N_11619);
xnor U12384 (N_12384,N_11627,N_11695);
and U12385 (N_12385,N_11796,N_11905);
xnor U12386 (N_12386,N_11940,N_11789);
nor U12387 (N_12387,N_11715,N_11737);
and U12388 (N_12388,N_11785,N_11636);
nor U12389 (N_12389,N_11701,N_11546);
and U12390 (N_12390,N_11892,N_11607);
xnor U12391 (N_12391,N_11842,N_11806);
or U12392 (N_12392,N_11718,N_11616);
nand U12393 (N_12393,N_11576,N_11912);
or U12394 (N_12394,N_11910,N_11920);
or U12395 (N_12395,N_11855,N_11929);
xnor U12396 (N_12396,N_11761,N_11986);
or U12397 (N_12397,N_11682,N_11818);
nor U12398 (N_12398,N_11584,N_11898);
nor U12399 (N_12399,N_11616,N_11586);
and U12400 (N_12400,N_11911,N_11706);
nor U12401 (N_12401,N_11815,N_11981);
nand U12402 (N_12402,N_11740,N_11965);
and U12403 (N_12403,N_11566,N_11661);
nor U12404 (N_12404,N_11569,N_11916);
nor U12405 (N_12405,N_11882,N_11962);
xnor U12406 (N_12406,N_11974,N_11995);
xnor U12407 (N_12407,N_11615,N_11570);
xor U12408 (N_12408,N_11794,N_11934);
nor U12409 (N_12409,N_11594,N_11646);
xor U12410 (N_12410,N_11673,N_11661);
or U12411 (N_12411,N_11883,N_11926);
nand U12412 (N_12412,N_11732,N_11847);
xor U12413 (N_12413,N_11861,N_11918);
or U12414 (N_12414,N_11546,N_11511);
and U12415 (N_12415,N_11591,N_11906);
nor U12416 (N_12416,N_11784,N_11585);
nor U12417 (N_12417,N_11667,N_11753);
and U12418 (N_12418,N_11615,N_11724);
nor U12419 (N_12419,N_11734,N_11802);
or U12420 (N_12420,N_11503,N_11969);
or U12421 (N_12421,N_11760,N_11719);
and U12422 (N_12422,N_11911,N_11568);
nor U12423 (N_12423,N_11767,N_11577);
nand U12424 (N_12424,N_11657,N_11527);
or U12425 (N_12425,N_11682,N_11656);
and U12426 (N_12426,N_11530,N_11749);
nand U12427 (N_12427,N_11710,N_11636);
nor U12428 (N_12428,N_11820,N_11853);
nor U12429 (N_12429,N_11543,N_11668);
nor U12430 (N_12430,N_11525,N_11553);
and U12431 (N_12431,N_11669,N_11946);
and U12432 (N_12432,N_11965,N_11694);
or U12433 (N_12433,N_11694,N_11783);
nand U12434 (N_12434,N_11530,N_11729);
and U12435 (N_12435,N_11771,N_11996);
xor U12436 (N_12436,N_11769,N_11589);
and U12437 (N_12437,N_11613,N_11593);
and U12438 (N_12438,N_11547,N_11951);
or U12439 (N_12439,N_11910,N_11979);
xor U12440 (N_12440,N_11652,N_11501);
or U12441 (N_12441,N_11876,N_11692);
nor U12442 (N_12442,N_11836,N_11581);
nor U12443 (N_12443,N_11990,N_11943);
nor U12444 (N_12444,N_11818,N_11972);
xor U12445 (N_12445,N_11934,N_11614);
nor U12446 (N_12446,N_11857,N_11660);
xnor U12447 (N_12447,N_11754,N_11654);
nand U12448 (N_12448,N_11589,N_11592);
xnor U12449 (N_12449,N_11637,N_11713);
or U12450 (N_12450,N_11529,N_11900);
nand U12451 (N_12451,N_11752,N_11706);
or U12452 (N_12452,N_11862,N_11957);
nor U12453 (N_12453,N_11632,N_11940);
or U12454 (N_12454,N_11797,N_11990);
xor U12455 (N_12455,N_11724,N_11623);
and U12456 (N_12456,N_11575,N_11981);
xnor U12457 (N_12457,N_11890,N_11510);
or U12458 (N_12458,N_11673,N_11651);
nor U12459 (N_12459,N_11984,N_11527);
and U12460 (N_12460,N_11655,N_11728);
or U12461 (N_12461,N_11568,N_11595);
nor U12462 (N_12462,N_11545,N_11644);
nor U12463 (N_12463,N_11739,N_11929);
xor U12464 (N_12464,N_11853,N_11977);
and U12465 (N_12465,N_11798,N_11864);
or U12466 (N_12466,N_11673,N_11746);
or U12467 (N_12467,N_11907,N_11862);
nor U12468 (N_12468,N_11847,N_11888);
nor U12469 (N_12469,N_11521,N_11834);
nand U12470 (N_12470,N_11563,N_11589);
or U12471 (N_12471,N_11693,N_11797);
nor U12472 (N_12472,N_11919,N_11647);
nand U12473 (N_12473,N_11696,N_11934);
xnor U12474 (N_12474,N_11542,N_11649);
nand U12475 (N_12475,N_11564,N_11912);
nand U12476 (N_12476,N_11941,N_11846);
nand U12477 (N_12477,N_11607,N_11543);
xnor U12478 (N_12478,N_11844,N_11848);
nor U12479 (N_12479,N_11522,N_11800);
nand U12480 (N_12480,N_11536,N_11737);
xnor U12481 (N_12481,N_11675,N_11511);
and U12482 (N_12482,N_11724,N_11717);
nor U12483 (N_12483,N_11873,N_11616);
nand U12484 (N_12484,N_11632,N_11900);
and U12485 (N_12485,N_11882,N_11573);
nand U12486 (N_12486,N_11786,N_11779);
nand U12487 (N_12487,N_11687,N_11728);
nand U12488 (N_12488,N_11974,N_11658);
xnor U12489 (N_12489,N_11744,N_11950);
or U12490 (N_12490,N_11645,N_11693);
nand U12491 (N_12491,N_11620,N_11910);
or U12492 (N_12492,N_11848,N_11561);
or U12493 (N_12493,N_11709,N_11525);
nor U12494 (N_12494,N_11868,N_11723);
nand U12495 (N_12495,N_11732,N_11600);
and U12496 (N_12496,N_11699,N_11723);
and U12497 (N_12497,N_11616,N_11843);
xnor U12498 (N_12498,N_11887,N_11538);
nand U12499 (N_12499,N_11589,N_11857);
nor U12500 (N_12500,N_12055,N_12020);
xnor U12501 (N_12501,N_12440,N_12271);
nor U12502 (N_12502,N_12322,N_12203);
or U12503 (N_12503,N_12135,N_12261);
or U12504 (N_12504,N_12302,N_12046);
or U12505 (N_12505,N_12007,N_12338);
or U12506 (N_12506,N_12009,N_12004);
or U12507 (N_12507,N_12354,N_12033);
nor U12508 (N_12508,N_12303,N_12433);
nand U12509 (N_12509,N_12325,N_12088);
nor U12510 (N_12510,N_12184,N_12052);
xor U12511 (N_12511,N_12437,N_12147);
xor U12512 (N_12512,N_12113,N_12213);
or U12513 (N_12513,N_12332,N_12152);
nand U12514 (N_12514,N_12132,N_12024);
or U12515 (N_12515,N_12498,N_12330);
or U12516 (N_12516,N_12427,N_12267);
nand U12517 (N_12517,N_12137,N_12171);
nand U12518 (N_12518,N_12413,N_12351);
xnor U12519 (N_12519,N_12443,N_12445);
nor U12520 (N_12520,N_12366,N_12396);
xnor U12521 (N_12521,N_12375,N_12476);
or U12522 (N_12522,N_12233,N_12090);
nand U12523 (N_12523,N_12238,N_12250);
xnor U12524 (N_12524,N_12352,N_12260);
and U12525 (N_12525,N_12000,N_12054);
nand U12526 (N_12526,N_12470,N_12160);
or U12527 (N_12527,N_12401,N_12071);
or U12528 (N_12528,N_12426,N_12157);
nand U12529 (N_12529,N_12166,N_12122);
nand U12530 (N_12530,N_12390,N_12191);
xor U12531 (N_12531,N_12008,N_12293);
and U12532 (N_12532,N_12156,N_12079);
or U12533 (N_12533,N_12255,N_12224);
nand U12534 (N_12534,N_12326,N_12223);
xor U12535 (N_12535,N_12386,N_12103);
xnor U12536 (N_12536,N_12339,N_12200);
or U12537 (N_12537,N_12497,N_12329);
and U12538 (N_12538,N_12111,N_12178);
or U12539 (N_12539,N_12116,N_12317);
or U12540 (N_12540,N_12406,N_12107);
xor U12541 (N_12541,N_12212,N_12381);
xnor U12542 (N_12542,N_12306,N_12202);
nor U12543 (N_12543,N_12370,N_12265);
xnor U12544 (N_12544,N_12123,N_12294);
xnor U12545 (N_12545,N_12006,N_12276);
xnor U12546 (N_12546,N_12320,N_12105);
nor U12547 (N_12547,N_12494,N_12448);
xor U12548 (N_12548,N_12488,N_12333);
xnor U12549 (N_12549,N_12242,N_12377);
nand U12550 (N_12550,N_12080,N_12095);
xor U12551 (N_12551,N_12419,N_12239);
xnor U12552 (N_12552,N_12415,N_12391);
or U12553 (N_12553,N_12279,N_12385);
nand U12554 (N_12554,N_12115,N_12049);
or U12555 (N_12555,N_12290,N_12272);
nand U12556 (N_12556,N_12145,N_12417);
and U12557 (N_12557,N_12360,N_12131);
nand U12558 (N_12558,N_12305,N_12268);
nor U12559 (N_12559,N_12134,N_12361);
nor U12560 (N_12560,N_12321,N_12349);
nand U12561 (N_12561,N_12138,N_12313);
nor U12562 (N_12562,N_12109,N_12291);
xnor U12563 (N_12563,N_12359,N_12042);
or U12564 (N_12564,N_12491,N_12379);
nor U12565 (N_12565,N_12258,N_12481);
xor U12566 (N_12566,N_12407,N_12136);
nand U12567 (N_12567,N_12285,N_12404);
nand U12568 (N_12568,N_12085,N_12344);
nor U12569 (N_12569,N_12314,N_12441);
and U12570 (N_12570,N_12382,N_12214);
xnor U12571 (N_12571,N_12167,N_12028);
nor U12572 (N_12572,N_12431,N_12133);
nand U12573 (N_12573,N_12193,N_12093);
and U12574 (N_12574,N_12014,N_12455);
xnor U12575 (N_12575,N_12101,N_12304);
and U12576 (N_12576,N_12149,N_12083);
nor U12577 (N_12577,N_12418,N_12402);
or U12578 (N_12578,N_12061,N_12403);
nand U12579 (N_12579,N_12310,N_12246);
and U12580 (N_12580,N_12438,N_12170);
and U12581 (N_12581,N_12034,N_12139);
xor U12582 (N_12582,N_12155,N_12192);
nor U12583 (N_12583,N_12266,N_12066);
xor U12584 (N_12584,N_12127,N_12311);
nand U12585 (N_12585,N_12281,N_12221);
or U12586 (N_12586,N_12289,N_12473);
nor U12587 (N_12587,N_12205,N_12493);
nand U12588 (N_12588,N_12274,N_12363);
nor U12589 (N_12589,N_12343,N_12197);
xnor U12590 (N_12590,N_12388,N_12462);
xnor U12591 (N_12591,N_12142,N_12432);
or U12592 (N_12592,N_12182,N_12451);
and U12593 (N_12593,N_12397,N_12316);
and U12594 (N_12594,N_12075,N_12183);
and U12595 (N_12595,N_12452,N_12172);
and U12596 (N_12596,N_12086,N_12056);
nor U12597 (N_12597,N_12236,N_12295);
xor U12598 (N_12598,N_12346,N_12496);
and U12599 (N_12599,N_12227,N_12120);
nand U12600 (N_12600,N_12015,N_12119);
nor U12601 (N_12601,N_12373,N_12057);
xor U12602 (N_12602,N_12051,N_12345);
and U12603 (N_12603,N_12082,N_12369);
nand U12604 (N_12604,N_12209,N_12254);
and U12605 (N_12605,N_12490,N_12199);
and U12606 (N_12606,N_12069,N_12282);
nand U12607 (N_12607,N_12169,N_12365);
or U12608 (N_12608,N_12424,N_12461);
or U12609 (N_12609,N_12472,N_12159);
or U12610 (N_12610,N_12060,N_12474);
xor U12611 (N_12611,N_12283,N_12237);
and U12612 (N_12612,N_12016,N_12168);
nand U12613 (N_12613,N_12031,N_12429);
nand U12614 (N_12614,N_12395,N_12226);
nand U12615 (N_12615,N_12298,N_12331);
nand U12616 (N_12616,N_12173,N_12324);
nand U12617 (N_12617,N_12252,N_12130);
or U12618 (N_12618,N_12161,N_12216);
and U12619 (N_12619,N_12464,N_12466);
xor U12620 (N_12620,N_12222,N_12175);
and U12621 (N_12621,N_12367,N_12078);
xnor U12622 (N_12622,N_12140,N_12450);
nand U12623 (N_12623,N_12334,N_12434);
nand U12624 (N_12624,N_12409,N_12231);
or U12625 (N_12625,N_12129,N_12019);
and U12626 (N_12626,N_12023,N_12387);
nand U12627 (N_12627,N_12411,N_12247);
xor U12628 (N_12628,N_12177,N_12074);
or U12629 (N_12629,N_12241,N_12341);
xnor U12630 (N_12630,N_12444,N_12243);
xnor U12631 (N_12631,N_12430,N_12297);
nand U12632 (N_12632,N_12483,N_12287);
nor U12633 (N_12633,N_12040,N_12368);
or U12634 (N_12634,N_12153,N_12005);
nand U12635 (N_12635,N_12141,N_12436);
nand U12636 (N_12636,N_12211,N_12220);
xnor U12637 (N_12637,N_12471,N_12463);
nor U12638 (N_12638,N_12479,N_12465);
nand U12639 (N_12639,N_12206,N_12357);
nor U12640 (N_12640,N_12154,N_12454);
nor U12641 (N_12641,N_12309,N_12301);
nand U12642 (N_12642,N_12335,N_12201);
nor U12643 (N_12643,N_12108,N_12414);
and U12644 (N_12644,N_12380,N_12067);
xor U12645 (N_12645,N_12245,N_12460);
xor U12646 (N_12646,N_12383,N_12398);
xnor U12647 (N_12647,N_12262,N_12084);
or U12648 (N_12648,N_12412,N_12050);
and U12649 (N_12649,N_12449,N_12356);
nand U12650 (N_12650,N_12013,N_12104);
nand U12651 (N_12651,N_12273,N_12043);
or U12652 (N_12652,N_12065,N_12002);
xor U12653 (N_12653,N_12336,N_12100);
nor U12654 (N_12654,N_12475,N_12277);
or U12655 (N_12655,N_12194,N_12208);
and U12656 (N_12656,N_12225,N_12076);
and U12657 (N_12657,N_12117,N_12143);
nand U12658 (N_12658,N_12393,N_12094);
or U12659 (N_12659,N_12089,N_12181);
and U12660 (N_12660,N_12376,N_12374);
and U12661 (N_12661,N_12392,N_12296);
and U12662 (N_12662,N_12469,N_12456);
nand U12663 (N_12663,N_12263,N_12187);
and U12664 (N_12664,N_12251,N_12045);
xor U12665 (N_12665,N_12308,N_12048);
xnor U12666 (N_12666,N_12499,N_12278);
or U12667 (N_12667,N_12106,N_12362);
nand U12668 (N_12668,N_12230,N_12328);
nand U12669 (N_12669,N_12010,N_12275);
xor U12670 (N_12670,N_12410,N_12102);
nand U12671 (N_12671,N_12228,N_12371);
xnor U12672 (N_12672,N_12022,N_12423);
and U12673 (N_12673,N_12240,N_12355);
and U12674 (N_12674,N_12389,N_12195);
and U12675 (N_12675,N_12124,N_12485);
or U12676 (N_12676,N_12098,N_12151);
xor U12677 (N_12677,N_12342,N_12063);
nor U12678 (N_12678,N_12235,N_12318);
xor U12679 (N_12679,N_12495,N_12315);
and U12680 (N_12680,N_12029,N_12215);
nor U12681 (N_12681,N_12092,N_12026);
or U12682 (N_12682,N_12378,N_12264);
nand U12683 (N_12683,N_12204,N_12164);
or U12684 (N_12684,N_12478,N_12259);
nor U12685 (N_12685,N_12112,N_12323);
nor U12686 (N_12686,N_12446,N_12358);
nand U12687 (N_12687,N_12190,N_12072);
nand U12688 (N_12688,N_12428,N_12299);
and U12689 (N_12689,N_12044,N_12425);
or U12690 (N_12690,N_12198,N_12058);
or U12691 (N_12691,N_12486,N_12070);
xor U12692 (N_12692,N_12421,N_12248);
nand U12693 (N_12693,N_12027,N_12091);
or U12694 (N_12694,N_12037,N_12165);
xor U12695 (N_12695,N_12280,N_12492);
or U12696 (N_12696,N_12096,N_12435);
nand U12697 (N_12697,N_12347,N_12229);
and U12698 (N_12698,N_12453,N_12257);
xor U12699 (N_12699,N_12081,N_12035);
nor U12700 (N_12700,N_12350,N_12219);
nor U12701 (N_12701,N_12300,N_12062);
or U12702 (N_12702,N_12482,N_12327);
or U12703 (N_12703,N_12128,N_12477);
xor U12704 (N_12704,N_12189,N_12348);
xor U12705 (N_12705,N_12353,N_12468);
xnor U12706 (N_12706,N_12041,N_12210);
and U12707 (N_12707,N_12185,N_12036);
nand U12708 (N_12708,N_12196,N_12244);
nand U12709 (N_12709,N_12012,N_12458);
nand U12710 (N_12710,N_12025,N_12207);
nor U12711 (N_12711,N_12001,N_12399);
nor U12712 (N_12712,N_12114,N_12087);
nand U12713 (N_12713,N_12121,N_12073);
nand U12714 (N_12714,N_12340,N_12186);
nor U12715 (N_12715,N_12144,N_12364);
xnor U12716 (N_12716,N_12234,N_12038);
nand U12717 (N_12717,N_12284,N_12394);
nor U12718 (N_12718,N_12480,N_12372);
nand U12719 (N_12719,N_12097,N_12148);
nor U12720 (N_12720,N_12408,N_12487);
xor U12721 (N_12721,N_12218,N_12188);
nor U12722 (N_12722,N_12126,N_12270);
xor U12723 (N_12723,N_12059,N_12253);
nor U12724 (N_12724,N_12146,N_12011);
xnor U12725 (N_12725,N_12439,N_12068);
and U12726 (N_12726,N_12099,N_12416);
and U12727 (N_12727,N_12420,N_12286);
nor U12728 (N_12728,N_12032,N_12489);
nor U12729 (N_12729,N_12180,N_12118);
xnor U12730 (N_12730,N_12158,N_12030);
and U12731 (N_12731,N_12174,N_12484);
nor U12732 (N_12732,N_12447,N_12053);
and U12733 (N_12733,N_12422,N_12307);
and U12734 (N_12734,N_12292,N_12459);
nand U12735 (N_12735,N_12249,N_12467);
nor U12736 (N_12736,N_12176,N_12288);
or U12737 (N_12737,N_12312,N_12232);
xor U12738 (N_12738,N_12110,N_12077);
nor U12739 (N_12739,N_12400,N_12064);
or U12740 (N_12740,N_12017,N_12018);
xor U12741 (N_12741,N_12256,N_12457);
nor U12742 (N_12742,N_12163,N_12442);
xor U12743 (N_12743,N_12125,N_12337);
and U12744 (N_12744,N_12269,N_12319);
nor U12745 (N_12745,N_12039,N_12003);
nand U12746 (N_12746,N_12217,N_12021);
or U12747 (N_12747,N_12047,N_12384);
xor U12748 (N_12748,N_12162,N_12179);
and U12749 (N_12749,N_12405,N_12150);
or U12750 (N_12750,N_12172,N_12215);
nand U12751 (N_12751,N_12368,N_12396);
xnor U12752 (N_12752,N_12009,N_12032);
nand U12753 (N_12753,N_12345,N_12314);
xor U12754 (N_12754,N_12175,N_12396);
and U12755 (N_12755,N_12470,N_12486);
nor U12756 (N_12756,N_12073,N_12189);
and U12757 (N_12757,N_12315,N_12293);
nor U12758 (N_12758,N_12278,N_12333);
nor U12759 (N_12759,N_12176,N_12436);
nand U12760 (N_12760,N_12299,N_12461);
nand U12761 (N_12761,N_12142,N_12269);
or U12762 (N_12762,N_12110,N_12146);
nand U12763 (N_12763,N_12442,N_12047);
nand U12764 (N_12764,N_12123,N_12356);
and U12765 (N_12765,N_12191,N_12100);
nand U12766 (N_12766,N_12049,N_12203);
nor U12767 (N_12767,N_12389,N_12224);
xnor U12768 (N_12768,N_12459,N_12332);
nor U12769 (N_12769,N_12386,N_12409);
nor U12770 (N_12770,N_12428,N_12350);
xnor U12771 (N_12771,N_12196,N_12093);
nand U12772 (N_12772,N_12097,N_12295);
xnor U12773 (N_12773,N_12266,N_12439);
and U12774 (N_12774,N_12469,N_12317);
nand U12775 (N_12775,N_12186,N_12245);
nor U12776 (N_12776,N_12218,N_12084);
nand U12777 (N_12777,N_12094,N_12344);
nand U12778 (N_12778,N_12134,N_12036);
and U12779 (N_12779,N_12030,N_12129);
xnor U12780 (N_12780,N_12358,N_12027);
or U12781 (N_12781,N_12133,N_12007);
or U12782 (N_12782,N_12485,N_12431);
xnor U12783 (N_12783,N_12352,N_12248);
nand U12784 (N_12784,N_12020,N_12056);
or U12785 (N_12785,N_12385,N_12081);
nor U12786 (N_12786,N_12102,N_12119);
and U12787 (N_12787,N_12088,N_12431);
xor U12788 (N_12788,N_12117,N_12199);
nor U12789 (N_12789,N_12178,N_12376);
nand U12790 (N_12790,N_12427,N_12319);
nand U12791 (N_12791,N_12212,N_12169);
nand U12792 (N_12792,N_12145,N_12148);
nor U12793 (N_12793,N_12329,N_12228);
nand U12794 (N_12794,N_12254,N_12042);
and U12795 (N_12795,N_12444,N_12165);
nand U12796 (N_12796,N_12423,N_12330);
nor U12797 (N_12797,N_12127,N_12197);
nor U12798 (N_12798,N_12222,N_12021);
and U12799 (N_12799,N_12056,N_12009);
and U12800 (N_12800,N_12134,N_12319);
and U12801 (N_12801,N_12155,N_12499);
and U12802 (N_12802,N_12305,N_12276);
xnor U12803 (N_12803,N_12065,N_12404);
xor U12804 (N_12804,N_12272,N_12209);
nand U12805 (N_12805,N_12133,N_12252);
xnor U12806 (N_12806,N_12420,N_12481);
and U12807 (N_12807,N_12355,N_12237);
or U12808 (N_12808,N_12081,N_12291);
or U12809 (N_12809,N_12378,N_12494);
and U12810 (N_12810,N_12249,N_12033);
or U12811 (N_12811,N_12135,N_12353);
nor U12812 (N_12812,N_12162,N_12381);
nor U12813 (N_12813,N_12395,N_12308);
or U12814 (N_12814,N_12131,N_12236);
xnor U12815 (N_12815,N_12164,N_12399);
nor U12816 (N_12816,N_12219,N_12077);
nor U12817 (N_12817,N_12020,N_12232);
xnor U12818 (N_12818,N_12222,N_12168);
or U12819 (N_12819,N_12096,N_12341);
xor U12820 (N_12820,N_12028,N_12372);
and U12821 (N_12821,N_12433,N_12281);
or U12822 (N_12822,N_12298,N_12122);
nand U12823 (N_12823,N_12301,N_12446);
nand U12824 (N_12824,N_12131,N_12167);
or U12825 (N_12825,N_12162,N_12425);
or U12826 (N_12826,N_12492,N_12122);
xor U12827 (N_12827,N_12434,N_12028);
nand U12828 (N_12828,N_12111,N_12052);
or U12829 (N_12829,N_12212,N_12133);
or U12830 (N_12830,N_12413,N_12393);
xor U12831 (N_12831,N_12378,N_12119);
nor U12832 (N_12832,N_12326,N_12439);
nor U12833 (N_12833,N_12292,N_12472);
or U12834 (N_12834,N_12166,N_12234);
xor U12835 (N_12835,N_12487,N_12373);
nor U12836 (N_12836,N_12417,N_12071);
xnor U12837 (N_12837,N_12339,N_12245);
xnor U12838 (N_12838,N_12101,N_12192);
nor U12839 (N_12839,N_12179,N_12114);
nand U12840 (N_12840,N_12470,N_12087);
or U12841 (N_12841,N_12174,N_12300);
nor U12842 (N_12842,N_12110,N_12182);
nand U12843 (N_12843,N_12184,N_12164);
nor U12844 (N_12844,N_12243,N_12357);
or U12845 (N_12845,N_12164,N_12394);
and U12846 (N_12846,N_12489,N_12279);
nand U12847 (N_12847,N_12358,N_12468);
and U12848 (N_12848,N_12461,N_12309);
xor U12849 (N_12849,N_12458,N_12348);
xor U12850 (N_12850,N_12014,N_12417);
xnor U12851 (N_12851,N_12077,N_12056);
xnor U12852 (N_12852,N_12157,N_12306);
nand U12853 (N_12853,N_12179,N_12489);
or U12854 (N_12854,N_12246,N_12250);
xnor U12855 (N_12855,N_12203,N_12149);
and U12856 (N_12856,N_12257,N_12305);
xnor U12857 (N_12857,N_12076,N_12455);
or U12858 (N_12858,N_12381,N_12404);
nor U12859 (N_12859,N_12391,N_12019);
nand U12860 (N_12860,N_12472,N_12064);
nand U12861 (N_12861,N_12055,N_12218);
nor U12862 (N_12862,N_12009,N_12489);
nand U12863 (N_12863,N_12127,N_12409);
and U12864 (N_12864,N_12391,N_12164);
and U12865 (N_12865,N_12371,N_12411);
nand U12866 (N_12866,N_12378,N_12099);
nand U12867 (N_12867,N_12139,N_12045);
or U12868 (N_12868,N_12408,N_12105);
and U12869 (N_12869,N_12050,N_12064);
xor U12870 (N_12870,N_12426,N_12302);
xnor U12871 (N_12871,N_12204,N_12251);
xor U12872 (N_12872,N_12200,N_12115);
and U12873 (N_12873,N_12344,N_12494);
xor U12874 (N_12874,N_12409,N_12418);
xor U12875 (N_12875,N_12286,N_12404);
and U12876 (N_12876,N_12338,N_12267);
and U12877 (N_12877,N_12016,N_12041);
nand U12878 (N_12878,N_12425,N_12458);
and U12879 (N_12879,N_12209,N_12243);
or U12880 (N_12880,N_12241,N_12396);
nand U12881 (N_12881,N_12388,N_12246);
xor U12882 (N_12882,N_12099,N_12496);
xnor U12883 (N_12883,N_12412,N_12293);
nand U12884 (N_12884,N_12464,N_12413);
and U12885 (N_12885,N_12289,N_12019);
or U12886 (N_12886,N_12132,N_12018);
and U12887 (N_12887,N_12297,N_12445);
nand U12888 (N_12888,N_12269,N_12099);
nand U12889 (N_12889,N_12175,N_12049);
nand U12890 (N_12890,N_12383,N_12411);
nand U12891 (N_12891,N_12078,N_12201);
and U12892 (N_12892,N_12226,N_12357);
nand U12893 (N_12893,N_12299,N_12080);
nor U12894 (N_12894,N_12162,N_12401);
and U12895 (N_12895,N_12046,N_12430);
nand U12896 (N_12896,N_12468,N_12458);
and U12897 (N_12897,N_12298,N_12074);
nand U12898 (N_12898,N_12224,N_12414);
nor U12899 (N_12899,N_12349,N_12037);
nand U12900 (N_12900,N_12424,N_12333);
nand U12901 (N_12901,N_12362,N_12313);
xnor U12902 (N_12902,N_12313,N_12422);
or U12903 (N_12903,N_12255,N_12003);
nor U12904 (N_12904,N_12475,N_12094);
xor U12905 (N_12905,N_12300,N_12490);
or U12906 (N_12906,N_12391,N_12485);
or U12907 (N_12907,N_12276,N_12108);
nand U12908 (N_12908,N_12069,N_12301);
and U12909 (N_12909,N_12299,N_12161);
nand U12910 (N_12910,N_12044,N_12310);
nand U12911 (N_12911,N_12037,N_12312);
and U12912 (N_12912,N_12450,N_12436);
xnor U12913 (N_12913,N_12355,N_12321);
nand U12914 (N_12914,N_12198,N_12229);
and U12915 (N_12915,N_12212,N_12225);
nor U12916 (N_12916,N_12375,N_12141);
nand U12917 (N_12917,N_12263,N_12226);
nand U12918 (N_12918,N_12227,N_12087);
or U12919 (N_12919,N_12319,N_12116);
and U12920 (N_12920,N_12428,N_12260);
nand U12921 (N_12921,N_12079,N_12084);
xnor U12922 (N_12922,N_12117,N_12029);
xor U12923 (N_12923,N_12370,N_12448);
nand U12924 (N_12924,N_12352,N_12202);
or U12925 (N_12925,N_12055,N_12115);
xor U12926 (N_12926,N_12243,N_12005);
nand U12927 (N_12927,N_12166,N_12236);
nor U12928 (N_12928,N_12035,N_12087);
nand U12929 (N_12929,N_12135,N_12093);
and U12930 (N_12930,N_12039,N_12392);
xnor U12931 (N_12931,N_12137,N_12118);
nand U12932 (N_12932,N_12164,N_12332);
nor U12933 (N_12933,N_12104,N_12497);
or U12934 (N_12934,N_12254,N_12194);
nor U12935 (N_12935,N_12171,N_12127);
nand U12936 (N_12936,N_12360,N_12287);
xor U12937 (N_12937,N_12369,N_12243);
nor U12938 (N_12938,N_12419,N_12335);
or U12939 (N_12939,N_12224,N_12259);
nand U12940 (N_12940,N_12264,N_12381);
xnor U12941 (N_12941,N_12394,N_12486);
or U12942 (N_12942,N_12111,N_12339);
nor U12943 (N_12943,N_12379,N_12011);
nand U12944 (N_12944,N_12378,N_12292);
nand U12945 (N_12945,N_12182,N_12307);
and U12946 (N_12946,N_12172,N_12047);
nor U12947 (N_12947,N_12181,N_12020);
or U12948 (N_12948,N_12175,N_12061);
nor U12949 (N_12949,N_12083,N_12250);
nand U12950 (N_12950,N_12138,N_12421);
or U12951 (N_12951,N_12049,N_12427);
and U12952 (N_12952,N_12441,N_12052);
nand U12953 (N_12953,N_12099,N_12022);
and U12954 (N_12954,N_12123,N_12000);
nor U12955 (N_12955,N_12424,N_12011);
or U12956 (N_12956,N_12262,N_12396);
nor U12957 (N_12957,N_12416,N_12227);
and U12958 (N_12958,N_12390,N_12088);
and U12959 (N_12959,N_12153,N_12074);
and U12960 (N_12960,N_12237,N_12111);
and U12961 (N_12961,N_12239,N_12300);
or U12962 (N_12962,N_12048,N_12294);
nor U12963 (N_12963,N_12300,N_12233);
nor U12964 (N_12964,N_12434,N_12100);
xnor U12965 (N_12965,N_12154,N_12360);
nand U12966 (N_12966,N_12338,N_12176);
nor U12967 (N_12967,N_12429,N_12150);
or U12968 (N_12968,N_12429,N_12048);
and U12969 (N_12969,N_12195,N_12452);
nor U12970 (N_12970,N_12153,N_12290);
nor U12971 (N_12971,N_12336,N_12117);
or U12972 (N_12972,N_12376,N_12352);
or U12973 (N_12973,N_12077,N_12407);
nand U12974 (N_12974,N_12437,N_12012);
or U12975 (N_12975,N_12296,N_12398);
nor U12976 (N_12976,N_12438,N_12216);
xnor U12977 (N_12977,N_12160,N_12330);
nor U12978 (N_12978,N_12354,N_12020);
or U12979 (N_12979,N_12158,N_12324);
nor U12980 (N_12980,N_12201,N_12120);
nand U12981 (N_12981,N_12041,N_12293);
nand U12982 (N_12982,N_12036,N_12076);
nor U12983 (N_12983,N_12399,N_12284);
and U12984 (N_12984,N_12337,N_12256);
nand U12985 (N_12985,N_12303,N_12464);
nand U12986 (N_12986,N_12435,N_12084);
and U12987 (N_12987,N_12367,N_12192);
nor U12988 (N_12988,N_12462,N_12342);
nand U12989 (N_12989,N_12312,N_12151);
xor U12990 (N_12990,N_12414,N_12170);
or U12991 (N_12991,N_12255,N_12445);
nor U12992 (N_12992,N_12409,N_12304);
and U12993 (N_12993,N_12019,N_12477);
nand U12994 (N_12994,N_12327,N_12065);
nor U12995 (N_12995,N_12477,N_12461);
xnor U12996 (N_12996,N_12026,N_12446);
xor U12997 (N_12997,N_12232,N_12098);
xor U12998 (N_12998,N_12004,N_12037);
or U12999 (N_12999,N_12104,N_12177);
and U13000 (N_13000,N_12676,N_12819);
xor U13001 (N_13001,N_12791,N_12995);
and U13002 (N_13002,N_12903,N_12952);
nand U13003 (N_13003,N_12810,N_12682);
nor U13004 (N_13004,N_12636,N_12932);
or U13005 (N_13005,N_12550,N_12823);
nor U13006 (N_13006,N_12941,N_12647);
nand U13007 (N_13007,N_12712,N_12699);
or U13008 (N_13008,N_12537,N_12643);
nor U13009 (N_13009,N_12911,N_12763);
xnor U13010 (N_13010,N_12985,N_12630);
and U13011 (N_13011,N_12695,N_12739);
or U13012 (N_13012,N_12981,N_12502);
and U13013 (N_13013,N_12626,N_12526);
and U13014 (N_13014,N_12917,N_12725);
or U13015 (N_13015,N_12849,N_12965);
and U13016 (N_13016,N_12582,N_12736);
and U13017 (N_13017,N_12871,N_12990);
or U13018 (N_13018,N_12873,N_12807);
xor U13019 (N_13019,N_12846,N_12548);
nand U13020 (N_13020,N_12616,N_12805);
nand U13021 (N_13021,N_12622,N_12832);
nor U13022 (N_13022,N_12910,N_12907);
xor U13023 (N_13023,N_12749,N_12930);
nand U13024 (N_13024,N_12727,N_12589);
nand U13025 (N_13025,N_12700,N_12926);
nand U13026 (N_13026,N_12912,N_12564);
xor U13027 (N_13027,N_12578,N_12742);
xor U13028 (N_13028,N_12728,N_12982);
or U13029 (N_13029,N_12558,N_12637);
nand U13030 (N_13030,N_12579,N_12828);
or U13031 (N_13031,N_12664,N_12519);
nor U13032 (N_13032,N_12938,N_12714);
and U13033 (N_13033,N_12734,N_12674);
nand U13034 (N_13034,N_12580,N_12959);
nand U13035 (N_13035,N_12600,N_12920);
and U13036 (N_13036,N_12639,N_12669);
nand U13037 (N_13037,N_12598,N_12603);
xor U13038 (N_13038,N_12748,N_12943);
or U13039 (N_13039,N_12833,N_12806);
xor U13040 (N_13040,N_12830,N_12535);
nor U13041 (N_13041,N_12989,N_12936);
xor U13042 (N_13042,N_12562,N_12593);
or U13043 (N_13043,N_12760,N_12796);
nand U13044 (N_13044,N_12500,N_12601);
or U13045 (N_13045,N_12688,N_12853);
xnor U13046 (N_13046,N_12949,N_12542);
and U13047 (N_13047,N_12776,N_12680);
nand U13048 (N_13048,N_12961,N_12569);
xnor U13049 (N_13049,N_12988,N_12673);
and U13050 (N_13050,N_12753,N_12511);
or U13051 (N_13051,N_12716,N_12528);
xnor U13052 (N_13052,N_12854,N_12824);
nor U13053 (N_13053,N_12861,N_12757);
xor U13054 (N_13054,N_12867,N_12623);
or U13055 (N_13055,N_12713,N_12890);
nand U13056 (N_13056,N_12545,N_12918);
nor U13057 (N_13057,N_12774,N_12969);
nand U13058 (N_13058,N_12521,N_12826);
or U13059 (N_13059,N_12976,N_12784);
nor U13060 (N_13060,N_12592,N_12966);
or U13061 (N_13061,N_12991,N_12983);
nand U13062 (N_13062,N_12841,N_12798);
xor U13063 (N_13063,N_12654,N_12914);
and U13064 (N_13064,N_12565,N_12708);
or U13065 (N_13065,N_12690,N_12684);
or U13066 (N_13066,N_12797,N_12892);
nor U13067 (N_13067,N_12642,N_12655);
and U13068 (N_13068,N_12978,N_12888);
or U13069 (N_13069,N_12720,N_12756);
xnor U13070 (N_13070,N_12663,N_12968);
or U13071 (N_13071,N_12813,N_12615);
nor U13072 (N_13072,N_12971,N_12617);
and U13073 (N_13073,N_12686,N_12808);
nand U13074 (N_13074,N_12577,N_12772);
xor U13075 (N_13075,N_12501,N_12886);
and U13076 (N_13076,N_12771,N_12998);
or U13077 (N_13077,N_12964,N_12814);
and U13078 (N_13078,N_12729,N_12840);
and U13079 (N_13079,N_12583,N_12707);
nor U13080 (N_13080,N_12765,N_12928);
xor U13081 (N_13081,N_12590,N_12546);
nor U13082 (N_13082,N_12747,N_12946);
xor U13083 (N_13083,N_12834,N_12818);
xnor U13084 (N_13084,N_12549,N_12882);
xor U13085 (N_13085,N_12665,N_12925);
nor U13086 (N_13086,N_12942,N_12605);
xor U13087 (N_13087,N_12934,N_12775);
and U13088 (N_13088,N_12524,N_12793);
nand U13089 (N_13089,N_12588,N_12611);
and U13090 (N_13090,N_12702,N_12878);
and U13091 (N_13091,N_12859,N_12954);
and U13092 (N_13092,N_12870,N_12721);
nand U13093 (N_13093,N_12513,N_12741);
and U13094 (N_13094,N_12717,N_12514);
xor U13095 (N_13095,N_12825,N_12602);
or U13096 (N_13096,N_12781,N_12661);
and U13097 (N_13097,N_12656,N_12566);
or U13098 (N_13098,N_12779,N_12599);
or U13099 (N_13099,N_12731,N_12575);
or U13100 (N_13100,N_12993,N_12881);
nor U13101 (N_13101,N_12539,N_12848);
and U13102 (N_13102,N_12745,N_12851);
nor U13103 (N_13103,N_12693,N_12666);
and U13104 (N_13104,N_12510,N_12672);
or U13105 (N_13105,N_12916,N_12758);
or U13106 (N_13106,N_12692,N_12940);
nand U13107 (N_13107,N_12865,N_12856);
nand U13108 (N_13108,N_12591,N_12785);
or U13109 (N_13109,N_12735,N_12863);
nand U13110 (N_13110,N_12746,N_12752);
and U13111 (N_13111,N_12627,N_12544);
xnor U13112 (N_13112,N_12653,N_12522);
xnor U13113 (N_13113,N_12670,N_12975);
nand U13114 (N_13114,N_12897,N_12921);
xor U13115 (N_13115,N_12773,N_12711);
or U13116 (N_13116,N_12860,N_12937);
nand U13117 (N_13117,N_12651,N_12766);
or U13118 (N_13118,N_12883,N_12821);
nand U13119 (N_13119,N_12827,N_12704);
nand U13120 (N_13120,N_12913,N_12970);
nor U13121 (N_13121,N_12650,N_12850);
nor U13122 (N_13122,N_12527,N_12900);
nand U13123 (N_13123,N_12847,N_12780);
xor U13124 (N_13124,N_12668,N_12646);
or U13125 (N_13125,N_12584,N_12563);
or U13126 (N_13126,N_12518,N_12640);
nor U13127 (N_13127,N_12905,N_12761);
nand U13128 (N_13128,N_12610,N_12788);
or U13129 (N_13129,N_12515,N_12869);
and U13130 (N_13130,N_12750,N_12629);
or U13131 (N_13131,N_12922,N_12703);
nor U13132 (N_13132,N_12614,N_12939);
or U13133 (N_13133,N_12767,N_12606);
xor U13134 (N_13134,N_12530,N_12738);
or U13135 (N_13135,N_12715,N_12898);
nand U13136 (N_13136,N_12845,N_12719);
nand U13137 (N_13137,N_12956,N_12868);
xor U13138 (N_13138,N_12657,N_12974);
xnor U13139 (N_13139,N_12768,N_12722);
or U13140 (N_13140,N_12523,N_12587);
or U13141 (N_13141,N_12586,N_12829);
nand U13142 (N_13142,N_12662,N_12759);
nor U13143 (N_13143,N_12876,N_12660);
xnor U13144 (N_13144,N_12594,N_12507);
nor U13145 (N_13145,N_12958,N_12885);
nand U13146 (N_13146,N_12604,N_12659);
and U13147 (N_13147,N_12732,N_12877);
xor U13148 (N_13148,N_12685,N_12538);
and U13149 (N_13149,N_12531,N_12764);
and U13150 (N_13150,N_12508,N_12996);
xnor U13151 (N_13151,N_12551,N_12979);
xnor U13152 (N_13152,N_12994,N_12635);
xnor U13153 (N_13153,N_12677,N_12815);
and U13154 (N_13154,N_12955,N_12908);
nor U13155 (N_13155,N_12572,N_12794);
xnor U13156 (N_13156,N_12787,N_12967);
nand U13157 (N_13157,N_12557,N_12778);
and U13158 (N_13158,N_12573,N_12632);
nor U13159 (N_13159,N_12864,N_12977);
nor U13160 (N_13160,N_12953,N_12570);
or U13161 (N_13161,N_12884,N_12691);
nor U13162 (N_13162,N_12540,N_12552);
nand U13163 (N_13163,N_12709,N_12844);
nand U13164 (N_13164,N_12574,N_12973);
and U13165 (N_13165,N_12895,N_12838);
nor U13166 (N_13166,N_12723,N_12596);
xor U13167 (N_13167,N_12987,N_12638);
xnor U13168 (N_13168,N_12901,N_12944);
nor U13169 (N_13169,N_12517,N_12618);
xor U13170 (N_13170,N_12836,N_12858);
xnor U13171 (N_13171,N_12678,N_12634);
xnor U13172 (N_13172,N_12963,N_12957);
nor U13173 (N_13173,N_12619,N_12960);
and U13174 (N_13174,N_12505,N_12751);
nor U13175 (N_13175,N_12857,N_12649);
and U13176 (N_13176,N_12997,N_12804);
or U13177 (N_13177,N_12929,N_12795);
nand U13178 (N_13178,N_12512,N_12831);
nand U13179 (N_13179,N_12769,N_12816);
nand U13180 (N_13180,N_12822,N_12644);
or U13181 (N_13181,N_12950,N_12803);
or U13182 (N_13182,N_12705,N_12710);
or U13183 (N_13183,N_12694,N_12697);
or U13184 (N_13184,N_12835,N_12924);
and U13185 (N_13185,N_12648,N_12812);
or U13186 (N_13186,N_12645,N_12624);
xor U13187 (N_13187,N_12631,N_12561);
xor U13188 (N_13188,N_12874,N_12899);
and U13189 (N_13189,N_12887,N_12609);
nor U13190 (N_13190,N_12532,N_12935);
and U13191 (N_13191,N_12658,N_12571);
nand U13192 (N_13192,N_12872,N_12945);
xnor U13193 (N_13193,N_12567,N_12792);
nand U13194 (N_13194,N_12679,N_12701);
and U13195 (N_13195,N_12724,N_12984);
or U13196 (N_13196,N_12799,N_12733);
nand U13197 (N_13197,N_12681,N_12726);
and U13198 (N_13198,N_12547,N_12754);
or U13199 (N_13199,N_12506,N_12948);
nand U13200 (N_13200,N_12811,N_12896);
nor U13201 (N_13201,N_12947,N_12889);
xor U13202 (N_13202,N_12559,N_12919);
nor U13203 (N_13203,N_12992,N_12875);
and U13204 (N_13204,N_12525,N_12891);
xor U13205 (N_13205,N_12743,N_12689);
nor U13206 (N_13206,N_12744,N_12633);
or U13207 (N_13207,N_12842,N_12931);
and U13208 (N_13208,N_12696,N_12855);
nand U13209 (N_13209,N_12843,N_12675);
nand U13210 (N_13210,N_12613,N_12698);
nor U13211 (N_13211,N_12556,N_12641);
nor U13212 (N_13212,N_12554,N_12608);
nand U13213 (N_13213,N_12628,N_12607);
or U13214 (N_13214,N_12516,N_12906);
or U13215 (N_13215,N_12621,N_12909);
xnor U13216 (N_13216,N_12800,N_12962);
nor U13217 (N_13217,N_12927,N_12576);
and U13218 (N_13218,N_12801,N_12687);
nor U13219 (N_13219,N_12762,N_12568);
and U13220 (N_13220,N_12770,N_12652);
and U13221 (N_13221,N_12625,N_12520);
nand U13222 (N_13222,N_12543,N_12999);
nor U13223 (N_13223,N_12783,N_12730);
xor U13224 (N_13224,N_12980,N_12820);
and U13225 (N_13225,N_12755,N_12683);
nand U13226 (N_13226,N_12972,N_12933);
xor U13227 (N_13227,N_12504,N_12560);
or U13228 (N_13228,N_12737,N_12866);
nor U13229 (N_13229,N_12789,N_12553);
and U13230 (N_13230,N_12718,N_12503);
and U13231 (N_13231,N_12536,N_12585);
and U13232 (N_13232,N_12777,N_12620);
nand U13233 (N_13233,N_12817,N_12534);
nand U13234 (N_13234,N_12902,N_12862);
and U13235 (N_13235,N_12893,N_12740);
or U13236 (N_13236,N_12671,N_12782);
and U13237 (N_13237,N_12852,N_12880);
xor U13238 (N_13238,N_12951,N_12555);
nor U13239 (N_13239,N_12529,N_12581);
xor U13240 (N_13240,N_12894,N_12533);
nand U13241 (N_13241,N_12923,N_12904);
nor U13242 (N_13242,N_12597,N_12790);
nand U13243 (N_13243,N_12667,N_12786);
nor U13244 (N_13244,N_12509,N_12802);
nand U13245 (N_13245,N_12986,N_12595);
and U13246 (N_13246,N_12612,N_12837);
nor U13247 (N_13247,N_12541,N_12809);
or U13248 (N_13248,N_12706,N_12839);
and U13249 (N_13249,N_12879,N_12915);
xnor U13250 (N_13250,N_12798,N_12863);
nor U13251 (N_13251,N_12741,N_12758);
nor U13252 (N_13252,N_12620,N_12854);
or U13253 (N_13253,N_12630,N_12999);
and U13254 (N_13254,N_12797,N_12550);
nor U13255 (N_13255,N_12782,N_12879);
xnor U13256 (N_13256,N_12990,N_12873);
nand U13257 (N_13257,N_12992,N_12823);
or U13258 (N_13258,N_12747,N_12995);
nand U13259 (N_13259,N_12702,N_12720);
and U13260 (N_13260,N_12776,N_12758);
nor U13261 (N_13261,N_12956,N_12660);
or U13262 (N_13262,N_12678,N_12872);
nand U13263 (N_13263,N_12529,N_12761);
or U13264 (N_13264,N_12779,N_12839);
xnor U13265 (N_13265,N_12987,N_12677);
or U13266 (N_13266,N_12804,N_12555);
and U13267 (N_13267,N_12781,N_12656);
nand U13268 (N_13268,N_12527,N_12971);
xnor U13269 (N_13269,N_12675,N_12570);
nand U13270 (N_13270,N_12897,N_12890);
or U13271 (N_13271,N_12717,N_12730);
xnor U13272 (N_13272,N_12961,N_12699);
or U13273 (N_13273,N_12506,N_12757);
and U13274 (N_13274,N_12639,N_12713);
or U13275 (N_13275,N_12638,N_12583);
nand U13276 (N_13276,N_12664,N_12693);
or U13277 (N_13277,N_12925,N_12544);
or U13278 (N_13278,N_12817,N_12566);
nand U13279 (N_13279,N_12570,N_12907);
and U13280 (N_13280,N_12780,N_12906);
nand U13281 (N_13281,N_12951,N_12728);
nand U13282 (N_13282,N_12801,N_12808);
and U13283 (N_13283,N_12754,N_12582);
xor U13284 (N_13284,N_12544,N_12591);
or U13285 (N_13285,N_12693,N_12740);
xor U13286 (N_13286,N_12651,N_12588);
nor U13287 (N_13287,N_12605,N_12860);
nand U13288 (N_13288,N_12784,N_12967);
and U13289 (N_13289,N_12554,N_12908);
or U13290 (N_13290,N_12592,N_12962);
or U13291 (N_13291,N_12602,N_12848);
nor U13292 (N_13292,N_12654,N_12709);
xnor U13293 (N_13293,N_12803,N_12527);
xnor U13294 (N_13294,N_12800,N_12820);
or U13295 (N_13295,N_12508,N_12928);
and U13296 (N_13296,N_12780,N_12675);
or U13297 (N_13297,N_12914,N_12962);
or U13298 (N_13298,N_12711,N_12687);
nand U13299 (N_13299,N_12850,N_12777);
xnor U13300 (N_13300,N_12999,N_12576);
xnor U13301 (N_13301,N_12631,N_12757);
or U13302 (N_13302,N_12519,N_12927);
xor U13303 (N_13303,N_12788,N_12903);
and U13304 (N_13304,N_12889,N_12886);
or U13305 (N_13305,N_12858,N_12636);
or U13306 (N_13306,N_12936,N_12973);
or U13307 (N_13307,N_12870,N_12689);
nand U13308 (N_13308,N_12740,N_12501);
xor U13309 (N_13309,N_12966,N_12894);
nor U13310 (N_13310,N_12840,N_12796);
xnor U13311 (N_13311,N_12861,N_12877);
nand U13312 (N_13312,N_12772,N_12823);
or U13313 (N_13313,N_12921,N_12765);
xnor U13314 (N_13314,N_12717,N_12640);
and U13315 (N_13315,N_12634,N_12648);
xnor U13316 (N_13316,N_12636,N_12609);
nand U13317 (N_13317,N_12769,N_12675);
or U13318 (N_13318,N_12639,N_12696);
nand U13319 (N_13319,N_12896,N_12943);
and U13320 (N_13320,N_12979,N_12674);
xor U13321 (N_13321,N_12658,N_12925);
and U13322 (N_13322,N_12813,N_12952);
or U13323 (N_13323,N_12597,N_12552);
and U13324 (N_13324,N_12668,N_12994);
and U13325 (N_13325,N_12846,N_12667);
xor U13326 (N_13326,N_12656,N_12680);
nor U13327 (N_13327,N_12723,N_12982);
xor U13328 (N_13328,N_12661,N_12707);
nand U13329 (N_13329,N_12602,N_12542);
or U13330 (N_13330,N_12594,N_12833);
nand U13331 (N_13331,N_12817,N_12933);
xnor U13332 (N_13332,N_12781,N_12765);
xnor U13333 (N_13333,N_12765,N_12533);
or U13334 (N_13334,N_12900,N_12586);
nor U13335 (N_13335,N_12993,N_12763);
nor U13336 (N_13336,N_12791,N_12973);
or U13337 (N_13337,N_12747,N_12897);
xor U13338 (N_13338,N_12828,N_12922);
nand U13339 (N_13339,N_12966,N_12620);
and U13340 (N_13340,N_12646,N_12895);
xnor U13341 (N_13341,N_12752,N_12754);
nor U13342 (N_13342,N_12500,N_12901);
xnor U13343 (N_13343,N_12887,N_12844);
xnor U13344 (N_13344,N_12651,N_12519);
or U13345 (N_13345,N_12742,N_12798);
or U13346 (N_13346,N_12664,N_12770);
or U13347 (N_13347,N_12782,N_12806);
xnor U13348 (N_13348,N_12942,N_12668);
nand U13349 (N_13349,N_12814,N_12638);
nor U13350 (N_13350,N_12766,N_12549);
nand U13351 (N_13351,N_12628,N_12700);
or U13352 (N_13352,N_12778,N_12776);
nor U13353 (N_13353,N_12985,N_12589);
or U13354 (N_13354,N_12587,N_12994);
and U13355 (N_13355,N_12893,N_12814);
xnor U13356 (N_13356,N_12846,N_12943);
and U13357 (N_13357,N_12712,N_12858);
or U13358 (N_13358,N_12666,N_12875);
nor U13359 (N_13359,N_12518,N_12992);
nand U13360 (N_13360,N_12983,N_12924);
xor U13361 (N_13361,N_12701,N_12578);
or U13362 (N_13362,N_12621,N_12907);
nand U13363 (N_13363,N_12865,N_12658);
xor U13364 (N_13364,N_12936,N_12693);
and U13365 (N_13365,N_12585,N_12719);
and U13366 (N_13366,N_12623,N_12725);
or U13367 (N_13367,N_12796,N_12815);
and U13368 (N_13368,N_12551,N_12735);
nand U13369 (N_13369,N_12596,N_12628);
xor U13370 (N_13370,N_12708,N_12769);
nor U13371 (N_13371,N_12610,N_12676);
xor U13372 (N_13372,N_12519,N_12734);
xnor U13373 (N_13373,N_12799,N_12604);
xor U13374 (N_13374,N_12797,N_12595);
xor U13375 (N_13375,N_12605,N_12596);
nand U13376 (N_13376,N_12584,N_12847);
nand U13377 (N_13377,N_12787,N_12706);
xor U13378 (N_13378,N_12655,N_12563);
nand U13379 (N_13379,N_12750,N_12930);
xor U13380 (N_13380,N_12907,N_12842);
nor U13381 (N_13381,N_12833,N_12990);
xor U13382 (N_13382,N_12910,N_12942);
or U13383 (N_13383,N_12535,N_12665);
xor U13384 (N_13384,N_12937,N_12820);
xor U13385 (N_13385,N_12924,N_12772);
xor U13386 (N_13386,N_12661,N_12566);
and U13387 (N_13387,N_12500,N_12973);
nor U13388 (N_13388,N_12637,N_12582);
nand U13389 (N_13389,N_12939,N_12803);
nand U13390 (N_13390,N_12854,N_12708);
or U13391 (N_13391,N_12859,N_12812);
xor U13392 (N_13392,N_12717,N_12851);
xor U13393 (N_13393,N_12503,N_12635);
nor U13394 (N_13394,N_12897,N_12693);
nor U13395 (N_13395,N_12892,N_12868);
and U13396 (N_13396,N_12841,N_12912);
nor U13397 (N_13397,N_12957,N_12563);
and U13398 (N_13398,N_12734,N_12706);
xor U13399 (N_13399,N_12698,N_12681);
nand U13400 (N_13400,N_12631,N_12733);
xor U13401 (N_13401,N_12833,N_12649);
nor U13402 (N_13402,N_12518,N_12547);
xor U13403 (N_13403,N_12798,N_12932);
xnor U13404 (N_13404,N_12706,N_12783);
nand U13405 (N_13405,N_12553,N_12809);
and U13406 (N_13406,N_12905,N_12614);
xor U13407 (N_13407,N_12950,N_12891);
nand U13408 (N_13408,N_12822,N_12987);
xnor U13409 (N_13409,N_12822,N_12899);
nor U13410 (N_13410,N_12697,N_12625);
and U13411 (N_13411,N_12856,N_12556);
xor U13412 (N_13412,N_12817,N_12582);
nand U13413 (N_13413,N_12806,N_12842);
nor U13414 (N_13414,N_12679,N_12939);
nor U13415 (N_13415,N_12586,N_12612);
nor U13416 (N_13416,N_12585,N_12881);
xor U13417 (N_13417,N_12994,N_12921);
nor U13418 (N_13418,N_12696,N_12815);
xor U13419 (N_13419,N_12876,N_12786);
nand U13420 (N_13420,N_12782,N_12812);
nand U13421 (N_13421,N_12572,N_12955);
xor U13422 (N_13422,N_12922,N_12931);
nand U13423 (N_13423,N_12732,N_12665);
xor U13424 (N_13424,N_12650,N_12686);
xor U13425 (N_13425,N_12747,N_12796);
nand U13426 (N_13426,N_12925,N_12908);
nor U13427 (N_13427,N_12693,N_12582);
nor U13428 (N_13428,N_12542,N_12856);
xnor U13429 (N_13429,N_12865,N_12681);
nand U13430 (N_13430,N_12553,N_12965);
xor U13431 (N_13431,N_12671,N_12588);
nand U13432 (N_13432,N_12520,N_12933);
nand U13433 (N_13433,N_12966,N_12977);
or U13434 (N_13434,N_12880,N_12922);
nand U13435 (N_13435,N_12817,N_12576);
nand U13436 (N_13436,N_12685,N_12771);
nand U13437 (N_13437,N_12933,N_12924);
and U13438 (N_13438,N_12564,N_12656);
xnor U13439 (N_13439,N_12528,N_12848);
and U13440 (N_13440,N_12982,N_12576);
nand U13441 (N_13441,N_12517,N_12823);
nand U13442 (N_13442,N_12984,N_12614);
nor U13443 (N_13443,N_12630,N_12746);
and U13444 (N_13444,N_12634,N_12868);
nor U13445 (N_13445,N_12947,N_12852);
and U13446 (N_13446,N_12905,N_12810);
nand U13447 (N_13447,N_12742,N_12991);
or U13448 (N_13448,N_12833,N_12702);
xor U13449 (N_13449,N_12730,N_12955);
xnor U13450 (N_13450,N_12512,N_12649);
xor U13451 (N_13451,N_12938,N_12776);
nor U13452 (N_13452,N_12536,N_12532);
nor U13453 (N_13453,N_12741,N_12744);
nor U13454 (N_13454,N_12616,N_12566);
or U13455 (N_13455,N_12926,N_12714);
and U13456 (N_13456,N_12856,N_12681);
nand U13457 (N_13457,N_12855,N_12940);
nor U13458 (N_13458,N_12589,N_12720);
nor U13459 (N_13459,N_12638,N_12624);
xnor U13460 (N_13460,N_12869,N_12855);
and U13461 (N_13461,N_12771,N_12939);
xnor U13462 (N_13462,N_12712,N_12653);
nor U13463 (N_13463,N_12924,N_12711);
nand U13464 (N_13464,N_12711,N_12925);
and U13465 (N_13465,N_12800,N_12763);
or U13466 (N_13466,N_12979,N_12873);
and U13467 (N_13467,N_12689,N_12942);
nand U13468 (N_13468,N_12502,N_12722);
and U13469 (N_13469,N_12585,N_12992);
nand U13470 (N_13470,N_12560,N_12517);
and U13471 (N_13471,N_12726,N_12504);
nand U13472 (N_13472,N_12747,N_12556);
nand U13473 (N_13473,N_12733,N_12717);
and U13474 (N_13474,N_12964,N_12855);
nand U13475 (N_13475,N_12960,N_12875);
nor U13476 (N_13476,N_12851,N_12824);
or U13477 (N_13477,N_12728,N_12751);
xnor U13478 (N_13478,N_12835,N_12878);
xor U13479 (N_13479,N_12833,N_12750);
or U13480 (N_13480,N_12740,N_12698);
xor U13481 (N_13481,N_12847,N_12854);
or U13482 (N_13482,N_12934,N_12667);
nor U13483 (N_13483,N_12955,N_12585);
xnor U13484 (N_13484,N_12836,N_12738);
or U13485 (N_13485,N_12621,N_12615);
nand U13486 (N_13486,N_12773,N_12677);
nor U13487 (N_13487,N_12974,N_12613);
or U13488 (N_13488,N_12503,N_12984);
nand U13489 (N_13489,N_12619,N_12850);
nand U13490 (N_13490,N_12744,N_12917);
and U13491 (N_13491,N_12711,N_12796);
nand U13492 (N_13492,N_12777,N_12724);
and U13493 (N_13493,N_12952,N_12979);
or U13494 (N_13494,N_12824,N_12652);
and U13495 (N_13495,N_12734,N_12715);
and U13496 (N_13496,N_12727,N_12534);
nor U13497 (N_13497,N_12627,N_12859);
or U13498 (N_13498,N_12937,N_12934);
nor U13499 (N_13499,N_12948,N_12795);
nand U13500 (N_13500,N_13125,N_13399);
xor U13501 (N_13501,N_13247,N_13212);
nand U13502 (N_13502,N_13191,N_13470);
nor U13503 (N_13503,N_13136,N_13021);
nand U13504 (N_13504,N_13152,N_13079);
or U13505 (N_13505,N_13359,N_13165);
or U13506 (N_13506,N_13181,N_13211);
xor U13507 (N_13507,N_13286,N_13010);
xnor U13508 (N_13508,N_13440,N_13043);
or U13509 (N_13509,N_13083,N_13184);
nand U13510 (N_13510,N_13108,N_13192);
nor U13511 (N_13511,N_13333,N_13237);
nand U13512 (N_13512,N_13213,N_13065);
nor U13513 (N_13513,N_13318,N_13174);
nor U13514 (N_13514,N_13419,N_13248);
nand U13515 (N_13515,N_13293,N_13154);
nor U13516 (N_13516,N_13497,N_13232);
xor U13517 (N_13517,N_13004,N_13009);
and U13518 (N_13518,N_13073,N_13473);
and U13519 (N_13519,N_13077,N_13026);
and U13520 (N_13520,N_13364,N_13283);
and U13521 (N_13521,N_13234,N_13469);
nor U13522 (N_13522,N_13229,N_13412);
nor U13523 (N_13523,N_13365,N_13219);
nor U13524 (N_13524,N_13096,N_13240);
xnor U13525 (N_13525,N_13171,N_13268);
and U13526 (N_13526,N_13341,N_13005);
nand U13527 (N_13527,N_13046,N_13047);
nand U13528 (N_13528,N_13263,N_13486);
nor U13529 (N_13529,N_13475,N_13415);
nand U13530 (N_13530,N_13159,N_13297);
xor U13531 (N_13531,N_13015,N_13353);
xor U13532 (N_13532,N_13081,N_13124);
nand U13533 (N_13533,N_13210,N_13214);
or U13534 (N_13534,N_13215,N_13205);
nand U13535 (N_13535,N_13106,N_13157);
and U13536 (N_13536,N_13455,N_13145);
nand U13537 (N_13537,N_13200,N_13345);
or U13538 (N_13538,N_13149,N_13404);
nand U13539 (N_13539,N_13334,N_13233);
or U13540 (N_13540,N_13355,N_13000);
or U13541 (N_13541,N_13044,N_13326);
or U13542 (N_13542,N_13180,N_13075);
xor U13543 (N_13543,N_13064,N_13493);
nand U13544 (N_13544,N_13447,N_13376);
nor U13545 (N_13545,N_13410,N_13480);
and U13546 (N_13546,N_13097,N_13262);
and U13547 (N_13547,N_13186,N_13499);
nand U13548 (N_13548,N_13199,N_13389);
xnor U13549 (N_13549,N_13319,N_13269);
or U13550 (N_13550,N_13142,N_13235);
nor U13551 (N_13551,N_13320,N_13148);
nand U13552 (N_13552,N_13312,N_13386);
or U13553 (N_13553,N_13035,N_13209);
or U13554 (N_13554,N_13462,N_13130);
and U13555 (N_13555,N_13280,N_13490);
and U13556 (N_13556,N_13056,N_13363);
nand U13557 (N_13557,N_13167,N_13024);
nand U13558 (N_13558,N_13337,N_13303);
nor U13559 (N_13559,N_13201,N_13471);
xor U13560 (N_13560,N_13298,N_13059);
nor U13561 (N_13561,N_13251,N_13485);
xor U13562 (N_13562,N_13383,N_13344);
and U13563 (N_13563,N_13394,N_13284);
nand U13564 (N_13564,N_13018,N_13484);
and U13565 (N_13565,N_13300,N_13008);
nand U13566 (N_13566,N_13395,N_13071);
xnor U13567 (N_13567,N_13443,N_13113);
nor U13568 (N_13568,N_13495,N_13374);
nor U13569 (N_13569,N_13141,N_13116);
or U13570 (N_13570,N_13218,N_13427);
nor U13571 (N_13571,N_13012,N_13267);
xor U13572 (N_13572,N_13225,N_13105);
or U13573 (N_13573,N_13132,N_13203);
and U13574 (N_13574,N_13007,N_13090);
and U13575 (N_13575,N_13445,N_13330);
or U13576 (N_13576,N_13328,N_13366);
xnor U13577 (N_13577,N_13336,N_13481);
nand U13578 (N_13578,N_13153,N_13245);
or U13579 (N_13579,N_13060,N_13243);
nand U13580 (N_13580,N_13204,N_13439);
nor U13581 (N_13581,N_13417,N_13092);
and U13582 (N_13582,N_13146,N_13372);
and U13583 (N_13583,N_13407,N_13143);
nor U13584 (N_13584,N_13054,N_13265);
or U13585 (N_13585,N_13465,N_13476);
or U13586 (N_13586,N_13117,N_13095);
nor U13587 (N_13587,N_13401,N_13451);
nor U13588 (N_13588,N_13102,N_13450);
or U13589 (N_13589,N_13348,N_13321);
or U13590 (N_13590,N_13368,N_13101);
nand U13591 (N_13591,N_13464,N_13400);
nand U13592 (N_13592,N_13128,N_13466);
xor U13593 (N_13593,N_13398,N_13271);
and U13594 (N_13594,N_13038,N_13133);
and U13595 (N_13595,N_13195,N_13340);
or U13596 (N_13596,N_13375,N_13429);
nand U13597 (N_13597,N_13226,N_13223);
nand U13598 (N_13598,N_13067,N_13162);
xnor U13599 (N_13599,N_13331,N_13411);
nor U13600 (N_13600,N_13260,N_13080);
and U13601 (N_13601,N_13311,N_13379);
and U13602 (N_13602,N_13356,N_13001);
and U13603 (N_13603,N_13266,N_13158);
nand U13604 (N_13604,N_13063,N_13289);
nor U13605 (N_13605,N_13335,N_13068);
or U13606 (N_13606,N_13388,N_13206);
nor U13607 (N_13607,N_13076,N_13244);
nand U13608 (N_13608,N_13129,N_13396);
nor U13609 (N_13609,N_13140,N_13479);
or U13610 (N_13610,N_13371,N_13058);
nor U13611 (N_13611,N_13357,N_13168);
or U13612 (N_13612,N_13224,N_13277);
nand U13613 (N_13613,N_13420,N_13037);
and U13614 (N_13614,N_13042,N_13343);
nor U13615 (N_13615,N_13072,N_13188);
xnor U13616 (N_13616,N_13441,N_13323);
nor U13617 (N_13617,N_13342,N_13314);
nor U13618 (N_13618,N_13431,N_13296);
xor U13619 (N_13619,N_13254,N_13208);
and U13620 (N_13620,N_13488,N_13178);
xor U13621 (N_13621,N_13099,N_13091);
nand U13622 (N_13622,N_13002,N_13170);
or U13623 (N_13623,N_13310,N_13442);
and U13624 (N_13624,N_13338,N_13309);
and U13625 (N_13625,N_13393,N_13422);
xnor U13626 (N_13626,N_13350,N_13084);
and U13627 (N_13627,N_13307,N_13425);
and U13628 (N_13628,N_13459,N_13222);
nor U13629 (N_13629,N_13161,N_13115);
and U13630 (N_13630,N_13169,N_13147);
xnor U13631 (N_13631,N_13182,N_13483);
xor U13632 (N_13632,N_13477,N_13332);
xor U13633 (N_13633,N_13238,N_13434);
xnor U13634 (N_13634,N_13373,N_13239);
xnor U13635 (N_13635,N_13272,N_13014);
and U13636 (N_13636,N_13019,N_13316);
nand U13637 (N_13637,N_13033,N_13457);
nand U13638 (N_13638,N_13246,N_13302);
and U13639 (N_13639,N_13492,N_13489);
or U13640 (N_13640,N_13382,N_13107);
xnor U13641 (N_13641,N_13045,N_13027);
or U13642 (N_13642,N_13156,N_13381);
or U13643 (N_13643,N_13144,N_13256);
and U13644 (N_13644,N_13322,N_13100);
nand U13645 (N_13645,N_13275,N_13327);
and U13646 (N_13646,N_13456,N_13406);
xnor U13647 (N_13647,N_13385,N_13351);
and U13648 (N_13648,N_13264,N_13250);
and U13649 (N_13649,N_13421,N_13408);
xnor U13650 (N_13650,N_13347,N_13216);
nor U13651 (N_13651,N_13409,N_13452);
nand U13652 (N_13652,N_13011,N_13236);
and U13653 (N_13653,N_13424,N_13114);
nand U13654 (N_13654,N_13025,N_13196);
xor U13655 (N_13655,N_13087,N_13362);
xnor U13656 (N_13656,N_13258,N_13110);
or U13657 (N_13657,N_13418,N_13472);
nor U13658 (N_13658,N_13463,N_13458);
xnor U13659 (N_13659,N_13402,N_13022);
and U13660 (N_13660,N_13428,N_13028);
nand U13661 (N_13661,N_13358,N_13313);
nand U13662 (N_13662,N_13164,N_13360);
and U13663 (N_13663,N_13066,N_13453);
and U13664 (N_13664,N_13029,N_13138);
nand U13665 (N_13665,N_13252,N_13467);
nor U13666 (N_13666,N_13187,N_13134);
xnor U13667 (N_13667,N_13403,N_13304);
xor U13668 (N_13668,N_13048,N_13448);
nor U13669 (N_13669,N_13020,N_13217);
nand U13670 (N_13670,N_13377,N_13207);
or U13671 (N_13671,N_13249,N_13131);
and U13672 (N_13672,N_13055,N_13185);
nor U13673 (N_13673,N_13384,N_13049);
nand U13674 (N_13674,N_13151,N_13098);
and U13675 (N_13675,N_13093,N_13416);
or U13676 (N_13676,N_13034,N_13104);
and U13677 (N_13677,N_13036,N_13139);
nand U13678 (N_13678,N_13498,N_13122);
nor U13679 (N_13679,N_13069,N_13436);
and U13680 (N_13680,N_13380,N_13198);
nor U13681 (N_13681,N_13190,N_13119);
or U13682 (N_13682,N_13039,N_13074);
and U13683 (N_13683,N_13414,N_13177);
nor U13684 (N_13684,N_13118,N_13040);
or U13685 (N_13685,N_13242,N_13294);
xor U13686 (N_13686,N_13163,N_13057);
nand U13687 (N_13687,N_13062,N_13306);
xnor U13688 (N_13688,N_13241,N_13017);
xnor U13689 (N_13689,N_13274,N_13354);
or U13690 (N_13690,N_13041,N_13287);
nor U13691 (N_13691,N_13423,N_13324);
nand U13692 (N_13692,N_13259,N_13491);
or U13693 (N_13693,N_13474,N_13120);
nand U13694 (N_13694,N_13288,N_13111);
xnor U13695 (N_13695,N_13449,N_13228);
and U13696 (N_13696,N_13050,N_13295);
or U13697 (N_13697,N_13231,N_13031);
nor U13698 (N_13698,N_13030,N_13227);
nor U13699 (N_13699,N_13278,N_13051);
xnor U13700 (N_13700,N_13285,N_13078);
or U13701 (N_13701,N_13305,N_13032);
or U13702 (N_13702,N_13397,N_13230);
or U13703 (N_13703,N_13430,N_13220);
and U13704 (N_13704,N_13325,N_13405);
nor U13705 (N_13705,N_13109,N_13183);
and U13706 (N_13706,N_13172,N_13179);
xnor U13707 (N_13707,N_13496,N_13487);
and U13708 (N_13708,N_13273,N_13085);
or U13709 (N_13709,N_13299,N_13454);
or U13710 (N_13710,N_13127,N_13468);
nor U13711 (N_13711,N_13494,N_13279);
nand U13712 (N_13712,N_13446,N_13482);
or U13713 (N_13713,N_13121,N_13221);
nand U13714 (N_13714,N_13061,N_13270);
or U13715 (N_13715,N_13282,N_13390);
nand U13716 (N_13716,N_13301,N_13166);
or U13717 (N_13717,N_13387,N_13253);
nand U13718 (N_13718,N_13352,N_13361);
nor U13719 (N_13719,N_13329,N_13094);
or U13720 (N_13720,N_13173,N_13437);
nor U13721 (N_13721,N_13392,N_13281);
xor U13722 (N_13722,N_13460,N_13367);
xor U13723 (N_13723,N_13082,N_13088);
and U13724 (N_13724,N_13276,N_13370);
and U13725 (N_13725,N_13013,N_13433);
and U13726 (N_13726,N_13176,N_13461);
and U13727 (N_13727,N_13053,N_13126);
xnor U13728 (N_13728,N_13378,N_13292);
nand U13729 (N_13729,N_13175,N_13255);
nand U13730 (N_13730,N_13086,N_13003);
or U13731 (N_13731,N_13016,N_13261);
and U13732 (N_13732,N_13315,N_13426);
nand U13733 (N_13733,N_13112,N_13308);
xnor U13734 (N_13734,N_13197,N_13257);
nand U13735 (N_13735,N_13052,N_13189);
or U13736 (N_13736,N_13202,N_13391);
nor U13737 (N_13737,N_13290,N_13339);
or U13738 (N_13738,N_13137,N_13089);
nor U13739 (N_13739,N_13070,N_13006);
or U13740 (N_13740,N_13478,N_13155);
nand U13741 (N_13741,N_13291,N_13413);
nand U13742 (N_13742,N_13444,N_13194);
nand U13743 (N_13743,N_13150,N_13193);
nor U13744 (N_13744,N_13103,N_13432);
xor U13745 (N_13745,N_13438,N_13369);
or U13746 (N_13746,N_13317,N_13435);
nor U13747 (N_13747,N_13123,N_13346);
xnor U13748 (N_13748,N_13160,N_13135);
or U13749 (N_13749,N_13349,N_13023);
or U13750 (N_13750,N_13045,N_13430);
xnor U13751 (N_13751,N_13386,N_13084);
xnor U13752 (N_13752,N_13192,N_13361);
xor U13753 (N_13753,N_13295,N_13016);
xor U13754 (N_13754,N_13310,N_13255);
nand U13755 (N_13755,N_13322,N_13359);
and U13756 (N_13756,N_13238,N_13390);
nand U13757 (N_13757,N_13020,N_13434);
and U13758 (N_13758,N_13007,N_13079);
xnor U13759 (N_13759,N_13348,N_13070);
xnor U13760 (N_13760,N_13076,N_13318);
nand U13761 (N_13761,N_13499,N_13335);
nor U13762 (N_13762,N_13300,N_13167);
or U13763 (N_13763,N_13318,N_13176);
nand U13764 (N_13764,N_13117,N_13364);
xnor U13765 (N_13765,N_13034,N_13386);
or U13766 (N_13766,N_13436,N_13116);
nand U13767 (N_13767,N_13346,N_13147);
xor U13768 (N_13768,N_13364,N_13053);
and U13769 (N_13769,N_13415,N_13328);
xnor U13770 (N_13770,N_13336,N_13309);
or U13771 (N_13771,N_13224,N_13143);
nand U13772 (N_13772,N_13223,N_13387);
xnor U13773 (N_13773,N_13465,N_13245);
nor U13774 (N_13774,N_13443,N_13117);
or U13775 (N_13775,N_13137,N_13054);
nand U13776 (N_13776,N_13044,N_13279);
and U13777 (N_13777,N_13262,N_13295);
or U13778 (N_13778,N_13381,N_13176);
nor U13779 (N_13779,N_13287,N_13284);
or U13780 (N_13780,N_13184,N_13195);
nor U13781 (N_13781,N_13392,N_13102);
or U13782 (N_13782,N_13012,N_13173);
xnor U13783 (N_13783,N_13013,N_13001);
xor U13784 (N_13784,N_13201,N_13460);
or U13785 (N_13785,N_13355,N_13377);
and U13786 (N_13786,N_13031,N_13471);
or U13787 (N_13787,N_13245,N_13080);
nor U13788 (N_13788,N_13290,N_13176);
or U13789 (N_13789,N_13359,N_13217);
or U13790 (N_13790,N_13360,N_13321);
or U13791 (N_13791,N_13473,N_13275);
nand U13792 (N_13792,N_13089,N_13224);
and U13793 (N_13793,N_13209,N_13340);
and U13794 (N_13794,N_13167,N_13032);
or U13795 (N_13795,N_13050,N_13247);
or U13796 (N_13796,N_13468,N_13120);
or U13797 (N_13797,N_13428,N_13218);
and U13798 (N_13798,N_13259,N_13355);
nand U13799 (N_13799,N_13420,N_13269);
xnor U13800 (N_13800,N_13154,N_13262);
or U13801 (N_13801,N_13057,N_13307);
and U13802 (N_13802,N_13416,N_13253);
or U13803 (N_13803,N_13228,N_13000);
nand U13804 (N_13804,N_13021,N_13023);
or U13805 (N_13805,N_13086,N_13461);
xor U13806 (N_13806,N_13305,N_13099);
and U13807 (N_13807,N_13395,N_13485);
nor U13808 (N_13808,N_13190,N_13344);
xnor U13809 (N_13809,N_13118,N_13347);
nand U13810 (N_13810,N_13160,N_13334);
and U13811 (N_13811,N_13124,N_13117);
xor U13812 (N_13812,N_13474,N_13342);
or U13813 (N_13813,N_13020,N_13039);
nor U13814 (N_13814,N_13422,N_13459);
xor U13815 (N_13815,N_13156,N_13089);
nor U13816 (N_13816,N_13172,N_13229);
nand U13817 (N_13817,N_13253,N_13355);
nand U13818 (N_13818,N_13368,N_13413);
nand U13819 (N_13819,N_13354,N_13342);
or U13820 (N_13820,N_13255,N_13344);
nand U13821 (N_13821,N_13276,N_13498);
nand U13822 (N_13822,N_13331,N_13001);
and U13823 (N_13823,N_13182,N_13180);
xor U13824 (N_13824,N_13003,N_13132);
or U13825 (N_13825,N_13322,N_13343);
xor U13826 (N_13826,N_13220,N_13230);
nor U13827 (N_13827,N_13175,N_13489);
nor U13828 (N_13828,N_13074,N_13396);
nand U13829 (N_13829,N_13281,N_13298);
xor U13830 (N_13830,N_13249,N_13366);
xor U13831 (N_13831,N_13287,N_13190);
and U13832 (N_13832,N_13356,N_13104);
xor U13833 (N_13833,N_13135,N_13481);
nor U13834 (N_13834,N_13142,N_13497);
and U13835 (N_13835,N_13276,N_13154);
nor U13836 (N_13836,N_13081,N_13330);
nand U13837 (N_13837,N_13472,N_13036);
nor U13838 (N_13838,N_13207,N_13076);
nor U13839 (N_13839,N_13213,N_13440);
xor U13840 (N_13840,N_13292,N_13269);
nand U13841 (N_13841,N_13161,N_13440);
or U13842 (N_13842,N_13093,N_13283);
nand U13843 (N_13843,N_13127,N_13319);
and U13844 (N_13844,N_13229,N_13494);
nand U13845 (N_13845,N_13072,N_13296);
nand U13846 (N_13846,N_13340,N_13084);
or U13847 (N_13847,N_13332,N_13162);
nand U13848 (N_13848,N_13315,N_13356);
nor U13849 (N_13849,N_13496,N_13424);
nor U13850 (N_13850,N_13389,N_13171);
nand U13851 (N_13851,N_13002,N_13387);
or U13852 (N_13852,N_13449,N_13246);
or U13853 (N_13853,N_13424,N_13201);
and U13854 (N_13854,N_13407,N_13311);
or U13855 (N_13855,N_13155,N_13086);
xnor U13856 (N_13856,N_13128,N_13142);
xor U13857 (N_13857,N_13045,N_13493);
xnor U13858 (N_13858,N_13233,N_13047);
nor U13859 (N_13859,N_13263,N_13243);
or U13860 (N_13860,N_13343,N_13250);
xor U13861 (N_13861,N_13394,N_13252);
nor U13862 (N_13862,N_13496,N_13112);
xor U13863 (N_13863,N_13205,N_13371);
nand U13864 (N_13864,N_13350,N_13449);
nand U13865 (N_13865,N_13366,N_13013);
nand U13866 (N_13866,N_13482,N_13298);
or U13867 (N_13867,N_13204,N_13440);
nand U13868 (N_13868,N_13088,N_13181);
or U13869 (N_13869,N_13078,N_13292);
nand U13870 (N_13870,N_13274,N_13241);
and U13871 (N_13871,N_13469,N_13184);
or U13872 (N_13872,N_13326,N_13161);
nand U13873 (N_13873,N_13179,N_13372);
nand U13874 (N_13874,N_13362,N_13184);
and U13875 (N_13875,N_13437,N_13266);
and U13876 (N_13876,N_13056,N_13427);
and U13877 (N_13877,N_13229,N_13187);
or U13878 (N_13878,N_13288,N_13002);
or U13879 (N_13879,N_13215,N_13258);
and U13880 (N_13880,N_13025,N_13170);
and U13881 (N_13881,N_13236,N_13268);
nand U13882 (N_13882,N_13088,N_13168);
and U13883 (N_13883,N_13472,N_13187);
nor U13884 (N_13884,N_13392,N_13095);
or U13885 (N_13885,N_13211,N_13193);
xor U13886 (N_13886,N_13253,N_13046);
nor U13887 (N_13887,N_13003,N_13163);
nand U13888 (N_13888,N_13293,N_13468);
xor U13889 (N_13889,N_13417,N_13051);
nor U13890 (N_13890,N_13286,N_13360);
xnor U13891 (N_13891,N_13087,N_13311);
or U13892 (N_13892,N_13350,N_13091);
or U13893 (N_13893,N_13194,N_13066);
nand U13894 (N_13894,N_13065,N_13027);
nand U13895 (N_13895,N_13004,N_13252);
nor U13896 (N_13896,N_13452,N_13439);
xor U13897 (N_13897,N_13175,N_13060);
or U13898 (N_13898,N_13224,N_13219);
xor U13899 (N_13899,N_13297,N_13408);
xnor U13900 (N_13900,N_13268,N_13402);
nor U13901 (N_13901,N_13112,N_13147);
nor U13902 (N_13902,N_13118,N_13492);
nor U13903 (N_13903,N_13213,N_13452);
or U13904 (N_13904,N_13060,N_13406);
xnor U13905 (N_13905,N_13456,N_13034);
nand U13906 (N_13906,N_13037,N_13201);
xor U13907 (N_13907,N_13117,N_13446);
or U13908 (N_13908,N_13293,N_13335);
and U13909 (N_13909,N_13391,N_13345);
nand U13910 (N_13910,N_13329,N_13328);
and U13911 (N_13911,N_13142,N_13380);
and U13912 (N_13912,N_13192,N_13057);
xnor U13913 (N_13913,N_13278,N_13381);
or U13914 (N_13914,N_13369,N_13054);
xor U13915 (N_13915,N_13464,N_13469);
and U13916 (N_13916,N_13153,N_13424);
xnor U13917 (N_13917,N_13154,N_13420);
or U13918 (N_13918,N_13159,N_13087);
or U13919 (N_13919,N_13201,N_13359);
and U13920 (N_13920,N_13412,N_13459);
xor U13921 (N_13921,N_13446,N_13196);
nand U13922 (N_13922,N_13354,N_13077);
nor U13923 (N_13923,N_13098,N_13139);
or U13924 (N_13924,N_13244,N_13411);
nor U13925 (N_13925,N_13477,N_13488);
xnor U13926 (N_13926,N_13400,N_13291);
nand U13927 (N_13927,N_13268,N_13226);
nor U13928 (N_13928,N_13366,N_13215);
and U13929 (N_13929,N_13362,N_13036);
nand U13930 (N_13930,N_13051,N_13455);
and U13931 (N_13931,N_13423,N_13373);
nand U13932 (N_13932,N_13307,N_13056);
or U13933 (N_13933,N_13332,N_13146);
xnor U13934 (N_13934,N_13113,N_13256);
or U13935 (N_13935,N_13327,N_13066);
nand U13936 (N_13936,N_13080,N_13464);
and U13937 (N_13937,N_13321,N_13236);
nand U13938 (N_13938,N_13070,N_13429);
or U13939 (N_13939,N_13336,N_13432);
nor U13940 (N_13940,N_13422,N_13242);
or U13941 (N_13941,N_13340,N_13409);
nand U13942 (N_13942,N_13322,N_13111);
xor U13943 (N_13943,N_13467,N_13190);
and U13944 (N_13944,N_13421,N_13146);
and U13945 (N_13945,N_13232,N_13479);
xnor U13946 (N_13946,N_13360,N_13028);
xor U13947 (N_13947,N_13230,N_13008);
nand U13948 (N_13948,N_13067,N_13473);
xnor U13949 (N_13949,N_13129,N_13094);
and U13950 (N_13950,N_13039,N_13494);
or U13951 (N_13951,N_13298,N_13137);
and U13952 (N_13952,N_13384,N_13142);
nor U13953 (N_13953,N_13164,N_13172);
nand U13954 (N_13954,N_13252,N_13436);
nor U13955 (N_13955,N_13059,N_13478);
xnor U13956 (N_13956,N_13235,N_13130);
nand U13957 (N_13957,N_13292,N_13129);
xnor U13958 (N_13958,N_13131,N_13165);
or U13959 (N_13959,N_13127,N_13461);
nor U13960 (N_13960,N_13147,N_13209);
xor U13961 (N_13961,N_13332,N_13234);
nand U13962 (N_13962,N_13488,N_13208);
nor U13963 (N_13963,N_13393,N_13007);
xor U13964 (N_13964,N_13362,N_13274);
xnor U13965 (N_13965,N_13119,N_13386);
nand U13966 (N_13966,N_13266,N_13378);
nand U13967 (N_13967,N_13297,N_13473);
nand U13968 (N_13968,N_13292,N_13418);
nor U13969 (N_13969,N_13241,N_13130);
nand U13970 (N_13970,N_13280,N_13110);
or U13971 (N_13971,N_13480,N_13070);
nand U13972 (N_13972,N_13237,N_13092);
nand U13973 (N_13973,N_13158,N_13074);
or U13974 (N_13974,N_13183,N_13218);
xnor U13975 (N_13975,N_13190,N_13483);
and U13976 (N_13976,N_13020,N_13260);
or U13977 (N_13977,N_13228,N_13039);
or U13978 (N_13978,N_13254,N_13150);
or U13979 (N_13979,N_13467,N_13203);
nand U13980 (N_13980,N_13099,N_13450);
nor U13981 (N_13981,N_13294,N_13302);
or U13982 (N_13982,N_13281,N_13261);
or U13983 (N_13983,N_13352,N_13495);
or U13984 (N_13984,N_13380,N_13265);
nand U13985 (N_13985,N_13299,N_13276);
or U13986 (N_13986,N_13459,N_13450);
or U13987 (N_13987,N_13445,N_13024);
nand U13988 (N_13988,N_13437,N_13263);
xor U13989 (N_13989,N_13319,N_13327);
nand U13990 (N_13990,N_13453,N_13336);
nor U13991 (N_13991,N_13357,N_13315);
nand U13992 (N_13992,N_13457,N_13055);
and U13993 (N_13993,N_13139,N_13124);
nor U13994 (N_13994,N_13191,N_13266);
and U13995 (N_13995,N_13020,N_13169);
nor U13996 (N_13996,N_13098,N_13346);
and U13997 (N_13997,N_13244,N_13395);
and U13998 (N_13998,N_13398,N_13087);
xnor U13999 (N_13999,N_13493,N_13219);
or U14000 (N_14000,N_13613,N_13911);
and U14001 (N_14001,N_13539,N_13526);
or U14002 (N_14002,N_13600,N_13980);
or U14003 (N_14003,N_13877,N_13651);
or U14004 (N_14004,N_13869,N_13700);
nand U14005 (N_14005,N_13833,N_13958);
xnor U14006 (N_14006,N_13992,N_13543);
and U14007 (N_14007,N_13918,N_13939);
nand U14008 (N_14008,N_13908,N_13741);
and U14009 (N_14009,N_13981,N_13919);
or U14010 (N_14010,N_13862,N_13948);
and U14011 (N_14011,N_13798,N_13786);
xnor U14012 (N_14012,N_13550,N_13610);
nand U14013 (N_14013,N_13721,N_13767);
nor U14014 (N_14014,N_13959,N_13515);
or U14015 (N_14015,N_13866,N_13743);
nand U14016 (N_14016,N_13556,N_13765);
and U14017 (N_14017,N_13787,N_13538);
or U14018 (N_14018,N_13520,N_13731);
nand U14019 (N_14019,N_13634,N_13923);
nor U14020 (N_14020,N_13548,N_13816);
nand U14021 (N_14021,N_13594,N_13847);
nand U14022 (N_14022,N_13977,N_13680);
and U14023 (N_14023,N_13702,N_13682);
nor U14024 (N_14024,N_13517,N_13739);
and U14025 (N_14025,N_13606,N_13684);
xnor U14026 (N_14026,N_13687,N_13521);
and U14027 (N_14027,N_13863,N_13542);
and U14028 (N_14028,N_13755,N_13834);
xor U14029 (N_14029,N_13635,N_13678);
nor U14030 (N_14030,N_13713,N_13857);
nor U14031 (N_14031,N_13621,N_13657);
xnor U14032 (N_14032,N_13936,N_13818);
xor U14033 (N_14033,N_13934,N_13507);
or U14034 (N_14034,N_13528,N_13845);
nor U14035 (N_14035,N_13750,N_13851);
nand U14036 (N_14036,N_13802,N_13576);
nand U14037 (N_14037,N_13852,N_13704);
and U14038 (N_14038,N_13985,N_13685);
nand U14039 (N_14039,N_13558,N_13940);
nand U14040 (N_14040,N_13695,N_13806);
or U14041 (N_14041,N_13995,N_13697);
or U14042 (N_14042,N_13575,N_13945);
nor U14043 (N_14043,N_13552,N_13503);
or U14044 (N_14044,N_13782,N_13585);
nand U14045 (N_14045,N_13873,N_13951);
nand U14046 (N_14046,N_13671,N_13547);
and U14047 (N_14047,N_13630,N_13904);
xor U14048 (N_14048,N_13691,N_13557);
nor U14049 (N_14049,N_13928,N_13997);
and U14050 (N_14050,N_13780,N_13648);
nor U14051 (N_14051,N_13701,N_13902);
or U14052 (N_14052,N_13579,N_13855);
xor U14053 (N_14053,N_13772,N_13778);
nand U14054 (N_14054,N_13795,N_13551);
nand U14055 (N_14055,N_13960,N_13819);
nand U14056 (N_14056,N_13588,N_13624);
and U14057 (N_14057,N_13903,N_13860);
and U14058 (N_14058,N_13897,N_13955);
nor U14059 (N_14059,N_13622,N_13712);
xnor U14060 (N_14060,N_13553,N_13783);
and U14061 (N_14061,N_13950,N_13896);
nand U14062 (N_14062,N_13753,N_13763);
and U14063 (N_14063,N_13616,N_13815);
xnor U14064 (N_14064,N_13524,N_13971);
or U14065 (N_14065,N_13728,N_13681);
nor U14066 (N_14066,N_13751,N_13830);
xor U14067 (N_14067,N_13650,N_13603);
nor U14068 (N_14068,N_13831,N_13566);
or U14069 (N_14069,N_13966,N_13676);
xor U14070 (N_14070,N_13722,N_13914);
or U14071 (N_14071,N_13719,N_13907);
or U14072 (N_14072,N_13703,N_13506);
or U14073 (N_14073,N_13508,N_13663);
or U14074 (N_14074,N_13848,N_13620);
nor U14075 (N_14075,N_13688,N_13867);
nand U14076 (N_14076,N_13589,N_13813);
nand U14077 (N_14077,N_13853,N_13698);
and U14078 (N_14078,N_13649,N_13623);
nor U14079 (N_14079,N_13692,N_13584);
xor U14080 (N_14080,N_13886,N_13673);
nor U14081 (N_14081,N_13826,N_13632);
or U14082 (N_14082,N_13982,N_13937);
and U14083 (N_14083,N_13799,N_13746);
xnor U14084 (N_14084,N_13920,N_13822);
or U14085 (N_14085,N_13514,N_13581);
nand U14086 (N_14086,N_13730,N_13757);
and U14087 (N_14087,N_13736,N_13762);
and U14088 (N_14088,N_13916,N_13724);
nand U14089 (N_14089,N_13626,N_13841);
or U14090 (N_14090,N_13737,N_13760);
and U14091 (N_14091,N_13643,N_13991);
xor U14092 (N_14092,N_13734,N_13609);
and U14093 (N_14093,N_13769,N_13509);
and U14094 (N_14094,N_13998,N_13775);
nand U14095 (N_14095,N_13582,N_13823);
or U14096 (N_14096,N_13935,N_13954);
and U14097 (N_14097,N_13619,N_13807);
and U14098 (N_14098,N_13779,N_13604);
nor U14099 (N_14099,N_13749,N_13870);
or U14100 (N_14100,N_13735,N_13773);
nand U14101 (N_14101,N_13549,N_13764);
and U14102 (N_14102,N_13989,N_13874);
nor U14103 (N_14103,N_13871,N_13617);
xor U14104 (N_14104,N_13797,N_13888);
xnor U14105 (N_14105,N_13597,N_13534);
nor U14106 (N_14106,N_13942,N_13660);
and U14107 (N_14107,N_13544,N_13518);
and U14108 (N_14108,N_13905,N_13710);
nand U14109 (N_14109,N_13522,N_13814);
and U14110 (N_14110,N_13525,N_13967);
or U14111 (N_14111,N_13884,N_13596);
nand U14112 (N_14112,N_13889,N_13652);
nor U14113 (N_14113,N_13562,N_13969);
nand U14114 (N_14114,N_13690,N_13745);
xnor U14115 (N_14115,N_13844,N_13975);
and U14116 (N_14116,N_13664,N_13835);
nand U14117 (N_14117,N_13895,N_13627);
xnor U14118 (N_14118,N_13591,N_13659);
nor U14119 (N_14119,N_13668,N_13832);
nand U14120 (N_14120,N_13513,N_13865);
or U14121 (N_14121,N_13718,N_13602);
xor U14122 (N_14122,N_13979,N_13666);
nand U14123 (N_14123,N_13973,N_13986);
nand U14124 (N_14124,N_13868,N_13561);
nand U14125 (N_14125,N_13727,N_13900);
or U14126 (N_14126,N_13983,N_13768);
nand U14127 (N_14127,N_13638,N_13527);
xnor U14128 (N_14128,N_13641,N_13824);
nor U14129 (N_14129,N_13829,N_13607);
or U14130 (N_14130,N_13988,N_13943);
xor U14131 (N_14131,N_13812,N_13825);
or U14132 (N_14132,N_13968,N_13742);
or U14133 (N_14133,N_13693,N_13500);
or U14134 (N_14134,N_13530,N_13628);
nand U14135 (N_14135,N_13744,N_13726);
and U14136 (N_14136,N_13661,N_13598);
nand U14137 (N_14137,N_13689,N_13752);
and U14138 (N_14138,N_13892,N_13861);
xnor U14139 (N_14139,N_13670,N_13696);
xnor U14140 (N_14140,N_13963,N_13910);
and U14141 (N_14141,N_13887,N_13647);
xor U14142 (N_14142,N_13504,N_13791);
nor U14143 (N_14143,N_13964,N_13839);
nand U14144 (N_14144,N_13974,N_13754);
and U14145 (N_14145,N_13707,N_13926);
nor U14146 (N_14146,N_13801,N_13850);
nor U14147 (N_14147,N_13972,N_13636);
and U14148 (N_14148,N_13578,N_13864);
nand U14149 (N_14149,N_13714,N_13587);
nand U14150 (N_14150,N_13876,N_13715);
nor U14151 (N_14151,N_13810,N_13674);
nand U14152 (N_14152,N_13859,N_13915);
xor U14153 (N_14153,N_13559,N_13747);
nand U14154 (N_14154,N_13709,N_13890);
nor U14155 (N_14155,N_13803,N_13932);
nand U14156 (N_14156,N_13523,N_13792);
nor U14157 (N_14157,N_13925,N_13879);
nor U14158 (N_14158,N_13679,N_13882);
and U14159 (N_14159,N_13796,N_13569);
nand U14160 (N_14160,N_13642,N_13574);
nand U14161 (N_14161,N_13501,N_13941);
or U14162 (N_14162,N_13637,N_13554);
xor U14163 (N_14163,N_13531,N_13804);
or U14164 (N_14164,N_13842,N_13567);
and U14165 (N_14165,N_13961,N_13725);
nor U14166 (N_14166,N_13706,N_13672);
and U14167 (N_14167,N_13683,N_13790);
nor U14168 (N_14168,N_13793,N_13808);
xor U14169 (N_14169,N_13717,N_13846);
nor U14170 (N_14170,N_13645,N_13956);
and U14171 (N_14171,N_13781,N_13921);
or U14172 (N_14172,N_13699,N_13629);
nor U14173 (N_14173,N_13608,N_13944);
nand U14174 (N_14174,N_13677,N_13540);
xnor U14175 (N_14175,N_13893,N_13733);
nand U14176 (N_14176,N_13878,N_13872);
nand U14177 (N_14177,N_13511,N_13720);
and U14178 (N_14178,N_13686,N_13883);
nand U14179 (N_14179,N_13563,N_13568);
xor U14180 (N_14180,N_13996,N_13560);
and U14181 (N_14181,N_13953,N_13922);
nand U14182 (N_14182,N_13512,N_13748);
or U14183 (N_14183,N_13555,N_13809);
nand U14184 (N_14184,N_13740,N_13827);
and U14185 (N_14185,N_13776,N_13811);
or U14186 (N_14186,N_13946,N_13618);
and U14187 (N_14187,N_13665,N_13800);
and U14188 (N_14188,N_13994,N_13881);
or U14189 (N_14189,N_13933,N_13631);
xor U14190 (N_14190,N_13510,N_13573);
and U14191 (N_14191,N_13614,N_13756);
nor U14192 (N_14192,N_13906,N_13858);
and U14193 (N_14193,N_13605,N_13894);
and U14194 (N_14194,N_13639,N_13952);
nand U14195 (N_14195,N_13820,N_13590);
nor U14196 (N_14196,N_13577,N_13532);
nor U14197 (N_14197,N_13794,N_13917);
and U14198 (N_14198,N_13962,N_13502);
nand U14199 (N_14199,N_13705,N_13817);
xnor U14200 (N_14200,N_13970,N_13976);
nand U14201 (N_14201,N_13729,N_13931);
xnor U14202 (N_14202,N_13732,N_13828);
xnor U14203 (N_14203,N_13565,N_13854);
and U14204 (N_14204,N_13947,N_13541);
and U14205 (N_14205,N_13761,N_13957);
nand U14206 (N_14206,N_13771,N_13837);
or U14207 (N_14207,N_13662,N_13535);
and U14208 (N_14208,N_13843,N_13993);
xor U14209 (N_14209,N_13564,N_13669);
nand U14210 (N_14210,N_13901,N_13949);
and U14211 (N_14211,N_13840,N_13533);
nand U14212 (N_14212,N_13653,N_13849);
and U14213 (N_14213,N_13880,N_13716);
or U14214 (N_14214,N_13675,N_13546);
nor U14215 (N_14215,N_13758,N_13536);
or U14216 (N_14216,N_13570,N_13938);
and U14217 (N_14217,N_13572,N_13519);
xor U14218 (N_14218,N_13978,N_13655);
or U14219 (N_14219,N_13708,N_13875);
and U14220 (N_14220,N_13785,N_13633);
or U14221 (N_14221,N_13601,N_13545);
or U14222 (N_14222,N_13821,N_13656);
nor U14223 (N_14223,N_13899,N_13836);
and U14224 (N_14224,N_13770,N_13580);
or U14225 (N_14225,N_13805,N_13738);
xnor U14226 (N_14226,N_13644,N_13723);
and U14227 (N_14227,N_13999,N_13583);
or U14228 (N_14228,N_13929,N_13891);
or U14229 (N_14229,N_13571,N_13927);
nand U14230 (N_14230,N_13856,N_13898);
xnor U14231 (N_14231,N_13586,N_13990);
nor U14232 (N_14232,N_13766,N_13611);
nand U14233 (N_14233,N_13838,N_13788);
and U14234 (N_14234,N_13930,N_13711);
or U14235 (N_14235,N_13615,N_13777);
xor U14236 (N_14236,N_13505,N_13759);
nor U14237 (N_14237,N_13599,N_13913);
and U14238 (N_14238,N_13984,N_13516);
and U14239 (N_14239,N_13592,N_13658);
nand U14240 (N_14240,N_13987,N_13965);
xnor U14241 (N_14241,N_13625,N_13646);
nor U14242 (N_14242,N_13640,N_13909);
nor U14243 (N_14243,N_13612,N_13885);
and U14244 (N_14244,N_13537,N_13784);
or U14245 (N_14245,N_13912,N_13595);
xnor U14246 (N_14246,N_13694,N_13529);
and U14247 (N_14247,N_13789,N_13924);
nand U14248 (N_14248,N_13654,N_13667);
or U14249 (N_14249,N_13774,N_13593);
xor U14250 (N_14250,N_13973,N_13953);
nand U14251 (N_14251,N_13906,N_13920);
xor U14252 (N_14252,N_13887,N_13724);
xnor U14253 (N_14253,N_13511,N_13703);
and U14254 (N_14254,N_13780,N_13875);
nand U14255 (N_14255,N_13952,N_13829);
and U14256 (N_14256,N_13949,N_13853);
and U14257 (N_14257,N_13583,N_13868);
and U14258 (N_14258,N_13524,N_13578);
and U14259 (N_14259,N_13518,N_13918);
or U14260 (N_14260,N_13712,N_13543);
nor U14261 (N_14261,N_13665,N_13650);
xnor U14262 (N_14262,N_13610,N_13618);
nor U14263 (N_14263,N_13698,N_13867);
or U14264 (N_14264,N_13631,N_13998);
or U14265 (N_14265,N_13511,N_13563);
and U14266 (N_14266,N_13730,N_13812);
nor U14267 (N_14267,N_13709,N_13942);
nand U14268 (N_14268,N_13749,N_13934);
and U14269 (N_14269,N_13949,N_13834);
or U14270 (N_14270,N_13678,N_13985);
and U14271 (N_14271,N_13817,N_13884);
or U14272 (N_14272,N_13576,N_13644);
and U14273 (N_14273,N_13787,N_13641);
nor U14274 (N_14274,N_13976,N_13511);
xor U14275 (N_14275,N_13988,N_13670);
nand U14276 (N_14276,N_13604,N_13990);
and U14277 (N_14277,N_13985,N_13550);
nor U14278 (N_14278,N_13753,N_13993);
xor U14279 (N_14279,N_13965,N_13898);
nor U14280 (N_14280,N_13594,N_13846);
and U14281 (N_14281,N_13647,N_13666);
and U14282 (N_14282,N_13913,N_13834);
xor U14283 (N_14283,N_13899,N_13620);
xnor U14284 (N_14284,N_13980,N_13603);
xor U14285 (N_14285,N_13523,N_13663);
or U14286 (N_14286,N_13586,N_13933);
nor U14287 (N_14287,N_13859,N_13870);
nand U14288 (N_14288,N_13781,N_13893);
or U14289 (N_14289,N_13970,N_13710);
or U14290 (N_14290,N_13559,N_13727);
nor U14291 (N_14291,N_13635,N_13862);
xor U14292 (N_14292,N_13562,N_13626);
nor U14293 (N_14293,N_13597,N_13991);
and U14294 (N_14294,N_13719,N_13935);
or U14295 (N_14295,N_13752,N_13796);
xnor U14296 (N_14296,N_13639,N_13991);
xnor U14297 (N_14297,N_13764,N_13789);
or U14298 (N_14298,N_13742,N_13791);
and U14299 (N_14299,N_13538,N_13500);
xnor U14300 (N_14300,N_13571,N_13670);
nor U14301 (N_14301,N_13964,N_13577);
nor U14302 (N_14302,N_13996,N_13729);
or U14303 (N_14303,N_13949,N_13771);
xnor U14304 (N_14304,N_13582,N_13765);
nor U14305 (N_14305,N_13533,N_13953);
nand U14306 (N_14306,N_13885,N_13870);
and U14307 (N_14307,N_13781,N_13522);
and U14308 (N_14308,N_13538,N_13603);
xor U14309 (N_14309,N_13680,N_13869);
nor U14310 (N_14310,N_13903,N_13610);
and U14311 (N_14311,N_13922,N_13568);
and U14312 (N_14312,N_13985,N_13799);
nand U14313 (N_14313,N_13965,N_13882);
nand U14314 (N_14314,N_13934,N_13944);
nand U14315 (N_14315,N_13572,N_13995);
nand U14316 (N_14316,N_13548,N_13692);
and U14317 (N_14317,N_13730,N_13844);
nand U14318 (N_14318,N_13520,N_13586);
and U14319 (N_14319,N_13960,N_13941);
and U14320 (N_14320,N_13939,N_13782);
nor U14321 (N_14321,N_13791,N_13527);
and U14322 (N_14322,N_13759,N_13735);
xor U14323 (N_14323,N_13834,N_13776);
and U14324 (N_14324,N_13524,N_13908);
and U14325 (N_14325,N_13630,N_13627);
nand U14326 (N_14326,N_13562,N_13726);
or U14327 (N_14327,N_13965,N_13577);
nor U14328 (N_14328,N_13730,N_13796);
nand U14329 (N_14329,N_13992,N_13759);
xnor U14330 (N_14330,N_13859,N_13744);
xor U14331 (N_14331,N_13524,N_13673);
or U14332 (N_14332,N_13748,N_13906);
xor U14333 (N_14333,N_13829,N_13675);
nor U14334 (N_14334,N_13735,N_13799);
or U14335 (N_14335,N_13883,N_13574);
and U14336 (N_14336,N_13763,N_13657);
and U14337 (N_14337,N_13701,N_13574);
nand U14338 (N_14338,N_13860,N_13864);
or U14339 (N_14339,N_13789,N_13830);
or U14340 (N_14340,N_13789,N_13808);
xnor U14341 (N_14341,N_13783,N_13752);
nor U14342 (N_14342,N_13717,N_13815);
xor U14343 (N_14343,N_13965,N_13779);
nand U14344 (N_14344,N_13797,N_13969);
nand U14345 (N_14345,N_13991,N_13910);
and U14346 (N_14346,N_13602,N_13553);
and U14347 (N_14347,N_13968,N_13558);
nand U14348 (N_14348,N_13655,N_13926);
or U14349 (N_14349,N_13883,N_13820);
and U14350 (N_14350,N_13885,N_13552);
nand U14351 (N_14351,N_13997,N_13809);
nand U14352 (N_14352,N_13907,N_13787);
xor U14353 (N_14353,N_13732,N_13907);
nand U14354 (N_14354,N_13905,N_13547);
nand U14355 (N_14355,N_13569,N_13721);
nor U14356 (N_14356,N_13933,N_13773);
and U14357 (N_14357,N_13803,N_13722);
nand U14358 (N_14358,N_13608,N_13751);
or U14359 (N_14359,N_13534,N_13754);
or U14360 (N_14360,N_13915,N_13842);
nand U14361 (N_14361,N_13762,N_13606);
nand U14362 (N_14362,N_13877,N_13766);
and U14363 (N_14363,N_13952,N_13828);
xnor U14364 (N_14364,N_13718,N_13502);
or U14365 (N_14365,N_13643,N_13912);
nand U14366 (N_14366,N_13693,N_13627);
and U14367 (N_14367,N_13603,N_13880);
and U14368 (N_14368,N_13583,N_13983);
and U14369 (N_14369,N_13666,N_13792);
and U14370 (N_14370,N_13797,N_13640);
nor U14371 (N_14371,N_13841,N_13931);
nand U14372 (N_14372,N_13542,N_13967);
xor U14373 (N_14373,N_13760,N_13949);
nor U14374 (N_14374,N_13801,N_13711);
nor U14375 (N_14375,N_13655,N_13640);
nor U14376 (N_14376,N_13990,N_13676);
and U14377 (N_14377,N_13615,N_13857);
xnor U14378 (N_14378,N_13737,N_13563);
and U14379 (N_14379,N_13692,N_13516);
and U14380 (N_14380,N_13989,N_13712);
or U14381 (N_14381,N_13951,N_13591);
nand U14382 (N_14382,N_13973,N_13510);
xor U14383 (N_14383,N_13515,N_13600);
or U14384 (N_14384,N_13608,N_13587);
and U14385 (N_14385,N_13793,N_13979);
nand U14386 (N_14386,N_13736,N_13668);
or U14387 (N_14387,N_13646,N_13576);
or U14388 (N_14388,N_13793,N_13710);
or U14389 (N_14389,N_13614,N_13846);
and U14390 (N_14390,N_13806,N_13732);
xnor U14391 (N_14391,N_13813,N_13766);
nor U14392 (N_14392,N_13764,N_13625);
nand U14393 (N_14393,N_13879,N_13687);
nor U14394 (N_14394,N_13588,N_13573);
nor U14395 (N_14395,N_13568,N_13952);
nor U14396 (N_14396,N_13924,N_13900);
nand U14397 (N_14397,N_13754,N_13897);
nor U14398 (N_14398,N_13713,N_13507);
nand U14399 (N_14399,N_13692,N_13794);
nand U14400 (N_14400,N_13922,N_13774);
nor U14401 (N_14401,N_13764,N_13893);
nor U14402 (N_14402,N_13501,N_13738);
or U14403 (N_14403,N_13596,N_13742);
and U14404 (N_14404,N_13940,N_13539);
nand U14405 (N_14405,N_13609,N_13611);
xnor U14406 (N_14406,N_13799,N_13995);
nand U14407 (N_14407,N_13906,N_13520);
xnor U14408 (N_14408,N_13714,N_13525);
and U14409 (N_14409,N_13841,N_13608);
nand U14410 (N_14410,N_13617,N_13544);
nand U14411 (N_14411,N_13953,N_13646);
nor U14412 (N_14412,N_13534,N_13675);
nor U14413 (N_14413,N_13776,N_13968);
nand U14414 (N_14414,N_13790,N_13518);
and U14415 (N_14415,N_13993,N_13740);
xor U14416 (N_14416,N_13600,N_13602);
or U14417 (N_14417,N_13727,N_13558);
nor U14418 (N_14418,N_13573,N_13774);
xor U14419 (N_14419,N_13946,N_13588);
and U14420 (N_14420,N_13813,N_13559);
nand U14421 (N_14421,N_13562,N_13896);
or U14422 (N_14422,N_13881,N_13739);
nand U14423 (N_14423,N_13843,N_13892);
and U14424 (N_14424,N_13529,N_13585);
xor U14425 (N_14425,N_13621,N_13968);
or U14426 (N_14426,N_13788,N_13823);
and U14427 (N_14427,N_13882,N_13732);
xnor U14428 (N_14428,N_13838,N_13982);
or U14429 (N_14429,N_13625,N_13876);
nor U14430 (N_14430,N_13793,N_13898);
nand U14431 (N_14431,N_13502,N_13571);
and U14432 (N_14432,N_13503,N_13642);
or U14433 (N_14433,N_13574,N_13977);
xnor U14434 (N_14434,N_13872,N_13634);
and U14435 (N_14435,N_13772,N_13975);
and U14436 (N_14436,N_13712,N_13754);
nor U14437 (N_14437,N_13540,N_13534);
nand U14438 (N_14438,N_13901,N_13583);
or U14439 (N_14439,N_13655,N_13589);
xnor U14440 (N_14440,N_13776,N_13795);
or U14441 (N_14441,N_13808,N_13605);
nand U14442 (N_14442,N_13817,N_13963);
xnor U14443 (N_14443,N_13941,N_13512);
and U14444 (N_14444,N_13551,N_13577);
xnor U14445 (N_14445,N_13578,N_13512);
or U14446 (N_14446,N_13960,N_13957);
nand U14447 (N_14447,N_13898,N_13598);
or U14448 (N_14448,N_13836,N_13614);
nor U14449 (N_14449,N_13633,N_13578);
xor U14450 (N_14450,N_13882,N_13557);
or U14451 (N_14451,N_13734,N_13708);
or U14452 (N_14452,N_13682,N_13958);
xor U14453 (N_14453,N_13637,N_13857);
or U14454 (N_14454,N_13767,N_13670);
nand U14455 (N_14455,N_13508,N_13611);
xnor U14456 (N_14456,N_13703,N_13587);
or U14457 (N_14457,N_13877,N_13789);
nor U14458 (N_14458,N_13585,N_13998);
nor U14459 (N_14459,N_13951,N_13732);
or U14460 (N_14460,N_13585,N_13663);
nand U14461 (N_14461,N_13700,N_13763);
xnor U14462 (N_14462,N_13773,N_13555);
xor U14463 (N_14463,N_13549,N_13506);
xnor U14464 (N_14464,N_13644,N_13796);
nor U14465 (N_14465,N_13779,N_13660);
and U14466 (N_14466,N_13786,N_13598);
xor U14467 (N_14467,N_13578,N_13931);
or U14468 (N_14468,N_13878,N_13657);
and U14469 (N_14469,N_13756,N_13543);
nor U14470 (N_14470,N_13944,N_13867);
or U14471 (N_14471,N_13659,N_13646);
nor U14472 (N_14472,N_13839,N_13907);
or U14473 (N_14473,N_13824,N_13687);
and U14474 (N_14474,N_13806,N_13713);
xor U14475 (N_14475,N_13815,N_13568);
nand U14476 (N_14476,N_13620,N_13832);
xor U14477 (N_14477,N_13547,N_13867);
nor U14478 (N_14478,N_13837,N_13738);
xor U14479 (N_14479,N_13588,N_13938);
nor U14480 (N_14480,N_13500,N_13864);
and U14481 (N_14481,N_13944,N_13732);
or U14482 (N_14482,N_13593,N_13860);
and U14483 (N_14483,N_13803,N_13541);
and U14484 (N_14484,N_13852,N_13562);
nand U14485 (N_14485,N_13705,N_13833);
and U14486 (N_14486,N_13987,N_13772);
and U14487 (N_14487,N_13557,N_13548);
and U14488 (N_14488,N_13637,N_13732);
nand U14489 (N_14489,N_13792,N_13737);
nand U14490 (N_14490,N_13674,N_13526);
or U14491 (N_14491,N_13971,N_13597);
xnor U14492 (N_14492,N_13857,N_13879);
or U14493 (N_14493,N_13971,N_13812);
nand U14494 (N_14494,N_13927,N_13561);
or U14495 (N_14495,N_13802,N_13932);
nand U14496 (N_14496,N_13793,N_13501);
nand U14497 (N_14497,N_13913,N_13888);
nand U14498 (N_14498,N_13998,N_13716);
or U14499 (N_14499,N_13515,N_13815);
nand U14500 (N_14500,N_14294,N_14168);
nand U14501 (N_14501,N_14326,N_14148);
and U14502 (N_14502,N_14440,N_14262);
and U14503 (N_14503,N_14385,N_14220);
nand U14504 (N_14504,N_14129,N_14467);
or U14505 (N_14505,N_14456,N_14119);
nand U14506 (N_14506,N_14007,N_14198);
nor U14507 (N_14507,N_14318,N_14425);
xor U14508 (N_14508,N_14340,N_14136);
xor U14509 (N_14509,N_14170,N_14342);
and U14510 (N_14510,N_14005,N_14265);
or U14511 (N_14511,N_14441,N_14354);
or U14512 (N_14512,N_14355,N_14317);
nor U14513 (N_14513,N_14033,N_14347);
xor U14514 (N_14514,N_14364,N_14161);
or U14515 (N_14515,N_14312,N_14057);
and U14516 (N_14516,N_14329,N_14357);
nor U14517 (N_14517,N_14348,N_14343);
nand U14518 (N_14518,N_14284,N_14041);
and U14519 (N_14519,N_14091,N_14038);
nor U14520 (N_14520,N_14472,N_14483);
nor U14521 (N_14521,N_14249,N_14020);
and U14522 (N_14522,N_14495,N_14200);
or U14523 (N_14523,N_14291,N_14131);
xnor U14524 (N_14524,N_14098,N_14463);
or U14525 (N_14525,N_14108,N_14388);
or U14526 (N_14526,N_14125,N_14071);
or U14527 (N_14527,N_14165,N_14345);
and U14528 (N_14528,N_14169,N_14195);
and U14529 (N_14529,N_14142,N_14427);
xnor U14530 (N_14530,N_14167,N_14060);
and U14531 (N_14531,N_14094,N_14276);
nand U14532 (N_14532,N_14448,N_14287);
and U14533 (N_14533,N_14277,N_14279);
nor U14534 (N_14534,N_14380,N_14303);
nor U14535 (N_14535,N_14429,N_14063);
or U14536 (N_14536,N_14360,N_14045);
nand U14537 (N_14537,N_14024,N_14036);
or U14538 (N_14538,N_14308,N_14025);
nor U14539 (N_14539,N_14133,N_14186);
and U14540 (N_14540,N_14451,N_14084);
or U14541 (N_14541,N_14235,N_14123);
xor U14542 (N_14542,N_14118,N_14029);
nand U14543 (N_14543,N_14367,N_14077);
xnor U14544 (N_14544,N_14092,N_14469);
nor U14545 (N_14545,N_14110,N_14002);
nor U14546 (N_14546,N_14274,N_14065);
or U14547 (N_14547,N_14461,N_14283);
and U14548 (N_14548,N_14246,N_14175);
nand U14549 (N_14549,N_14420,N_14115);
nand U14550 (N_14550,N_14327,N_14212);
nor U14551 (N_14551,N_14482,N_14059);
or U14552 (N_14552,N_14035,N_14245);
or U14553 (N_14553,N_14134,N_14358);
xor U14554 (N_14554,N_14229,N_14314);
and U14555 (N_14555,N_14346,N_14078);
nand U14556 (N_14556,N_14371,N_14064);
nand U14557 (N_14557,N_14137,N_14275);
or U14558 (N_14558,N_14412,N_14491);
or U14559 (N_14559,N_14408,N_14179);
nand U14560 (N_14560,N_14122,N_14386);
and U14561 (N_14561,N_14419,N_14426);
xnor U14562 (N_14562,N_14185,N_14101);
nor U14563 (N_14563,N_14076,N_14389);
nor U14564 (N_14564,N_14305,N_14428);
xor U14565 (N_14565,N_14183,N_14117);
and U14566 (N_14566,N_14485,N_14295);
nor U14567 (N_14567,N_14434,N_14010);
nor U14568 (N_14568,N_14039,N_14356);
xnor U14569 (N_14569,N_14376,N_14177);
nand U14570 (N_14570,N_14104,N_14166);
xor U14571 (N_14571,N_14404,N_14266);
xnor U14572 (N_14572,N_14079,N_14192);
or U14573 (N_14573,N_14339,N_14324);
nand U14574 (N_14574,N_14344,N_14350);
nand U14575 (N_14575,N_14099,N_14213);
nand U14576 (N_14576,N_14333,N_14152);
and U14577 (N_14577,N_14302,N_14218);
nor U14578 (N_14578,N_14151,N_14121);
or U14579 (N_14579,N_14251,N_14013);
or U14580 (N_14580,N_14335,N_14257);
or U14581 (N_14581,N_14297,N_14252);
nor U14582 (N_14582,N_14256,N_14062);
nor U14583 (N_14583,N_14146,N_14163);
nor U14584 (N_14584,N_14489,N_14442);
nand U14585 (N_14585,N_14199,N_14113);
xor U14586 (N_14586,N_14263,N_14362);
xnor U14587 (N_14587,N_14226,N_14431);
xnor U14588 (N_14588,N_14225,N_14160);
nor U14589 (N_14589,N_14400,N_14074);
and U14590 (N_14590,N_14103,N_14202);
nand U14591 (N_14591,N_14444,N_14234);
nand U14592 (N_14592,N_14407,N_14219);
nor U14593 (N_14593,N_14468,N_14178);
nand U14594 (N_14594,N_14487,N_14349);
or U14595 (N_14595,N_14466,N_14374);
xnor U14596 (N_14596,N_14452,N_14158);
nor U14597 (N_14597,N_14492,N_14015);
nor U14598 (N_14598,N_14174,N_14301);
nor U14599 (N_14599,N_14311,N_14053);
and U14600 (N_14600,N_14424,N_14187);
nand U14601 (N_14601,N_14260,N_14361);
and U14602 (N_14602,N_14410,N_14352);
nor U14603 (N_14603,N_14116,N_14109);
and U14604 (N_14604,N_14465,N_14061);
nor U14605 (N_14605,N_14201,N_14164);
xnor U14606 (N_14606,N_14056,N_14089);
nor U14607 (N_14607,N_14173,N_14268);
nor U14608 (N_14608,N_14379,N_14027);
xnor U14609 (N_14609,N_14189,N_14250);
and U14610 (N_14610,N_14338,N_14460);
or U14611 (N_14611,N_14241,N_14406);
xnor U14612 (N_14612,N_14032,N_14224);
nand U14613 (N_14613,N_14414,N_14139);
or U14614 (N_14614,N_14204,N_14100);
and U14615 (N_14615,N_14484,N_14377);
or U14616 (N_14616,N_14264,N_14070);
nand U14617 (N_14617,N_14395,N_14332);
xnor U14618 (N_14618,N_14272,N_14000);
xor U14619 (N_14619,N_14023,N_14363);
or U14620 (N_14620,N_14267,N_14402);
nand U14621 (N_14621,N_14067,N_14081);
and U14622 (N_14622,N_14331,N_14088);
or U14623 (N_14623,N_14285,N_14316);
xnor U14624 (N_14624,N_14097,N_14221);
nor U14625 (N_14625,N_14227,N_14017);
and U14626 (N_14626,N_14366,N_14243);
or U14627 (N_14627,N_14474,N_14396);
and U14628 (N_14628,N_14135,N_14240);
nor U14629 (N_14629,N_14397,N_14281);
xnor U14630 (N_14630,N_14073,N_14269);
nand U14631 (N_14631,N_14341,N_14421);
nor U14632 (N_14632,N_14498,N_14323);
nand U14633 (N_14633,N_14141,N_14058);
nor U14634 (N_14634,N_14019,N_14009);
or U14635 (N_14635,N_14066,N_14403);
or U14636 (N_14636,N_14171,N_14215);
nor U14637 (N_14637,N_14370,N_14181);
or U14638 (N_14638,N_14014,N_14155);
nand U14639 (N_14639,N_14315,N_14083);
and U14640 (N_14640,N_14239,N_14493);
nand U14641 (N_14641,N_14449,N_14399);
xor U14642 (N_14642,N_14184,N_14191);
or U14643 (N_14643,N_14042,N_14196);
xnor U14644 (N_14644,N_14411,N_14209);
nand U14645 (N_14645,N_14445,N_14143);
nor U14646 (N_14646,N_14154,N_14499);
or U14647 (N_14647,N_14496,N_14401);
xor U14648 (N_14648,N_14475,N_14417);
nand U14649 (N_14649,N_14398,N_14270);
nor U14650 (N_14650,N_14222,N_14373);
nor U14651 (N_14651,N_14443,N_14180);
and U14652 (N_14652,N_14273,N_14040);
or U14653 (N_14653,N_14409,N_14255);
and U14654 (N_14654,N_14150,N_14383);
and U14655 (N_14655,N_14248,N_14216);
nor U14656 (N_14656,N_14018,N_14437);
xor U14657 (N_14657,N_14390,N_14320);
or U14658 (N_14658,N_14494,N_14028);
nor U14659 (N_14659,N_14394,N_14086);
nand U14660 (N_14660,N_14147,N_14309);
and U14661 (N_14661,N_14423,N_14415);
nor U14662 (N_14662,N_14378,N_14021);
nor U14663 (N_14663,N_14242,N_14111);
nor U14664 (N_14664,N_14286,N_14391);
xor U14665 (N_14665,N_14322,N_14405);
nor U14666 (N_14666,N_14034,N_14247);
xor U14667 (N_14667,N_14048,N_14051);
xnor U14668 (N_14668,N_14006,N_14353);
or U14669 (N_14669,N_14497,N_14016);
xnor U14670 (N_14670,N_14278,N_14128);
or U14671 (N_14671,N_14476,N_14430);
or U14672 (N_14672,N_14011,N_14080);
and U14673 (N_14673,N_14293,N_14223);
nand U14674 (N_14674,N_14127,N_14193);
nor U14675 (N_14675,N_14176,N_14208);
or U14676 (N_14676,N_14190,N_14043);
and U14677 (N_14677,N_14030,N_14436);
and U14678 (N_14678,N_14313,N_14351);
xnor U14679 (N_14679,N_14069,N_14244);
xor U14680 (N_14680,N_14207,N_14289);
or U14681 (N_14681,N_14464,N_14182);
or U14682 (N_14682,N_14159,N_14282);
xnor U14683 (N_14683,N_14157,N_14306);
xnor U14684 (N_14684,N_14261,N_14228);
or U14685 (N_14685,N_14149,N_14112);
xnor U14686 (N_14686,N_14138,N_14130);
xor U14687 (N_14687,N_14001,N_14479);
nand U14688 (N_14688,N_14416,N_14049);
xor U14689 (N_14689,N_14156,N_14457);
or U14690 (N_14690,N_14299,N_14037);
or U14691 (N_14691,N_14292,N_14140);
or U14692 (N_14692,N_14231,N_14392);
or U14693 (N_14693,N_14438,N_14298);
and U14694 (N_14694,N_14258,N_14336);
nor U14695 (N_14695,N_14307,N_14459);
xor U14696 (N_14696,N_14393,N_14003);
and U14697 (N_14697,N_14325,N_14254);
or U14698 (N_14698,N_14106,N_14233);
xor U14699 (N_14699,N_14271,N_14422);
and U14700 (N_14700,N_14031,N_14238);
nand U14701 (N_14701,N_14330,N_14114);
xor U14702 (N_14702,N_14280,N_14087);
nand U14703 (N_14703,N_14359,N_14082);
and U14704 (N_14704,N_14085,N_14418);
or U14705 (N_14705,N_14290,N_14205);
or U14706 (N_14706,N_14477,N_14488);
and U14707 (N_14707,N_14105,N_14046);
xnor U14708 (N_14708,N_14300,N_14090);
and U14709 (N_14709,N_14236,N_14044);
nor U14710 (N_14710,N_14230,N_14481);
xor U14711 (N_14711,N_14026,N_14217);
nor U14712 (N_14712,N_14450,N_14197);
or U14713 (N_14713,N_14054,N_14486);
or U14714 (N_14714,N_14453,N_14210);
nand U14715 (N_14715,N_14153,N_14206);
xor U14716 (N_14716,N_14432,N_14194);
or U14717 (N_14717,N_14075,N_14433);
and U14718 (N_14718,N_14068,N_14480);
nor U14719 (N_14719,N_14337,N_14369);
or U14720 (N_14720,N_14296,N_14446);
or U14721 (N_14721,N_14047,N_14132);
nand U14722 (N_14722,N_14372,N_14203);
nand U14723 (N_14723,N_14470,N_14120);
xnor U14724 (N_14724,N_14102,N_14439);
and U14725 (N_14725,N_14162,N_14310);
nor U14726 (N_14726,N_14055,N_14328);
or U14727 (N_14727,N_14126,N_14237);
or U14728 (N_14728,N_14471,N_14304);
nand U14729 (N_14729,N_14321,N_14107);
or U14730 (N_14730,N_14012,N_14455);
and U14731 (N_14731,N_14259,N_14435);
nand U14732 (N_14732,N_14447,N_14145);
or U14733 (N_14733,N_14144,N_14384);
xor U14734 (N_14734,N_14253,N_14072);
xnor U14735 (N_14735,N_14188,N_14387);
and U14736 (N_14736,N_14004,N_14093);
and U14737 (N_14737,N_14211,N_14462);
or U14738 (N_14738,N_14478,N_14381);
xnor U14739 (N_14739,N_14232,N_14052);
or U14740 (N_14740,N_14008,N_14490);
xor U14741 (N_14741,N_14214,N_14172);
and U14742 (N_14742,N_14413,N_14473);
nor U14743 (N_14743,N_14365,N_14375);
nor U14744 (N_14744,N_14288,N_14454);
xnor U14745 (N_14745,N_14124,N_14458);
nand U14746 (N_14746,N_14382,N_14022);
nor U14747 (N_14747,N_14334,N_14096);
and U14748 (N_14748,N_14368,N_14095);
or U14749 (N_14749,N_14319,N_14050);
and U14750 (N_14750,N_14354,N_14206);
nor U14751 (N_14751,N_14115,N_14162);
nor U14752 (N_14752,N_14442,N_14209);
or U14753 (N_14753,N_14011,N_14496);
nor U14754 (N_14754,N_14098,N_14203);
nor U14755 (N_14755,N_14399,N_14153);
xor U14756 (N_14756,N_14315,N_14011);
or U14757 (N_14757,N_14090,N_14403);
or U14758 (N_14758,N_14026,N_14025);
nor U14759 (N_14759,N_14051,N_14001);
xnor U14760 (N_14760,N_14229,N_14479);
and U14761 (N_14761,N_14306,N_14040);
and U14762 (N_14762,N_14150,N_14270);
xor U14763 (N_14763,N_14019,N_14482);
nand U14764 (N_14764,N_14366,N_14433);
and U14765 (N_14765,N_14010,N_14312);
or U14766 (N_14766,N_14387,N_14165);
xor U14767 (N_14767,N_14441,N_14332);
xnor U14768 (N_14768,N_14430,N_14358);
nor U14769 (N_14769,N_14145,N_14490);
or U14770 (N_14770,N_14317,N_14468);
nand U14771 (N_14771,N_14307,N_14148);
and U14772 (N_14772,N_14060,N_14023);
nand U14773 (N_14773,N_14195,N_14412);
nor U14774 (N_14774,N_14405,N_14153);
or U14775 (N_14775,N_14010,N_14163);
and U14776 (N_14776,N_14337,N_14120);
or U14777 (N_14777,N_14242,N_14308);
nor U14778 (N_14778,N_14223,N_14336);
or U14779 (N_14779,N_14364,N_14351);
and U14780 (N_14780,N_14067,N_14078);
and U14781 (N_14781,N_14298,N_14414);
and U14782 (N_14782,N_14185,N_14488);
nand U14783 (N_14783,N_14383,N_14242);
xnor U14784 (N_14784,N_14376,N_14296);
xor U14785 (N_14785,N_14110,N_14163);
xnor U14786 (N_14786,N_14461,N_14113);
nor U14787 (N_14787,N_14201,N_14334);
nor U14788 (N_14788,N_14152,N_14185);
xor U14789 (N_14789,N_14249,N_14212);
nor U14790 (N_14790,N_14418,N_14051);
and U14791 (N_14791,N_14186,N_14351);
nand U14792 (N_14792,N_14254,N_14467);
nor U14793 (N_14793,N_14066,N_14467);
and U14794 (N_14794,N_14051,N_14432);
xor U14795 (N_14795,N_14088,N_14043);
nand U14796 (N_14796,N_14469,N_14330);
nand U14797 (N_14797,N_14060,N_14196);
nand U14798 (N_14798,N_14436,N_14195);
xnor U14799 (N_14799,N_14158,N_14274);
or U14800 (N_14800,N_14468,N_14131);
or U14801 (N_14801,N_14001,N_14029);
nand U14802 (N_14802,N_14442,N_14122);
xor U14803 (N_14803,N_14086,N_14342);
and U14804 (N_14804,N_14484,N_14187);
and U14805 (N_14805,N_14244,N_14231);
or U14806 (N_14806,N_14419,N_14034);
and U14807 (N_14807,N_14301,N_14322);
or U14808 (N_14808,N_14261,N_14100);
nor U14809 (N_14809,N_14298,N_14464);
xnor U14810 (N_14810,N_14082,N_14067);
and U14811 (N_14811,N_14145,N_14032);
and U14812 (N_14812,N_14041,N_14355);
nand U14813 (N_14813,N_14354,N_14113);
and U14814 (N_14814,N_14272,N_14102);
nor U14815 (N_14815,N_14429,N_14059);
nand U14816 (N_14816,N_14467,N_14341);
and U14817 (N_14817,N_14400,N_14371);
nor U14818 (N_14818,N_14194,N_14341);
xor U14819 (N_14819,N_14425,N_14015);
nand U14820 (N_14820,N_14259,N_14343);
and U14821 (N_14821,N_14093,N_14115);
xnor U14822 (N_14822,N_14304,N_14455);
nand U14823 (N_14823,N_14288,N_14042);
and U14824 (N_14824,N_14288,N_14209);
nor U14825 (N_14825,N_14443,N_14102);
nor U14826 (N_14826,N_14338,N_14362);
nor U14827 (N_14827,N_14351,N_14334);
or U14828 (N_14828,N_14461,N_14181);
nand U14829 (N_14829,N_14045,N_14015);
and U14830 (N_14830,N_14452,N_14274);
xor U14831 (N_14831,N_14168,N_14394);
and U14832 (N_14832,N_14465,N_14020);
xor U14833 (N_14833,N_14058,N_14181);
nand U14834 (N_14834,N_14024,N_14207);
xnor U14835 (N_14835,N_14065,N_14352);
or U14836 (N_14836,N_14020,N_14316);
xor U14837 (N_14837,N_14071,N_14422);
xnor U14838 (N_14838,N_14393,N_14459);
or U14839 (N_14839,N_14493,N_14366);
and U14840 (N_14840,N_14416,N_14220);
and U14841 (N_14841,N_14185,N_14390);
nor U14842 (N_14842,N_14166,N_14037);
nor U14843 (N_14843,N_14144,N_14475);
or U14844 (N_14844,N_14497,N_14012);
or U14845 (N_14845,N_14362,N_14229);
or U14846 (N_14846,N_14175,N_14318);
xnor U14847 (N_14847,N_14043,N_14306);
nand U14848 (N_14848,N_14437,N_14220);
nor U14849 (N_14849,N_14441,N_14081);
nand U14850 (N_14850,N_14292,N_14037);
nor U14851 (N_14851,N_14318,N_14459);
xnor U14852 (N_14852,N_14224,N_14272);
nor U14853 (N_14853,N_14149,N_14456);
nand U14854 (N_14854,N_14333,N_14047);
xor U14855 (N_14855,N_14426,N_14409);
and U14856 (N_14856,N_14289,N_14153);
nor U14857 (N_14857,N_14218,N_14313);
nor U14858 (N_14858,N_14284,N_14253);
nand U14859 (N_14859,N_14281,N_14127);
nor U14860 (N_14860,N_14194,N_14307);
or U14861 (N_14861,N_14142,N_14040);
xor U14862 (N_14862,N_14022,N_14296);
or U14863 (N_14863,N_14495,N_14001);
or U14864 (N_14864,N_14017,N_14136);
nor U14865 (N_14865,N_14307,N_14300);
and U14866 (N_14866,N_14487,N_14016);
and U14867 (N_14867,N_14413,N_14094);
and U14868 (N_14868,N_14283,N_14235);
and U14869 (N_14869,N_14097,N_14472);
xnor U14870 (N_14870,N_14365,N_14064);
or U14871 (N_14871,N_14338,N_14340);
xnor U14872 (N_14872,N_14221,N_14176);
nor U14873 (N_14873,N_14371,N_14092);
xor U14874 (N_14874,N_14430,N_14235);
or U14875 (N_14875,N_14339,N_14318);
nor U14876 (N_14876,N_14035,N_14133);
nand U14877 (N_14877,N_14278,N_14086);
and U14878 (N_14878,N_14437,N_14181);
nor U14879 (N_14879,N_14090,N_14204);
nand U14880 (N_14880,N_14010,N_14362);
nor U14881 (N_14881,N_14255,N_14237);
nand U14882 (N_14882,N_14273,N_14447);
nor U14883 (N_14883,N_14256,N_14210);
or U14884 (N_14884,N_14309,N_14241);
or U14885 (N_14885,N_14144,N_14260);
or U14886 (N_14886,N_14477,N_14456);
or U14887 (N_14887,N_14190,N_14337);
and U14888 (N_14888,N_14180,N_14238);
xnor U14889 (N_14889,N_14247,N_14456);
or U14890 (N_14890,N_14126,N_14378);
nand U14891 (N_14891,N_14309,N_14230);
and U14892 (N_14892,N_14216,N_14250);
or U14893 (N_14893,N_14275,N_14053);
xor U14894 (N_14894,N_14444,N_14327);
and U14895 (N_14895,N_14402,N_14089);
nor U14896 (N_14896,N_14239,N_14322);
xor U14897 (N_14897,N_14058,N_14067);
nor U14898 (N_14898,N_14343,N_14351);
or U14899 (N_14899,N_14115,N_14281);
or U14900 (N_14900,N_14450,N_14460);
nand U14901 (N_14901,N_14139,N_14482);
nor U14902 (N_14902,N_14020,N_14042);
or U14903 (N_14903,N_14360,N_14452);
nand U14904 (N_14904,N_14250,N_14338);
xnor U14905 (N_14905,N_14490,N_14174);
and U14906 (N_14906,N_14170,N_14302);
and U14907 (N_14907,N_14368,N_14234);
nor U14908 (N_14908,N_14310,N_14495);
nor U14909 (N_14909,N_14294,N_14265);
xnor U14910 (N_14910,N_14316,N_14305);
nand U14911 (N_14911,N_14391,N_14261);
and U14912 (N_14912,N_14450,N_14280);
xor U14913 (N_14913,N_14136,N_14290);
and U14914 (N_14914,N_14391,N_14175);
xor U14915 (N_14915,N_14111,N_14247);
or U14916 (N_14916,N_14277,N_14106);
or U14917 (N_14917,N_14119,N_14452);
or U14918 (N_14918,N_14198,N_14019);
nand U14919 (N_14919,N_14096,N_14379);
nor U14920 (N_14920,N_14186,N_14289);
and U14921 (N_14921,N_14411,N_14319);
nand U14922 (N_14922,N_14108,N_14039);
or U14923 (N_14923,N_14055,N_14377);
and U14924 (N_14924,N_14400,N_14104);
or U14925 (N_14925,N_14175,N_14277);
or U14926 (N_14926,N_14262,N_14169);
and U14927 (N_14927,N_14394,N_14002);
or U14928 (N_14928,N_14129,N_14261);
xor U14929 (N_14929,N_14349,N_14068);
xnor U14930 (N_14930,N_14196,N_14032);
nor U14931 (N_14931,N_14416,N_14267);
nand U14932 (N_14932,N_14137,N_14293);
or U14933 (N_14933,N_14250,N_14442);
xnor U14934 (N_14934,N_14035,N_14088);
nand U14935 (N_14935,N_14191,N_14204);
and U14936 (N_14936,N_14321,N_14326);
and U14937 (N_14937,N_14436,N_14010);
or U14938 (N_14938,N_14045,N_14055);
nand U14939 (N_14939,N_14159,N_14091);
nor U14940 (N_14940,N_14066,N_14038);
nand U14941 (N_14941,N_14284,N_14063);
and U14942 (N_14942,N_14486,N_14068);
xnor U14943 (N_14943,N_14326,N_14128);
xnor U14944 (N_14944,N_14006,N_14013);
xnor U14945 (N_14945,N_14034,N_14255);
or U14946 (N_14946,N_14203,N_14076);
or U14947 (N_14947,N_14307,N_14112);
nor U14948 (N_14948,N_14035,N_14137);
xnor U14949 (N_14949,N_14015,N_14369);
nand U14950 (N_14950,N_14354,N_14428);
nand U14951 (N_14951,N_14370,N_14154);
xor U14952 (N_14952,N_14049,N_14220);
nand U14953 (N_14953,N_14235,N_14490);
or U14954 (N_14954,N_14042,N_14382);
nand U14955 (N_14955,N_14254,N_14438);
nand U14956 (N_14956,N_14004,N_14380);
nand U14957 (N_14957,N_14187,N_14420);
or U14958 (N_14958,N_14272,N_14009);
xnor U14959 (N_14959,N_14060,N_14352);
nor U14960 (N_14960,N_14133,N_14185);
or U14961 (N_14961,N_14203,N_14303);
or U14962 (N_14962,N_14209,N_14277);
nand U14963 (N_14963,N_14060,N_14030);
nor U14964 (N_14964,N_14400,N_14276);
or U14965 (N_14965,N_14055,N_14400);
or U14966 (N_14966,N_14308,N_14142);
nor U14967 (N_14967,N_14278,N_14487);
nand U14968 (N_14968,N_14035,N_14201);
nand U14969 (N_14969,N_14249,N_14175);
and U14970 (N_14970,N_14254,N_14346);
nand U14971 (N_14971,N_14080,N_14064);
nand U14972 (N_14972,N_14323,N_14359);
xor U14973 (N_14973,N_14422,N_14110);
and U14974 (N_14974,N_14321,N_14153);
or U14975 (N_14975,N_14383,N_14020);
xor U14976 (N_14976,N_14035,N_14320);
nor U14977 (N_14977,N_14282,N_14448);
or U14978 (N_14978,N_14472,N_14467);
xor U14979 (N_14979,N_14219,N_14015);
and U14980 (N_14980,N_14205,N_14185);
nand U14981 (N_14981,N_14399,N_14233);
or U14982 (N_14982,N_14195,N_14091);
nor U14983 (N_14983,N_14078,N_14441);
nor U14984 (N_14984,N_14494,N_14419);
xor U14985 (N_14985,N_14136,N_14022);
nor U14986 (N_14986,N_14098,N_14089);
nand U14987 (N_14987,N_14262,N_14186);
nor U14988 (N_14988,N_14009,N_14408);
and U14989 (N_14989,N_14198,N_14446);
nor U14990 (N_14990,N_14425,N_14256);
xnor U14991 (N_14991,N_14188,N_14480);
xnor U14992 (N_14992,N_14211,N_14281);
nor U14993 (N_14993,N_14013,N_14412);
nand U14994 (N_14994,N_14326,N_14487);
xor U14995 (N_14995,N_14307,N_14303);
nor U14996 (N_14996,N_14109,N_14391);
nor U14997 (N_14997,N_14126,N_14035);
nor U14998 (N_14998,N_14462,N_14217);
nand U14999 (N_14999,N_14189,N_14329);
or U15000 (N_15000,N_14718,N_14590);
nand U15001 (N_15001,N_14772,N_14706);
nand U15002 (N_15002,N_14974,N_14702);
nor U15003 (N_15003,N_14555,N_14569);
and U15004 (N_15004,N_14519,N_14707);
or U15005 (N_15005,N_14563,N_14808);
and U15006 (N_15006,N_14885,N_14870);
nor U15007 (N_15007,N_14814,N_14995);
nand U15008 (N_15008,N_14527,N_14534);
or U15009 (N_15009,N_14780,N_14861);
xor U15010 (N_15010,N_14990,N_14753);
xnor U15011 (N_15011,N_14533,N_14865);
xor U15012 (N_15012,N_14605,N_14608);
xor U15013 (N_15013,N_14757,N_14786);
nand U15014 (N_15014,N_14629,N_14970);
xor U15015 (N_15015,N_14602,N_14871);
xor U15016 (N_15016,N_14846,N_14604);
nand U15017 (N_15017,N_14679,N_14875);
and U15018 (N_15018,N_14804,N_14665);
and U15019 (N_15019,N_14614,N_14709);
xnor U15020 (N_15020,N_14637,N_14802);
or U15021 (N_15021,N_14963,N_14518);
and U15022 (N_15022,N_14984,N_14971);
and U15023 (N_15023,N_14944,N_14580);
nand U15024 (N_15024,N_14838,N_14742);
xnor U15025 (N_15025,N_14503,N_14728);
nand U15026 (N_15026,N_14909,N_14557);
xor U15027 (N_15027,N_14986,N_14594);
xnor U15028 (N_15028,N_14523,N_14920);
nor U15029 (N_15029,N_14953,N_14933);
or U15030 (N_15030,N_14685,N_14627);
nand U15031 (N_15031,N_14784,N_14715);
nand U15032 (N_15032,N_14847,N_14688);
and U15033 (N_15033,N_14811,N_14979);
nand U15034 (N_15034,N_14782,N_14731);
and U15035 (N_15035,N_14776,N_14897);
nor U15036 (N_15036,N_14734,N_14807);
xor U15037 (N_15037,N_14929,N_14854);
or U15038 (N_15038,N_14573,N_14544);
and U15039 (N_15039,N_14672,N_14740);
nand U15040 (N_15040,N_14789,N_14524);
nand U15041 (N_15041,N_14801,N_14714);
and U15042 (N_15042,N_14930,N_14531);
nor U15043 (N_15043,N_14769,N_14717);
nand U15044 (N_15044,N_14904,N_14556);
xnor U15045 (N_15045,N_14517,N_14975);
and U15046 (N_15046,N_14873,N_14547);
or U15047 (N_15047,N_14997,N_14673);
and U15048 (N_15048,N_14813,N_14546);
nor U15049 (N_15049,N_14908,N_14638);
xor U15050 (N_15050,N_14691,N_14586);
nor U15051 (N_15051,N_14856,N_14515);
or U15052 (N_15052,N_14831,N_14790);
nor U15053 (N_15053,N_14644,N_14643);
nor U15054 (N_15054,N_14570,N_14677);
nand U15055 (N_15055,N_14712,N_14658);
or U15056 (N_15056,N_14833,N_14919);
nand U15057 (N_15057,N_14800,N_14899);
nor U15058 (N_15058,N_14934,N_14835);
nor U15059 (N_15059,N_14987,N_14575);
nand U15060 (N_15060,N_14701,N_14616);
xor U15061 (N_15061,N_14922,N_14945);
xnor U15062 (N_15062,N_14678,N_14798);
and U15063 (N_15063,N_14656,N_14795);
nand U15064 (N_15064,N_14659,N_14724);
nor U15065 (N_15065,N_14585,N_14763);
xor U15066 (N_15066,N_14579,N_14628);
or U15067 (N_15067,N_14642,N_14552);
nand U15068 (N_15068,N_14852,N_14827);
or U15069 (N_15069,N_14821,N_14617);
or U15070 (N_15070,N_14771,N_14501);
xor U15071 (N_15071,N_14905,N_14635);
xor U15072 (N_15072,N_14747,N_14526);
and U15073 (N_15073,N_14752,N_14983);
and U15074 (N_15074,N_14777,N_14946);
and U15075 (N_15075,N_14924,N_14916);
nor U15076 (N_15076,N_14516,N_14948);
xnor U15077 (N_15077,N_14849,N_14826);
or U15078 (N_15078,N_14610,N_14957);
and U15079 (N_15079,N_14779,N_14887);
and U15080 (N_15080,N_14622,N_14834);
nand U15081 (N_15081,N_14906,N_14907);
nand U15082 (N_15082,N_14860,N_14620);
nor U15083 (N_15083,N_14660,N_14674);
or U15084 (N_15084,N_14538,N_14978);
nand U15085 (N_15085,N_14896,N_14976);
nor U15086 (N_15086,N_14537,N_14699);
and U15087 (N_15087,N_14964,N_14894);
xnor U15088 (N_15088,N_14525,N_14867);
or U15089 (N_15089,N_14554,N_14598);
or U15090 (N_15090,N_14650,N_14618);
nand U15091 (N_15091,N_14597,N_14545);
nor U15092 (N_15092,N_14609,N_14893);
or U15093 (N_15093,N_14912,N_14961);
and U15094 (N_15094,N_14773,N_14584);
xnor U15095 (N_15095,N_14695,N_14500);
nand U15096 (N_15096,N_14532,N_14631);
and U15097 (N_15097,N_14721,N_14550);
nor U15098 (N_15098,N_14915,N_14733);
nor U15099 (N_15099,N_14823,N_14993);
nor U15100 (N_15100,N_14596,N_14632);
xor U15101 (N_15101,N_14931,N_14536);
nor U15102 (N_15102,N_14935,N_14541);
or U15103 (N_15103,N_14704,N_14992);
or U15104 (N_15104,N_14938,N_14864);
xnor U15105 (N_15105,N_14874,N_14880);
and U15106 (N_15106,N_14589,N_14921);
nor U15107 (N_15107,N_14886,N_14535);
and U15108 (N_15108,N_14843,N_14566);
xnor U15109 (N_15109,N_14661,N_14850);
nor U15110 (N_15110,N_14510,N_14781);
xor U15111 (N_15111,N_14505,N_14741);
nand U15112 (N_15112,N_14509,N_14792);
or U15113 (N_15113,N_14810,N_14560);
and U15114 (N_15114,N_14900,N_14568);
or U15115 (N_15115,N_14895,N_14687);
nor U15116 (N_15116,N_14967,N_14954);
or U15117 (N_15117,N_14806,N_14889);
or U15118 (N_15118,N_14748,N_14891);
and U15119 (N_15119,N_14832,N_14882);
xnor U15120 (N_15120,N_14950,N_14996);
or U15121 (N_15121,N_14949,N_14751);
xnor U15122 (N_15122,N_14606,N_14947);
nand U15123 (N_15123,N_14540,N_14654);
nor U15124 (N_15124,N_14711,N_14825);
nand U15125 (N_15125,N_14514,N_14582);
nor U15126 (N_15126,N_14663,N_14567);
or U15127 (N_15127,N_14593,N_14793);
or U15128 (N_15128,N_14926,N_14778);
or U15129 (N_15129,N_14812,N_14743);
xor U15130 (N_15130,N_14574,N_14783);
nand U15131 (N_15131,N_14646,N_14888);
nor U15132 (N_15132,N_14937,N_14508);
and U15133 (N_15133,N_14700,N_14732);
nor U15134 (N_15134,N_14766,N_14543);
xnor U15135 (N_15135,N_14729,N_14991);
and U15136 (N_15136,N_14939,N_14840);
xor U15137 (N_15137,N_14667,N_14940);
or U15138 (N_15138,N_14710,N_14746);
xor U15139 (N_15139,N_14565,N_14866);
and U15140 (N_15140,N_14855,N_14841);
nor U15141 (N_15141,N_14858,N_14853);
nand U15142 (N_15142,N_14848,N_14819);
nor U15143 (N_15143,N_14966,N_14542);
xnor U15144 (N_15144,N_14977,N_14621);
and U15145 (N_15145,N_14839,N_14910);
or U15146 (N_15146,N_14951,N_14558);
and U15147 (N_15147,N_14881,N_14539);
nor U15148 (N_15148,N_14564,N_14581);
and U15149 (N_15149,N_14911,N_14863);
or U15150 (N_15150,N_14980,N_14682);
nor U15151 (N_15151,N_14805,N_14817);
or U15152 (N_15152,N_14928,N_14754);
xnor U15153 (N_15153,N_14969,N_14903);
xor U15154 (N_15154,N_14762,N_14859);
nor U15155 (N_15155,N_14836,N_14942);
and U15156 (N_15156,N_14681,N_14730);
or U15157 (N_15157,N_14723,N_14719);
nor U15158 (N_15158,N_14657,N_14703);
and U15159 (N_15159,N_14521,N_14561);
nor U15160 (N_15160,N_14818,N_14872);
and U15161 (N_15161,N_14630,N_14520);
and U15162 (N_15162,N_14932,N_14759);
xnor U15163 (N_15163,N_14998,N_14761);
xor U15164 (N_15164,N_14815,N_14739);
and U15165 (N_15165,N_14767,N_14645);
and U15166 (N_15166,N_14698,N_14973);
xnor U15167 (N_15167,N_14655,N_14612);
or U15168 (N_15168,N_14716,N_14744);
nor U15169 (N_15169,N_14883,N_14725);
or U15170 (N_15170,N_14830,N_14576);
or U15171 (N_15171,N_14670,N_14624);
and U15172 (N_15172,N_14512,N_14914);
nand U15173 (N_15173,N_14749,N_14962);
nand U15174 (N_15174,N_14756,N_14708);
nand U15175 (N_15175,N_14693,N_14528);
nor U15176 (N_15176,N_14513,N_14676);
nor U15177 (N_15177,N_14822,N_14694);
xnor U15178 (N_15178,N_14799,N_14797);
nand U15179 (N_15179,N_14738,N_14684);
nor U15180 (N_15180,N_14842,N_14634);
xnor U15181 (N_15181,N_14941,N_14879);
or U15182 (N_15182,N_14913,N_14619);
or U15183 (N_15183,N_14599,N_14760);
and U15184 (N_15184,N_14726,N_14690);
xnor U15185 (N_15185,N_14653,N_14648);
or U15186 (N_15186,N_14623,N_14775);
or U15187 (N_15187,N_14768,N_14958);
nor U15188 (N_15188,N_14803,N_14918);
xor U15189 (N_15189,N_14662,N_14960);
xnor U15190 (N_15190,N_14669,N_14943);
and U15191 (N_15191,N_14615,N_14705);
or U15192 (N_15192,N_14745,N_14588);
and U15193 (N_15193,N_14972,N_14549);
nor U15194 (N_15194,N_14595,N_14758);
xor U15195 (N_15195,N_14591,N_14868);
and U15196 (N_15196,N_14664,N_14816);
or U15197 (N_15197,N_14553,N_14529);
nand U15198 (N_15198,N_14857,N_14727);
xor U15199 (N_15199,N_14692,N_14956);
nand U15200 (N_15200,N_14828,N_14666);
and U15201 (N_15201,N_14869,N_14809);
nand U15202 (N_15202,N_14820,N_14844);
nor U15203 (N_15203,N_14876,N_14936);
and U15204 (N_15204,N_14583,N_14927);
xnor U15205 (N_15205,N_14720,N_14735);
nand U15206 (N_15206,N_14603,N_14671);
or U15207 (N_15207,N_14755,N_14994);
and U15208 (N_15208,N_14639,N_14901);
nand U15209 (N_15209,N_14686,N_14788);
nand U15210 (N_15210,N_14774,N_14737);
or U15211 (N_15211,N_14794,N_14504);
or U15212 (N_15212,N_14791,N_14592);
nor U15213 (N_15213,N_14765,N_14502);
and U15214 (N_15214,N_14633,N_14571);
xnor U15215 (N_15215,N_14925,N_14965);
or U15216 (N_15216,N_14988,N_14506);
nor U15217 (N_15217,N_14649,N_14507);
and U15218 (N_15218,N_14952,N_14985);
or U15219 (N_15219,N_14736,N_14917);
or U15220 (N_15220,N_14968,N_14625);
nor U15221 (N_15221,N_14764,N_14607);
and U15222 (N_15222,N_14522,N_14902);
nor U15223 (N_15223,N_14837,N_14551);
nor U15224 (N_15224,N_14548,N_14611);
nand U15225 (N_15225,N_14511,N_14878);
and U15226 (N_15226,N_14577,N_14884);
xor U15227 (N_15227,N_14578,N_14770);
nand U15228 (N_15228,N_14572,N_14923);
nand U15229 (N_15229,N_14982,N_14640);
xor U15230 (N_15230,N_14862,N_14668);
xor U15231 (N_15231,N_14829,N_14824);
xor U15232 (N_15232,N_14722,N_14999);
and U15233 (N_15233,N_14796,N_14636);
or U15234 (N_15234,N_14787,N_14562);
or U15235 (N_15235,N_14587,N_14559);
nor U15236 (N_15236,N_14981,N_14898);
nand U15237 (N_15237,N_14750,N_14601);
xor U15238 (N_15238,N_14959,N_14851);
xor U15239 (N_15239,N_14890,N_14641);
xor U15240 (N_15240,N_14713,N_14683);
xnor U15241 (N_15241,N_14845,N_14652);
nand U15242 (N_15242,N_14697,N_14785);
nand U15243 (N_15243,N_14651,N_14600);
or U15244 (N_15244,N_14892,N_14696);
or U15245 (N_15245,N_14675,N_14877);
nor U15246 (N_15246,N_14626,N_14680);
nor U15247 (N_15247,N_14689,N_14989);
xnor U15248 (N_15248,N_14955,N_14530);
and U15249 (N_15249,N_14647,N_14613);
nor U15250 (N_15250,N_14542,N_14907);
nor U15251 (N_15251,N_14981,N_14934);
nand U15252 (N_15252,N_14531,N_14634);
xor U15253 (N_15253,N_14718,N_14780);
or U15254 (N_15254,N_14507,N_14594);
nor U15255 (N_15255,N_14509,N_14736);
or U15256 (N_15256,N_14987,N_14578);
xor U15257 (N_15257,N_14733,N_14983);
nand U15258 (N_15258,N_14524,N_14625);
nor U15259 (N_15259,N_14528,N_14741);
nand U15260 (N_15260,N_14538,N_14560);
nor U15261 (N_15261,N_14619,N_14939);
nor U15262 (N_15262,N_14734,N_14607);
and U15263 (N_15263,N_14730,N_14657);
xnor U15264 (N_15264,N_14542,N_14820);
nor U15265 (N_15265,N_14605,N_14693);
and U15266 (N_15266,N_14569,N_14937);
nand U15267 (N_15267,N_14733,N_14777);
nand U15268 (N_15268,N_14925,N_14500);
and U15269 (N_15269,N_14518,N_14796);
and U15270 (N_15270,N_14727,N_14910);
or U15271 (N_15271,N_14680,N_14950);
xnor U15272 (N_15272,N_14866,N_14815);
nor U15273 (N_15273,N_14717,N_14910);
or U15274 (N_15274,N_14547,N_14554);
xnor U15275 (N_15275,N_14705,N_14777);
xnor U15276 (N_15276,N_14720,N_14973);
nor U15277 (N_15277,N_14673,N_14963);
nand U15278 (N_15278,N_14908,N_14600);
nand U15279 (N_15279,N_14607,N_14577);
nand U15280 (N_15280,N_14657,N_14529);
or U15281 (N_15281,N_14519,N_14868);
xnor U15282 (N_15282,N_14646,N_14988);
nor U15283 (N_15283,N_14555,N_14812);
or U15284 (N_15284,N_14776,N_14668);
or U15285 (N_15285,N_14926,N_14893);
nand U15286 (N_15286,N_14824,N_14896);
and U15287 (N_15287,N_14720,N_14897);
or U15288 (N_15288,N_14757,N_14686);
or U15289 (N_15289,N_14825,N_14681);
and U15290 (N_15290,N_14589,N_14798);
or U15291 (N_15291,N_14930,N_14634);
and U15292 (N_15292,N_14668,N_14731);
or U15293 (N_15293,N_14861,N_14836);
nor U15294 (N_15294,N_14903,N_14725);
or U15295 (N_15295,N_14543,N_14933);
or U15296 (N_15296,N_14777,N_14698);
xnor U15297 (N_15297,N_14892,N_14705);
and U15298 (N_15298,N_14961,N_14830);
or U15299 (N_15299,N_14845,N_14550);
xnor U15300 (N_15300,N_14741,N_14814);
nor U15301 (N_15301,N_14894,N_14881);
xor U15302 (N_15302,N_14536,N_14967);
nand U15303 (N_15303,N_14704,N_14741);
or U15304 (N_15304,N_14845,N_14617);
and U15305 (N_15305,N_14976,N_14813);
xnor U15306 (N_15306,N_14984,N_14918);
xor U15307 (N_15307,N_14910,N_14943);
and U15308 (N_15308,N_14929,N_14732);
nand U15309 (N_15309,N_14691,N_14551);
and U15310 (N_15310,N_14734,N_14510);
or U15311 (N_15311,N_14814,N_14878);
nand U15312 (N_15312,N_14990,N_14989);
nand U15313 (N_15313,N_14717,N_14852);
or U15314 (N_15314,N_14772,N_14982);
and U15315 (N_15315,N_14507,N_14756);
xnor U15316 (N_15316,N_14560,N_14946);
and U15317 (N_15317,N_14519,N_14736);
or U15318 (N_15318,N_14715,N_14891);
or U15319 (N_15319,N_14923,N_14505);
nand U15320 (N_15320,N_14910,N_14754);
xnor U15321 (N_15321,N_14692,N_14544);
xnor U15322 (N_15322,N_14833,N_14892);
nor U15323 (N_15323,N_14640,N_14902);
and U15324 (N_15324,N_14730,N_14509);
xnor U15325 (N_15325,N_14689,N_14636);
xor U15326 (N_15326,N_14762,N_14577);
or U15327 (N_15327,N_14890,N_14849);
nand U15328 (N_15328,N_14572,N_14714);
or U15329 (N_15329,N_14614,N_14923);
nand U15330 (N_15330,N_14659,N_14518);
or U15331 (N_15331,N_14885,N_14670);
and U15332 (N_15332,N_14642,N_14637);
nand U15333 (N_15333,N_14822,N_14795);
and U15334 (N_15334,N_14521,N_14736);
nand U15335 (N_15335,N_14680,N_14989);
xor U15336 (N_15336,N_14946,N_14666);
xnor U15337 (N_15337,N_14579,N_14923);
or U15338 (N_15338,N_14955,N_14502);
or U15339 (N_15339,N_14625,N_14559);
and U15340 (N_15340,N_14563,N_14920);
nand U15341 (N_15341,N_14574,N_14674);
nand U15342 (N_15342,N_14958,N_14881);
nor U15343 (N_15343,N_14613,N_14984);
nand U15344 (N_15344,N_14957,N_14896);
nand U15345 (N_15345,N_14870,N_14719);
xnor U15346 (N_15346,N_14803,N_14783);
nor U15347 (N_15347,N_14813,N_14547);
nor U15348 (N_15348,N_14672,N_14957);
xor U15349 (N_15349,N_14551,N_14847);
nand U15350 (N_15350,N_14817,N_14511);
or U15351 (N_15351,N_14530,N_14753);
xnor U15352 (N_15352,N_14858,N_14712);
xnor U15353 (N_15353,N_14945,N_14594);
nor U15354 (N_15354,N_14522,N_14735);
and U15355 (N_15355,N_14945,N_14999);
nand U15356 (N_15356,N_14811,N_14789);
nor U15357 (N_15357,N_14875,N_14576);
xor U15358 (N_15358,N_14950,N_14808);
or U15359 (N_15359,N_14612,N_14816);
nand U15360 (N_15360,N_14716,N_14726);
or U15361 (N_15361,N_14924,N_14968);
xnor U15362 (N_15362,N_14752,N_14877);
xnor U15363 (N_15363,N_14578,N_14843);
nand U15364 (N_15364,N_14825,N_14635);
and U15365 (N_15365,N_14877,N_14985);
nor U15366 (N_15366,N_14707,N_14591);
nor U15367 (N_15367,N_14872,N_14617);
nand U15368 (N_15368,N_14633,N_14570);
xor U15369 (N_15369,N_14998,N_14692);
nand U15370 (N_15370,N_14546,N_14862);
and U15371 (N_15371,N_14745,N_14551);
or U15372 (N_15372,N_14580,N_14689);
or U15373 (N_15373,N_14738,N_14831);
and U15374 (N_15374,N_14521,N_14560);
nor U15375 (N_15375,N_14693,N_14760);
nand U15376 (N_15376,N_14633,N_14949);
and U15377 (N_15377,N_14670,N_14571);
and U15378 (N_15378,N_14847,N_14955);
xnor U15379 (N_15379,N_14864,N_14577);
nor U15380 (N_15380,N_14856,N_14774);
and U15381 (N_15381,N_14783,N_14615);
nand U15382 (N_15382,N_14931,N_14738);
and U15383 (N_15383,N_14666,N_14824);
nand U15384 (N_15384,N_14919,N_14716);
nor U15385 (N_15385,N_14866,N_14982);
xor U15386 (N_15386,N_14500,N_14952);
nand U15387 (N_15387,N_14753,N_14888);
xnor U15388 (N_15388,N_14588,N_14865);
xor U15389 (N_15389,N_14887,N_14900);
and U15390 (N_15390,N_14845,N_14781);
nor U15391 (N_15391,N_14781,N_14613);
and U15392 (N_15392,N_14909,N_14713);
nand U15393 (N_15393,N_14811,N_14985);
nor U15394 (N_15394,N_14995,N_14985);
and U15395 (N_15395,N_14670,N_14788);
nand U15396 (N_15396,N_14575,N_14816);
xor U15397 (N_15397,N_14653,N_14791);
or U15398 (N_15398,N_14799,N_14935);
or U15399 (N_15399,N_14837,N_14504);
nor U15400 (N_15400,N_14889,N_14737);
nor U15401 (N_15401,N_14870,N_14791);
xnor U15402 (N_15402,N_14689,N_14598);
nand U15403 (N_15403,N_14511,N_14619);
nand U15404 (N_15404,N_14727,N_14577);
and U15405 (N_15405,N_14867,N_14537);
nor U15406 (N_15406,N_14979,N_14807);
nor U15407 (N_15407,N_14654,N_14843);
nand U15408 (N_15408,N_14904,N_14769);
nand U15409 (N_15409,N_14880,N_14604);
nor U15410 (N_15410,N_14646,N_14890);
or U15411 (N_15411,N_14720,N_14779);
nand U15412 (N_15412,N_14679,N_14654);
xnor U15413 (N_15413,N_14887,N_14838);
xor U15414 (N_15414,N_14710,N_14655);
and U15415 (N_15415,N_14811,N_14761);
or U15416 (N_15416,N_14644,N_14632);
and U15417 (N_15417,N_14609,N_14879);
xor U15418 (N_15418,N_14948,N_14933);
and U15419 (N_15419,N_14925,N_14666);
and U15420 (N_15420,N_14930,N_14501);
and U15421 (N_15421,N_14562,N_14832);
and U15422 (N_15422,N_14919,N_14845);
nand U15423 (N_15423,N_14796,N_14526);
or U15424 (N_15424,N_14672,N_14983);
nor U15425 (N_15425,N_14728,N_14501);
and U15426 (N_15426,N_14744,N_14940);
xor U15427 (N_15427,N_14629,N_14962);
xnor U15428 (N_15428,N_14514,N_14852);
or U15429 (N_15429,N_14906,N_14545);
xor U15430 (N_15430,N_14593,N_14625);
nand U15431 (N_15431,N_14871,N_14837);
nor U15432 (N_15432,N_14773,N_14532);
xor U15433 (N_15433,N_14986,N_14708);
nand U15434 (N_15434,N_14962,N_14570);
nand U15435 (N_15435,N_14661,N_14609);
and U15436 (N_15436,N_14857,N_14594);
or U15437 (N_15437,N_14918,N_14582);
and U15438 (N_15438,N_14898,N_14913);
nor U15439 (N_15439,N_14662,N_14861);
nor U15440 (N_15440,N_14687,N_14984);
nand U15441 (N_15441,N_14750,N_14843);
nand U15442 (N_15442,N_14743,N_14909);
or U15443 (N_15443,N_14544,N_14567);
or U15444 (N_15444,N_14655,N_14630);
xor U15445 (N_15445,N_14502,N_14906);
and U15446 (N_15446,N_14527,N_14831);
xor U15447 (N_15447,N_14717,N_14728);
or U15448 (N_15448,N_14918,N_14500);
nor U15449 (N_15449,N_14768,N_14788);
nand U15450 (N_15450,N_14647,N_14600);
nor U15451 (N_15451,N_14767,N_14779);
or U15452 (N_15452,N_14809,N_14854);
or U15453 (N_15453,N_14611,N_14680);
xnor U15454 (N_15454,N_14942,N_14920);
xor U15455 (N_15455,N_14924,N_14950);
xnor U15456 (N_15456,N_14726,N_14919);
nand U15457 (N_15457,N_14763,N_14989);
and U15458 (N_15458,N_14552,N_14806);
and U15459 (N_15459,N_14906,N_14558);
nand U15460 (N_15460,N_14552,N_14759);
nand U15461 (N_15461,N_14954,N_14833);
and U15462 (N_15462,N_14527,N_14772);
or U15463 (N_15463,N_14745,N_14765);
xnor U15464 (N_15464,N_14992,N_14841);
nand U15465 (N_15465,N_14531,N_14991);
or U15466 (N_15466,N_14778,N_14966);
nand U15467 (N_15467,N_14624,N_14575);
xor U15468 (N_15468,N_14943,N_14889);
or U15469 (N_15469,N_14843,N_14777);
xor U15470 (N_15470,N_14588,N_14527);
and U15471 (N_15471,N_14572,N_14762);
nor U15472 (N_15472,N_14633,N_14867);
and U15473 (N_15473,N_14905,N_14654);
and U15474 (N_15474,N_14634,N_14795);
and U15475 (N_15475,N_14893,N_14788);
or U15476 (N_15476,N_14559,N_14868);
nor U15477 (N_15477,N_14910,N_14680);
and U15478 (N_15478,N_14698,N_14655);
xor U15479 (N_15479,N_14651,N_14841);
xnor U15480 (N_15480,N_14795,N_14798);
or U15481 (N_15481,N_14809,N_14882);
nand U15482 (N_15482,N_14818,N_14765);
and U15483 (N_15483,N_14567,N_14757);
nor U15484 (N_15484,N_14508,N_14590);
and U15485 (N_15485,N_14796,N_14578);
or U15486 (N_15486,N_14578,N_14933);
nor U15487 (N_15487,N_14765,N_14573);
and U15488 (N_15488,N_14570,N_14675);
and U15489 (N_15489,N_14745,N_14859);
and U15490 (N_15490,N_14581,N_14990);
or U15491 (N_15491,N_14669,N_14966);
nor U15492 (N_15492,N_14914,N_14849);
xnor U15493 (N_15493,N_14759,N_14845);
or U15494 (N_15494,N_14931,N_14599);
xnor U15495 (N_15495,N_14973,N_14968);
nor U15496 (N_15496,N_14694,N_14518);
xnor U15497 (N_15497,N_14745,N_14779);
nor U15498 (N_15498,N_14710,N_14941);
or U15499 (N_15499,N_14519,N_14827);
nor U15500 (N_15500,N_15178,N_15064);
or U15501 (N_15501,N_15108,N_15391);
or U15502 (N_15502,N_15125,N_15021);
nor U15503 (N_15503,N_15033,N_15310);
or U15504 (N_15504,N_15198,N_15373);
or U15505 (N_15505,N_15397,N_15182);
nand U15506 (N_15506,N_15496,N_15118);
xor U15507 (N_15507,N_15499,N_15435);
nor U15508 (N_15508,N_15038,N_15274);
or U15509 (N_15509,N_15461,N_15066);
xor U15510 (N_15510,N_15112,N_15234);
nand U15511 (N_15511,N_15138,N_15255);
nor U15512 (N_15512,N_15277,N_15464);
and U15513 (N_15513,N_15074,N_15212);
nor U15514 (N_15514,N_15290,N_15229);
xor U15515 (N_15515,N_15406,N_15478);
nand U15516 (N_15516,N_15437,N_15413);
and U15517 (N_15517,N_15246,N_15408);
and U15518 (N_15518,N_15150,N_15367);
xor U15519 (N_15519,N_15484,N_15339);
xnor U15520 (N_15520,N_15011,N_15265);
nand U15521 (N_15521,N_15051,N_15284);
and U15522 (N_15522,N_15134,N_15090);
nand U15523 (N_15523,N_15026,N_15126);
and U15524 (N_15524,N_15457,N_15318);
nand U15525 (N_15525,N_15216,N_15482);
or U15526 (N_15526,N_15106,N_15231);
or U15527 (N_15527,N_15470,N_15130);
or U15528 (N_15528,N_15189,N_15131);
nor U15529 (N_15529,N_15202,N_15114);
nor U15530 (N_15530,N_15084,N_15225);
nor U15531 (N_15531,N_15077,N_15195);
and U15532 (N_15532,N_15151,N_15230);
nor U15533 (N_15533,N_15203,N_15096);
and U15534 (N_15534,N_15219,N_15013);
or U15535 (N_15535,N_15376,N_15141);
nand U15536 (N_15536,N_15241,N_15043);
xor U15537 (N_15537,N_15271,N_15117);
xnor U15538 (N_15538,N_15083,N_15172);
or U15539 (N_15539,N_15379,N_15440);
nand U15540 (N_15540,N_15162,N_15489);
xor U15541 (N_15541,N_15344,N_15049);
and U15542 (N_15542,N_15208,N_15433);
nor U15543 (N_15543,N_15067,N_15065);
nand U15544 (N_15544,N_15341,N_15334);
nor U15545 (N_15545,N_15307,N_15417);
and U15546 (N_15546,N_15314,N_15005);
nor U15547 (N_15547,N_15153,N_15110);
xnor U15548 (N_15548,N_15159,N_15034);
and U15549 (N_15549,N_15010,N_15474);
nand U15550 (N_15550,N_15115,N_15177);
or U15551 (N_15551,N_15263,N_15302);
and U15552 (N_15552,N_15031,N_15042);
nand U15553 (N_15553,N_15393,N_15317);
and U15554 (N_15554,N_15381,N_15235);
or U15555 (N_15555,N_15335,N_15168);
nor U15556 (N_15556,N_15135,N_15346);
xnor U15557 (N_15557,N_15097,N_15261);
nand U15558 (N_15558,N_15188,N_15295);
xnor U15559 (N_15559,N_15256,N_15259);
and U15560 (N_15560,N_15293,N_15094);
or U15561 (N_15561,N_15415,N_15392);
xor U15562 (N_15562,N_15477,N_15194);
or U15563 (N_15563,N_15137,N_15384);
nand U15564 (N_15564,N_15213,N_15401);
nor U15565 (N_15565,N_15060,N_15411);
nor U15566 (N_15566,N_15000,N_15347);
nor U15567 (N_15567,N_15087,N_15113);
nand U15568 (N_15568,N_15073,N_15220);
xor U15569 (N_15569,N_15398,N_15123);
nand U15570 (N_15570,N_15364,N_15396);
or U15571 (N_15571,N_15463,N_15248);
nor U15572 (N_15572,N_15244,N_15175);
or U15573 (N_15573,N_15306,N_15085);
xor U15574 (N_15574,N_15047,N_15018);
xor U15575 (N_15575,N_15210,N_15345);
or U15576 (N_15576,N_15350,N_15154);
nor U15577 (N_15577,N_15360,N_15405);
nand U15578 (N_15578,N_15163,N_15080);
and U15579 (N_15579,N_15170,N_15395);
xor U15580 (N_15580,N_15236,N_15326);
or U15581 (N_15581,N_15322,N_15429);
or U15582 (N_15582,N_15497,N_15289);
nor U15583 (N_15583,N_15127,N_15380);
nor U15584 (N_15584,N_15280,N_15491);
or U15585 (N_15585,N_15253,N_15467);
or U15586 (N_15586,N_15129,N_15264);
and U15587 (N_15587,N_15423,N_15100);
nand U15588 (N_15588,N_15340,N_15283);
nand U15589 (N_15589,N_15431,N_15057);
nand U15590 (N_15590,N_15351,N_15173);
and U15591 (N_15591,N_15382,N_15328);
xor U15592 (N_15592,N_15040,N_15358);
or U15593 (N_15593,N_15363,N_15139);
nor U15594 (N_15594,N_15069,N_15086);
nand U15595 (N_15595,N_15451,N_15362);
and U15596 (N_15596,N_15458,N_15032);
or U15597 (N_15597,N_15309,N_15070);
nand U15598 (N_15598,N_15399,N_15389);
nand U15599 (N_15599,N_15015,N_15166);
xnor U15600 (N_15600,N_15472,N_15352);
and U15601 (N_15601,N_15121,N_15357);
xor U15602 (N_15602,N_15479,N_15494);
xor U15603 (N_15603,N_15454,N_15174);
nand U15604 (N_15604,N_15483,N_15098);
and U15605 (N_15605,N_15120,N_15331);
and U15606 (N_15606,N_15157,N_15002);
xor U15607 (N_15607,N_15407,N_15250);
or U15608 (N_15608,N_15209,N_15095);
xor U15609 (N_15609,N_15416,N_15387);
and U15610 (N_15610,N_15238,N_15281);
and U15611 (N_15611,N_15003,N_15204);
xor U15612 (N_15612,N_15019,N_15372);
nor U15613 (N_15613,N_15434,N_15430);
and U15614 (N_15614,N_15428,N_15036);
xnor U15615 (N_15615,N_15354,N_15320);
xor U15616 (N_15616,N_15426,N_15254);
or U15617 (N_15617,N_15155,N_15240);
nand U15618 (N_15618,N_15388,N_15185);
nor U15619 (N_15619,N_15432,N_15409);
or U15620 (N_15620,N_15303,N_15124);
nor U15621 (N_15621,N_15349,N_15298);
nand U15622 (N_15622,N_15232,N_15245);
xor U15623 (N_15623,N_15315,N_15498);
nand U15624 (N_15624,N_15152,N_15279);
or U15625 (N_15625,N_15156,N_15160);
xnor U15626 (N_15626,N_15378,N_15128);
nand U15627 (N_15627,N_15319,N_15275);
xor U15628 (N_15628,N_15308,N_15476);
nor U15629 (N_15629,N_15329,N_15390);
nand U15630 (N_15630,N_15111,N_15148);
xor U15631 (N_15631,N_15471,N_15348);
xnor U15632 (N_15632,N_15427,N_15078);
xor U15633 (N_15633,N_15055,N_15361);
nand U15634 (N_15634,N_15022,N_15400);
nand U15635 (N_15635,N_15207,N_15278);
or U15636 (N_15636,N_15375,N_15059);
xnor U15637 (N_15637,N_15251,N_15233);
nor U15638 (N_15638,N_15054,N_15495);
xnor U15639 (N_15639,N_15455,N_15422);
nor U15640 (N_15640,N_15146,N_15030);
xnor U15641 (N_15641,N_15099,N_15468);
and U15642 (N_15642,N_15136,N_15014);
or U15643 (N_15643,N_15191,N_15368);
nand U15644 (N_15644,N_15291,N_15149);
xnor U15645 (N_15645,N_15052,N_15039);
or U15646 (N_15646,N_15205,N_15460);
nor U15647 (N_15647,N_15420,N_15325);
or U15648 (N_15648,N_15243,N_15488);
nand U15649 (N_15649,N_15142,N_15321);
xor U15650 (N_15650,N_15075,N_15029);
nor U15651 (N_15651,N_15092,N_15201);
nor U15652 (N_15652,N_15176,N_15404);
nor U15653 (N_15653,N_15490,N_15300);
nor U15654 (N_15654,N_15342,N_15072);
nand U15655 (N_15655,N_15273,N_15020);
and U15656 (N_15656,N_15343,N_15403);
or U15657 (N_15657,N_15260,N_15025);
xnor U15658 (N_15658,N_15140,N_15359);
xor U15659 (N_15659,N_15053,N_15383);
and U15660 (N_15660,N_15266,N_15410);
or U15661 (N_15661,N_15105,N_15184);
and U15662 (N_15662,N_15007,N_15103);
nor U15663 (N_15663,N_15102,N_15257);
nand U15664 (N_15664,N_15439,N_15324);
and U15665 (N_15665,N_15061,N_15171);
xor U15666 (N_15666,N_15267,N_15164);
and U15667 (N_15667,N_15370,N_15045);
xnor U15668 (N_15668,N_15414,N_15436);
and U15669 (N_15669,N_15145,N_15465);
xor U15670 (N_15670,N_15167,N_15028);
xnor U15671 (N_15671,N_15452,N_15487);
nor U15672 (N_15672,N_15187,N_15402);
and U15673 (N_15673,N_15356,N_15093);
and U15674 (N_15674,N_15200,N_15023);
nor U15675 (N_15675,N_15050,N_15247);
and U15676 (N_15676,N_15444,N_15056);
nor U15677 (N_15677,N_15355,N_15425);
nor U15678 (N_15678,N_15206,N_15285);
nand U15679 (N_15679,N_15089,N_15294);
xor U15680 (N_15680,N_15377,N_15268);
or U15681 (N_15681,N_15332,N_15012);
xnor U15682 (N_15682,N_15492,N_15104);
nor U15683 (N_15683,N_15453,N_15211);
nor U15684 (N_15684,N_15116,N_15443);
and U15685 (N_15685,N_15469,N_15386);
or U15686 (N_15686,N_15282,N_15249);
nand U15687 (N_15687,N_15486,N_15299);
xor U15688 (N_15688,N_15296,N_15223);
and U15689 (N_15689,N_15199,N_15009);
nor U15690 (N_15690,N_15165,N_15044);
xnor U15691 (N_15691,N_15224,N_15197);
nor U15692 (N_15692,N_15161,N_15237);
or U15693 (N_15693,N_15001,N_15107);
nor U15694 (N_15694,N_15221,N_15071);
nand U15695 (N_15695,N_15101,N_15186);
or U15696 (N_15696,N_15217,N_15081);
nor U15697 (N_15697,N_15466,N_15313);
nand U15698 (N_15698,N_15462,N_15035);
xnor U15699 (N_15699,N_15369,N_15133);
and U15700 (N_15700,N_15017,N_15258);
and U15701 (N_15701,N_15196,N_15447);
xnor U15702 (N_15702,N_15180,N_15063);
or U15703 (N_15703,N_15330,N_15424);
and U15704 (N_15704,N_15024,N_15132);
and U15705 (N_15705,N_15048,N_15305);
xor U15706 (N_15706,N_15008,N_15493);
or U15707 (N_15707,N_15158,N_15288);
nand U15708 (N_15708,N_15179,N_15336);
and U15709 (N_15709,N_15448,N_15269);
and U15710 (N_15710,N_15252,N_15169);
and U15711 (N_15711,N_15006,N_15181);
nor U15712 (N_15712,N_15337,N_15016);
xor U15713 (N_15713,N_15475,N_15192);
nor U15714 (N_15714,N_15365,N_15473);
nand U15715 (N_15715,N_15449,N_15147);
or U15716 (N_15716,N_15333,N_15286);
nor U15717 (N_15717,N_15144,N_15076);
or U15718 (N_15718,N_15027,N_15218);
or U15719 (N_15719,N_15366,N_15292);
and U15720 (N_15720,N_15394,N_15419);
nor U15721 (N_15721,N_15323,N_15371);
and U15722 (N_15722,N_15190,N_15304);
xor U15723 (N_15723,N_15480,N_15215);
xnor U15724 (N_15724,N_15004,N_15421);
nor U15725 (N_15725,N_15270,N_15459);
nand U15726 (N_15726,N_15262,N_15214);
xnor U15727 (N_15727,N_15119,N_15046);
and U15728 (N_15728,N_15438,N_15485);
or U15729 (N_15729,N_15418,N_15088);
and U15730 (N_15730,N_15228,N_15338);
xnor U15731 (N_15731,N_15327,N_15412);
and U15732 (N_15732,N_15297,N_15442);
or U15733 (N_15733,N_15082,N_15276);
xor U15734 (N_15734,N_15079,N_15450);
nor U15735 (N_15735,N_15109,N_15239);
nor U15736 (N_15736,N_15353,N_15287);
nor U15737 (N_15737,N_15068,N_15374);
nor U15738 (N_15738,N_15441,N_15062);
nor U15739 (N_15739,N_15446,N_15311);
nand U15740 (N_15740,N_15272,N_15301);
nor U15741 (N_15741,N_15041,N_15226);
nand U15742 (N_15742,N_15385,N_15456);
nor U15743 (N_15743,N_15037,N_15193);
nor U15744 (N_15744,N_15312,N_15222);
nand U15745 (N_15745,N_15058,N_15091);
and U15746 (N_15746,N_15122,N_15242);
xnor U15747 (N_15747,N_15227,N_15143);
nand U15748 (N_15748,N_15183,N_15481);
and U15749 (N_15749,N_15445,N_15316);
and U15750 (N_15750,N_15006,N_15419);
or U15751 (N_15751,N_15170,N_15463);
xor U15752 (N_15752,N_15392,N_15206);
xnor U15753 (N_15753,N_15295,N_15331);
or U15754 (N_15754,N_15183,N_15164);
or U15755 (N_15755,N_15287,N_15037);
or U15756 (N_15756,N_15253,N_15489);
xnor U15757 (N_15757,N_15229,N_15342);
nor U15758 (N_15758,N_15187,N_15026);
and U15759 (N_15759,N_15138,N_15306);
and U15760 (N_15760,N_15272,N_15378);
and U15761 (N_15761,N_15330,N_15327);
and U15762 (N_15762,N_15013,N_15256);
or U15763 (N_15763,N_15329,N_15228);
or U15764 (N_15764,N_15225,N_15249);
xor U15765 (N_15765,N_15053,N_15002);
and U15766 (N_15766,N_15042,N_15371);
xor U15767 (N_15767,N_15378,N_15309);
nor U15768 (N_15768,N_15254,N_15198);
nand U15769 (N_15769,N_15121,N_15313);
xor U15770 (N_15770,N_15227,N_15075);
or U15771 (N_15771,N_15294,N_15034);
nor U15772 (N_15772,N_15154,N_15224);
nor U15773 (N_15773,N_15260,N_15301);
nand U15774 (N_15774,N_15422,N_15354);
nand U15775 (N_15775,N_15421,N_15139);
nand U15776 (N_15776,N_15093,N_15126);
nand U15777 (N_15777,N_15117,N_15237);
or U15778 (N_15778,N_15130,N_15076);
nor U15779 (N_15779,N_15332,N_15111);
xor U15780 (N_15780,N_15049,N_15083);
or U15781 (N_15781,N_15396,N_15262);
nor U15782 (N_15782,N_15211,N_15499);
nand U15783 (N_15783,N_15207,N_15001);
or U15784 (N_15784,N_15186,N_15225);
or U15785 (N_15785,N_15092,N_15030);
nor U15786 (N_15786,N_15493,N_15145);
or U15787 (N_15787,N_15402,N_15274);
nand U15788 (N_15788,N_15330,N_15204);
and U15789 (N_15789,N_15485,N_15487);
nor U15790 (N_15790,N_15321,N_15145);
nor U15791 (N_15791,N_15322,N_15117);
nand U15792 (N_15792,N_15005,N_15254);
nor U15793 (N_15793,N_15026,N_15390);
nand U15794 (N_15794,N_15142,N_15044);
and U15795 (N_15795,N_15138,N_15473);
xor U15796 (N_15796,N_15304,N_15383);
nor U15797 (N_15797,N_15005,N_15430);
xor U15798 (N_15798,N_15003,N_15290);
and U15799 (N_15799,N_15417,N_15141);
nand U15800 (N_15800,N_15483,N_15484);
xnor U15801 (N_15801,N_15011,N_15395);
or U15802 (N_15802,N_15389,N_15346);
nand U15803 (N_15803,N_15251,N_15446);
nand U15804 (N_15804,N_15137,N_15390);
xnor U15805 (N_15805,N_15045,N_15049);
xor U15806 (N_15806,N_15451,N_15452);
xnor U15807 (N_15807,N_15187,N_15443);
nand U15808 (N_15808,N_15060,N_15320);
nand U15809 (N_15809,N_15222,N_15109);
xnor U15810 (N_15810,N_15445,N_15034);
xor U15811 (N_15811,N_15101,N_15117);
nor U15812 (N_15812,N_15333,N_15150);
nor U15813 (N_15813,N_15015,N_15423);
or U15814 (N_15814,N_15418,N_15040);
or U15815 (N_15815,N_15456,N_15163);
nor U15816 (N_15816,N_15102,N_15099);
nor U15817 (N_15817,N_15416,N_15449);
or U15818 (N_15818,N_15222,N_15330);
and U15819 (N_15819,N_15296,N_15117);
xor U15820 (N_15820,N_15104,N_15059);
and U15821 (N_15821,N_15162,N_15023);
and U15822 (N_15822,N_15390,N_15192);
or U15823 (N_15823,N_15306,N_15190);
nand U15824 (N_15824,N_15495,N_15194);
and U15825 (N_15825,N_15228,N_15472);
nand U15826 (N_15826,N_15300,N_15134);
nand U15827 (N_15827,N_15001,N_15310);
nor U15828 (N_15828,N_15215,N_15095);
nor U15829 (N_15829,N_15148,N_15079);
nand U15830 (N_15830,N_15164,N_15381);
nand U15831 (N_15831,N_15354,N_15334);
and U15832 (N_15832,N_15144,N_15058);
or U15833 (N_15833,N_15432,N_15340);
xnor U15834 (N_15834,N_15181,N_15473);
or U15835 (N_15835,N_15453,N_15255);
nand U15836 (N_15836,N_15119,N_15409);
and U15837 (N_15837,N_15402,N_15310);
nor U15838 (N_15838,N_15431,N_15252);
and U15839 (N_15839,N_15463,N_15315);
or U15840 (N_15840,N_15203,N_15319);
nand U15841 (N_15841,N_15317,N_15401);
xor U15842 (N_15842,N_15176,N_15093);
or U15843 (N_15843,N_15275,N_15332);
xnor U15844 (N_15844,N_15060,N_15407);
nand U15845 (N_15845,N_15350,N_15189);
nand U15846 (N_15846,N_15481,N_15206);
and U15847 (N_15847,N_15296,N_15065);
nor U15848 (N_15848,N_15169,N_15388);
and U15849 (N_15849,N_15329,N_15430);
xnor U15850 (N_15850,N_15325,N_15109);
or U15851 (N_15851,N_15464,N_15415);
or U15852 (N_15852,N_15165,N_15239);
or U15853 (N_15853,N_15101,N_15137);
nor U15854 (N_15854,N_15017,N_15216);
nand U15855 (N_15855,N_15411,N_15499);
or U15856 (N_15856,N_15124,N_15335);
nor U15857 (N_15857,N_15031,N_15138);
xor U15858 (N_15858,N_15329,N_15265);
nor U15859 (N_15859,N_15384,N_15236);
nor U15860 (N_15860,N_15019,N_15006);
xor U15861 (N_15861,N_15109,N_15352);
xor U15862 (N_15862,N_15256,N_15176);
xor U15863 (N_15863,N_15359,N_15273);
or U15864 (N_15864,N_15281,N_15335);
nand U15865 (N_15865,N_15428,N_15066);
nor U15866 (N_15866,N_15252,N_15005);
nor U15867 (N_15867,N_15052,N_15432);
xnor U15868 (N_15868,N_15123,N_15136);
or U15869 (N_15869,N_15479,N_15440);
or U15870 (N_15870,N_15433,N_15249);
nor U15871 (N_15871,N_15171,N_15055);
nand U15872 (N_15872,N_15461,N_15028);
and U15873 (N_15873,N_15365,N_15446);
or U15874 (N_15874,N_15435,N_15195);
and U15875 (N_15875,N_15490,N_15462);
or U15876 (N_15876,N_15062,N_15393);
and U15877 (N_15877,N_15217,N_15010);
nand U15878 (N_15878,N_15276,N_15026);
nand U15879 (N_15879,N_15319,N_15338);
xnor U15880 (N_15880,N_15489,N_15067);
and U15881 (N_15881,N_15031,N_15100);
or U15882 (N_15882,N_15144,N_15275);
and U15883 (N_15883,N_15402,N_15429);
xnor U15884 (N_15884,N_15385,N_15107);
nor U15885 (N_15885,N_15074,N_15004);
and U15886 (N_15886,N_15271,N_15438);
nor U15887 (N_15887,N_15236,N_15064);
nor U15888 (N_15888,N_15214,N_15058);
or U15889 (N_15889,N_15106,N_15490);
xor U15890 (N_15890,N_15246,N_15373);
and U15891 (N_15891,N_15405,N_15490);
and U15892 (N_15892,N_15017,N_15267);
and U15893 (N_15893,N_15097,N_15099);
nand U15894 (N_15894,N_15393,N_15058);
nand U15895 (N_15895,N_15020,N_15475);
or U15896 (N_15896,N_15328,N_15239);
and U15897 (N_15897,N_15010,N_15260);
nor U15898 (N_15898,N_15181,N_15359);
xor U15899 (N_15899,N_15310,N_15333);
and U15900 (N_15900,N_15174,N_15357);
nand U15901 (N_15901,N_15168,N_15282);
xor U15902 (N_15902,N_15183,N_15358);
and U15903 (N_15903,N_15365,N_15441);
or U15904 (N_15904,N_15115,N_15439);
xnor U15905 (N_15905,N_15201,N_15422);
and U15906 (N_15906,N_15275,N_15401);
nor U15907 (N_15907,N_15333,N_15161);
nor U15908 (N_15908,N_15275,N_15222);
nor U15909 (N_15909,N_15369,N_15349);
or U15910 (N_15910,N_15213,N_15239);
xnor U15911 (N_15911,N_15042,N_15387);
and U15912 (N_15912,N_15361,N_15455);
nand U15913 (N_15913,N_15285,N_15341);
and U15914 (N_15914,N_15343,N_15138);
xnor U15915 (N_15915,N_15299,N_15021);
or U15916 (N_15916,N_15069,N_15481);
nand U15917 (N_15917,N_15086,N_15342);
or U15918 (N_15918,N_15447,N_15450);
and U15919 (N_15919,N_15307,N_15073);
and U15920 (N_15920,N_15445,N_15188);
xnor U15921 (N_15921,N_15104,N_15261);
and U15922 (N_15922,N_15433,N_15288);
nor U15923 (N_15923,N_15031,N_15143);
xor U15924 (N_15924,N_15180,N_15122);
or U15925 (N_15925,N_15332,N_15274);
xor U15926 (N_15926,N_15041,N_15042);
or U15927 (N_15927,N_15117,N_15228);
nand U15928 (N_15928,N_15078,N_15442);
or U15929 (N_15929,N_15087,N_15403);
or U15930 (N_15930,N_15017,N_15201);
or U15931 (N_15931,N_15212,N_15142);
nand U15932 (N_15932,N_15116,N_15331);
xnor U15933 (N_15933,N_15290,N_15240);
nand U15934 (N_15934,N_15117,N_15308);
or U15935 (N_15935,N_15372,N_15339);
nor U15936 (N_15936,N_15063,N_15083);
and U15937 (N_15937,N_15306,N_15498);
or U15938 (N_15938,N_15164,N_15083);
and U15939 (N_15939,N_15200,N_15002);
xor U15940 (N_15940,N_15057,N_15387);
and U15941 (N_15941,N_15373,N_15472);
xor U15942 (N_15942,N_15410,N_15217);
nand U15943 (N_15943,N_15099,N_15267);
or U15944 (N_15944,N_15004,N_15220);
xor U15945 (N_15945,N_15152,N_15316);
and U15946 (N_15946,N_15343,N_15208);
xnor U15947 (N_15947,N_15324,N_15054);
nor U15948 (N_15948,N_15239,N_15362);
nor U15949 (N_15949,N_15280,N_15180);
nand U15950 (N_15950,N_15466,N_15124);
nor U15951 (N_15951,N_15470,N_15186);
xnor U15952 (N_15952,N_15074,N_15116);
nand U15953 (N_15953,N_15128,N_15275);
or U15954 (N_15954,N_15179,N_15497);
nor U15955 (N_15955,N_15205,N_15439);
or U15956 (N_15956,N_15404,N_15332);
or U15957 (N_15957,N_15268,N_15101);
xnor U15958 (N_15958,N_15279,N_15027);
nor U15959 (N_15959,N_15416,N_15329);
or U15960 (N_15960,N_15142,N_15201);
nand U15961 (N_15961,N_15280,N_15315);
nand U15962 (N_15962,N_15077,N_15256);
xor U15963 (N_15963,N_15355,N_15385);
and U15964 (N_15964,N_15423,N_15051);
and U15965 (N_15965,N_15164,N_15283);
nand U15966 (N_15966,N_15003,N_15378);
and U15967 (N_15967,N_15387,N_15338);
xor U15968 (N_15968,N_15065,N_15009);
xor U15969 (N_15969,N_15111,N_15456);
nand U15970 (N_15970,N_15389,N_15149);
or U15971 (N_15971,N_15029,N_15247);
and U15972 (N_15972,N_15091,N_15252);
xor U15973 (N_15973,N_15224,N_15275);
or U15974 (N_15974,N_15421,N_15394);
xnor U15975 (N_15975,N_15361,N_15464);
or U15976 (N_15976,N_15179,N_15031);
and U15977 (N_15977,N_15005,N_15429);
nand U15978 (N_15978,N_15138,N_15283);
xnor U15979 (N_15979,N_15462,N_15008);
or U15980 (N_15980,N_15065,N_15339);
or U15981 (N_15981,N_15494,N_15327);
nand U15982 (N_15982,N_15298,N_15418);
nand U15983 (N_15983,N_15487,N_15222);
or U15984 (N_15984,N_15200,N_15079);
or U15985 (N_15985,N_15122,N_15438);
xnor U15986 (N_15986,N_15006,N_15313);
nor U15987 (N_15987,N_15257,N_15088);
or U15988 (N_15988,N_15293,N_15499);
or U15989 (N_15989,N_15276,N_15084);
xor U15990 (N_15990,N_15396,N_15025);
or U15991 (N_15991,N_15048,N_15275);
or U15992 (N_15992,N_15139,N_15462);
and U15993 (N_15993,N_15164,N_15209);
xnor U15994 (N_15994,N_15321,N_15066);
and U15995 (N_15995,N_15198,N_15331);
nor U15996 (N_15996,N_15050,N_15001);
nand U15997 (N_15997,N_15033,N_15308);
nand U15998 (N_15998,N_15173,N_15003);
nor U15999 (N_15999,N_15007,N_15205);
and U16000 (N_16000,N_15817,N_15745);
nor U16001 (N_16001,N_15731,N_15901);
xnor U16002 (N_16002,N_15961,N_15809);
and U16003 (N_16003,N_15791,N_15523);
xor U16004 (N_16004,N_15606,N_15579);
and U16005 (N_16005,N_15870,N_15859);
nor U16006 (N_16006,N_15630,N_15504);
xnor U16007 (N_16007,N_15705,N_15522);
nor U16008 (N_16008,N_15852,N_15920);
xor U16009 (N_16009,N_15932,N_15605);
xnor U16010 (N_16010,N_15615,N_15595);
xor U16011 (N_16011,N_15729,N_15542);
xor U16012 (N_16012,N_15805,N_15984);
and U16013 (N_16013,N_15535,N_15891);
xnor U16014 (N_16014,N_15767,N_15665);
or U16015 (N_16015,N_15916,N_15617);
xnor U16016 (N_16016,N_15872,N_15879);
nand U16017 (N_16017,N_15570,N_15746);
and U16018 (N_16018,N_15765,N_15759);
xnor U16019 (N_16019,N_15744,N_15720);
or U16020 (N_16020,N_15868,N_15700);
xor U16021 (N_16021,N_15703,N_15904);
nor U16022 (N_16022,N_15930,N_15592);
and U16023 (N_16023,N_15661,N_15926);
xor U16024 (N_16024,N_15892,N_15575);
nor U16025 (N_16025,N_15913,N_15540);
nand U16026 (N_16026,N_15781,N_15794);
xor U16027 (N_16027,N_15969,N_15616);
and U16028 (N_16028,N_15629,N_15977);
nor U16029 (N_16029,N_15826,N_15847);
nand U16030 (N_16030,N_15712,N_15797);
xnor U16031 (N_16031,N_15866,N_15845);
xor U16032 (N_16032,N_15931,N_15771);
xor U16033 (N_16033,N_15632,N_15896);
nor U16034 (N_16034,N_15530,N_15514);
nand U16035 (N_16035,N_15688,N_15580);
and U16036 (N_16036,N_15832,N_15560);
nand U16037 (N_16037,N_15853,N_15676);
nor U16038 (N_16038,N_15707,N_15704);
and U16039 (N_16039,N_15634,N_15571);
xor U16040 (N_16040,N_15858,N_15666);
or U16041 (N_16041,N_15785,N_15644);
or U16042 (N_16042,N_15730,N_15633);
xor U16043 (N_16043,N_15878,N_15719);
and U16044 (N_16044,N_15573,N_15925);
xnor U16045 (N_16045,N_15821,N_15923);
nor U16046 (N_16046,N_15658,N_15854);
or U16047 (N_16047,N_15671,N_15871);
and U16048 (N_16048,N_15724,N_15699);
or U16049 (N_16049,N_15763,N_15538);
or U16050 (N_16050,N_15792,N_15812);
nor U16051 (N_16051,N_15897,N_15820);
and U16052 (N_16052,N_15622,N_15902);
nand U16053 (N_16053,N_15987,N_15788);
nand U16054 (N_16054,N_15681,N_15774);
nand U16055 (N_16055,N_15947,N_15756);
nor U16056 (N_16056,N_15950,N_15548);
nand U16057 (N_16057,N_15793,N_15803);
nand U16058 (N_16058,N_15670,N_15577);
xor U16059 (N_16059,N_15851,N_15928);
nand U16060 (N_16060,N_15698,N_15856);
or U16061 (N_16061,N_15784,N_15786);
xnor U16062 (N_16062,N_15808,N_15985);
nand U16063 (N_16063,N_15914,N_15515);
xor U16064 (N_16064,N_15869,N_15567);
nor U16065 (N_16065,N_15513,N_15819);
or U16066 (N_16066,N_15960,N_15751);
or U16067 (N_16067,N_15741,N_15789);
and U16068 (N_16068,N_15899,N_15663);
nor U16069 (N_16069,N_15804,N_15941);
or U16070 (N_16070,N_15511,N_15546);
and U16071 (N_16071,N_15843,N_15625);
nor U16072 (N_16072,N_15938,N_15922);
and U16073 (N_16073,N_15999,N_15718);
nand U16074 (N_16074,N_15628,N_15900);
nor U16075 (N_16075,N_15848,N_15773);
nor U16076 (N_16076,N_15728,N_15710);
xor U16077 (N_16077,N_15850,N_15591);
xnor U16078 (N_16078,N_15754,N_15768);
or U16079 (N_16079,N_15687,N_15971);
nor U16080 (N_16080,N_15825,N_15711);
nor U16081 (N_16081,N_15715,N_15647);
nor U16082 (N_16082,N_15508,N_15838);
xnor U16083 (N_16083,N_15936,N_15701);
and U16084 (N_16084,N_15709,N_15737);
xnor U16085 (N_16085,N_15586,N_15653);
and U16086 (N_16086,N_15713,N_15702);
or U16087 (N_16087,N_15637,N_15951);
nor U16088 (N_16088,N_15520,N_15877);
xor U16089 (N_16089,N_15956,N_15506);
xor U16090 (N_16090,N_15888,N_15993);
or U16091 (N_16091,N_15883,N_15937);
nand U16092 (N_16092,N_15684,N_15988);
or U16093 (N_16093,N_15994,N_15584);
and U16094 (N_16094,N_15662,N_15991);
nor U16095 (N_16095,N_15749,N_15549);
xnor U16096 (N_16096,N_15837,N_15777);
or U16097 (N_16097,N_15618,N_15521);
nor U16098 (N_16098,N_15559,N_15551);
xnor U16099 (N_16099,N_15680,N_15898);
xnor U16100 (N_16100,N_15933,N_15917);
or U16101 (N_16101,N_15693,N_15802);
nand U16102 (N_16102,N_15553,N_15833);
or U16103 (N_16103,N_15959,N_15949);
and U16104 (N_16104,N_15816,N_15695);
xnor U16105 (N_16105,N_15641,N_15624);
nand U16106 (N_16106,N_15613,N_15772);
or U16107 (N_16107,N_15849,N_15566);
nand U16108 (N_16108,N_15750,N_15536);
or U16109 (N_16109,N_15799,N_15547);
and U16110 (N_16110,N_15528,N_15865);
nand U16111 (N_16111,N_15979,N_15503);
nor U16112 (N_16112,N_15942,N_15939);
and U16113 (N_16113,N_15642,N_15968);
or U16114 (N_16114,N_15690,N_15655);
and U16115 (N_16115,N_15708,N_15783);
or U16116 (N_16116,N_15611,N_15518);
nand U16117 (N_16117,N_15934,N_15534);
and U16118 (N_16118,N_15552,N_15921);
and U16119 (N_16119,N_15512,N_15955);
nor U16120 (N_16120,N_15685,N_15940);
or U16121 (N_16121,N_15667,N_15829);
nor U16122 (N_16122,N_15590,N_15723);
and U16123 (N_16123,N_15556,N_15758);
nor U16124 (N_16124,N_15964,N_15970);
xnor U16125 (N_16125,N_15810,N_15760);
nand U16126 (N_16126,N_15906,N_15656);
xor U16127 (N_16127,N_15526,N_15814);
nor U16128 (N_16128,N_15717,N_15974);
xor U16129 (N_16129,N_15766,N_15739);
or U16130 (N_16130,N_15948,N_15885);
and U16131 (N_16131,N_15908,N_15596);
nor U16132 (N_16132,N_15735,N_15679);
xor U16133 (N_16133,N_15747,N_15568);
or U16134 (N_16134,N_15981,N_15697);
nand U16135 (N_16135,N_15539,N_15953);
xnor U16136 (N_16136,N_15895,N_15813);
or U16137 (N_16137,N_15998,N_15909);
nor U16138 (N_16138,N_15675,N_15578);
or U16139 (N_16139,N_15686,N_15725);
or U16140 (N_16140,N_15927,N_15753);
nor U16141 (N_16141,N_15780,N_15738);
xor U16142 (N_16142,N_15995,N_15664);
nor U16143 (N_16143,N_15643,N_15529);
and U16144 (N_16144,N_15588,N_15654);
nor U16145 (N_16145,N_15574,N_15516);
xnor U16146 (N_16146,N_15841,N_15620);
xor U16147 (N_16147,N_15593,N_15798);
and U16148 (N_16148,N_15648,N_15980);
xnor U16149 (N_16149,N_15764,N_15603);
xor U16150 (N_16150,N_15646,N_15752);
or U16151 (N_16151,N_15517,N_15945);
nor U16152 (N_16152,N_15696,N_15682);
nand U16153 (N_16153,N_15842,N_15597);
xnor U16154 (N_16154,N_15860,N_15770);
or U16155 (N_16155,N_15828,N_15801);
xor U16156 (N_16156,N_15594,N_15935);
xor U16157 (N_16157,N_15972,N_15543);
nor U16158 (N_16158,N_15533,N_15608);
xnor U16159 (N_16159,N_15835,N_15544);
xor U16160 (N_16160,N_15598,N_15507);
xnor U16161 (N_16161,N_15692,N_15732);
nor U16162 (N_16162,N_15963,N_15557);
xnor U16163 (N_16163,N_15525,N_15903);
nor U16164 (N_16164,N_15880,N_15857);
nand U16165 (N_16165,N_15874,N_15527);
nand U16166 (N_16166,N_15531,N_15776);
nand U16167 (N_16167,N_15631,N_15996);
xnor U16168 (N_16168,N_15722,N_15524);
and U16169 (N_16169,N_15790,N_15855);
and U16170 (N_16170,N_15602,N_15502);
nand U16171 (N_16171,N_15743,N_15623);
nand U16172 (N_16172,N_15861,N_15886);
xor U16173 (N_16173,N_15876,N_15889);
nor U16174 (N_16174,N_15796,N_15569);
and U16175 (N_16175,N_15600,N_15550);
nor U16176 (N_16176,N_15541,N_15678);
nand U16177 (N_16177,N_15965,N_15867);
xnor U16178 (N_16178,N_15609,N_15582);
and U16179 (N_16179,N_15882,N_15831);
and U16180 (N_16180,N_15839,N_15887);
xor U16181 (N_16181,N_15986,N_15672);
nor U16182 (N_16182,N_15510,N_15893);
and U16183 (N_16183,N_15558,N_15599);
and U16184 (N_16184,N_15782,N_15554);
xnor U16185 (N_16185,N_15601,N_15500);
nand U16186 (N_16186,N_15827,N_15762);
xnor U16187 (N_16187,N_15505,N_15537);
xor U16188 (N_16188,N_15881,N_15966);
nand U16189 (N_16189,N_15824,N_15587);
xor U16190 (N_16190,N_15915,N_15565);
and U16191 (N_16191,N_15519,N_15585);
nand U16192 (N_16192,N_15651,N_15946);
nand U16193 (N_16193,N_15627,N_15564);
nand U16194 (N_16194,N_15983,N_15757);
nor U16195 (N_16195,N_15639,N_15962);
nor U16196 (N_16196,N_15677,N_15614);
and U16197 (N_16197,N_15576,N_15561);
and U16198 (N_16198,N_15822,N_15674);
nor U16199 (N_16199,N_15742,N_15555);
or U16200 (N_16200,N_15673,N_15836);
or U16201 (N_16201,N_15716,N_15807);
xnor U16202 (N_16202,N_15612,N_15795);
nor U16203 (N_16203,N_15668,N_15989);
nand U16204 (N_16204,N_15740,N_15875);
nor U16205 (N_16205,N_15636,N_15638);
xnor U16206 (N_16206,N_15572,N_15929);
or U16207 (N_16207,N_15944,N_15604);
xor U16208 (N_16208,N_15919,N_15645);
nand U16209 (N_16209,N_15806,N_15918);
or U16210 (N_16210,N_15992,N_15683);
or U16211 (N_16211,N_15894,N_15726);
xor U16212 (N_16212,N_15652,N_15973);
xnor U16213 (N_16213,N_15581,N_15583);
or U16214 (N_16214,N_15621,N_15501);
nor U16215 (N_16215,N_15610,N_15976);
xor U16216 (N_16216,N_15840,N_15924);
nand U16217 (N_16217,N_15863,N_15650);
or U16218 (N_16218,N_15689,N_15635);
or U16219 (N_16219,N_15748,N_15657);
xnor U16220 (N_16220,N_15706,N_15967);
and U16221 (N_16221,N_15818,N_15830);
nor U16222 (N_16222,N_15990,N_15659);
nand U16223 (N_16223,N_15911,N_15978);
nand U16224 (N_16224,N_15734,N_15815);
xnor U16225 (N_16225,N_15787,N_15761);
xnor U16226 (N_16226,N_15912,N_15714);
nand U16227 (N_16227,N_15952,N_15864);
xor U16228 (N_16228,N_15982,N_15873);
xnor U16229 (N_16229,N_15957,N_15779);
or U16230 (N_16230,N_15669,N_15640);
and U16231 (N_16231,N_15562,N_15954);
nor U16232 (N_16232,N_15619,N_15532);
and U16233 (N_16233,N_15721,N_15626);
nand U16234 (N_16234,N_15755,N_15509);
or U16235 (N_16235,N_15890,N_15884);
xor U16236 (N_16236,N_15727,N_15660);
or U16237 (N_16237,N_15862,N_15778);
nor U16238 (N_16238,N_15775,N_15607);
nor U16239 (N_16239,N_15563,N_15844);
and U16240 (N_16240,N_15846,N_15545);
nor U16241 (N_16241,N_15800,N_15910);
or U16242 (N_16242,N_15649,N_15958);
xnor U16243 (N_16243,N_15907,N_15733);
xnor U16244 (N_16244,N_15736,N_15769);
xor U16245 (N_16245,N_15589,N_15811);
xor U16246 (N_16246,N_15691,N_15823);
and U16247 (N_16247,N_15905,N_15943);
nor U16248 (N_16248,N_15834,N_15997);
xnor U16249 (N_16249,N_15975,N_15694);
nand U16250 (N_16250,N_15998,N_15794);
nand U16251 (N_16251,N_15936,N_15693);
xnor U16252 (N_16252,N_15809,N_15626);
and U16253 (N_16253,N_15932,N_15624);
nand U16254 (N_16254,N_15773,N_15559);
nand U16255 (N_16255,N_15930,N_15826);
or U16256 (N_16256,N_15546,N_15798);
and U16257 (N_16257,N_15707,N_15615);
nor U16258 (N_16258,N_15592,N_15582);
and U16259 (N_16259,N_15631,N_15605);
nor U16260 (N_16260,N_15982,N_15949);
and U16261 (N_16261,N_15654,N_15889);
nand U16262 (N_16262,N_15713,N_15920);
or U16263 (N_16263,N_15893,N_15601);
nor U16264 (N_16264,N_15841,N_15586);
or U16265 (N_16265,N_15585,N_15624);
nor U16266 (N_16266,N_15690,N_15841);
or U16267 (N_16267,N_15620,N_15849);
xor U16268 (N_16268,N_15860,N_15590);
and U16269 (N_16269,N_15793,N_15939);
xnor U16270 (N_16270,N_15509,N_15779);
nand U16271 (N_16271,N_15885,N_15855);
nand U16272 (N_16272,N_15548,N_15961);
nand U16273 (N_16273,N_15840,N_15992);
xor U16274 (N_16274,N_15520,N_15566);
xor U16275 (N_16275,N_15631,N_15946);
nor U16276 (N_16276,N_15863,N_15564);
xor U16277 (N_16277,N_15665,N_15746);
and U16278 (N_16278,N_15999,N_15553);
and U16279 (N_16279,N_15847,N_15933);
nor U16280 (N_16280,N_15527,N_15790);
nor U16281 (N_16281,N_15743,N_15914);
nor U16282 (N_16282,N_15913,N_15641);
nand U16283 (N_16283,N_15628,N_15994);
nor U16284 (N_16284,N_15957,N_15922);
nand U16285 (N_16285,N_15875,N_15908);
nor U16286 (N_16286,N_15587,N_15747);
and U16287 (N_16287,N_15578,N_15663);
xor U16288 (N_16288,N_15890,N_15592);
nor U16289 (N_16289,N_15561,N_15807);
and U16290 (N_16290,N_15671,N_15530);
nand U16291 (N_16291,N_15947,N_15933);
nor U16292 (N_16292,N_15948,N_15919);
nor U16293 (N_16293,N_15563,N_15984);
xor U16294 (N_16294,N_15720,N_15965);
xnor U16295 (N_16295,N_15929,N_15911);
and U16296 (N_16296,N_15781,N_15662);
or U16297 (N_16297,N_15769,N_15742);
nor U16298 (N_16298,N_15877,N_15584);
and U16299 (N_16299,N_15877,N_15920);
nor U16300 (N_16300,N_15820,N_15638);
or U16301 (N_16301,N_15578,N_15690);
nor U16302 (N_16302,N_15662,N_15892);
and U16303 (N_16303,N_15587,N_15965);
nor U16304 (N_16304,N_15630,N_15989);
or U16305 (N_16305,N_15991,N_15648);
or U16306 (N_16306,N_15561,N_15885);
xor U16307 (N_16307,N_15660,N_15993);
or U16308 (N_16308,N_15596,N_15984);
or U16309 (N_16309,N_15538,N_15635);
nand U16310 (N_16310,N_15695,N_15904);
xnor U16311 (N_16311,N_15659,N_15756);
and U16312 (N_16312,N_15582,N_15872);
xnor U16313 (N_16313,N_15604,N_15755);
nor U16314 (N_16314,N_15808,N_15884);
nand U16315 (N_16315,N_15538,N_15784);
xnor U16316 (N_16316,N_15900,N_15699);
xor U16317 (N_16317,N_15778,N_15586);
xor U16318 (N_16318,N_15754,N_15968);
or U16319 (N_16319,N_15587,N_15868);
or U16320 (N_16320,N_15506,N_15821);
xor U16321 (N_16321,N_15949,N_15545);
xor U16322 (N_16322,N_15607,N_15964);
xor U16323 (N_16323,N_15712,N_15710);
xor U16324 (N_16324,N_15820,N_15667);
or U16325 (N_16325,N_15624,N_15991);
xnor U16326 (N_16326,N_15872,N_15677);
nand U16327 (N_16327,N_15809,N_15610);
and U16328 (N_16328,N_15838,N_15724);
nand U16329 (N_16329,N_15830,N_15973);
or U16330 (N_16330,N_15766,N_15546);
or U16331 (N_16331,N_15547,N_15948);
nor U16332 (N_16332,N_15519,N_15610);
xor U16333 (N_16333,N_15590,N_15631);
nor U16334 (N_16334,N_15666,N_15517);
or U16335 (N_16335,N_15952,N_15557);
and U16336 (N_16336,N_15730,N_15775);
or U16337 (N_16337,N_15522,N_15643);
or U16338 (N_16338,N_15635,N_15945);
nor U16339 (N_16339,N_15691,N_15821);
nor U16340 (N_16340,N_15644,N_15676);
or U16341 (N_16341,N_15987,N_15722);
xor U16342 (N_16342,N_15738,N_15646);
xor U16343 (N_16343,N_15601,N_15550);
and U16344 (N_16344,N_15518,N_15765);
nand U16345 (N_16345,N_15883,N_15552);
nor U16346 (N_16346,N_15877,N_15730);
or U16347 (N_16347,N_15544,N_15913);
nand U16348 (N_16348,N_15568,N_15676);
xnor U16349 (N_16349,N_15614,N_15645);
nor U16350 (N_16350,N_15755,N_15618);
nand U16351 (N_16351,N_15538,N_15948);
nand U16352 (N_16352,N_15694,N_15844);
or U16353 (N_16353,N_15985,N_15711);
and U16354 (N_16354,N_15698,N_15614);
xor U16355 (N_16355,N_15852,N_15735);
nand U16356 (N_16356,N_15501,N_15736);
nor U16357 (N_16357,N_15931,N_15908);
or U16358 (N_16358,N_15770,N_15522);
or U16359 (N_16359,N_15589,N_15941);
nor U16360 (N_16360,N_15804,N_15884);
nand U16361 (N_16361,N_15770,N_15596);
nor U16362 (N_16362,N_15908,N_15735);
and U16363 (N_16363,N_15804,N_15636);
xor U16364 (N_16364,N_15641,N_15671);
and U16365 (N_16365,N_15898,N_15904);
or U16366 (N_16366,N_15859,N_15821);
or U16367 (N_16367,N_15820,N_15804);
xnor U16368 (N_16368,N_15714,N_15552);
or U16369 (N_16369,N_15795,N_15802);
nor U16370 (N_16370,N_15919,N_15503);
nor U16371 (N_16371,N_15552,N_15736);
nor U16372 (N_16372,N_15600,N_15853);
nor U16373 (N_16373,N_15786,N_15605);
xnor U16374 (N_16374,N_15695,N_15811);
xnor U16375 (N_16375,N_15614,N_15730);
nor U16376 (N_16376,N_15744,N_15569);
nand U16377 (N_16377,N_15980,N_15789);
or U16378 (N_16378,N_15825,N_15699);
and U16379 (N_16379,N_15987,N_15592);
and U16380 (N_16380,N_15593,N_15532);
or U16381 (N_16381,N_15991,N_15841);
nand U16382 (N_16382,N_15990,N_15825);
nor U16383 (N_16383,N_15906,N_15529);
and U16384 (N_16384,N_15987,N_15529);
nor U16385 (N_16385,N_15900,N_15939);
and U16386 (N_16386,N_15697,N_15712);
nor U16387 (N_16387,N_15541,N_15577);
nand U16388 (N_16388,N_15745,N_15897);
xnor U16389 (N_16389,N_15952,N_15526);
nand U16390 (N_16390,N_15520,N_15568);
nand U16391 (N_16391,N_15782,N_15600);
nor U16392 (N_16392,N_15584,N_15975);
and U16393 (N_16393,N_15982,N_15725);
or U16394 (N_16394,N_15726,N_15515);
nand U16395 (N_16395,N_15744,N_15585);
nor U16396 (N_16396,N_15861,N_15954);
nor U16397 (N_16397,N_15967,N_15586);
or U16398 (N_16398,N_15599,N_15885);
xnor U16399 (N_16399,N_15585,N_15735);
xnor U16400 (N_16400,N_15707,N_15786);
nand U16401 (N_16401,N_15624,N_15718);
nor U16402 (N_16402,N_15984,N_15698);
xnor U16403 (N_16403,N_15723,N_15540);
nand U16404 (N_16404,N_15691,N_15543);
or U16405 (N_16405,N_15509,N_15717);
and U16406 (N_16406,N_15798,N_15547);
and U16407 (N_16407,N_15904,N_15957);
and U16408 (N_16408,N_15520,N_15885);
nor U16409 (N_16409,N_15625,N_15643);
nand U16410 (N_16410,N_15699,N_15562);
or U16411 (N_16411,N_15711,N_15730);
and U16412 (N_16412,N_15590,N_15845);
and U16413 (N_16413,N_15901,N_15778);
and U16414 (N_16414,N_15584,N_15967);
or U16415 (N_16415,N_15981,N_15567);
nand U16416 (N_16416,N_15525,N_15530);
xor U16417 (N_16417,N_15590,N_15551);
nor U16418 (N_16418,N_15646,N_15802);
or U16419 (N_16419,N_15556,N_15838);
nor U16420 (N_16420,N_15536,N_15607);
nand U16421 (N_16421,N_15925,N_15822);
xor U16422 (N_16422,N_15959,N_15658);
or U16423 (N_16423,N_15779,N_15869);
nand U16424 (N_16424,N_15961,N_15654);
and U16425 (N_16425,N_15565,N_15962);
nor U16426 (N_16426,N_15766,N_15883);
nor U16427 (N_16427,N_15574,N_15972);
and U16428 (N_16428,N_15947,N_15818);
nand U16429 (N_16429,N_15629,N_15917);
nand U16430 (N_16430,N_15517,N_15915);
or U16431 (N_16431,N_15977,N_15791);
nand U16432 (N_16432,N_15514,N_15764);
and U16433 (N_16433,N_15527,N_15546);
nand U16434 (N_16434,N_15671,N_15690);
nor U16435 (N_16435,N_15626,N_15786);
nand U16436 (N_16436,N_15601,N_15703);
or U16437 (N_16437,N_15564,N_15535);
nor U16438 (N_16438,N_15529,N_15870);
or U16439 (N_16439,N_15730,N_15896);
nand U16440 (N_16440,N_15901,N_15670);
nand U16441 (N_16441,N_15800,N_15595);
nor U16442 (N_16442,N_15818,N_15756);
or U16443 (N_16443,N_15992,N_15741);
nor U16444 (N_16444,N_15796,N_15826);
or U16445 (N_16445,N_15992,N_15963);
nor U16446 (N_16446,N_15518,N_15618);
or U16447 (N_16447,N_15786,N_15680);
or U16448 (N_16448,N_15543,N_15638);
nor U16449 (N_16449,N_15540,N_15533);
nand U16450 (N_16450,N_15957,N_15689);
nand U16451 (N_16451,N_15549,N_15504);
xor U16452 (N_16452,N_15715,N_15721);
nor U16453 (N_16453,N_15745,N_15513);
or U16454 (N_16454,N_15682,N_15524);
nor U16455 (N_16455,N_15821,N_15738);
and U16456 (N_16456,N_15789,N_15819);
nor U16457 (N_16457,N_15822,N_15537);
nand U16458 (N_16458,N_15709,N_15874);
or U16459 (N_16459,N_15579,N_15920);
or U16460 (N_16460,N_15835,N_15754);
xor U16461 (N_16461,N_15789,N_15972);
xor U16462 (N_16462,N_15816,N_15972);
or U16463 (N_16463,N_15797,N_15767);
xor U16464 (N_16464,N_15835,N_15605);
nand U16465 (N_16465,N_15722,N_15577);
nor U16466 (N_16466,N_15605,N_15968);
or U16467 (N_16467,N_15518,N_15871);
xor U16468 (N_16468,N_15739,N_15728);
and U16469 (N_16469,N_15946,N_15654);
nand U16470 (N_16470,N_15519,N_15854);
and U16471 (N_16471,N_15614,N_15889);
nand U16472 (N_16472,N_15638,N_15936);
xor U16473 (N_16473,N_15732,N_15561);
nand U16474 (N_16474,N_15903,N_15865);
or U16475 (N_16475,N_15883,N_15732);
nor U16476 (N_16476,N_15640,N_15845);
nand U16477 (N_16477,N_15587,N_15724);
and U16478 (N_16478,N_15754,N_15593);
nor U16479 (N_16479,N_15605,N_15751);
and U16480 (N_16480,N_15567,N_15934);
nand U16481 (N_16481,N_15905,N_15785);
nand U16482 (N_16482,N_15852,N_15583);
or U16483 (N_16483,N_15568,N_15523);
xor U16484 (N_16484,N_15794,N_15846);
or U16485 (N_16485,N_15824,N_15562);
or U16486 (N_16486,N_15544,N_15684);
or U16487 (N_16487,N_15961,N_15705);
nor U16488 (N_16488,N_15903,N_15973);
or U16489 (N_16489,N_15662,N_15852);
nand U16490 (N_16490,N_15696,N_15675);
and U16491 (N_16491,N_15721,N_15990);
xor U16492 (N_16492,N_15831,N_15566);
nand U16493 (N_16493,N_15518,N_15823);
nand U16494 (N_16494,N_15970,N_15887);
nand U16495 (N_16495,N_15688,N_15657);
or U16496 (N_16496,N_15766,N_15618);
nand U16497 (N_16497,N_15905,N_15815);
or U16498 (N_16498,N_15912,N_15556);
and U16499 (N_16499,N_15569,N_15587);
or U16500 (N_16500,N_16298,N_16492);
xnor U16501 (N_16501,N_16238,N_16170);
and U16502 (N_16502,N_16416,N_16200);
or U16503 (N_16503,N_16001,N_16141);
nor U16504 (N_16504,N_16305,N_16084);
xnor U16505 (N_16505,N_16035,N_16257);
or U16506 (N_16506,N_16380,N_16253);
xnor U16507 (N_16507,N_16112,N_16366);
nand U16508 (N_16508,N_16296,N_16307);
nand U16509 (N_16509,N_16326,N_16198);
and U16510 (N_16510,N_16462,N_16418);
nor U16511 (N_16511,N_16343,N_16099);
xnor U16512 (N_16512,N_16496,N_16093);
or U16513 (N_16513,N_16105,N_16102);
or U16514 (N_16514,N_16373,N_16053);
xor U16515 (N_16515,N_16031,N_16321);
nor U16516 (N_16516,N_16166,N_16284);
and U16517 (N_16517,N_16362,N_16458);
or U16518 (N_16518,N_16176,N_16056);
nand U16519 (N_16519,N_16493,N_16452);
and U16520 (N_16520,N_16333,N_16008);
and U16521 (N_16521,N_16441,N_16218);
xnor U16522 (N_16522,N_16219,N_16303);
or U16523 (N_16523,N_16354,N_16325);
nand U16524 (N_16524,N_16036,N_16071);
or U16525 (N_16525,N_16454,N_16486);
nor U16526 (N_16526,N_16385,N_16087);
and U16527 (N_16527,N_16327,N_16291);
or U16528 (N_16528,N_16227,N_16448);
xor U16529 (N_16529,N_16187,N_16329);
nand U16530 (N_16530,N_16078,N_16247);
nand U16531 (N_16531,N_16269,N_16421);
nand U16532 (N_16532,N_16406,N_16183);
and U16533 (N_16533,N_16092,N_16022);
nor U16534 (N_16534,N_16383,N_16018);
xnor U16535 (N_16535,N_16480,N_16419);
nor U16536 (N_16536,N_16415,N_16049);
nor U16537 (N_16537,N_16094,N_16216);
nor U16538 (N_16538,N_16317,N_16185);
nor U16539 (N_16539,N_16498,N_16080);
nor U16540 (N_16540,N_16289,N_16365);
xnor U16541 (N_16541,N_16372,N_16217);
nor U16542 (N_16542,N_16434,N_16360);
and U16543 (N_16543,N_16339,N_16275);
and U16544 (N_16544,N_16260,N_16456);
and U16545 (N_16545,N_16075,N_16435);
or U16546 (N_16546,N_16125,N_16029);
and U16547 (N_16547,N_16174,N_16015);
or U16548 (N_16548,N_16083,N_16330);
or U16549 (N_16549,N_16020,N_16004);
xnor U16550 (N_16550,N_16427,N_16204);
nor U16551 (N_16551,N_16489,N_16107);
and U16552 (N_16552,N_16194,N_16320);
nor U16553 (N_16553,N_16256,N_16258);
or U16554 (N_16554,N_16450,N_16195);
or U16555 (N_16555,N_16390,N_16313);
or U16556 (N_16556,N_16440,N_16143);
xnor U16557 (N_16557,N_16046,N_16072);
and U16558 (N_16558,N_16173,N_16285);
nor U16559 (N_16559,N_16495,N_16229);
or U16560 (N_16560,N_16283,N_16106);
and U16561 (N_16561,N_16199,N_16158);
nand U16562 (N_16562,N_16070,N_16108);
xnor U16563 (N_16563,N_16381,N_16153);
or U16564 (N_16564,N_16426,N_16074);
or U16565 (N_16565,N_16213,N_16119);
nor U16566 (N_16566,N_16451,N_16379);
nor U16567 (N_16567,N_16266,N_16484);
xor U16568 (N_16568,N_16287,N_16364);
or U16569 (N_16569,N_16398,N_16466);
xnor U16570 (N_16570,N_16005,N_16461);
nand U16571 (N_16571,N_16475,N_16323);
nor U16572 (N_16572,N_16089,N_16393);
xor U16573 (N_16573,N_16446,N_16161);
nor U16574 (N_16574,N_16397,N_16344);
nand U16575 (N_16575,N_16282,N_16206);
and U16576 (N_16576,N_16130,N_16131);
and U16577 (N_16577,N_16164,N_16394);
xor U16578 (N_16578,N_16134,N_16288);
nand U16579 (N_16579,N_16403,N_16026);
or U16580 (N_16580,N_16097,N_16154);
xor U16581 (N_16581,N_16472,N_16473);
xnor U16582 (N_16582,N_16028,N_16384);
nor U16583 (N_16583,N_16483,N_16007);
xor U16584 (N_16584,N_16274,N_16359);
nor U16585 (N_16585,N_16220,N_16011);
nor U16586 (N_16586,N_16024,N_16202);
or U16587 (N_16587,N_16363,N_16042);
xor U16588 (N_16588,N_16404,N_16271);
nand U16589 (N_16589,N_16273,N_16293);
and U16590 (N_16590,N_16044,N_16335);
and U16591 (N_16591,N_16348,N_16414);
nor U16592 (N_16592,N_16150,N_16355);
and U16593 (N_16593,N_16090,N_16180);
xor U16594 (N_16594,N_16063,N_16244);
nand U16595 (N_16595,N_16405,N_16332);
xnor U16596 (N_16596,N_16336,N_16442);
xor U16597 (N_16597,N_16010,N_16371);
nand U16598 (N_16598,N_16347,N_16225);
nor U16599 (N_16599,N_16148,N_16133);
xor U16600 (N_16600,N_16351,N_16230);
xor U16601 (N_16601,N_16369,N_16478);
nor U16602 (N_16602,N_16037,N_16226);
nor U16603 (N_16603,N_16016,N_16444);
or U16604 (N_16604,N_16453,N_16062);
or U16605 (N_16605,N_16312,N_16252);
nor U16606 (N_16606,N_16413,N_16115);
and U16607 (N_16607,N_16157,N_16254);
nand U16608 (N_16608,N_16168,N_16025);
xor U16609 (N_16609,N_16428,N_16278);
or U16610 (N_16610,N_16245,N_16349);
nand U16611 (N_16611,N_16165,N_16377);
xnor U16612 (N_16612,N_16051,N_16255);
and U16613 (N_16613,N_16128,N_16346);
or U16614 (N_16614,N_16100,N_16449);
or U16615 (N_16615,N_16203,N_16400);
nor U16616 (N_16616,N_16251,N_16032);
nand U16617 (N_16617,N_16048,N_16306);
xor U16618 (N_16618,N_16171,N_16027);
or U16619 (N_16619,N_16311,N_16436);
xnor U16620 (N_16620,N_16116,N_16239);
or U16621 (N_16621,N_16182,N_16152);
xor U16622 (N_16622,N_16276,N_16352);
and U16623 (N_16623,N_16370,N_16350);
nor U16624 (N_16624,N_16002,N_16212);
or U16625 (N_16625,N_16392,N_16375);
xnor U16626 (N_16626,N_16043,N_16345);
xor U16627 (N_16627,N_16468,N_16232);
and U16628 (N_16628,N_16262,N_16412);
or U16629 (N_16629,N_16302,N_16184);
xnor U16630 (N_16630,N_16163,N_16211);
and U16631 (N_16631,N_16270,N_16124);
nor U16632 (N_16632,N_16109,N_16110);
or U16633 (N_16633,N_16013,N_16367);
nor U16634 (N_16634,N_16067,N_16017);
or U16635 (N_16635,N_16021,N_16139);
or U16636 (N_16636,N_16420,N_16309);
nor U16637 (N_16637,N_16012,N_16060);
and U16638 (N_16638,N_16019,N_16085);
or U16639 (N_16639,N_16300,N_16417);
nor U16640 (N_16640,N_16210,N_16374);
nor U16641 (N_16641,N_16234,N_16151);
nand U16642 (N_16642,N_16272,N_16052);
nand U16643 (N_16643,N_16463,N_16140);
or U16644 (N_16644,N_16459,N_16353);
nand U16645 (N_16645,N_16358,N_16438);
and U16646 (N_16646,N_16248,N_16069);
nand U16647 (N_16647,N_16224,N_16485);
and U16648 (N_16648,N_16117,N_16259);
nand U16649 (N_16649,N_16009,N_16395);
xor U16650 (N_16650,N_16445,N_16160);
nand U16651 (N_16651,N_16177,N_16261);
nand U16652 (N_16652,N_16433,N_16214);
nand U16653 (N_16653,N_16465,N_16066);
or U16654 (N_16654,N_16250,N_16341);
and U16655 (N_16655,N_16030,N_16023);
or U16656 (N_16656,N_16491,N_16429);
and U16657 (N_16657,N_16172,N_16249);
nand U16658 (N_16658,N_16129,N_16127);
xnor U16659 (N_16659,N_16361,N_16233);
nor U16660 (N_16660,N_16146,N_16231);
nand U16661 (N_16661,N_16156,N_16136);
and U16662 (N_16662,N_16041,N_16082);
xor U16663 (N_16663,N_16142,N_16470);
and U16664 (N_16664,N_16378,N_16208);
or U16665 (N_16665,N_16264,N_16101);
nand U16666 (N_16666,N_16310,N_16304);
or U16667 (N_16667,N_16457,N_16081);
or U16668 (N_16668,N_16482,N_16215);
and U16669 (N_16669,N_16389,N_16149);
xnor U16670 (N_16670,N_16123,N_16111);
nor U16671 (N_16671,N_16467,N_16396);
nand U16672 (N_16672,N_16207,N_16401);
nand U16673 (N_16673,N_16314,N_16235);
or U16674 (N_16674,N_16205,N_16159);
xnor U16675 (N_16675,N_16086,N_16447);
nand U16676 (N_16676,N_16096,N_16196);
and U16677 (N_16677,N_16280,N_16263);
and U16678 (N_16678,N_16479,N_16223);
nand U16679 (N_16679,N_16034,N_16337);
nand U16680 (N_16680,N_16064,N_16286);
nor U16681 (N_16681,N_16430,N_16126);
nand U16682 (N_16682,N_16399,N_16464);
nand U16683 (N_16683,N_16324,N_16281);
and U16684 (N_16684,N_16228,N_16181);
nor U16685 (N_16685,N_16382,N_16144);
or U16686 (N_16686,N_16192,N_16190);
and U16687 (N_16687,N_16033,N_16167);
xnor U16688 (N_16688,N_16193,N_16474);
or U16689 (N_16689,N_16318,N_16014);
and U16690 (N_16690,N_16240,N_16424);
and U16691 (N_16691,N_16422,N_16055);
or U16692 (N_16692,N_16179,N_16073);
or U16693 (N_16693,N_16301,N_16000);
nand U16694 (N_16694,N_16471,N_16357);
and U16695 (N_16695,N_16045,N_16460);
xor U16696 (N_16696,N_16050,N_16294);
nor U16697 (N_16697,N_16186,N_16040);
and U16698 (N_16698,N_16342,N_16308);
and U16699 (N_16699,N_16267,N_16494);
nand U16700 (N_16700,N_16065,N_16038);
nor U16701 (N_16701,N_16221,N_16118);
nor U16702 (N_16702,N_16003,N_16237);
nor U16703 (N_16703,N_16423,N_16432);
xor U16704 (N_16704,N_16376,N_16091);
or U16705 (N_16705,N_16408,N_16391);
xor U16706 (N_16706,N_16322,N_16425);
xnor U16707 (N_16707,N_16297,N_16277);
xor U16708 (N_16708,N_16409,N_16431);
xnor U16709 (N_16709,N_16114,N_16411);
or U16710 (N_16710,N_16061,N_16059);
or U16711 (N_16711,N_16334,N_16487);
nor U16712 (N_16712,N_16299,N_16079);
or U16713 (N_16713,N_16145,N_16169);
xnor U16714 (N_16714,N_16132,N_16175);
nor U16715 (N_16715,N_16356,N_16120);
and U16716 (N_16716,N_16138,N_16242);
nor U16717 (N_16717,N_16315,N_16490);
xnor U16718 (N_16718,N_16387,N_16054);
or U16719 (N_16719,N_16499,N_16188);
xnor U16720 (N_16720,N_16077,N_16095);
xor U16721 (N_16721,N_16047,N_16488);
nor U16722 (N_16722,N_16068,N_16135);
nand U16723 (N_16723,N_16189,N_16279);
and U16724 (N_16724,N_16340,N_16104);
and U16725 (N_16725,N_16147,N_16410);
nand U16726 (N_16726,N_16455,N_16290);
xnor U16727 (N_16727,N_16209,N_16331);
xnor U16728 (N_16728,N_16469,N_16477);
nor U16729 (N_16729,N_16197,N_16088);
nor U16730 (N_16730,N_16319,N_16098);
and U16731 (N_16731,N_16076,N_16338);
nor U16732 (N_16732,N_16201,N_16316);
nor U16733 (N_16733,N_16121,N_16368);
nand U16734 (N_16734,N_16295,N_16006);
and U16735 (N_16735,N_16268,N_16155);
and U16736 (N_16736,N_16407,N_16058);
nor U16737 (N_16737,N_16386,N_16328);
xnor U16738 (N_16738,N_16497,N_16113);
nor U16739 (N_16739,N_16265,N_16439);
nand U16740 (N_16740,N_16481,N_16402);
or U16741 (N_16741,N_16443,N_16191);
or U16742 (N_16742,N_16437,N_16246);
nand U16743 (N_16743,N_16162,N_16222);
nor U16744 (N_16744,N_16137,N_16039);
and U16745 (N_16745,N_16292,N_16103);
xor U16746 (N_16746,N_16243,N_16236);
and U16747 (N_16747,N_16388,N_16178);
xnor U16748 (N_16748,N_16057,N_16241);
nand U16749 (N_16749,N_16122,N_16476);
or U16750 (N_16750,N_16428,N_16063);
nand U16751 (N_16751,N_16221,N_16115);
or U16752 (N_16752,N_16187,N_16140);
xnor U16753 (N_16753,N_16247,N_16293);
nor U16754 (N_16754,N_16443,N_16420);
xnor U16755 (N_16755,N_16291,N_16391);
xnor U16756 (N_16756,N_16010,N_16328);
nor U16757 (N_16757,N_16484,N_16409);
nor U16758 (N_16758,N_16004,N_16320);
nand U16759 (N_16759,N_16196,N_16419);
or U16760 (N_16760,N_16188,N_16334);
or U16761 (N_16761,N_16445,N_16191);
and U16762 (N_16762,N_16186,N_16434);
or U16763 (N_16763,N_16292,N_16150);
nand U16764 (N_16764,N_16383,N_16455);
and U16765 (N_16765,N_16347,N_16111);
nand U16766 (N_16766,N_16003,N_16208);
xnor U16767 (N_16767,N_16429,N_16430);
and U16768 (N_16768,N_16220,N_16425);
xor U16769 (N_16769,N_16172,N_16400);
nor U16770 (N_16770,N_16188,N_16028);
and U16771 (N_16771,N_16017,N_16458);
xnor U16772 (N_16772,N_16174,N_16256);
and U16773 (N_16773,N_16140,N_16155);
nor U16774 (N_16774,N_16392,N_16468);
or U16775 (N_16775,N_16267,N_16444);
xnor U16776 (N_16776,N_16438,N_16123);
and U16777 (N_16777,N_16350,N_16470);
and U16778 (N_16778,N_16370,N_16311);
and U16779 (N_16779,N_16080,N_16215);
nor U16780 (N_16780,N_16018,N_16107);
nor U16781 (N_16781,N_16474,N_16382);
xnor U16782 (N_16782,N_16171,N_16284);
xnor U16783 (N_16783,N_16055,N_16168);
nor U16784 (N_16784,N_16483,N_16144);
xnor U16785 (N_16785,N_16006,N_16127);
and U16786 (N_16786,N_16031,N_16444);
nor U16787 (N_16787,N_16295,N_16340);
xor U16788 (N_16788,N_16120,N_16108);
nand U16789 (N_16789,N_16331,N_16076);
and U16790 (N_16790,N_16090,N_16033);
and U16791 (N_16791,N_16203,N_16416);
and U16792 (N_16792,N_16279,N_16305);
or U16793 (N_16793,N_16070,N_16082);
and U16794 (N_16794,N_16010,N_16230);
nand U16795 (N_16795,N_16419,N_16181);
nand U16796 (N_16796,N_16399,N_16402);
and U16797 (N_16797,N_16000,N_16384);
nand U16798 (N_16798,N_16097,N_16456);
nor U16799 (N_16799,N_16099,N_16009);
or U16800 (N_16800,N_16220,N_16467);
and U16801 (N_16801,N_16073,N_16173);
nor U16802 (N_16802,N_16016,N_16163);
xnor U16803 (N_16803,N_16398,N_16495);
xnor U16804 (N_16804,N_16076,N_16089);
nand U16805 (N_16805,N_16417,N_16343);
nor U16806 (N_16806,N_16129,N_16144);
xor U16807 (N_16807,N_16333,N_16089);
nor U16808 (N_16808,N_16447,N_16112);
nand U16809 (N_16809,N_16052,N_16021);
nand U16810 (N_16810,N_16043,N_16053);
nor U16811 (N_16811,N_16312,N_16417);
nor U16812 (N_16812,N_16058,N_16419);
xnor U16813 (N_16813,N_16273,N_16336);
nand U16814 (N_16814,N_16425,N_16146);
nand U16815 (N_16815,N_16328,N_16478);
and U16816 (N_16816,N_16136,N_16196);
xor U16817 (N_16817,N_16070,N_16086);
or U16818 (N_16818,N_16197,N_16201);
or U16819 (N_16819,N_16045,N_16495);
nor U16820 (N_16820,N_16466,N_16050);
nand U16821 (N_16821,N_16304,N_16207);
or U16822 (N_16822,N_16024,N_16087);
xnor U16823 (N_16823,N_16222,N_16150);
or U16824 (N_16824,N_16157,N_16027);
nor U16825 (N_16825,N_16317,N_16458);
nor U16826 (N_16826,N_16056,N_16159);
xor U16827 (N_16827,N_16311,N_16494);
or U16828 (N_16828,N_16018,N_16032);
or U16829 (N_16829,N_16251,N_16242);
xnor U16830 (N_16830,N_16219,N_16404);
and U16831 (N_16831,N_16474,N_16303);
nor U16832 (N_16832,N_16248,N_16202);
nor U16833 (N_16833,N_16406,N_16038);
xnor U16834 (N_16834,N_16280,N_16304);
nor U16835 (N_16835,N_16222,N_16142);
xor U16836 (N_16836,N_16182,N_16146);
and U16837 (N_16837,N_16114,N_16487);
nand U16838 (N_16838,N_16040,N_16192);
nand U16839 (N_16839,N_16224,N_16213);
and U16840 (N_16840,N_16031,N_16308);
xor U16841 (N_16841,N_16468,N_16092);
nor U16842 (N_16842,N_16362,N_16341);
and U16843 (N_16843,N_16486,N_16094);
or U16844 (N_16844,N_16131,N_16116);
nand U16845 (N_16845,N_16248,N_16066);
xnor U16846 (N_16846,N_16494,N_16284);
nor U16847 (N_16847,N_16264,N_16216);
xor U16848 (N_16848,N_16241,N_16006);
or U16849 (N_16849,N_16113,N_16197);
nand U16850 (N_16850,N_16293,N_16376);
or U16851 (N_16851,N_16493,N_16368);
and U16852 (N_16852,N_16343,N_16477);
nor U16853 (N_16853,N_16496,N_16261);
nand U16854 (N_16854,N_16408,N_16099);
nor U16855 (N_16855,N_16127,N_16097);
and U16856 (N_16856,N_16445,N_16078);
nand U16857 (N_16857,N_16351,N_16310);
nand U16858 (N_16858,N_16488,N_16348);
xnor U16859 (N_16859,N_16008,N_16281);
nand U16860 (N_16860,N_16347,N_16429);
xor U16861 (N_16861,N_16151,N_16060);
and U16862 (N_16862,N_16003,N_16394);
nor U16863 (N_16863,N_16117,N_16095);
or U16864 (N_16864,N_16123,N_16105);
and U16865 (N_16865,N_16218,N_16426);
xnor U16866 (N_16866,N_16149,N_16184);
and U16867 (N_16867,N_16345,N_16497);
and U16868 (N_16868,N_16099,N_16222);
or U16869 (N_16869,N_16229,N_16010);
and U16870 (N_16870,N_16492,N_16396);
and U16871 (N_16871,N_16021,N_16117);
nor U16872 (N_16872,N_16016,N_16474);
nand U16873 (N_16873,N_16021,N_16151);
nor U16874 (N_16874,N_16132,N_16128);
xor U16875 (N_16875,N_16181,N_16418);
and U16876 (N_16876,N_16145,N_16305);
nor U16877 (N_16877,N_16148,N_16486);
xnor U16878 (N_16878,N_16495,N_16131);
xnor U16879 (N_16879,N_16100,N_16413);
xor U16880 (N_16880,N_16013,N_16445);
or U16881 (N_16881,N_16199,N_16212);
nand U16882 (N_16882,N_16493,N_16202);
and U16883 (N_16883,N_16452,N_16200);
nor U16884 (N_16884,N_16421,N_16028);
or U16885 (N_16885,N_16398,N_16197);
nor U16886 (N_16886,N_16000,N_16263);
nor U16887 (N_16887,N_16130,N_16319);
xor U16888 (N_16888,N_16082,N_16053);
nor U16889 (N_16889,N_16357,N_16393);
or U16890 (N_16890,N_16101,N_16281);
nor U16891 (N_16891,N_16215,N_16433);
xnor U16892 (N_16892,N_16283,N_16276);
nand U16893 (N_16893,N_16458,N_16020);
xor U16894 (N_16894,N_16333,N_16345);
xor U16895 (N_16895,N_16243,N_16381);
nor U16896 (N_16896,N_16325,N_16429);
or U16897 (N_16897,N_16401,N_16410);
nor U16898 (N_16898,N_16371,N_16226);
nor U16899 (N_16899,N_16011,N_16390);
xor U16900 (N_16900,N_16292,N_16078);
and U16901 (N_16901,N_16080,N_16081);
and U16902 (N_16902,N_16229,N_16092);
xnor U16903 (N_16903,N_16330,N_16399);
or U16904 (N_16904,N_16302,N_16412);
and U16905 (N_16905,N_16437,N_16215);
nand U16906 (N_16906,N_16050,N_16344);
xor U16907 (N_16907,N_16499,N_16279);
xor U16908 (N_16908,N_16006,N_16044);
nor U16909 (N_16909,N_16199,N_16311);
or U16910 (N_16910,N_16218,N_16325);
nor U16911 (N_16911,N_16462,N_16291);
or U16912 (N_16912,N_16177,N_16052);
nor U16913 (N_16913,N_16120,N_16225);
or U16914 (N_16914,N_16254,N_16229);
or U16915 (N_16915,N_16264,N_16417);
xnor U16916 (N_16916,N_16482,N_16408);
and U16917 (N_16917,N_16257,N_16416);
xor U16918 (N_16918,N_16421,N_16447);
nand U16919 (N_16919,N_16413,N_16340);
xnor U16920 (N_16920,N_16248,N_16135);
and U16921 (N_16921,N_16124,N_16475);
xor U16922 (N_16922,N_16115,N_16030);
and U16923 (N_16923,N_16181,N_16465);
nor U16924 (N_16924,N_16179,N_16449);
nand U16925 (N_16925,N_16141,N_16170);
nand U16926 (N_16926,N_16391,N_16397);
and U16927 (N_16927,N_16383,N_16407);
xor U16928 (N_16928,N_16036,N_16102);
nor U16929 (N_16929,N_16177,N_16394);
and U16930 (N_16930,N_16120,N_16124);
nor U16931 (N_16931,N_16405,N_16499);
and U16932 (N_16932,N_16499,N_16059);
nand U16933 (N_16933,N_16325,N_16216);
nor U16934 (N_16934,N_16311,N_16117);
or U16935 (N_16935,N_16323,N_16175);
and U16936 (N_16936,N_16327,N_16115);
nand U16937 (N_16937,N_16020,N_16005);
nand U16938 (N_16938,N_16267,N_16270);
nor U16939 (N_16939,N_16348,N_16482);
xnor U16940 (N_16940,N_16388,N_16163);
and U16941 (N_16941,N_16494,N_16003);
and U16942 (N_16942,N_16050,N_16102);
and U16943 (N_16943,N_16335,N_16222);
nor U16944 (N_16944,N_16198,N_16357);
nor U16945 (N_16945,N_16077,N_16123);
xor U16946 (N_16946,N_16102,N_16150);
nand U16947 (N_16947,N_16202,N_16298);
and U16948 (N_16948,N_16303,N_16398);
xor U16949 (N_16949,N_16415,N_16301);
or U16950 (N_16950,N_16443,N_16481);
xor U16951 (N_16951,N_16268,N_16047);
nor U16952 (N_16952,N_16074,N_16164);
nor U16953 (N_16953,N_16412,N_16333);
or U16954 (N_16954,N_16045,N_16200);
and U16955 (N_16955,N_16025,N_16032);
nor U16956 (N_16956,N_16312,N_16296);
nand U16957 (N_16957,N_16009,N_16200);
or U16958 (N_16958,N_16321,N_16403);
xor U16959 (N_16959,N_16163,N_16343);
or U16960 (N_16960,N_16233,N_16285);
nor U16961 (N_16961,N_16226,N_16435);
xor U16962 (N_16962,N_16424,N_16494);
nor U16963 (N_16963,N_16422,N_16430);
nand U16964 (N_16964,N_16217,N_16425);
and U16965 (N_16965,N_16393,N_16136);
or U16966 (N_16966,N_16435,N_16294);
nor U16967 (N_16967,N_16299,N_16038);
xor U16968 (N_16968,N_16003,N_16064);
nor U16969 (N_16969,N_16345,N_16089);
or U16970 (N_16970,N_16278,N_16165);
and U16971 (N_16971,N_16237,N_16093);
xnor U16972 (N_16972,N_16011,N_16292);
nor U16973 (N_16973,N_16361,N_16262);
nor U16974 (N_16974,N_16163,N_16437);
and U16975 (N_16975,N_16447,N_16364);
nand U16976 (N_16976,N_16269,N_16112);
nand U16977 (N_16977,N_16298,N_16106);
xor U16978 (N_16978,N_16164,N_16374);
nand U16979 (N_16979,N_16279,N_16459);
xor U16980 (N_16980,N_16046,N_16320);
xnor U16981 (N_16981,N_16375,N_16094);
xnor U16982 (N_16982,N_16094,N_16265);
xnor U16983 (N_16983,N_16498,N_16369);
xor U16984 (N_16984,N_16286,N_16261);
nand U16985 (N_16985,N_16208,N_16449);
nor U16986 (N_16986,N_16217,N_16428);
nor U16987 (N_16987,N_16455,N_16421);
or U16988 (N_16988,N_16393,N_16238);
nand U16989 (N_16989,N_16013,N_16119);
nor U16990 (N_16990,N_16468,N_16193);
or U16991 (N_16991,N_16252,N_16089);
nand U16992 (N_16992,N_16414,N_16156);
nor U16993 (N_16993,N_16497,N_16221);
nor U16994 (N_16994,N_16361,N_16305);
or U16995 (N_16995,N_16018,N_16013);
or U16996 (N_16996,N_16007,N_16333);
and U16997 (N_16997,N_16486,N_16350);
and U16998 (N_16998,N_16281,N_16052);
xor U16999 (N_16999,N_16279,N_16264);
nand U17000 (N_17000,N_16589,N_16907);
or U17001 (N_17001,N_16980,N_16902);
nand U17002 (N_17002,N_16716,N_16765);
nor U17003 (N_17003,N_16813,N_16603);
nand U17004 (N_17004,N_16837,N_16674);
and U17005 (N_17005,N_16804,N_16541);
or U17006 (N_17006,N_16672,N_16618);
or U17007 (N_17007,N_16789,N_16905);
or U17008 (N_17008,N_16525,N_16664);
nor U17009 (N_17009,N_16501,N_16788);
and U17010 (N_17010,N_16536,N_16696);
and U17011 (N_17011,N_16998,N_16706);
nand U17012 (N_17012,N_16947,N_16909);
nor U17013 (N_17013,N_16744,N_16683);
or U17014 (N_17014,N_16883,N_16671);
and U17015 (N_17015,N_16967,N_16896);
nor U17016 (N_17016,N_16955,N_16577);
or U17017 (N_17017,N_16820,N_16818);
nor U17018 (N_17018,N_16926,N_16780);
nand U17019 (N_17019,N_16686,N_16502);
nand U17020 (N_17020,N_16522,N_16785);
xor U17021 (N_17021,N_16509,N_16771);
or U17022 (N_17022,N_16638,N_16935);
nand U17023 (N_17023,N_16931,N_16613);
and U17024 (N_17024,N_16971,N_16985);
or U17025 (N_17025,N_16938,N_16793);
or U17026 (N_17026,N_16977,N_16772);
and U17027 (N_17027,N_16611,N_16957);
and U17028 (N_17028,N_16619,N_16946);
nor U17029 (N_17029,N_16500,N_16911);
nand U17030 (N_17030,N_16861,N_16827);
nor U17031 (N_17031,N_16572,N_16960);
nor U17032 (N_17032,N_16973,N_16610);
xnor U17033 (N_17033,N_16524,N_16503);
or U17034 (N_17034,N_16505,N_16677);
or U17035 (N_17035,N_16760,N_16699);
nand U17036 (N_17036,N_16682,N_16615);
nor U17037 (N_17037,N_16836,N_16616);
xnor U17038 (N_17038,N_16758,N_16568);
xor U17039 (N_17039,N_16727,N_16679);
and U17040 (N_17040,N_16890,N_16702);
xor U17041 (N_17041,N_16959,N_16596);
nand U17042 (N_17042,N_16571,N_16825);
xor U17043 (N_17043,N_16995,N_16845);
and U17044 (N_17044,N_16885,N_16529);
or U17045 (N_17045,N_16752,N_16792);
nand U17046 (N_17046,N_16592,N_16530);
nand U17047 (N_17047,N_16652,N_16533);
nand U17048 (N_17048,N_16757,N_16940);
nor U17049 (N_17049,N_16704,N_16745);
nor U17050 (N_17050,N_16711,N_16715);
or U17051 (N_17051,N_16848,N_16874);
xnor U17052 (N_17052,N_16846,N_16988);
or U17053 (N_17053,N_16520,N_16647);
nand U17054 (N_17054,N_16733,N_16554);
nand U17055 (N_17055,N_16510,N_16979);
nand U17056 (N_17056,N_16651,N_16630);
or U17057 (N_17057,N_16976,N_16857);
or U17058 (N_17058,N_16910,N_16504);
nand U17059 (N_17059,N_16642,N_16769);
nor U17060 (N_17060,N_16653,N_16763);
nor U17061 (N_17061,N_16969,N_16599);
and U17062 (N_17062,N_16670,N_16643);
xnor U17063 (N_17063,N_16790,N_16594);
nand U17064 (N_17064,N_16842,N_16843);
xnor U17065 (N_17065,N_16767,N_16717);
nand U17066 (N_17066,N_16739,N_16864);
nor U17067 (N_17067,N_16514,N_16564);
xor U17068 (N_17068,N_16741,N_16990);
xnor U17069 (N_17069,N_16644,N_16560);
or U17070 (N_17070,N_16558,N_16597);
or U17071 (N_17071,N_16802,N_16863);
nand U17072 (N_17072,N_16736,N_16889);
and U17073 (N_17073,N_16588,N_16662);
and U17074 (N_17074,N_16943,N_16878);
nor U17075 (N_17075,N_16847,N_16828);
xnor U17076 (N_17076,N_16612,N_16581);
xnor U17077 (N_17077,N_16856,N_16685);
nand U17078 (N_17078,N_16915,N_16567);
nand U17079 (N_17079,N_16726,N_16645);
and U17080 (N_17080,N_16707,N_16838);
and U17081 (N_17081,N_16557,N_16867);
or U17082 (N_17082,N_16584,N_16556);
nor U17083 (N_17083,N_16582,N_16776);
nand U17084 (N_17084,N_16703,N_16797);
or U17085 (N_17085,N_16851,N_16900);
xor U17086 (N_17086,N_16994,N_16839);
xor U17087 (N_17087,N_16562,N_16724);
and U17088 (N_17088,N_16552,N_16928);
xnor U17089 (N_17089,N_16812,N_16869);
nand U17090 (N_17090,N_16698,N_16866);
nor U17091 (N_17091,N_16929,N_16640);
nor U17092 (N_17092,N_16508,N_16690);
xnor U17093 (N_17093,N_16840,N_16538);
nand U17094 (N_17094,N_16543,N_16519);
nor U17095 (N_17095,N_16748,N_16873);
or U17096 (N_17096,N_16849,N_16753);
xor U17097 (N_17097,N_16799,N_16852);
or U17098 (N_17098,N_16815,N_16806);
nand U17099 (N_17099,N_16924,N_16937);
and U17100 (N_17100,N_16854,N_16553);
and U17101 (N_17101,N_16656,N_16999);
and U17102 (N_17102,N_16563,N_16834);
or U17103 (N_17103,N_16921,N_16949);
nand U17104 (N_17104,N_16676,N_16775);
nor U17105 (N_17105,N_16578,N_16574);
or U17106 (N_17106,N_16822,N_16819);
and U17107 (N_17107,N_16648,N_16930);
nand U17108 (N_17108,N_16958,N_16824);
nand U17109 (N_17109,N_16646,N_16660);
xnor U17110 (N_17110,N_16996,N_16912);
xor U17111 (N_17111,N_16963,N_16617);
nand U17112 (N_17112,N_16579,N_16983);
nor U17113 (N_17113,N_16532,N_16941);
xor U17114 (N_17114,N_16901,N_16925);
xor U17115 (N_17115,N_16576,N_16721);
nand U17116 (N_17116,N_16986,N_16922);
nand U17117 (N_17117,N_16665,N_16629);
xnor U17118 (N_17118,N_16991,N_16535);
xor U17119 (N_17119,N_16904,N_16876);
nor U17120 (N_17120,N_16942,N_16561);
and U17121 (N_17121,N_16808,N_16787);
nor U17122 (N_17122,N_16580,N_16691);
xnor U17123 (N_17123,N_16607,N_16829);
nand U17124 (N_17124,N_16573,N_16962);
nor U17125 (N_17125,N_16987,N_16666);
or U17126 (N_17126,N_16518,N_16527);
nor U17127 (N_17127,N_16766,N_16654);
and U17128 (N_17128,N_16540,N_16982);
or U17129 (N_17129,N_16583,N_16626);
nand U17130 (N_17130,N_16981,N_16749);
nand U17131 (N_17131,N_16585,N_16517);
or U17132 (N_17132,N_16868,N_16590);
xnor U17133 (N_17133,N_16528,N_16779);
nand U17134 (N_17134,N_16534,N_16545);
xor U17135 (N_17135,N_16693,N_16650);
and U17136 (N_17136,N_16547,N_16521);
or U17137 (N_17137,N_16742,N_16855);
nor U17138 (N_17138,N_16669,N_16860);
nor U17139 (N_17139,N_16784,N_16743);
and U17140 (N_17140,N_16723,N_16841);
nor U17141 (N_17141,N_16953,N_16768);
nor U17142 (N_17142,N_16516,N_16734);
or U17143 (N_17143,N_16908,N_16796);
xor U17144 (N_17144,N_16906,N_16968);
xnor U17145 (N_17145,N_16695,N_16884);
nand U17146 (N_17146,N_16718,N_16531);
nand U17147 (N_17147,N_16526,N_16899);
or U17148 (N_17148,N_16879,N_16978);
or U17149 (N_17149,N_16635,N_16692);
xor U17150 (N_17150,N_16798,N_16800);
xnor U17151 (N_17151,N_16762,N_16606);
nand U17152 (N_17152,N_16759,N_16895);
nand U17153 (N_17153,N_16725,N_16892);
xor U17154 (N_17154,N_16663,N_16515);
nor U17155 (N_17155,N_16903,N_16546);
nand U17156 (N_17156,N_16641,N_16891);
nor U17157 (N_17157,N_16795,N_16777);
and U17158 (N_17158,N_16713,N_16786);
nor U17159 (N_17159,N_16731,N_16810);
and U17160 (N_17160,N_16507,N_16627);
nor U17161 (N_17161,N_16701,N_16913);
and U17162 (N_17162,N_16887,N_16655);
nor U17163 (N_17163,N_16992,N_16625);
nand U17164 (N_17164,N_16551,N_16659);
or U17165 (N_17165,N_16951,N_16512);
or U17166 (N_17166,N_16565,N_16722);
nand U17167 (N_17167,N_16623,N_16523);
and U17168 (N_17168,N_16897,N_16833);
or U17169 (N_17169,N_16729,N_16542);
nor U17170 (N_17170,N_16694,N_16712);
nor U17171 (N_17171,N_16673,N_16948);
or U17172 (N_17172,N_16865,N_16681);
nand U17173 (N_17173,N_16614,N_16919);
nand U17174 (N_17174,N_16939,N_16700);
nor U17175 (N_17175,N_16956,N_16756);
and U17176 (N_17176,N_16816,N_16705);
or U17177 (N_17177,N_16680,N_16972);
or U17178 (N_17178,N_16950,N_16595);
and U17179 (N_17179,N_16550,N_16933);
and U17180 (N_17180,N_16805,N_16920);
or U17181 (N_17181,N_16738,N_16831);
nor U17182 (N_17182,N_16608,N_16661);
nor U17183 (N_17183,N_16945,N_16587);
nor U17184 (N_17184,N_16778,N_16811);
and U17185 (N_17185,N_16728,N_16675);
and U17186 (N_17186,N_16814,N_16888);
and U17187 (N_17187,N_16932,N_16821);
and U17188 (N_17188,N_16601,N_16761);
or U17189 (N_17189,N_16871,N_16850);
or U17190 (N_17190,N_16886,N_16853);
xor U17191 (N_17191,N_16602,N_16894);
and U17192 (N_17192,N_16774,N_16559);
xor U17193 (N_17193,N_16997,N_16737);
xor U17194 (N_17194,N_16624,N_16746);
xor U17195 (N_17195,N_16605,N_16586);
nand U17196 (N_17196,N_16993,N_16506);
and U17197 (N_17197,N_16549,N_16697);
nand U17198 (N_17198,N_16591,N_16604);
xnor U17199 (N_17199,N_16791,N_16730);
and U17200 (N_17200,N_16575,N_16844);
or U17201 (N_17201,N_16639,N_16667);
nand U17202 (N_17202,N_16832,N_16794);
nand U17203 (N_17203,N_16875,N_16764);
xor U17204 (N_17204,N_16881,N_16633);
and U17205 (N_17205,N_16918,N_16637);
and U17206 (N_17206,N_16750,N_16513);
or U17207 (N_17207,N_16877,N_16593);
or U17208 (N_17208,N_16975,N_16747);
xor U17209 (N_17209,N_16803,N_16740);
nor U17210 (N_17210,N_16966,N_16658);
or U17211 (N_17211,N_16773,N_16751);
and U17212 (N_17212,N_16898,N_16684);
nor U17213 (N_17213,N_16688,N_16830);
nand U17214 (N_17214,N_16555,N_16870);
and U17215 (N_17215,N_16923,N_16936);
xnor U17216 (N_17216,N_16916,N_16801);
or U17217 (N_17217,N_16719,N_16754);
xnor U17218 (N_17218,N_16622,N_16539);
nor U17219 (N_17219,N_16970,N_16961);
nand U17220 (N_17220,N_16974,N_16710);
or U17221 (N_17221,N_16632,N_16954);
nor U17222 (N_17222,N_16755,N_16634);
nand U17223 (N_17223,N_16649,N_16783);
xnor U17224 (N_17224,N_16735,N_16858);
or U17225 (N_17225,N_16770,N_16859);
and U17226 (N_17226,N_16678,N_16708);
or U17227 (N_17227,N_16823,N_16570);
xor U17228 (N_17228,N_16984,N_16989);
xnor U17229 (N_17229,N_16620,N_16668);
nand U17230 (N_17230,N_16826,N_16598);
nand U17231 (N_17231,N_16809,N_16714);
xnor U17232 (N_17232,N_16709,N_16927);
nor U17233 (N_17233,N_16537,N_16862);
and U17234 (N_17234,N_16817,N_16781);
or U17235 (N_17235,N_16566,N_16934);
nand U17236 (N_17236,N_16511,N_16569);
and U17237 (N_17237,N_16600,N_16882);
and U17238 (N_17238,N_16628,N_16544);
xnor U17239 (N_17239,N_16621,N_16631);
xnor U17240 (N_17240,N_16893,N_16689);
xor U17241 (N_17241,N_16636,N_16687);
xor U17242 (N_17242,N_16917,N_16880);
or U17243 (N_17243,N_16964,N_16657);
and U17244 (N_17244,N_16872,N_16835);
or U17245 (N_17245,N_16914,N_16548);
nand U17246 (N_17246,N_16965,N_16720);
xor U17247 (N_17247,N_16952,N_16609);
and U17248 (N_17248,N_16944,N_16732);
or U17249 (N_17249,N_16782,N_16807);
nor U17250 (N_17250,N_16788,N_16953);
and U17251 (N_17251,N_16804,N_16671);
nand U17252 (N_17252,N_16960,N_16659);
or U17253 (N_17253,N_16605,N_16634);
and U17254 (N_17254,N_16665,N_16792);
or U17255 (N_17255,N_16907,N_16597);
and U17256 (N_17256,N_16821,N_16777);
nor U17257 (N_17257,N_16755,N_16808);
or U17258 (N_17258,N_16844,N_16559);
or U17259 (N_17259,N_16838,N_16976);
nor U17260 (N_17260,N_16520,N_16755);
and U17261 (N_17261,N_16802,N_16522);
xnor U17262 (N_17262,N_16689,N_16592);
and U17263 (N_17263,N_16548,N_16858);
nor U17264 (N_17264,N_16974,N_16625);
nor U17265 (N_17265,N_16969,N_16638);
nand U17266 (N_17266,N_16716,N_16766);
nand U17267 (N_17267,N_16980,N_16604);
nand U17268 (N_17268,N_16558,N_16514);
xnor U17269 (N_17269,N_16924,N_16984);
nor U17270 (N_17270,N_16937,N_16779);
or U17271 (N_17271,N_16528,N_16751);
or U17272 (N_17272,N_16771,N_16715);
nor U17273 (N_17273,N_16727,N_16925);
nor U17274 (N_17274,N_16613,N_16903);
nor U17275 (N_17275,N_16883,N_16913);
nand U17276 (N_17276,N_16770,N_16881);
or U17277 (N_17277,N_16814,N_16809);
xnor U17278 (N_17278,N_16545,N_16838);
and U17279 (N_17279,N_16825,N_16900);
xnor U17280 (N_17280,N_16541,N_16713);
or U17281 (N_17281,N_16572,N_16529);
and U17282 (N_17282,N_16822,N_16717);
nand U17283 (N_17283,N_16600,N_16990);
nand U17284 (N_17284,N_16893,N_16557);
nor U17285 (N_17285,N_16966,N_16994);
or U17286 (N_17286,N_16959,N_16576);
nand U17287 (N_17287,N_16725,N_16872);
or U17288 (N_17288,N_16944,N_16733);
nand U17289 (N_17289,N_16684,N_16899);
xor U17290 (N_17290,N_16753,N_16630);
nor U17291 (N_17291,N_16527,N_16510);
nand U17292 (N_17292,N_16991,N_16560);
xor U17293 (N_17293,N_16762,N_16580);
xor U17294 (N_17294,N_16596,N_16551);
nand U17295 (N_17295,N_16611,N_16884);
xnor U17296 (N_17296,N_16782,N_16942);
nand U17297 (N_17297,N_16515,N_16753);
and U17298 (N_17298,N_16739,N_16894);
and U17299 (N_17299,N_16609,N_16655);
nor U17300 (N_17300,N_16757,N_16881);
nand U17301 (N_17301,N_16992,N_16785);
nand U17302 (N_17302,N_16660,N_16708);
nor U17303 (N_17303,N_16993,N_16521);
nand U17304 (N_17304,N_16544,N_16807);
and U17305 (N_17305,N_16946,N_16577);
xnor U17306 (N_17306,N_16522,N_16929);
xor U17307 (N_17307,N_16948,N_16983);
nand U17308 (N_17308,N_16776,N_16688);
nor U17309 (N_17309,N_16607,N_16990);
nor U17310 (N_17310,N_16648,N_16762);
xnor U17311 (N_17311,N_16543,N_16629);
nor U17312 (N_17312,N_16798,N_16563);
nor U17313 (N_17313,N_16923,N_16586);
nand U17314 (N_17314,N_16752,N_16797);
nor U17315 (N_17315,N_16849,N_16515);
xnor U17316 (N_17316,N_16541,N_16526);
or U17317 (N_17317,N_16696,N_16719);
nand U17318 (N_17318,N_16889,N_16765);
or U17319 (N_17319,N_16588,N_16759);
and U17320 (N_17320,N_16877,N_16545);
and U17321 (N_17321,N_16614,N_16672);
nand U17322 (N_17322,N_16822,N_16646);
nand U17323 (N_17323,N_16740,N_16884);
nand U17324 (N_17324,N_16794,N_16667);
and U17325 (N_17325,N_16931,N_16520);
nand U17326 (N_17326,N_16911,N_16920);
nand U17327 (N_17327,N_16752,N_16836);
or U17328 (N_17328,N_16654,N_16845);
or U17329 (N_17329,N_16811,N_16921);
and U17330 (N_17330,N_16965,N_16685);
and U17331 (N_17331,N_16653,N_16966);
nor U17332 (N_17332,N_16950,N_16547);
xor U17333 (N_17333,N_16891,N_16876);
and U17334 (N_17334,N_16968,N_16639);
xnor U17335 (N_17335,N_16645,N_16800);
nand U17336 (N_17336,N_16537,N_16770);
xnor U17337 (N_17337,N_16719,N_16665);
and U17338 (N_17338,N_16976,N_16681);
nand U17339 (N_17339,N_16537,N_16779);
or U17340 (N_17340,N_16647,N_16758);
or U17341 (N_17341,N_16640,N_16889);
nor U17342 (N_17342,N_16815,N_16833);
xor U17343 (N_17343,N_16507,N_16630);
nor U17344 (N_17344,N_16855,N_16941);
and U17345 (N_17345,N_16536,N_16669);
and U17346 (N_17346,N_16778,N_16700);
nand U17347 (N_17347,N_16696,N_16695);
and U17348 (N_17348,N_16832,N_16583);
or U17349 (N_17349,N_16726,N_16997);
or U17350 (N_17350,N_16823,N_16995);
nand U17351 (N_17351,N_16766,N_16872);
nand U17352 (N_17352,N_16771,N_16746);
nand U17353 (N_17353,N_16999,N_16623);
nor U17354 (N_17354,N_16908,N_16640);
nor U17355 (N_17355,N_16703,N_16806);
or U17356 (N_17356,N_16953,N_16824);
nand U17357 (N_17357,N_16571,N_16525);
or U17358 (N_17358,N_16893,N_16994);
xor U17359 (N_17359,N_16560,N_16879);
and U17360 (N_17360,N_16985,N_16633);
xnor U17361 (N_17361,N_16821,N_16957);
and U17362 (N_17362,N_16757,N_16761);
and U17363 (N_17363,N_16717,N_16814);
xor U17364 (N_17364,N_16675,N_16961);
or U17365 (N_17365,N_16909,N_16632);
and U17366 (N_17366,N_16771,N_16902);
and U17367 (N_17367,N_16861,N_16790);
nand U17368 (N_17368,N_16860,N_16986);
nor U17369 (N_17369,N_16889,N_16993);
xor U17370 (N_17370,N_16855,N_16817);
nand U17371 (N_17371,N_16641,N_16572);
and U17372 (N_17372,N_16695,N_16527);
and U17373 (N_17373,N_16957,N_16999);
nand U17374 (N_17374,N_16723,N_16960);
and U17375 (N_17375,N_16539,N_16925);
nor U17376 (N_17376,N_16900,N_16910);
xor U17377 (N_17377,N_16648,N_16622);
or U17378 (N_17378,N_16924,N_16918);
nand U17379 (N_17379,N_16593,N_16867);
xor U17380 (N_17380,N_16875,N_16549);
and U17381 (N_17381,N_16853,N_16594);
or U17382 (N_17382,N_16662,N_16674);
and U17383 (N_17383,N_16649,N_16534);
nor U17384 (N_17384,N_16836,N_16604);
nor U17385 (N_17385,N_16871,N_16949);
and U17386 (N_17386,N_16530,N_16765);
nand U17387 (N_17387,N_16650,N_16648);
nand U17388 (N_17388,N_16845,N_16738);
or U17389 (N_17389,N_16528,N_16594);
xnor U17390 (N_17390,N_16589,N_16675);
or U17391 (N_17391,N_16559,N_16824);
or U17392 (N_17392,N_16959,N_16758);
nand U17393 (N_17393,N_16684,N_16783);
xor U17394 (N_17394,N_16986,N_16534);
xor U17395 (N_17395,N_16963,N_16769);
nor U17396 (N_17396,N_16578,N_16559);
and U17397 (N_17397,N_16782,N_16509);
or U17398 (N_17398,N_16615,N_16873);
or U17399 (N_17399,N_16811,N_16838);
and U17400 (N_17400,N_16755,N_16751);
or U17401 (N_17401,N_16530,N_16782);
and U17402 (N_17402,N_16839,N_16734);
and U17403 (N_17403,N_16621,N_16629);
or U17404 (N_17404,N_16882,N_16834);
or U17405 (N_17405,N_16971,N_16759);
xnor U17406 (N_17406,N_16555,N_16517);
nor U17407 (N_17407,N_16717,N_16771);
nor U17408 (N_17408,N_16660,N_16964);
xor U17409 (N_17409,N_16799,N_16921);
nor U17410 (N_17410,N_16863,N_16762);
and U17411 (N_17411,N_16907,N_16660);
nor U17412 (N_17412,N_16584,N_16948);
and U17413 (N_17413,N_16965,N_16795);
nor U17414 (N_17414,N_16754,N_16730);
nand U17415 (N_17415,N_16725,N_16705);
nor U17416 (N_17416,N_16809,N_16668);
nor U17417 (N_17417,N_16805,N_16739);
and U17418 (N_17418,N_16706,N_16982);
and U17419 (N_17419,N_16637,N_16816);
or U17420 (N_17420,N_16565,N_16979);
and U17421 (N_17421,N_16851,N_16847);
nor U17422 (N_17422,N_16756,N_16777);
xor U17423 (N_17423,N_16508,N_16975);
nor U17424 (N_17424,N_16977,N_16849);
xor U17425 (N_17425,N_16686,N_16997);
nor U17426 (N_17426,N_16589,N_16781);
and U17427 (N_17427,N_16537,N_16906);
xor U17428 (N_17428,N_16772,N_16928);
xor U17429 (N_17429,N_16678,N_16734);
or U17430 (N_17430,N_16680,N_16744);
and U17431 (N_17431,N_16943,N_16968);
nor U17432 (N_17432,N_16790,N_16989);
nand U17433 (N_17433,N_16574,N_16776);
nand U17434 (N_17434,N_16893,N_16861);
nor U17435 (N_17435,N_16867,N_16828);
and U17436 (N_17436,N_16890,N_16620);
or U17437 (N_17437,N_16651,N_16922);
or U17438 (N_17438,N_16699,N_16987);
nor U17439 (N_17439,N_16518,N_16844);
nand U17440 (N_17440,N_16600,N_16608);
xor U17441 (N_17441,N_16559,N_16511);
and U17442 (N_17442,N_16794,N_16886);
nor U17443 (N_17443,N_16693,N_16801);
and U17444 (N_17444,N_16988,N_16665);
xor U17445 (N_17445,N_16559,N_16847);
nand U17446 (N_17446,N_16829,N_16837);
nor U17447 (N_17447,N_16804,N_16877);
and U17448 (N_17448,N_16938,N_16883);
nand U17449 (N_17449,N_16900,N_16911);
and U17450 (N_17450,N_16701,N_16667);
or U17451 (N_17451,N_16869,N_16737);
and U17452 (N_17452,N_16552,N_16749);
xnor U17453 (N_17453,N_16670,N_16523);
and U17454 (N_17454,N_16920,N_16643);
or U17455 (N_17455,N_16653,N_16993);
or U17456 (N_17456,N_16787,N_16819);
xnor U17457 (N_17457,N_16626,N_16836);
nor U17458 (N_17458,N_16791,N_16660);
and U17459 (N_17459,N_16811,N_16973);
or U17460 (N_17460,N_16979,N_16555);
nor U17461 (N_17461,N_16759,N_16808);
nand U17462 (N_17462,N_16521,N_16833);
nand U17463 (N_17463,N_16505,N_16881);
or U17464 (N_17464,N_16923,N_16549);
and U17465 (N_17465,N_16875,N_16767);
nand U17466 (N_17466,N_16800,N_16937);
nor U17467 (N_17467,N_16853,N_16739);
nor U17468 (N_17468,N_16603,N_16664);
nand U17469 (N_17469,N_16821,N_16810);
xor U17470 (N_17470,N_16790,N_16715);
nand U17471 (N_17471,N_16900,N_16891);
or U17472 (N_17472,N_16561,N_16771);
nand U17473 (N_17473,N_16863,N_16645);
nand U17474 (N_17474,N_16584,N_16676);
and U17475 (N_17475,N_16503,N_16975);
or U17476 (N_17476,N_16654,N_16815);
nand U17477 (N_17477,N_16813,N_16533);
and U17478 (N_17478,N_16995,N_16980);
nor U17479 (N_17479,N_16810,N_16596);
and U17480 (N_17480,N_16969,N_16653);
nand U17481 (N_17481,N_16698,N_16918);
nor U17482 (N_17482,N_16950,N_16518);
and U17483 (N_17483,N_16505,N_16613);
and U17484 (N_17484,N_16618,N_16581);
nand U17485 (N_17485,N_16869,N_16521);
nor U17486 (N_17486,N_16712,N_16613);
or U17487 (N_17487,N_16999,N_16969);
nor U17488 (N_17488,N_16907,N_16812);
or U17489 (N_17489,N_16562,N_16515);
nand U17490 (N_17490,N_16697,N_16698);
and U17491 (N_17491,N_16803,N_16917);
xnor U17492 (N_17492,N_16696,N_16679);
nand U17493 (N_17493,N_16574,N_16559);
xor U17494 (N_17494,N_16619,N_16705);
xnor U17495 (N_17495,N_16664,N_16887);
and U17496 (N_17496,N_16875,N_16652);
xor U17497 (N_17497,N_16678,N_16526);
and U17498 (N_17498,N_16893,N_16826);
or U17499 (N_17499,N_16720,N_16962);
xnor U17500 (N_17500,N_17072,N_17071);
nand U17501 (N_17501,N_17094,N_17223);
and U17502 (N_17502,N_17300,N_17386);
xor U17503 (N_17503,N_17265,N_17290);
nand U17504 (N_17504,N_17384,N_17417);
and U17505 (N_17505,N_17325,N_17160);
and U17506 (N_17506,N_17061,N_17497);
nand U17507 (N_17507,N_17331,N_17237);
xor U17508 (N_17508,N_17430,N_17239);
nand U17509 (N_17509,N_17316,N_17016);
or U17510 (N_17510,N_17208,N_17057);
and U17511 (N_17511,N_17197,N_17367);
nand U17512 (N_17512,N_17264,N_17204);
xnor U17513 (N_17513,N_17083,N_17442);
xor U17514 (N_17514,N_17099,N_17104);
nor U17515 (N_17515,N_17284,N_17117);
or U17516 (N_17516,N_17110,N_17196);
nand U17517 (N_17517,N_17076,N_17496);
xor U17518 (N_17518,N_17470,N_17089);
or U17519 (N_17519,N_17073,N_17093);
and U17520 (N_17520,N_17411,N_17010);
xnor U17521 (N_17521,N_17182,N_17238);
or U17522 (N_17522,N_17378,N_17092);
and U17523 (N_17523,N_17233,N_17294);
nand U17524 (N_17524,N_17306,N_17123);
nor U17525 (N_17525,N_17224,N_17003);
nand U17526 (N_17526,N_17486,N_17293);
nor U17527 (N_17527,N_17419,N_17254);
nand U17528 (N_17528,N_17203,N_17102);
or U17529 (N_17529,N_17198,N_17079);
xnor U17530 (N_17530,N_17312,N_17049);
nor U17531 (N_17531,N_17370,N_17122);
or U17532 (N_17532,N_17002,N_17267);
nor U17533 (N_17533,N_17303,N_17052);
and U17534 (N_17534,N_17460,N_17200);
or U17535 (N_17535,N_17206,N_17188);
or U17536 (N_17536,N_17077,N_17458);
nand U17537 (N_17537,N_17229,N_17056);
and U17538 (N_17538,N_17462,N_17365);
or U17539 (N_17539,N_17402,N_17322);
nand U17540 (N_17540,N_17245,N_17205);
xnor U17541 (N_17541,N_17334,N_17115);
and U17542 (N_17542,N_17226,N_17431);
nand U17543 (N_17543,N_17218,N_17336);
nand U17544 (N_17544,N_17338,N_17440);
nor U17545 (N_17545,N_17219,N_17022);
and U17546 (N_17546,N_17166,N_17328);
nor U17547 (N_17547,N_17078,N_17211);
nor U17548 (N_17548,N_17351,N_17189);
nor U17549 (N_17549,N_17429,N_17080);
nor U17550 (N_17550,N_17362,N_17291);
nand U17551 (N_17551,N_17120,N_17344);
and U17552 (N_17552,N_17054,N_17042);
nand U17553 (N_17553,N_17481,N_17221);
and U17554 (N_17554,N_17405,N_17318);
or U17555 (N_17555,N_17454,N_17064);
nand U17556 (N_17556,N_17070,N_17187);
and U17557 (N_17557,N_17013,N_17461);
or U17558 (N_17558,N_17485,N_17395);
xor U17559 (N_17559,N_17051,N_17382);
nor U17560 (N_17560,N_17305,N_17296);
nand U17561 (N_17561,N_17260,N_17242);
and U17562 (N_17562,N_17114,N_17340);
nor U17563 (N_17563,N_17287,N_17032);
xor U17564 (N_17564,N_17292,N_17048);
xnor U17565 (N_17565,N_17310,N_17379);
nor U17566 (N_17566,N_17220,N_17225);
nor U17567 (N_17567,N_17084,N_17317);
and U17568 (N_17568,N_17154,N_17261);
xor U17569 (N_17569,N_17007,N_17158);
and U17570 (N_17570,N_17424,N_17493);
xor U17571 (N_17571,N_17029,N_17358);
and U17572 (N_17572,N_17031,N_17190);
xor U17573 (N_17573,N_17184,N_17162);
nor U17574 (N_17574,N_17345,N_17451);
and U17575 (N_17575,N_17088,N_17389);
nor U17576 (N_17576,N_17183,N_17157);
and U17577 (N_17577,N_17422,N_17464);
or U17578 (N_17578,N_17376,N_17450);
nand U17579 (N_17579,N_17034,N_17255);
xnor U17580 (N_17580,N_17369,N_17217);
and U17581 (N_17581,N_17240,N_17323);
nand U17582 (N_17582,N_17398,N_17373);
and U17583 (N_17583,N_17339,N_17280);
and U17584 (N_17584,N_17106,N_17215);
xor U17585 (N_17585,N_17437,N_17314);
or U17586 (N_17586,N_17281,N_17046);
nor U17587 (N_17587,N_17037,N_17447);
nand U17588 (N_17588,N_17155,N_17130);
and U17589 (N_17589,N_17385,N_17014);
xor U17590 (N_17590,N_17026,N_17000);
nand U17591 (N_17591,N_17194,N_17480);
nor U17592 (N_17592,N_17116,N_17343);
nand U17593 (N_17593,N_17179,N_17435);
and U17594 (N_17594,N_17019,N_17308);
nor U17595 (N_17595,N_17085,N_17065);
nand U17596 (N_17596,N_17145,N_17474);
or U17597 (N_17597,N_17324,N_17494);
or U17598 (N_17598,N_17439,N_17359);
nor U17599 (N_17599,N_17035,N_17403);
xor U17600 (N_17600,N_17258,N_17018);
nand U17601 (N_17601,N_17274,N_17231);
nand U17602 (N_17602,N_17364,N_17138);
or U17603 (N_17603,N_17406,N_17086);
and U17604 (N_17604,N_17272,N_17456);
or U17605 (N_17605,N_17087,N_17298);
nand U17606 (N_17606,N_17443,N_17361);
or U17607 (N_17607,N_17477,N_17167);
and U17608 (N_17608,N_17191,N_17315);
and U17609 (N_17609,N_17235,N_17243);
or U17610 (N_17610,N_17269,N_17069);
nand U17611 (N_17611,N_17449,N_17387);
xor U17612 (N_17612,N_17353,N_17326);
nor U17613 (N_17613,N_17473,N_17377);
nand U17614 (N_17614,N_17289,N_17043);
or U17615 (N_17615,N_17036,N_17445);
nand U17616 (N_17616,N_17113,N_17128);
or U17617 (N_17617,N_17201,N_17025);
and U17618 (N_17618,N_17047,N_17136);
nand U17619 (N_17619,N_17108,N_17408);
xor U17620 (N_17620,N_17333,N_17251);
xnor U17621 (N_17621,N_17416,N_17023);
nand U17622 (N_17622,N_17309,N_17392);
or U17623 (N_17623,N_17476,N_17144);
and U17624 (N_17624,N_17030,N_17412);
or U17625 (N_17625,N_17495,N_17250);
nand U17626 (N_17626,N_17012,N_17161);
nand U17627 (N_17627,N_17060,N_17380);
nor U17628 (N_17628,N_17181,N_17105);
nand U17629 (N_17629,N_17368,N_17095);
or U17630 (N_17630,N_17172,N_17366);
xnor U17631 (N_17631,N_17302,N_17349);
xnor U17632 (N_17632,N_17174,N_17468);
and U17633 (N_17633,N_17170,N_17109);
nand U17634 (N_17634,N_17149,N_17283);
nor U17635 (N_17635,N_17180,N_17058);
or U17636 (N_17636,N_17410,N_17301);
nand U17637 (N_17637,N_17150,N_17295);
and U17638 (N_17638,N_17396,N_17210);
nor U17639 (N_17639,N_17207,N_17414);
xor U17640 (N_17640,N_17173,N_17271);
nand U17641 (N_17641,N_17313,N_17241);
nor U17642 (N_17642,N_17348,N_17492);
nand U17643 (N_17643,N_17459,N_17471);
nor U17644 (N_17644,N_17090,N_17121);
nand U17645 (N_17645,N_17275,N_17137);
or U17646 (N_17646,N_17466,N_17399);
xor U17647 (N_17647,N_17270,N_17354);
and U17648 (N_17648,N_17488,N_17011);
xnor U17649 (N_17649,N_17125,N_17244);
xnor U17650 (N_17650,N_17001,N_17247);
or U17651 (N_17651,N_17214,N_17222);
or U17652 (N_17652,N_17268,N_17409);
nand U17653 (N_17653,N_17304,N_17118);
nand U17654 (N_17654,N_17028,N_17383);
or U17655 (N_17655,N_17252,N_17371);
xor U17656 (N_17656,N_17446,N_17352);
or U17657 (N_17657,N_17276,N_17393);
nand U17658 (N_17658,N_17327,N_17050);
or U17659 (N_17659,N_17165,N_17024);
or U17660 (N_17660,N_17487,N_17127);
or U17661 (N_17661,N_17259,N_17401);
nand U17662 (N_17662,N_17132,N_17067);
nand U17663 (N_17663,N_17146,N_17151);
or U17664 (N_17664,N_17212,N_17273);
xnor U17665 (N_17665,N_17335,N_17282);
or U17666 (N_17666,N_17257,N_17178);
and U17667 (N_17667,N_17465,N_17311);
and U17668 (N_17668,N_17248,N_17341);
xnor U17669 (N_17669,N_17143,N_17498);
xor U17670 (N_17670,N_17027,N_17469);
nand U17671 (N_17671,N_17482,N_17297);
and U17672 (N_17672,N_17062,N_17319);
xnor U17673 (N_17673,N_17216,N_17472);
nand U17674 (N_17674,N_17418,N_17156);
xnor U17675 (N_17675,N_17213,N_17192);
xnor U17676 (N_17676,N_17285,N_17433);
nand U17677 (N_17677,N_17420,N_17041);
and U17678 (N_17678,N_17288,N_17101);
xnor U17679 (N_17679,N_17236,N_17074);
xor U17680 (N_17680,N_17129,N_17263);
nor U17681 (N_17681,N_17091,N_17186);
or U17682 (N_17682,N_17195,N_17453);
nand U17683 (N_17683,N_17434,N_17490);
nand U17684 (N_17684,N_17478,N_17008);
xor U17685 (N_17685,N_17484,N_17400);
nand U17686 (N_17686,N_17425,N_17081);
xnor U17687 (N_17687,N_17278,N_17082);
nor U17688 (N_17688,N_17467,N_17234);
xor U17689 (N_17689,N_17499,N_17164);
nor U17690 (N_17690,N_17098,N_17111);
xor U17691 (N_17691,N_17483,N_17045);
and U17692 (N_17692,N_17112,N_17253);
xnor U17693 (N_17693,N_17141,N_17246);
nor U17694 (N_17694,N_17413,N_17388);
and U17695 (N_17695,N_17142,N_17038);
nand U17696 (N_17696,N_17040,N_17332);
xor U17697 (N_17697,N_17159,N_17330);
or U17698 (N_17698,N_17202,N_17321);
nor U17699 (N_17699,N_17004,N_17124);
and U17700 (N_17700,N_17153,N_17139);
nand U17701 (N_17701,N_17126,N_17438);
and U17702 (N_17702,N_17059,N_17404);
or U17703 (N_17703,N_17033,N_17426);
xnor U17704 (N_17704,N_17185,N_17475);
xor U17705 (N_17705,N_17177,N_17249);
and U17706 (N_17706,N_17209,N_17346);
nand U17707 (N_17707,N_17448,N_17415);
and U17708 (N_17708,N_17075,N_17147);
nand U17709 (N_17709,N_17053,N_17097);
nand U17710 (N_17710,N_17452,N_17163);
nor U17711 (N_17711,N_17381,N_17175);
nand U17712 (N_17712,N_17394,N_17407);
and U17713 (N_17713,N_17140,N_17021);
and U17714 (N_17714,N_17360,N_17279);
or U17715 (N_17715,N_17457,N_17491);
or U17716 (N_17716,N_17390,N_17299);
nand U17717 (N_17717,N_17307,N_17427);
xnor U17718 (N_17718,N_17350,N_17286);
nand U17719 (N_17719,N_17355,N_17227);
or U17720 (N_17720,N_17017,N_17055);
nand U17721 (N_17721,N_17133,N_17009);
xor U17722 (N_17722,N_17171,N_17169);
nor U17723 (N_17723,N_17372,N_17363);
xnor U17724 (N_17724,N_17066,N_17228);
nand U17725 (N_17725,N_17397,N_17100);
or U17726 (N_17726,N_17444,N_17262);
xnor U17727 (N_17727,N_17096,N_17391);
nor U17728 (N_17728,N_17119,N_17428);
nand U17729 (N_17729,N_17421,N_17479);
nor U17730 (N_17730,N_17103,N_17193);
xnor U17731 (N_17731,N_17232,N_17005);
or U17732 (N_17732,N_17375,N_17356);
xor U17733 (N_17733,N_17168,N_17266);
or U17734 (N_17734,N_17230,N_17337);
and U17735 (N_17735,N_17131,N_17347);
xor U17736 (N_17736,N_17152,N_17423);
or U17737 (N_17737,N_17176,N_17342);
nand U17738 (N_17738,N_17134,N_17357);
nand U17739 (N_17739,N_17463,N_17374);
nand U17740 (N_17740,N_17436,N_17015);
nor U17741 (N_17741,N_17063,N_17135);
or U17742 (N_17742,N_17006,N_17148);
and U17743 (N_17743,N_17320,N_17329);
nor U17744 (N_17744,N_17199,N_17277);
or U17745 (N_17745,N_17441,N_17039);
nor U17746 (N_17746,N_17432,N_17256);
and U17747 (N_17747,N_17068,N_17020);
nor U17748 (N_17748,N_17489,N_17455);
and U17749 (N_17749,N_17107,N_17044);
nand U17750 (N_17750,N_17204,N_17248);
nand U17751 (N_17751,N_17064,N_17106);
xnor U17752 (N_17752,N_17227,N_17186);
xor U17753 (N_17753,N_17027,N_17006);
and U17754 (N_17754,N_17435,N_17053);
and U17755 (N_17755,N_17295,N_17380);
or U17756 (N_17756,N_17151,N_17271);
xor U17757 (N_17757,N_17173,N_17324);
nand U17758 (N_17758,N_17498,N_17199);
or U17759 (N_17759,N_17319,N_17441);
xnor U17760 (N_17760,N_17482,N_17099);
nor U17761 (N_17761,N_17339,N_17244);
nor U17762 (N_17762,N_17450,N_17341);
nand U17763 (N_17763,N_17411,N_17311);
nor U17764 (N_17764,N_17048,N_17030);
nor U17765 (N_17765,N_17360,N_17465);
xor U17766 (N_17766,N_17239,N_17231);
and U17767 (N_17767,N_17075,N_17401);
xor U17768 (N_17768,N_17211,N_17103);
or U17769 (N_17769,N_17143,N_17295);
and U17770 (N_17770,N_17349,N_17471);
nor U17771 (N_17771,N_17168,N_17075);
nand U17772 (N_17772,N_17427,N_17100);
and U17773 (N_17773,N_17058,N_17279);
and U17774 (N_17774,N_17070,N_17277);
and U17775 (N_17775,N_17447,N_17164);
xor U17776 (N_17776,N_17463,N_17355);
and U17777 (N_17777,N_17380,N_17119);
nor U17778 (N_17778,N_17084,N_17276);
or U17779 (N_17779,N_17124,N_17342);
xor U17780 (N_17780,N_17086,N_17208);
nand U17781 (N_17781,N_17015,N_17058);
nor U17782 (N_17782,N_17212,N_17230);
nand U17783 (N_17783,N_17322,N_17319);
nand U17784 (N_17784,N_17117,N_17254);
nor U17785 (N_17785,N_17097,N_17041);
nor U17786 (N_17786,N_17381,N_17196);
xor U17787 (N_17787,N_17404,N_17018);
and U17788 (N_17788,N_17194,N_17311);
xor U17789 (N_17789,N_17194,N_17326);
and U17790 (N_17790,N_17281,N_17490);
and U17791 (N_17791,N_17304,N_17171);
nor U17792 (N_17792,N_17402,N_17092);
nand U17793 (N_17793,N_17004,N_17266);
nor U17794 (N_17794,N_17145,N_17156);
or U17795 (N_17795,N_17226,N_17182);
or U17796 (N_17796,N_17313,N_17460);
and U17797 (N_17797,N_17165,N_17145);
xnor U17798 (N_17798,N_17396,N_17125);
or U17799 (N_17799,N_17075,N_17173);
nor U17800 (N_17800,N_17471,N_17321);
or U17801 (N_17801,N_17469,N_17254);
and U17802 (N_17802,N_17187,N_17092);
or U17803 (N_17803,N_17347,N_17484);
nor U17804 (N_17804,N_17134,N_17019);
and U17805 (N_17805,N_17383,N_17274);
nand U17806 (N_17806,N_17488,N_17063);
nand U17807 (N_17807,N_17034,N_17195);
and U17808 (N_17808,N_17424,N_17082);
nor U17809 (N_17809,N_17494,N_17131);
and U17810 (N_17810,N_17485,N_17496);
nand U17811 (N_17811,N_17080,N_17172);
xor U17812 (N_17812,N_17374,N_17399);
nand U17813 (N_17813,N_17227,N_17279);
nor U17814 (N_17814,N_17429,N_17181);
nand U17815 (N_17815,N_17083,N_17236);
xor U17816 (N_17816,N_17411,N_17078);
xor U17817 (N_17817,N_17454,N_17422);
xnor U17818 (N_17818,N_17305,N_17048);
and U17819 (N_17819,N_17492,N_17159);
nor U17820 (N_17820,N_17196,N_17342);
xnor U17821 (N_17821,N_17332,N_17494);
nor U17822 (N_17822,N_17084,N_17370);
nand U17823 (N_17823,N_17274,N_17013);
or U17824 (N_17824,N_17002,N_17411);
and U17825 (N_17825,N_17425,N_17274);
nor U17826 (N_17826,N_17427,N_17120);
nand U17827 (N_17827,N_17361,N_17327);
and U17828 (N_17828,N_17489,N_17272);
nor U17829 (N_17829,N_17340,N_17443);
and U17830 (N_17830,N_17466,N_17241);
and U17831 (N_17831,N_17103,N_17375);
xor U17832 (N_17832,N_17161,N_17221);
or U17833 (N_17833,N_17115,N_17134);
nand U17834 (N_17834,N_17305,N_17198);
or U17835 (N_17835,N_17263,N_17469);
and U17836 (N_17836,N_17145,N_17316);
and U17837 (N_17837,N_17272,N_17468);
nand U17838 (N_17838,N_17482,N_17314);
nand U17839 (N_17839,N_17263,N_17390);
xnor U17840 (N_17840,N_17084,N_17442);
nand U17841 (N_17841,N_17340,N_17086);
nand U17842 (N_17842,N_17467,N_17424);
and U17843 (N_17843,N_17411,N_17001);
or U17844 (N_17844,N_17100,N_17273);
or U17845 (N_17845,N_17298,N_17449);
and U17846 (N_17846,N_17376,N_17059);
xnor U17847 (N_17847,N_17461,N_17480);
or U17848 (N_17848,N_17358,N_17339);
nor U17849 (N_17849,N_17418,N_17076);
nor U17850 (N_17850,N_17198,N_17480);
xnor U17851 (N_17851,N_17438,N_17012);
nor U17852 (N_17852,N_17486,N_17104);
and U17853 (N_17853,N_17197,N_17348);
xnor U17854 (N_17854,N_17199,N_17324);
or U17855 (N_17855,N_17140,N_17390);
xor U17856 (N_17856,N_17150,N_17305);
nor U17857 (N_17857,N_17006,N_17290);
xor U17858 (N_17858,N_17050,N_17174);
nand U17859 (N_17859,N_17067,N_17148);
or U17860 (N_17860,N_17058,N_17027);
and U17861 (N_17861,N_17445,N_17355);
and U17862 (N_17862,N_17273,N_17063);
nor U17863 (N_17863,N_17153,N_17058);
nor U17864 (N_17864,N_17420,N_17059);
and U17865 (N_17865,N_17315,N_17186);
or U17866 (N_17866,N_17144,N_17214);
and U17867 (N_17867,N_17016,N_17306);
nor U17868 (N_17868,N_17298,N_17075);
or U17869 (N_17869,N_17041,N_17287);
and U17870 (N_17870,N_17143,N_17228);
xor U17871 (N_17871,N_17025,N_17387);
xnor U17872 (N_17872,N_17184,N_17384);
xor U17873 (N_17873,N_17111,N_17196);
xnor U17874 (N_17874,N_17008,N_17280);
or U17875 (N_17875,N_17006,N_17024);
or U17876 (N_17876,N_17031,N_17084);
or U17877 (N_17877,N_17201,N_17067);
or U17878 (N_17878,N_17262,N_17047);
or U17879 (N_17879,N_17188,N_17498);
xor U17880 (N_17880,N_17203,N_17310);
or U17881 (N_17881,N_17498,N_17479);
nand U17882 (N_17882,N_17359,N_17411);
or U17883 (N_17883,N_17445,N_17314);
nor U17884 (N_17884,N_17346,N_17369);
and U17885 (N_17885,N_17403,N_17073);
and U17886 (N_17886,N_17355,N_17453);
nand U17887 (N_17887,N_17271,N_17177);
and U17888 (N_17888,N_17171,N_17118);
xor U17889 (N_17889,N_17171,N_17355);
nor U17890 (N_17890,N_17197,N_17109);
xnor U17891 (N_17891,N_17203,N_17369);
nor U17892 (N_17892,N_17027,N_17335);
xor U17893 (N_17893,N_17467,N_17263);
nand U17894 (N_17894,N_17155,N_17314);
xor U17895 (N_17895,N_17433,N_17073);
nand U17896 (N_17896,N_17222,N_17051);
and U17897 (N_17897,N_17088,N_17461);
nor U17898 (N_17898,N_17260,N_17142);
nor U17899 (N_17899,N_17086,N_17381);
or U17900 (N_17900,N_17426,N_17322);
and U17901 (N_17901,N_17089,N_17246);
nand U17902 (N_17902,N_17088,N_17350);
nand U17903 (N_17903,N_17359,N_17026);
or U17904 (N_17904,N_17461,N_17355);
xnor U17905 (N_17905,N_17107,N_17148);
and U17906 (N_17906,N_17067,N_17159);
and U17907 (N_17907,N_17029,N_17122);
and U17908 (N_17908,N_17381,N_17014);
and U17909 (N_17909,N_17134,N_17327);
or U17910 (N_17910,N_17305,N_17267);
and U17911 (N_17911,N_17011,N_17081);
nand U17912 (N_17912,N_17493,N_17274);
nand U17913 (N_17913,N_17425,N_17481);
and U17914 (N_17914,N_17083,N_17352);
nor U17915 (N_17915,N_17036,N_17131);
nor U17916 (N_17916,N_17242,N_17228);
or U17917 (N_17917,N_17259,N_17465);
xor U17918 (N_17918,N_17062,N_17031);
and U17919 (N_17919,N_17409,N_17100);
and U17920 (N_17920,N_17127,N_17201);
nor U17921 (N_17921,N_17095,N_17089);
xnor U17922 (N_17922,N_17021,N_17404);
and U17923 (N_17923,N_17006,N_17476);
or U17924 (N_17924,N_17027,N_17255);
and U17925 (N_17925,N_17339,N_17102);
xnor U17926 (N_17926,N_17178,N_17101);
xnor U17927 (N_17927,N_17476,N_17032);
nor U17928 (N_17928,N_17297,N_17423);
or U17929 (N_17929,N_17490,N_17087);
nor U17930 (N_17930,N_17245,N_17350);
or U17931 (N_17931,N_17125,N_17385);
nand U17932 (N_17932,N_17303,N_17089);
xnor U17933 (N_17933,N_17096,N_17306);
or U17934 (N_17934,N_17256,N_17499);
nor U17935 (N_17935,N_17329,N_17131);
and U17936 (N_17936,N_17000,N_17044);
xnor U17937 (N_17937,N_17240,N_17038);
and U17938 (N_17938,N_17318,N_17252);
xnor U17939 (N_17939,N_17275,N_17296);
nand U17940 (N_17940,N_17493,N_17211);
xor U17941 (N_17941,N_17206,N_17432);
or U17942 (N_17942,N_17110,N_17270);
xor U17943 (N_17943,N_17404,N_17237);
and U17944 (N_17944,N_17163,N_17210);
nand U17945 (N_17945,N_17399,N_17451);
or U17946 (N_17946,N_17428,N_17115);
and U17947 (N_17947,N_17081,N_17427);
and U17948 (N_17948,N_17206,N_17078);
or U17949 (N_17949,N_17496,N_17098);
and U17950 (N_17950,N_17301,N_17201);
and U17951 (N_17951,N_17079,N_17326);
nand U17952 (N_17952,N_17456,N_17031);
or U17953 (N_17953,N_17107,N_17362);
xnor U17954 (N_17954,N_17213,N_17087);
and U17955 (N_17955,N_17459,N_17261);
and U17956 (N_17956,N_17144,N_17194);
nand U17957 (N_17957,N_17347,N_17262);
xnor U17958 (N_17958,N_17412,N_17236);
xnor U17959 (N_17959,N_17013,N_17462);
and U17960 (N_17960,N_17232,N_17330);
nor U17961 (N_17961,N_17246,N_17043);
nand U17962 (N_17962,N_17006,N_17259);
nor U17963 (N_17963,N_17270,N_17499);
xnor U17964 (N_17964,N_17032,N_17236);
or U17965 (N_17965,N_17123,N_17271);
nand U17966 (N_17966,N_17150,N_17440);
xnor U17967 (N_17967,N_17062,N_17388);
xor U17968 (N_17968,N_17116,N_17191);
nand U17969 (N_17969,N_17431,N_17206);
xnor U17970 (N_17970,N_17096,N_17195);
xor U17971 (N_17971,N_17026,N_17062);
nand U17972 (N_17972,N_17002,N_17402);
and U17973 (N_17973,N_17155,N_17019);
nand U17974 (N_17974,N_17222,N_17463);
nand U17975 (N_17975,N_17078,N_17091);
nor U17976 (N_17976,N_17454,N_17089);
nor U17977 (N_17977,N_17037,N_17462);
nand U17978 (N_17978,N_17218,N_17223);
xor U17979 (N_17979,N_17185,N_17219);
and U17980 (N_17980,N_17116,N_17411);
nand U17981 (N_17981,N_17197,N_17340);
xnor U17982 (N_17982,N_17282,N_17289);
and U17983 (N_17983,N_17458,N_17001);
xnor U17984 (N_17984,N_17428,N_17363);
or U17985 (N_17985,N_17438,N_17401);
or U17986 (N_17986,N_17399,N_17059);
nor U17987 (N_17987,N_17442,N_17369);
nor U17988 (N_17988,N_17436,N_17090);
nor U17989 (N_17989,N_17036,N_17042);
xnor U17990 (N_17990,N_17256,N_17442);
nor U17991 (N_17991,N_17287,N_17232);
nand U17992 (N_17992,N_17325,N_17432);
nand U17993 (N_17993,N_17336,N_17372);
or U17994 (N_17994,N_17331,N_17004);
xnor U17995 (N_17995,N_17351,N_17075);
or U17996 (N_17996,N_17123,N_17272);
xor U17997 (N_17997,N_17240,N_17445);
xnor U17998 (N_17998,N_17158,N_17246);
or U17999 (N_17999,N_17441,N_17432);
or U18000 (N_18000,N_17584,N_17821);
xnor U18001 (N_18001,N_17915,N_17740);
or U18002 (N_18002,N_17678,N_17531);
nor U18003 (N_18003,N_17566,N_17646);
nor U18004 (N_18004,N_17642,N_17693);
xor U18005 (N_18005,N_17792,N_17551);
or U18006 (N_18006,N_17541,N_17501);
and U18007 (N_18007,N_17809,N_17935);
nand U18008 (N_18008,N_17718,N_17976);
and U18009 (N_18009,N_17909,N_17567);
or U18010 (N_18010,N_17638,N_17800);
nor U18011 (N_18011,N_17712,N_17635);
or U18012 (N_18012,N_17947,N_17794);
and U18013 (N_18013,N_17630,N_17980);
nor U18014 (N_18014,N_17985,N_17589);
xor U18015 (N_18015,N_17723,N_17746);
or U18016 (N_18016,N_17580,N_17953);
nand U18017 (N_18017,N_17708,N_17899);
nor U18018 (N_18018,N_17941,N_17609);
nand U18019 (N_18019,N_17908,N_17592);
nor U18020 (N_18020,N_17905,N_17857);
and U18021 (N_18021,N_17859,N_17563);
nor U18022 (N_18022,N_17679,N_17841);
and U18023 (N_18023,N_17731,N_17513);
nor U18024 (N_18024,N_17863,N_17872);
and U18025 (N_18025,N_17690,N_17578);
and U18026 (N_18026,N_17697,N_17839);
and U18027 (N_18027,N_17738,N_17576);
and U18028 (N_18028,N_17787,N_17572);
or U18029 (N_18029,N_17665,N_17916);
nor U18030 (N_18030,N_17827,N_17819);
nand U18031 (N_18031,N_17922,N_17610);
nor U18032 (N_18032,N_17571,N_17733);
xor U18033 (N_18033,N_17755,N_17856);
nand U18034 (N_18034,N_17993,N_17885);
nor U18035 (N_18035,N_17730,N_17932);
nand U18036 (N_18036,N_17979,N_17546);
nand U18037 (N_18037,N_17761,N_17648);
nand U18038 (N_18038,N_17754,N_17945);
nand U18039 (N_18039,N_17777,N_17954);
nor U18040 (N_18040,N_17978,N_17785);
nor U18041 (N_18041,N_17688,N_17711);
xor U18042 (N_18042,N_17503,N_17561);
or U18043 (N_18043,N_17948,N_17673);
or U18044 (N_18044,N_17997,N_17533);
nor U18045 (N_18045,N_17637,N_17525);
xor U18046 (N_18046,N_17903,N_17694);
nor U18047 (N_18047,N_17601,N_17766);
xor U18048 (N_18048,N_17747,N_17611);
xnor U18049 (N_18049,N_17682,N_17986);
and U18050 (N_18050,N_17790,N_17606);
xor U18051 (N_18051,N_17502,N_17547);
nand U18052 (N_18052,N_17880,N_17901);
and U18053 (N_18053,N_17581,N_17799);
nor U18054 (N_18054,N_17701,N_17649);
nor U18055 (N_18055,N_17864,N_17894);
and U18056 (N_18056,N_17600,N_17770);
or U18057 (N_18057,N_17728,N_17861);
nand U18058 (N_18058,N_17680,N_17812);
nor U18059 (N_18059,N_17805,N_17781);
nor U18060 (N_18060,N_17512,N_17904);
nand U18061 (N_18061,N_17780,N_17644);
nor U18062 (N_18062,N_17760,N_17921);
xor U18063 (N_18063,N_17564,N_17815);
and U18064 (N_18064,N_17764,N_17726);
nand U18065 (N_18065,N_17869,N_17789);
nand U18066 (N_18066,N_17706,N_17984);
xor U18067 (N_18067,N_17801,N_17772);
and U18068 (N_18068,N_17749,N_17778);
and U18069 (N_18069,N_17962,N_17539);
nor U18070 (N_18070,N_17897,N_17931);
xnor U18071 (N_18071,N_17937,N_17517);
and U18072 (N_18072,N_17753,N_17602);
and U18073 (N_18073,N_17959,N_17739);
and U18074 (N_18074,N_17737,N_17720);
and U18075 (N_18075,N_17520,N_17519);
and U18076 (N_18076,N_17586,N_17994);
or U18077 (N_18077,N_17656,N_17703);
nand U18078 (N_18078,N_17875,N_17615);
and U18079 (N_18079,N_17585,N_17717);
xor U18080 (N_18080,N_17988,N_17906);
xnor U18081 (N_18081,N_17583,N_17775);
nand U18082 (N_18082,N_17573,N_17873);
and U18083 (N_18083,N_17970,N_17716);
and U18084 (N_18084,N_17672,N_17537);
nand U18085 (N_18085,N_17536,N_17882);
xnor U18086 (N_18086,N_17612,N_17829);
nand U18087 (N_18087,N_17868,N_17808);
nand U18088 (N_18088,N_17913,N_17735);
or U18089 (N_18089,N_17555,N_17732);
xor U18090 (N_18090,N_17964,N_17917);
xnor U18091 (N_18091,N_17556,N_17876);
nor U18092 (N_18092,N_17846,N_17991);
xnor U18093 (N_18093,N_17524,N_17834);
and U18094 (N_18094,N_17620,N_17751);
nor U18095 (N_18095,N_17927,N_17558);
xnor U18096 (N_18096,N_17643,N_17527);
xor U18097 (N_18097,N_17830,N_17532);
xor U18098 (N_18098,N_17858,N_17614);
nand U18099 (N_18099,N_17709,N_17568);
and U18100 (N_18100,N_17878,N_17824);
and U18101 (N_18101,N_17847,N_17587);
and U18102 (N_18102,N_17996,N_17695);
or U18103 (N_18103,N_17641,N_17943);
or U18104 (N_18104,N_17798,N_17992);
xor U18105 (N_18105,N_17837,N_17776);
xnor U18106 (N_18106,N_17514,N_17553);
or U18107 (N_18107,N_17627,N_17759);
xnor U18108 (N_18108,N_17895,N_17851);
or U18109 (N_18109,N_17636,N_17548);
nor U18110 (N_18110,N_17534,N_17683);
xor U18111 (N_18111,N_17845,N_17686);
xor U18112 (N_18112,N_17590,N_17862);
nand U18113 (N_18113,N_17719,N_17955);
or U18114 (N_18114,N_17657,N_17811);
nor U18115 (N_18115,N_17804,N_17818);
and U18116 (N_18116,N_17890,N_17763);
and U18117 (N_18117,N_17950,N_17866);
xnor U18118 (N_18118,N_17783,N_17704);
and U18119 (N_18119,N_17743,N_17826);
or U18120 (N_18120,N_17757,N_17727);
nand U18121 (N_18121,N_17762,N_17545);
nor U18122 (N_18122,N_17983,N_17628);
xnor U18123 (N_18123,N_17971,N_17653);
and U18124 (N_18124,N_17510,N_17516);
nor U18125 (N_18125,N_17651,N_17791);
or U18126 (N_18126,N_17544,N_17562);
xor U18127 (N_18127,N_17575,N_17752);
nand U18128 (N_18128,N_17807,N_17956);
nand U18129 (N_18129,N_17919,N_17676);
xnor U18130 (N_18130,N_17634,N_17797);
and U18131 (N_18131,N_17893,N_17960);
or U18132 (N_18132,N_17666,N_17670);
xor U18133 (N_18133,N_17820,N_17618);
and U18134 (N_18134,N_17987,N_17542);
nor U18135 (N_18135,N_17814,N_17940);
xnor U18136 (N_18136,N_17639,N_17700);
nand U18137 (N_18137,N_17570,N_17967);
nand U18138 (N_18138,N_17707,N_17603);
nor U18139 (N_18139,N_17881,N_17828);
and U18140 (N_18140,N_17745,N_17902);
nor U18141 (N_18141,N_17806,N_17961);
xor U18142 (N_18142,N_17848,N_17944);
xnor U18143 (N_18143,N_17816,N_17802);
or U18144 (N_18144,N_17810,N_17850);
and U18145 (N_18145,N_17741,N_17951);
nor U18146 (N_18146,N_17929,N_17599);
and U18147 (N_18147,N_17604,N_17684);
xor U18148 (N_18148,N_17977,N_17822);
nand U18149 (N_18149,N_17692,N_17938);
and U18150 (N_18150,N_17557,N_17958);
xor U18151 (N_18151,N_17623,N_17912);
and U18152 (N_18152,N_17849,N_17650);
xnor U18153 (N_18153,N_17926,N_17825);
nor U18154 (N_18154,N_17963,N_17803);
xnor U18155 (N_18155,N_17663,N_17925);
or U18156 (N_18156,N_17874,N_17687);
nand U18157 (N_18157,N_17668,N_17647);
nor U18158 (N_18158,N_17854,N_17594);
nor U18159 (N_18159,N_17619,N_17523);
nor U18160 (N_18160,N_17898,N_17867);
xnor U18161 (N_18161,N_17538,N_17833);
nand U18162 (N_18162,N_17793,N_17625);
nand U18163 (N_18163,N_17871,N_17598);
nor U18164 (N_18164,N_17914,N_17549);
nand U18165 (N_18165,N_17933,N_17840);
nand U18166 (N_18166,N_17522,N_17559);
xnor U18167 (N_18167,N_17710,N_17595);
xor U18168 (N_18168,N_17744,N_17729);
nor U18169 (N_18169,N_17907,N_17702);
or U18170 (N_18170,N_17528,N_17569);
xor U18171 (N_18171,N_17633,N_17645);
and U18172 (N_18172,N_17530,N_17565);
nand U18173 (N_18173,N_17714,N_17588);
nand U18174 (N_18174,N_17835,N_17554);
nor U18175 (N_18175,N_17928,N_17577);
nor U18176 (N_18176,N_17966,N_17934);
and U18177 (N_18177,N_17973,N_17795);
nor U18178 (N_18178,N_17608,N_17574);
or U18179 (N_18179,N_17505,N_17844);
and U18180 (N_18180,N_17838,N_17667);
or U18181 (N_18181,N_17836,N_17796);
and U18182 (N_18182,N_17734,N_17842);
nand U18183 (N_18183,N_17560,N_17788);
xnor U18184 (N_18184,N_17918,N_17952);
xor U18185 (N_18185,N_17617,N_17957);
nand U18186 (N_18186,N_17689,N_17853);
or U18187 (N_18187,N_17831,N_17660);
nand U18188 (N_18188,N_17661,N_17884);
nand U18189 (N_18189,N_17591,N_17865);
nand U18190 (N_18190,N_17896,N_17936);
nor U18191 (N_18191,N_17974,N_17900);
or U18192 (N_18192,N_17924,N_17879);
or U18193 (N_18193,N_17771,N_17626);
nand U18194 (N_18194,N_17892,N_17658);
nand U18195 (N_18195,N_17705,N_17671);
xor U18196 (N_18196,N_17540,N_17677);
xor U18197 (N_18197,N_17886,N_17631);
or U18198 (N_18198,N_17972,N_17742);
or U18199 (N_18199,N_17998,N_17655);
nand U18200 (N_18200,N_17664,N_17995);
and U18201 (N_18201,N_17817,N_17508);
xnor U18202 (N_18202,N_17725,N_17765);
xnor U18203 (N_18203,N_17681,N_17507);
nor U18204 (N_18204,N_17999,N_17813);
and U18205 (N_18205,N_17981,N_17659);
nor U18206 (N_18206,N_17939,N_17942);
and U18207 (N_18207,N_17911,N_17515);
and U18208 (N_18208,N_17654,N_17552);
nor U18209 (N_18209,N_17969,N_17923);
nand U18210 (N_18210,N_17989,N_17843);
xnor U18211 (N_18211,N_17509,N_17975);
xor U18212 (N_18212,N_17621,N_17550);
nand U18213 (N_18213,N_17782,N_17773);
xnor U18214 (N_18214,N_17860,N_17582);
xor U18215 (N_18215,N_17887,N_17696);
xor U18216 (N_18216,N_17691,N_17500);
and U18217 (N_18217,N_17504,N_17715);
xnor U18218 (N_18218,N_17767,N_17669);
or U18219 (N_18219,N_17748,N_17889);
nand U18220 (N_18220,N_17698,N_17624);
nor U18221 (N_18221,N_17662,N_17852);
or U18222 (N_18222,N_17768,N_17632);
nor U18223 (N_18223,N_17910,N_17769);
xor U18224 (N_18224,N_17675,N_17736);
or U18225 (N_18225,N_17883,N_17526);
xor U18226 (N_18226,N_17949,N_17786);
and U18227 (N_18227,N_17756,N_17506);
xor U18228 (N_18228,N_17888,N_17629);
nor U18229 (N_18229,N_17832,N_17870);
xor U18230 (N_18230,N_17990,N_17779);
nand U18231 (N_18231,N_17982,N_17674);
or U18232 (N_18232,N_17784,N_17652);
nor U18233 (N_18233,N_17518,N_17685);
xor U18234 (N_18234,N_17521,N_17607);
nand U18235 (N_18235,N_17721,N_17597);
nand U18236 (N_18236,N_17640,N_17758);
nand U18237 (N_18237,N_17946,N_17920);
nor U18238 (N_18238,N_17877,N_17891);
or U18239 (N_18239,N_17593,N_17579);
nor U18240 (N_18240,N_17713,N_17774);
and U18241 (N_18241,N_17596,N_17529);
nand U18242 (N_18242,N_17965,N_17968);
nand U18243 (N_18243,N_17722,N_17930);
or U18244 (N_18244,N_17543,N_17535);
nand U18245 (N_18245,N_17724,N_17613);
nand U18246 (N_18246,N_17823,N_17605);
xor U18247 (N_18247,N_17750,N_17616);
xor U18248 (N_18248,N_17511,N_17699);
xnor U18249 (N_18249,N_17622,N_17855);
or U18250 (N_18250,N_17891,N_17823);
nand U18251 (N_18251,N_17519,N_17547);
and U18252 (N_18252,N_17547,N_17812);
and U18253 (N_18253,N_17711,N_17873);
xnor U18254 (N_18254,N_17777,N_17699);
xnor U18255 (N_18255,N_17790,N_17692);
nand U18256 (N_18256,N_17865,N_17531);
nand U18257 (N_18257,N_17656,N_17945);
xnor U18258 (N_18258,N_17686,N_17776);
or U18259 (N_18259,N_17866,N_17796);
and U18260 (N_18260,N_17589,N_17635);
and U18261 (N_18261,N_17684,N_17898);
and U18262 (N_18262,N_17590,N_17893);
xnor U18263 (N_18263,N_17580,N_17633);
xnor U18264 (N_18264,N_17726,N_17576);
and U18265 (N_18265,N_17956,N_17589);
nand U18266 (N_18266,N_17816,N_17528);
nor U18267 (N_18267,N_17787,N_17995);
nor U18268 (N_18268,N_17946,N_17841);
or U18269 (N_18269,N_17601,N_17865);
or U18270 (N_18270,N_17878,N_17993);
nor U18271 (N_18271,N_17618,N_17958);
xnor U18272 (N_18272,N_17851,N_17898);
nand U18273 (N_18273,N_17951,N_17836);
xor U18274 (N_18274,N_17954,N_17510);
nand U18275 (N_18275,N_17897,N_17763);
xnor U18276 (N_18276,N_17523,N_17658);
xor U18277 (N_18277,N_17562,N_17676);
nor U18278 (N_18278,N_17819,N_17767);
xor U18279 (N_18279,N_17647,N_17783);
and U18280 (N_18280,N_17790,N_17971);
nand U18281 (N_18281,N_17790,N_17701);
nor U18282 (N_18282,N_17799,N_17670);
xor U18283 (N_18283,N_17522,N_17872);
nand U18284 (N_18284,N_17931,N_17775);
nor U18285 (N_18285,N_17815,N_17778);
nor U18286 (N_18286,N_17847,N_17666);
xor U18287 (N_18287,N_17907,N_17682);
or U18288 (N_18288,N_17939,N_17670);
xnor U18289 (N_18289,N_17949,N_17967);
nor U18290 (N_18290,N_17754,N_17692);
or U18291 (N_18291,N_17791,N_17749);
nand U18292 (N_18292,N_17752,N_17979);
or U18293 (N_18293,N_17693,N_17906);
nand U18294 (N_18294,N_17760,N_17898);
and U18295 (N_18295,N_17766,N_17742);
or U18296 (N_18296,N_17716,N_17918);
or U18297 (N_18297,N_17526,N_17855);
or U18298 (N_18298,N_17636,N_17951);
or U18299 (N_18299,N_17733,N_17800);
or U18300 (N_18300,N_17627,N_17862);
nor U18301 (N_18301,N_17622,N_17801);
and U18302 (N_18302,N_17973,N_17847);
and U18303 (N_18303,N_17950,N_17552);
and U18304 (N_18304,N_17559,N_17633);
nand U18305 (N_18305,N_17896,N_17672);
xnor U18306 (N_18306,N_17942,N_17595);
or U18307 (N_18307,N_17764,N_17530);
nor U18308 (N_18308,N_17952,N_17731);
and U18309 (N_18309,N_17866,N_17969);
nand U18310 (N_18310,N_17545,N_17903);
and U18311 (N_18311,N_17650,N_17804);
and U18312 (N_18312,N_17770,N_17505);
nand U18313 (N_18313,N_17844,N_17920);
nor U18314 (N_18314,N_17965,N_17978);
nand U18315 (N_18315,N_17716,N_17526);
or U18316 (N_18316,N_17831,N_17858);
or U18317 (N_18317,N_17515,N_17926);
nor U18318 (N_18318,N_17785,N_17853);
nand U18319 (N_18319,N_17874,N_17693);
or U18320 (N_18320,N_17612,N_17524);
nand U18321 (N_18321,N_17638,N_17823);
nand U18322 (N_18322,N_17707,N_17674);
xnor U18323 (N_18323,N_17821,N_17870);
nor U18324 (N_18324,N_17783,N_17616);
nor U18325 (N_18325,N_17950,N_17660);
nor U18326 (N_18326,N_17888,N_17563);
nand U18327 (N_18327,N_17635,N_17734);
or U18328 (N_18328,N_17920,N_17704);
nor U18329 (N_18329,N_17847,N_17501);
nand U18330 (N_18330,N_17702,N_17869);
nor U18331 (N_18331,N_17994,N_17732);
nand U18332 (N_18332,N_17510,N_17752);
or U18333 (N_18333,N_17580,N_17724);
and U18334 (N_18334,N_17875,N_17690);
nor U18335 (N_18335,N_17908,N_17925);
nand U18336 (N_18336,N_17642,N_17834);
nor U18337 (N_18337,N_17948,N_17836);
nand U18338 (N_18338,N_17607,N_17968);
nor U18339 (N_18339,N_17962,N_17824);
nand U18340 (N_18340,N_17944,N_17850);
and U18341 (N_18341,N_17881,N_17707);
xor U18342 (N_18342,N_17755,N_17788);
xor U18343 (N_18343,N_17581,N_17722);
and U18344 (N_18344,N_17596,N_17836);
and U18345 (N_18345,N_17835,N_17826);
or U18346 (N_18346,N_17521,N_17634);
nor U18347 (N_18347,N_17578,N_17995);
nand U18348 (N_18348,N_17566,N_17586);
xor U18349 (N_18349,N_17600,N_17759);
nor U18350 (N_18350,N_17670,N_17989);
nand U18351 (N_18351,N_17731,N_17887);
and U18352 (N_18352,N_17518,N_17574);
nor U18353 (N_18353,N_17918,N_17688);
nor U18354 (N_18354,N_17685,N_17883);
or U18355 (N_18355,N_17661,N_17718);
or U18356 (N_18356,N_17981,N_17801);
and U18357 (N_18357,N_17620,N_17955);
and U18358 (N_18358,N_17790,N_17728);
nor U18359 (N_18359,N_17803,N_17510);
and U18360 (N_18360,N_17920,N_17977);
nand U18361 (N_18361,N_17571,N_17979);
and U18362 (N_18362,N_17712,N_17586);
xor U18363 (N_18363,N_17740,N_17644);
and U18364 (N_18364,N_17519,N_17569);
nor U18365 (N_18365,N_17630,N_17531);
and U18366 (N_18366,N_17532,N_17779);
and U18367 (N_18367,N_17690,N_17819);
xor U18368 (N_18368,N_17755,N_17676);
nor U18369 (N_18369,N_17715,N_17916);
or U18370 (N_18370,N_17972,N_17868);
or U18371 (N_18371,N_17634,N_17658);
and U18372 (N_18372,N_17861,N_17929);
or U18373 (N_18373,N_17653,N_17770);
or U18374 (N_18374,N_17753,N_17655);
and U18375 (N_18375,N_17667,N_17666);
xnor U18376 (N_18376,N_17916,N_17864);
nor U18377 (N_18377,N_17898,N_17638);
nor U18378 (N_18378,N_17847,N_17880);
and U18379 (N_18379,N_17628,N_17552);
nor U18380 (N_18380,N_17800,N_17582);
nor U18381 (N_18381,N_17808,N_17919);
or U18382 (N_18382,N_17502,N_17749);
xnor U18383 (N_18383,N_17567,N_17826);
or U18384 (N_18384,N_17984,N_17971);
or U18385 (N_18385,N_17576,N_17581);
and U18386 (N_18386,N_17618,N_17737);
or U18387 (N_18387,N_17571,N_17877);
nand U18388 (N_18388,N_17859,N_17834);
or U18389 (N_18389,N_17579,N_17692);
xnor U18390 (N_18390,N_17865,N_17911);
xnor U18391 (N_18391,N_17927,N_17787);
or U18392 (N_18392,N_17558,N_17755);
or U18393 (N_18393,N_17678,N_17774);
xnor U18394 (N_18394,N_17787,N_17867);
or U18395 (N_18395,N_17631,N_17632);
nor U18396 (N_18396,N_17935,N_17825);
nand U18397 (N_18397,N_17883,N_17627);
or U18398 (N_18398,N_17618,N_17756);
or U18399 (N_18399,N_17608,N_17922);
and U18400 (N_18400,N_17552,N_17666);
nand U18401 (N_18401,N_17866,N_17701);
and U18402 (N_18402,N_17708,N_17714);
nor U18403 (N_18403,N_17892,N_17593);
xnor U18404 (N_18404,N_17821,N_17636);
or U18405 (N_18405,N_17554,N_17816);
nand U18406 (N_18406,N_17900,N_17573);
nor U18407 (N_18407,N_17614,N_17516);
nand U18408 (N_18408,N_17761,N_17557);
xnor U18409 (N_18409,N_17587,N_17648);
nand U18410 (N_18410,N_17592,N_17931);
xor U18411 (N_18411,N_17559,N_17723);
xnor U18412 (N_18412,N_17559,N_17776);
nor U18413 (N_18413,N_17519,N_17639);
xor U18414 (N_18414,N_17585,N_17681);
or U18415 (N_18415,N_17520,N_17528);
xnor U18416 (N_18416,N_17884,N_17635);
or U18417 (N_18417,N_17883,N_17916);
nand U18418 (N_18418,N_17679,N_17727);
nor U18419 (N_18419,N_17517,N_17535);
nor U18420 (N_18420,N_17632,N_17999);
xor U18421 (N_18421,N_17614,N_17696);
nand U18422 (N_18422,N_17739,N_17910);
or U18423 (N_18423,N_17763,N_17709);
and U18424 (N_18424,N_17513,N_17785);
and U18425 (N_18425,N_17613,N_17519);
and U18426 (N_18426,N_17641,N_17754);
nor U18427 (N_18427,N_17928,N_17812);
xnor U18428 (N_18428,N_17537,N_17884);
and U18429 (N_18429,N_17911,N_17976);
xnor U18430 (N_18430,N_17559,N_17569);
nor U18431 (N_18431,N_17744,N_17732);
or U18432 (N_18432,N_17772,N_17576);
and U18433 (N_18433,N_17945,N_17995);
nand U18434 (N_18434,N_17861,N_17554);
xnor U18435 (N_18435,N_17886,N_17508);
nand U18436 (N_18436,N_17861,N_17720);
nor U18437 (N_18437,N_17539,N_17883);
xor U18438 (N_18438,N_17600,N_17567);
nor U18439 (N_18439,N_17756,N_17953);
nand U18440 (N_18440,N_17601,N_17623);
xnor U18441 (N_18441,N_17645,N_17624);
xnor U18442 (N_18442,N_17562,N_17633);
xor U18443 (N_18443,N_17570,N_17700);
and U18444 (N_18444,N_17946,N_17829);
or U18445 (N_18445,N_17665,N_17542);
and U18446 (N_18446,N_17695,N_17738);
and U18447 (N_18447,N_17823,N_17630);
xnor U18448 (N_18448,N_17509,N_17640);
xor U18449 (N_18449,N_17598,N_17540);
or U18450 (N_18450,N_17966,N_17739);
xor U18451 (N_18451,N_17637,N_17700);
nor U18452 (N_18452,N_17755,N_17638);
nand U18453 (N_18453,N_17808,N_17817);
and U18454 (N_18454,N_17811,N_17560);
nor U18455 (N_18455,N_17506,N_17659);
xnor U18456 (N_18456,N_17741,N_17524);
nor U18457 (N_18457,N_17944,N_17846);
and U18458 (N_18458,N_17506,N_17507);
nor U18459 (N_18459,N_17756,N_17788);
xor U18460 (N_18460,N_17519,N_17574);
or U18461 (N_18461,N_17713,N_17797);
nand U18462 (N_18462,N_17717,N_17518);
or U18463 (N_18463,N_17581,N_17648);
or U18464 (N_18464,N_17813,N_17905);
or U18465 (N_18465,N_17515,N_17715);
xnor U18466 (N_18466,N_17955,N_17823);
nand U18467 (N_18467,N_17855,N_17505);
and U18468 (N_18468,N_17747,N_17983);
and U18469 (N_18469,N_17920,N_17560);
or U18470 (N_18470,N_17741,N_17776);
xnor U18471 (N_18471,N_17646,N_17884);
or U18472 (N_18472,N_17510,N_17938);
nand U18473 (N_18473,N_17825,N_17586);
nor U18474 (N_18474,N_17883,N_17558);
and U18475 (N_18475,N_17954,N_17902);
nor U18476 (N_18476,N_17547,N_17784);
xnor U18477 (N_18477,N_17671,N_17973);
or U18478 (N_18478,N_17519,N_17916);
and U18479 (N_18479,N_17687,N_17926);
nand U18480 (N_18480,N_17730,N_17979);
and U18481 (N_18481,N_17886,N_17691);
nor U18482 (N_18482,N_17712,N_17866);
or U18483 (N_18483,N_17585,N_17702);
and U18484 (N_18484,N_17793,N_17509);
xnor U18485 (N_18485,N_17766,N_17728);
and U18486 (N_18486,N_17976,N_17772);
nor U18487 (N_18487,N_17636,N_17836);
or U18488 (N_18488,N_17715,N_17588);
xor U18489 (N_18489,N_17683,N_17855);
xnor U18490 (N_18490,N_17500,N_17694);
xnor U18491 (N_18491,N_17684,N_17615);
or U18492 (N_18492,N_17779,N_17579);
nand U18493 (N_18493,N_17516,N_17942);
or U18494 (N_18494,N_17618,N_17531);
or U18495 (N_18495,N_17667,N_17536);
nor U18496 (N_18496,N_17544,N_17629);
or U18497 (N_18497,N_17975,N_17591);
nand U18498 (N_18498,N_17571,N_17633);
nand U18499 (N_18499,N_17601,N_17618);
nor U18500 (N_18500,N_18210,N_18051);
nand U18501 (N_18501,N_18413,N_18009);
xor U18502 (N_18502,N_18481,N_18011);
and U18503 (N_18503,N_18108,N_18468);
nor U18504 (N_18504,N_18129,N_18118);
nand U18505 (N_18505,N_18078,N_18279);
nand U18506 (N_18506,N_18286,N_18484);
xnor U18507 (N_18507,N_18347,N_18115);
nor U18508 (N_18508,N_18159,N_18213);
nand U18509 (N_18509,N_18191,N_18330);
nor U18510 (N_18510,N_18201,N_18271);
nand U18511 (N_18511,N_18250,N_18217);
nand U18512 (N_18512,N_18483,N_18243);
and U18513 (N_18513,N_18200,N_18339);
xor U18514 (N_18514,N_18153,N_18454);
nor U18515 (N_18515,N_18099,N_18391);
xnor U18516 (N_18516,N_18486,N_18378);
or U18517 (N_18517,N_18329,N_18182);
nand U18518 (N_18518,N_18066,N_18097);
or U18519 (N_18519,N_18179,N_18125);
and U18520 (N_18520,N_18290,N_18475);
and U18521 (N_18521,N_18253,N_18448);
nor U18522 (N_18522,N_18398,N_18270);
or U18523 (N_18523,N_18312,N_18462);
and U18524 (N_18524,N_18176,N_18023);
and U18525 (N_18525,N_18084,N_18429);
or U18526 (N_18526,N_18377,N_18111);
xnor U18527 (N_18527,N_18070,N_18300);
xnor U18528 (N_18528,N_18180,N_18247);
and U18529 (N_18529,N_18292,N_18198);
or U18530 (N_18530,N_18225,N_18054);
xnor U18531 (N_18531,N_18249,N_18203);
nand U18532 (N_18532,N_18216,N_18166);
and U18533 (N_18533,N_18031,N_18058);
nand U18534 (N_18534,N_18173,N_18049);
xor U18535 (N_18535,N_18068,N_18245);
nand U18536 (N_18536,N_18367,N_18388);
nand U18537 (N_18537,N_18012,N_18387);
nand U18538 (N_18538,N_18220,N_18206);
and U18539 (N_18539,N_18352,N_18294);
or U18540 (N_18540,N_18114,N_18473);
or U18541 (N_18541,N_18187,N_18440);
or U18542 (N_18542,N_18291,N_18426);
or U18543 (N_18543,N_18053,N_18465);
or U18544 (N_18544,N_18328,N_18326);
nand U18545 (N_18545,N_18255,N_18446);
and U18546 (N_18546,N_18062,N_18241);
or U18547 (N_18547,N_18124,N_18267);
and U18548 (N_18548,N_18237,N_18445);
nor U18549 (N_18549,N_18458,N_18252);
xnor U18550 (N_18550,N_18162,N_18441);
nor U18551 (N_18551,N_18299,N_18412);
nand U18552 (N_18552,N_18007,N_18067);
xnor U18553 (N_18553,N_18197,N_18359);
nor U18554 (N_18554,N_18401,N_18364);
xor U18555 (N_18555,N_18288,N_18490);
and U18556 (N_18556,N_18019,N_18365);
nand U18557 (N_18557,N_18323,N_18382);
or U18558 (N_18558,N_18296,N_18383);
nor U18559 (N_18559,N_18427,N_18144);
or U18560 (N_18560,N_18061,N_18017);
nand U18561 (N_18561,N_18302,N_18374);
nor U18562 (N_18562,N_18188,N_18319);
and U18563 (N_18563,N_18466,N_18244);
nor U18564 (N_18564,N_18010,N_18022);
and U18565 (N_18565,N_18327,N_18452);
xor U18566 (N_18566,N_18029,N_18100);
and U18567 (N_18567,N_18467,N_18492);
xor U18568 (N_18568,N_18306,N_18167);
nor U18569 (N_18569,N_18417,N_18092);
nor U18570 (N_18570,N_18331,N_18334);
xor U18571 (N_18571,N_18231,N_18322);
nand U18572 (N_18572,N_18212,N_18280);
and U18573 (N_18573,N_18154,N_18227);
or U18574 (N_18574,N_18041,N_18254);
nand U18575 (N_18575,N_18433,N_18172);
xor U18576 (N_18576,N_18119,N_18344);
xor U18577 (N_18577,N_18015,N_18464);
and U18578 (N_18578,N_18091,N_18222);
xor U18579 (N_18579,N_18209,N_18480);
nor U18580 (N_18580,N_18397,N_18205);
and U18581 (N_18581,N_18149,N_18236);
or U18582 (N_18582,N_18190,N_18263);
nand U18583 (N_18583,N_18341,N_18335);
or U18584 (N_18584,N_18064,N_18207);
nand U18585 (N_18585,N_18076,N_18265);
and U18586 (N_18586,N_18143,N_18351);
and U18587 (N_18587,N_18109,N_18141);
xor U18588 (N_18588,N_18314,N_18379);
xor U18589 (N_18589,N_18059,N_18419);
and U18590 (N_18590,N_18275,N_18434);
nand U18591 (N_18591,N_18442,N_18407);
nor U18592 (N_18592,N_18333,N_18194);
or U18593 (N_18593,N_18324,N_18251);
xnor U18594 (N_18594,N_18080,N_18307);
and U18595 (N_18595,N_18455,N_18376);
or U18596 (N_18596,N_18199,N_18134);
or U18597 (N_18597,N_18140,N_18348);
nor U18598 (N_18598,N_18037,N_18077);
or U18599 (N_18599,N_18408,N_18082);
xor U18600 (N_18600,N_18242,N_18380);
nor U18601 (N_18601,N_18152,N_18355);
and U18602 (N_18602,N_18024,N_18073);
or U18603 (N_18603,N_18298,N_18156);
nand U18604 (N_18604,N_18132,N_18451);
nor U18605 (N_18605,N_18420,N_18346);
and U18606 (N_18606,N_18121,N_18219);
and U18607 (N_18607,N_18120,N_18033);
and U18608 (N_18608,N_18470,N_18342);
and U18609 (N_18609,N_18192,N_18488);
nor U18610 (N_18610,N_18196,N_18360);
and U18611 (N_18611,N_18297,N_18085);
and U18612 (N_18612,N_18142,N_18357);
nor U18613 (N_18613,N_18261,N_18487);
or U18614 (N_18614,N_18040,N_18272);
and U18615 (N_18615,N_18406,N_18095);
and U18616 (N_18616,N_18349,N_18164);
nor U18617 (N_18617,N_18148,N_18060);
and U18618 (N_18618,N_18226,N_18287);
nand U18619 (N_18619,N_18447,N_18093);
or U18620 (N_18620,N_18424,N_18425);
xor U18621 (N_18621,N_18276,N_18128);
or U18622 (N_18622,N_18138,N_18171);
or U18623 (N_18623,N_18453,N_18087);
nand U18624 (N_18624,N_18285,N_18145);
xnor U18625 (N_18625,N_18014,N_18256);
nand U18626 (N_18626,N_18423,N_18411);
xor U18627 (N_18627,N_18289,N_18325);
and U18628 (N_18628,N_18358,N_18135);
xor U18629 (N_18629,N_18083,N_18372);
and U18630 (N_18630,N_18421,N_18257);
or U18631 (N_18631,N_18018,N_18338);
or U18632 (N_18632,N_18089,N_18384);
nand U18633 (N_18633,N_18160,N_18181);
and U18634 (N_18634,N_18146,N_18394);
xor U18635 (N_18635,N_18479,N_18110);
nand U18636 (N_18636,N_18238,N_18195);
and U18637 (N_18637,N_18021,N_18337);
nand U18638 (N_18638,N_18170,N_18090);
nand U18639 (N_18639,N_18034,N_18248);
or U18640 (N_18640,N_18370,N_18165);
nand U18641 (N_18641,N_18386,N_18320);
and U18642 (N_18642,N_18321,N_18476);
or U18643 (N_18643,N_18042,N_18035);
or U18644 (N_18644,N_18028,N_18472);
or U18645 (N_18645,N_18268,N_18079);
and U18646 (N_18646,N_18157,N_18178);
nand U18647 (N_18647,N_18431,N_18032);
xor U18648 (N_18648,N_18202,N_18013);
and U18649 (N_18649,N_18390,N_18381);
xor U18650 (N_18650,N_18074,N_18046);
nand U18651 (N_18651,N_18311,N_18027);
or U18652 (N_18652,N_18150,N_18282);
nor U18653 (N_18653,N_18277,N_18036);
xor U18654 (N_18654,N_18395,N_18436);
or U18655 (N_18655,N_18356,N_18163);
or U18656 (N_18656,N_18112,N_18235);
nor U18657 (N_18657,N_18402,N_18315);
and U18658 (N_18658,N_18052,N_18081);
or U18659 (N_18659,N_18204,N_18189);
or U18660 (N_18660,N_18432,N_18185);
and U18661 (N_18661,N_18169,N_18489);
nor U18662 (N_18662,N_18416,N_18496);
nor U18663 (N_18663,N_18105,N_18404);
or U18664 (N_18664,N_18044,N_18385);
nor U18665 (N_18665,N_18158,N_18422);
and U18666 (N_18666,N_18233,N_18403);
nor U18667 (N_18667,N_18008,N_18177);
or U18668 (N_18668,N_18332,N_18350);
nor U18669 (N_18669,N_18122,N_18269);
or U18670 (N_18670,N_18369,N_18246);
or U18671 (N_18671,N_18495,N_18025);
or U18672 (N_18672,N_18450,N_18086);
or U18673 (N_18673,N_18463,N_18001);
or U18674 (N_18674,N_18497,N_18006);
and U18675 (N_18675,N_18396,N_18106);
nand U18676 (N_18676,N_18469,N_18107);
or U18677 (N_18677,N_18284,N_18224);
or U18678 (N_18678,N_18435,N_18499);
and U18679 (N_18679,N_18259,N_18116);
and U18680 (N_18680,N_18439,N_18030);
xnor U18681 (N_18681,N_18096,N_18260);
or U18682 (N_18682,N_18047,N_18234);
nand U18683 (N_18683,N_18309,N_18283);
nand U18684 (N_18684,N_18437,N_18399);
xnor U18685 (N_18685,N_18005,N_18461);
nand U18686 (N_18686,N_18045,N_18123);
or U18687 (N_18687,N_18147,N_18211);
xnor U18688 (N_18688,N_18186,N_18175);
xor U18689 (N_18689,N_18354,N_18094);
nor U18690 (N_18690,N_18183,N_18214);
and U18691 (N_18691,N_18155,N_18151);
xor U18692 (N_18692,N_18363,N_18438);
nor U18693 (N_18693,N_18418,N_18343);
xor U18694 (N_18694,N_18498,N_18477);
xnor U18695 (N_18695,N_18471,N_18136);
or U18696 (N_18696,N_18139,N_18003);
or U18697 (N_18697,N_18016,N_18168);
or U18698 (N_18698,N_18117,N_18460);
or U18699 (N_18699,N_18230,N_18184);
nand U18700 (N_18700,N_18273,N_18295);
and U18701 (N_18701,N_18056,N_18389);
xor U18702 (N_18702,N_18494,N_18039);
or U18703 (N_18703,N_18137,N_18414);
or U18704 (N_18704,N_18057,N_18362);
and U18705 (N_18705,N_18101,N_18050);
nand U18706 (N_18706,N_18308,N_18443);
or U18707 (N_18707,N_18239,N_18072);
nand U18708 (N_18708,N_18313,N_18310);
nor U18709 (N_18709,N_18258,N_18336);
nand U18710 (N_18710,N_18459,N_18221);
nand U18711 (N_18711,N_18223,N_18065);
and U18712 (N_18712,N_18228,N_18069);
or U18713 (N_18713,N_18161,N_18055);
nor U18714 (N_18714,N_18405,N_18174);
xnor U18715 (N_18715,N_18215,N_18102);
nand U18716 (N_18716,N_18491,N_18126);
nor U18717 (N_18717,N_18193,N_18368);
nor U18718 (N_18718,N_18127,N_18361);
and U18719 (N_18719,N_18043,N_18371);
xor U18720 (N_18720,N_18305,N_18318);
and U18721 (N_18721,N_18493,N_18340);
or U18722 (N_18722,N_18232,N_18410);
xor U18723 (N_18723,N_18345,N_18373);
nand U18724 (N_18724,N_18104,N_18000);
nand U18725 (N_18725,N_18485,N_18366);
nand U18726 (N_18726,N_18444,N_18088);
nand U18727 (N_18727,N_18278,N_18304);
and U18728 (N_18728,N_18415,N_18474);
nor U18729 (N_18729,N_18482,N_18301);
nor U18730 (N_18730,N_18038,N_18020);
xnor U18731 (N_18731,N_18430,N_18208);
or U18732 (N_18732,N_18375,N_18130);
xnor U18733 (N_18733,N_18002,N_18457);
nor U18734 (N_18734,N_18264,N_18478);
xnor U18735 (N_18735,N_18133,N_18131);
nand U18736 (N_18736,N_18048,N_18303);
and U18737 (N_18737,N_18240,N_18393);
xor U18738 (N_18738,N_18317,N_18428);
and U18739 (N_18739,N_18281,N_18071);
xnor U18740 (N_18740,N_18075,N_18392);
or U18741 (N_18741,N_18449,N_18113);
nor U18742 (N_18742,N_18229,N_18103);
xnor U18743 (N_18743,N_18353,N_18266);
nand U18744 (N_18744,N_18293,N_18316);
nor U18745 (N_18745,N_18098,N_18274);
or U18746 (N_18746,N_18400,N_18456);
or U18747 (N_18747,N_18262,N_18409);
nor U18748 (N_18748,N_18026,N_18218);
or U18749 (N_18749,N_18063,N_18004);
nand U18750 (N_18750,N_18383,N_18386);
nor U18751 (N_18751,N_18245,N_18180);
or U18752 (N_18752,N_18021,N_18463);
or U18753 (N_18753,N_18257,N_18243);
or U18754 (N_18754,N_18324,N_18309);
and U18755 (N_18755,N_18140,N_18351);
xnor U18756 (N_18756,N_18028,N_18306);
nand U18757 (N_18757,N_18174,N_18427);
or U18758 (N_18758,N_18308,N_18284);
and U18759 (N_18759,N_18389,N_18483);
nor U18760 (N_18760,N_18404,N_18463);
or U18761 (N_18761,N_18403,N_18162);
xor U18762 (N_18762,N_18487,N_18358);
nor U18763 (N_18763,N_18249,N_18379);
nand U18764 (N_18764,N_18218,N_18113);
and U18765 (N_18765,N_18312,N_18390);
nand U18766 (N_18766,N_18489,N_18443);
nand U18767 (N_18767,N_18133,N_18474);
and U18768 (N_18768,N_18365,N_18067);
xor U18769 (N_18769,N_18499,N_18450);
nand U18770 (N_18770,N_18294,N_18435);
or U18771 (N_18771,N_18319,N_18068);
nand U18772 (N_18772,N_18463,N_18212);
or U18773 (N_18773,N_18383,N_18488);
nand U18774 (N_18774,N_18466,N_18431);
or U18775 (N_18775,N_18029,N_18432);
or U18776 (N_18776,N_18375,N_18188);
xor U18777 (N_18777,N_18125,N_18007);
nand U18778 (N_18778,N_18202,N_18201);
nor U18779 (N_18779,N_18255,N_18427);
and U18780 (N_18780,N_18139,N_18434);
or U18781 (N_18781,N_18255,N_18284);
or U18782 (N_18782,N_18117,N_18105);
xor U18783 (N_18783,N_18495,N_18402);
and U18784 (N_18784,N_18060,N_18469);
xor U18785 (N_18785,N_18323,N_18156);
nor U18786 (N_18786,N_18248,N_18008);
nand U18787 (N_18787,N_18480,N_18456);
nand U18788 (N_18788,N_18384,N_18288);
nand U18789 (N_18789,N_18152,N_18047);
xnor U18790 (N_18790,N_18316,N_18087);
and U18791 (N_18791,N_18032,N_18158);
nor U18792 (N_18792,N_18397,N_18498);
nor U18793 (N_18793,N_18142,N_18171);
or U18794 (N_18794,N_18466,N_18051);
xor U18795 (N_18795,N_18150,N_18309);
or U18796 (N_18796,N_18258,N_18459);
and U18797 (N_18797,N_18325,N_18424);
or U18798 (N_18798,N_18063,N_18054);
xor U18799 (N_18799,N_18099,N_18223);
nand U18800 (N_18800,N_18441,N_18145);
nor U18801 (N_18801,N_18277,N_18147);
or U18802 (N_18802,N_18057,N_18385);
nand U18803 (N_18803,N_18160,N_18123);
and U18804 (N_18804,N_18401,N_18499);
and U18805 (N_18805,N_18336,N_18182);
or U18806 (N_18806,N_18157,N_18334);
nor U18807 (N_18807,N_18266,N_18470);
nand U18808 (N_18808,N_18091,N_18340);
nor U18809 (N_18809,N_18458,N_18439);
nand U18810 (N_18810,N_18419,N_18167);
nand U18811 (N_18811,N_18006,N_18218);
or U18812 (N_18812,N_18172,N_18168);
nand U18813 (N_18813,N_18362,N_18062);
and U18814 (N_18814,N_18059,N_18266);
nor U18815 (N_18815,N_18116,N_18114);
nand U18816 (N_18816,N_18297,N_18469);
nand U18817 (N_18817,N_18144,N_18214);
or U18818 (N_18818,N_18184,N_18003);
and U18819 (N_18819,N_18219,N_18499);
nand U18820 (N_18820,N_18265,N_18274);
nor U18821 (N_18821,N_18141,N_18308);
nand U18822 (N_18822,N_18236,N_18273);
xor U18823 (N_18823,N_18056,N_18013);
xnor U18824 (N_18824,N_18018,N_18448);
nand U18825 (N_18825,N_18048,N_18381);
nor U18826 (N_18826,N_18132,N_18035);
and U18827 (N_18827,N_18026,N_18163);
xnor U18828 (N_18828,N_18055,N_18331);
or U18829 (N_18829,N_18256,N_18054);
nand U18830 (N_18830,N_18355,N_18123);
nor U18831 (N_18831,N_18316,N_18010);
nor U18832 (N_18832,N_18059,N_18064);
and U18833 (N_18833,N_18216,N_18459);
nor U18834 (N_18834,N_18296,N_18293);
nor U18835 (N_18835,N_18018,N_18284);
nor U18836 (N_18836,N_18306,N_18257);
nand U18837 (N_18837,N_18393,N_18208);
and U18838 (N_18838,N_18295,N_18105);
and U18839 (N_18839,N_18197,N_18098);
or U18840 (N_18840,N_18441,N_18361);
or U18841 (N_18841,N_18023,N_18369);
nand U18842 (N_18842,N_18414,N_18486);
xor U18843 (N_18843,N_18292,N_18117);
nor U18844 (N_18844,N_18402,N_18181);
nor U18845 (N_18845,N_18377,N_18423);
nand U18846 (N_18846,N_18100,N_18308);
and U18847 (N_18847,N_18101,N_18366);
nand U18848 (N_18848,N_18343,N_18279);
nor U18849 (N_18849,N_18226,N_18080);
and U18850 (N_18850,N_18041,N_18169);
xor U18851 (N_18851,N_18174,N_18299);
and U18852 (N_18852,N_18022,N_18119);
and U18853 (N_18853,N_18424,N_18176);
and U18854 (N_18854,N_18017,N_18132);
nor U18855 (N_18855,N_18008,N_18457);
nor U18856 (N_18856,N_18027,N_18151);
xor U18857 (N_18857,N_18157,N_18395);
or U18858 (N_18858,N_18047,N_18008);
nand U18859 (N_18859,N_18171,N_18192);
nor U18860 (N_18860,N_18175,N_18345);
and U18861 (N_18861,N_18269,N_18375);
xnor U18862 (N_18862,N_18101,N_18294);
and U18863 (N_18863,N_18388,N_18211);
or U18864 (N_18864,N_18307,N_18051);
or U18865 (N_18865,N_18229,N_18248);
nor U18866 (N_18866,N_18034,N_18009);
nand U18867 (N_18867,N_18317,N_18144);
nand U18868 (N_18868,N_18310,N_18316);
or U18869 (N_18869,N_18332,N_18413);
and U18870 (N_18870,N_18096,N_18421);
and U18871 (N_18871,N_18077,N_18176);
or U18872 (N_18872,N_18084,N_18400);
nand U18873 (N_18873,N_18286,N_18280);
nor U18874 (N_18874,N_18318,N_18307);
xor U18875 (N_18875,N_18416,N_18305);
nor U18876 (N_18876,N_18494,N_18242);
nor U18877 (N_18877,N_18031,N_18137);
nand U18878 (N_18878,N_18042,N_18370);
xor U18879 (N_18879,N_18364,N_18142);
nor U18880 (N_18880,N_18068,N_18394);
nand U18881 (N_18881,N_18106,N_18198);
nand U18882 (N_18882,N_18460,N_18471);
and U18883 (N_18883,N_18393,N_18295);
nor U18884 (N_18884,N_18083,N_18381);
nor U18885 (N_18885,N_18165,N_18288);
or U18886 (N_18886,N_18204,N_18499);
nand U18887 (N_18887,N_18021,N_18179);
or U18888 (N_18888,N_18160,N_18024);
xor U18889 (N_18889,N_18115,N_18038);
or U18890 (N_18890,N_18221,N_18416);
nor U18891 (N_18891,N_18169,N_18252);
or U18892 (N_18892,N_18346,N_18392);
or U18893 (N_18893,N_18435,N_18448);
or U18894 (N_18894,N_18132,N_18099);
nand U18895 (N_18895,N_18459,N_18450);
nor U18896 (N_18896,N_18069,N_18473);
and U18897 (N_18897,N_18108,N_18044);
xnor U18898 (N_18898,N_18195,N_18026);
nand U18899 (N_18899,N_18190,N_18230);
or U18900 (N_18900,N_18462,N_18466);
nand U18901 (N_18901,N_18146,N_18177);
xor U18902 (N_18902,N_18153,N_18162);
nor U18903 (N_18903,N_18215,N_18194);
nor U18904 (N_18904,N_18435,N_18322);
nand U18905 (N_18905,N_18199,N_18174);
nand U18906 (N_18906,N_18086,N_18132);
and U18907 (N_18907,N_18049,N_18315);
nor U18908 (N_18908,N_18413,N_18103);
nand U18909 (N_18909,N_18321,N_18414);
or U18910 (N_18910,N_18346,N_18250);
nand U18911 (N_18911,N_18042,N_18464);
or U18912 (N_18912,N_18381,N_18349);
and U18913 (N_18913,N_18267,N_18297);
nor U18914 (N_18914,N_18499,N_18283);
nand U18915 (N_18915,N_18399,N_18192);
xor U18916 (N_18916,N_18281,N_18373);
nand U18917 (N_18917,N_18044,N_18226);
nor U18918 (N_18918,N_18447,N_18470);
xnor U18919 (N_18919,N_18133,N_18141);
and U18920 (N_18920,N_18473,N_18403);
xnor U18921 (N_18921,N_18098,N_18434);
and U18922 (N_18922,N_18254,N_18042);
nand U18923 (N_18923,N_18075,N_18491);
or U18924 (N_18924,N_18181,N_18150);
nand U18925 (N_18925,N_18196,N_18118);
and U18926 (N_18926,N_18156,N_18458);
and U18927 (N_18927,N_18155,N_18427);
nand U18928 (N_18928,N_18417,N_18038);
nor U18929 (N_18929,N_18313,N_18162);
and U18930 (N_18930,N_18062,N_18153);
xor U18931 (N_18931,N_18038,N_18268);
xnor U18932 (N_18932,N_18199,N_18293);
and U18933 (N_18933,N_18311,N_18443);
nand U18934 (N_18934,N_18183,N_18472);
and U18935 (N_18935,N_18330,N_18458);
nor U18936 (N_18936,N_18481,N_18293);
and U18937 (N_18937,N_18239,N_18383);
and U18938 (N_18938,N_18116,N_18278);
nand U18939 (N_18939,N_18186,N_18166);
and U18940 (N_18940,N_18377,N_18339);
nand U18941 (N_18941,N_18186,N_18436);
or U18942 (N_18942,N_18444,N_18000);
xor U18943 (N_18943,N_18344,N_18289);
nand U18944 (N_18944,N_18346,N_18344);
and U18945 (N_18945,N_18155,N_18470);
or U18946 (N_18946,N_18346,N_18257);
xor U18947 (N_18947,N_18216,N_18205);
or U18948 (N_18948,N_18417,N_18303);
xor U18949 (N_18949,N_18126,N_18314);
nor U18950 (N_18950,N_18361,N_18072);
xor U18951 (N_18951,N_18252,N_18488);
nor U18952 (N_18952,N_18062,N_18277);
or U18953 (N_18953,N_18450,N_18331);
and U18954 (N_18954,N_18311,N_18037);
nor U18955 (N_18955,N_18478,N_18300);
or U18956 (N_18956,N_18034,N_18276);
and U18957 (N_18957,N_18395,N_18099);
nor U18958 (N_18958,N_18209,N_18271);
and U18959 (N_18959,N_18009,N_18398);
nor U18960 (N_18960,N_18239,N_18250);
xnor U18961 (N_18961,N_18035,N_18423);
and U18962 (N_18962,N_18199,N_18300);
nand U18963 (N_18963,N_18167,N_18185);
nand U18964 (N_18964,N_18315,N_18196);
xor U18965 (N_18965,N_18137,N_18053);
nor U18966 (N_18966,N_18401,N_18417);
or U18967 (N_18967,N_18055,N_18044);
nand U18968 (N_18968,N_18153,N_18202);
and U18969 (N_18969,N_18471,N_18475);
xor U18970 (N_18970,N_18410,N_18458);
and U18971 (N_18971,N_18222,N_18423);
xor U18972 (N_18972,N_18348,N_18003);
or U18973 (N_18973,N_18090,N_18001);
nand U18974 (N_18974,N_18457,N_18365);
nor U18975 (N_18975,N_18418,N_18414);
xnor U18976 (N_18976,N_18119,N_18116);
nand U18977 (N_18977,N_18041,N_18399);
xor U18978 (N_18978,N_18335,N_18125);
xnor U18979 (N_18979,N_18042,N_18465);
or U18980 (N_18980,N_18140,N_18035);
or U18981 (N_18981,N_18309,N_18357);
and U18982 (N_18982,N_18256,N_18286);
nand U18983 (N_18983,N_18447,N_18326);
xnor U18984 (N_18984,N_18339,N_18353);
nor U18985 (N_18985,N_18398,N_18090);
and U18986 (N_18986,N_18405,N_18236);
or U18987 (N_18987,N_18210,N_18402);
nor U18988 (N_18988,N_18483,N_18414);
xor U18989 (N_18989,N_18118,N_18097);
and U18990 (N_18990,N_18234,N_18185);
or U18991 (N_18991,N_18120,N_18012);
nand U18992 (N_18992,N_18217,N_18293);
and U18993 (N_18993,N_18426,N_18270);
nand U18994 (N_18994,N_18325,N_18316);
xnor U18995 (N_18995,N_18048,N_18424);
or U18996 (N_18996,N_18085,N_18219);
and U18997 (N_18997,N_18449,N_18326);
nor U18998 (N_18998,N_18452,N_18473);
nand U18999 (N_18999,N_18252,N_18198);
nand U19000 (N_19000,N_18960,N_18621);
and U19001 (N_19001,N_18702,N_18793);
nor U19002 (N_19002,N_18779,N_18601);
or U19003 (N_19003,N_18772,N_18656);
xnor U19004 (N_19004,N_18883,N_18941);
or U19005 (N_19005,N_18928,N_18874);
xnor U19006 (N_19006,N_18940,N_18629);
or U19007 (N_19007,N_18857,N_18548);
xnor U19008 (N_19008,N_18682,N_18972);
nand U19009 (N_19009,N_18732,N_18627);
or U19010 (N_19010,N_18892,N_18692);
or U19011 (N_19011,N_18937,N_18908);
and U19012 (N_19012,N_18554,N_18983);
or U19013 (N_19013,N_18582,N_18947);
and U19014 (N_19014,N_18865,N_18859);
xnor U19015 (N_19015,N_18804,N_18596);
xnor U19016 (N_19016,N_18815,N_18673);
nand U19017 (N_19017,N_18752,N_18990);
nor U19018 (N_19018,N_18574,N_18878);
nand U19019 (N_19019,N_18899,N_18800);
xnor U19020 (N_19020,N_18630,N_18733);
nand U19021 (N_19021,N_18560,N_18696);
nor U19022 (N_19022,N_18666,N_18506);
and U19023 (N_19023,N_18740,N_18712);
nand U19024 (N_19024,N_18739,N_18890);
and U19025 (N_19025,N_18715,N_18895);
nand U19026 (N_19026,N_18515,N_18557);
and U19027 (N_19027,N_18658,N_18994);
nor U19028 (N_19028,N_18597,N_18897);
nand U19029 (N_19029,N_18681,N_18575);
nand U19030 (N_19030,N_18829,N_18588);
nand U19031 (N_19031,N_18850,N_18900);
or U19032 (N_19032,N_18759,N_18765);
and U19033 (N_19033,N_18573,N_18884);
nor U19034 (N_19034,N_18813,N_18507);
xnor U19035 (N_19035,N_18531,N_18710);
xnor U19036 (N_19036,N_18678,N_18611);
xor U19037 (N_19037,N_18959,N_18663);
xnor U19038 (N_19038,N_18585,N_18555);
or U19039 (N_19039,N_18768,N_18542);
and U19040 (N_19040,N_18709,N_18769);
nor U19041 (N_19041,N_18910,N_18721);
nand U19042 (N_19042,N_18571,N_18838);
nand U19043 (N_19043,N_18747,N_18835);
or U19044 (N_19044,N_18978,N_18816);
nand U19045 (N_19045,N_18840,N_18902);
xnor U19046 (N_19046,N_18823,N_18610);
or U19047 (N_19047,N_18862,N_18876);
nor U19048 (N_19048,N_18618,N_18736);
or U19049 (N_19049,N_18967,N_18684);
and U19050 (N_19050,N_18975,N_18837);
xor U19051 (N_19051,N_18523,N_18821);
xor U19052 (N_19052,N_18955,N_18671);
xor U19053 (N_19053,N_18849,N_18676);
xor U19054 (N_19054,N_18638,N_18964);
or U19055 (N_19055,N_18672,N_18654);
nor U19056 (N_19056,N_18894,N_18547);
xor U19057 (N_19057,N_18784,N_18819);
xnor U19058 (N_19058,N_18510,N_18737);
and U19059 (N_19059,N_18650,N_18980);
or U19060 (N_19060,N_18754,N_18688);
or U19061 (N_19061,N_18750,N_18742);
or U19062 (N_19062,N_18636,N_18807);
nor U19063 (N_19063,N_18956,N_18581);
or U19064 (N_19064,N_18648,N_18877);
or U19065 (N_19065,N_18624,N_18602);
and U19066 (N_19066,N_18701,N_18860);
nand U19067 (N_19067,N_18896,N_18934);
or U19068 (N_19068,N_18679,N_18616);
xnor U19069 (N_19069,N_18628,N_18834);
or U19070 (N_19070,N_18758,N_18801);
and U19071 (N_19071,N_18609,N_18786);
xor U19072 (N_19072,N_18851,N_18643);
nor U19073 (N_19073,N_18642,N_18566);
or U19074 (N_19074,N_18761,N_18968);
nand U19075 (N_19075,N_18722,N_18870);
nand U19076 (N_19076,N_18619,N_18848);
or U19077 (N_19077,N_18526,N_18683);
or U19078 (N_19078,N_18923,N_18993);
and U19079 (N_19079,N_18977,N_18519);
xnor U19080 (N_19080,N_18952,N_18522);
nor U19081 (N_19081,N_18958,N_18949);
xor U19082 (N_19082,N_18824,N_18713);
nand U19083 (N_19083,N_18961,N_18505);
nor U19084 (N_19084,N_18562,N_18511);
and U19085 (N_19085,N_18795,N_18707);
nand U19086 (N_19086,N_18518,N_18527);
and U19087 (N_19087,N_18730,N_18734);
nor U19088 (N_19088,N_18844,N_18647);
nor U19089 (N_19089,N_18625,N_18659);
nor U19090 (N_19090,N_18741,N_18728);
xnor U19091 (N_19091,N_18589,N_18533);
or U19092 (N_19092,N_18942,N_18861);
xor U19093 (N_19093,N_18568,N_18864);
nand U19094 (N_19094,N_18953,N_18546);
nand U19095 (N_19095,N_18782,N_18595);
or U19096 (N_19096,N_18916,N_18974);
nor U19097 (N_19097,N_18693,N_18988);
and U19098 (N_19098,N_18564,N_18634);
or U19099 (N_19099,N_18969,N_18987);
or U19100 (N_19100,N_18704,N_18528);
and U19101 (N_19101,N_18986,N_18996);
nand U19102 (N_19102,N_18637,N_18600);
and U19103 (N_19103,N_18748,N_18918);
or U19104 (N_19104,N_18976,N_18592);
nand U19105 (N_19105,N_18871,N_18852);
and U19106 (N_19106,N_18911,N_18771);
nor U19107 (N_19107,N_18500,N_18605);
xor U19108 (N_19108,N_18863,N_18646);
xor U19109 (N_19109,N_18965,N_18790);
nand U19110 (N_19110,N_18622,N_18989);
and U19111 (N_19111,N_18762,N_18567);
nor U19112 (N_19112,N_18898,N_18788);
xnor U19113 (N_19113,N_18590,N_18887);
and U19114 (N_19114,N_18924,N_18631);
nor U19115 (N_19115,N_18919,N_18775);
or U19116 (N_19116,N_18751,N_18945);
nand U19117 (N_19117,N_18708,N_18579);
or U19118 (N_19118,N_18551,N_18591);
xor U19119 (N_19119,N_18984,N_18660);
and U19120 (N_19120,N_18901,N_18735);
nor U19121 (N_19121,N_18723,N_18904);
nor U19122 (N_19122,N_18820,N_18925);
xor U19123 (N_19123,N_18729,N_18513);
and U19124 (N_19124,N_18879,N_18839);
nand U19125 (N_19125,N_18875,N_18830);
nor U19126 (N_19126,N_18806,N_18537);
and U19127 (N_19127,N_18530,N_18770);
xnor U19128 (N_19128,N_18661,N_18933);
nand U19129 (N_19129,N_18749,N_18694);
or U19130 (N_19130,N_18586,N_18503);
and U19131 (N_19131,N_18517,N_18615);
xor U19132 (N_19132,N_18556,N_18799);
xor U19133 (N_19133,N_18843,N_18936);
or U19134 (N_19134,N_18598,N_18787);
nor U19135 (N_19135,N_18954,N_18827);
or U19136 (N_19136,N_18982,N_18664);
nor U19137 (N_19137,N_18550,N_18690);
or U19138 (N_19138,N_18998,N_18726);
nor U19139 (N_19139,N_18888,N_18791);
xor U19140 (N_19140,N_18535,N_18508);
and U19141 (N_19141,N_18979,N_18842);
nand U19142 (N_19142,N_18691,N_18521);
and U19143 (N_19143,N_18803,N_18716);
nand U19144 (N_19144,N_18536,N_18767);
nand U19145 (N_19145,N_18962,N_18623);
nor U19146 (N_19146,N_18633,N_18549);
and U19147 (N_19147,N_18774,N_18826);
xnor U19148 (N_19148,N_18603,N_18810);
nand U19149 (N_19149,N_18680,N_18565);
nand U19150 (N_19150,N_18607,N_18699);
and U19151 (N_19151,N_18669,N_18753);
nand U19152 (N_19152,N_18698,N_18563);
xor U19153 (N_19153,N_18612,N_18572);
nor U19154 (N_19154,N_18997,N_18743);
or U19155 (N_19155,N_18685,N_18697);
nor U19156 (N_19156,N_18948,N_18662);
nor U19157 (N_19157,N_18912,N_18906);
nor U19158 (N_19158,N_18532,N_18525);
or U19159 (N_19159,N_18738,N_18516);
nor U19160 (N_19160,N_18655,N_18846);
or U19161 (N_19161,N_18921,N_18985);
nand U19162 (N_19162,N_18881,N_18893);
or U19163 (N_19163,N_18845,N_18794);
nand U19164 (N_19164,N_18746,N_18577);
or U19165 (N_19165,N_18913,N_18653);
nand U19166 (N_19166,N_18886,N_18825);
nand U19167 (N_19167,N_18544,N_18995);
and U19168 (N_19168,N_18926,N_18635);
nor U19169 (N_19169,N_18714,N_18868);
nand U19170 (N_19170,N_18543,N_18727);
and U19171 (N_19171,N_18812,N_18882);
or U19172 (N_19172,N_18966,N_18781);
nor U19173 (N_19173,N_18731,N_18760);
and U19174 (N_19174,N_18785,N_18814);
xor U19175 (N_19175,N_18764,N_18705);
or U19176 (N_19176,N_18808,N_18855);
or U19177 (N_19177,N_18944,N_18687);
nand U19178 (N_19178,N_18614,N_18796);
and U19179 (N_19179,N_18719,N_18501);
nor U19180 (N_19180,N_18540,N_18641);
or U19181 (N_19181,N_18724,N_18828);
and U19182 (N_19182,N_18670,N_18700);
and U19183 (N_19183,N_18689,N_18970);
or U19184 (N_19184,N_18817,N_18584);
xor U19185 (N_19185,N_18880,N_18915);
nor U19186 (N_19186,N_18538,N_18905);
or U19187 (N_19187,N_18873,N_18939);
nand U19188 (N_19188,N_18756,N_18657);
xnor U19189 (N_19189,N_18576,N_18599);
nand U19190 (N_19190,N_18668,N_18539);
xor U19191 (N_19191,N_18512,N_18504);
or U19192 (N_19192,N_18578,N_18640);
and U19193 (N_19193,N_18755,N_18675);
and U19194 (N_19194,N_18608,N_18836);
or U19195 (N_19195,N_18792,N_18797);
and U19196 (N_19196,N_18502,N_18514);
nor U19197 (N_19197,N_18951,N_18541);
nand U19198 (N_19198,N_18667,N_18917);
xor U19199 (N_19199,N_18773,N_18626);
and U19200 (N_19200,N_18776,N_18822);
and U19201 (N_19201,N_18811,N_18981);
nand U19202 (N_19202,N_18652,N_18674);
or U19203 (N_19203,N_18718,N_18677);
nand U19204 (N_19204,N_18922,N_18867);
or U19205 (N_19205,N_18720,N_18620);
xnor U19206 (N_19206,N_18927,N_18903);
and U19207 (N_19207,N_18999,N_18725);
xnor U19208 (N_19208,N_18963,N_18858);
or U19209 (N_19209,N_18766,N_18569);
and U19210 (N_19210,N_18872,N_18931);
xnor U19211 (N_19211,N_18920,N_18534);
xor U19212 (N_19212,N_18606,N_18932);
nand U19213 (N_19213,N_18891,N_18703);
nor U19214 (N_19214,N_18744,N_18950);
xor U19215 (N_19215,N_18545,N_18798);
or U19216 (N_19216,N_18757,N_18853);
or U19217 (N_19217,N_18587,N_18909);
nor U19218 (N_19218,N_18706,N_18869);
nand U19219 (N_19219,N_18973,N_18789);
or U19220 (N_19220,N_18818,N_18866);
xnor U19221 (N_19221,N_18552,N_18559);
or U19222 (N_19222,N_18717,N_18832);
nor U19223 (N_19223,N_18971,N_18778);
nand U19224 (N_19224,N_18847,N_18889);
and U19225 (N_19225,N_18617,N_18763);
nor U19226 (N_19226,N_18929,N_18651);
nand U19227 (N_19227,N_18529,N_18802);
or U19228 (N_19228,N_18558,N_18854);
nand U19229 (N_19229,N_18780,N_18809);
or U19230 (N_19230,N_18841,N_18649);
and U19231 (N_19231,N_18520,N_18665);
and U19232 (N_19232,N_18686,N_18524);
xnor U19233 (N_19233,N_18580,N_18935);
nor U19234 (N_19234,N_18644,N_18938);
and U19235 (N_19235,N_18561,N_18946);
nor U19236 (N_19236,N_18833,N_18632);
xnor U19237 (N_19237,N_18594,N_18613);
nor U19238 (N_19238,N_18509,N_18570);
or U19239 (N_19239,N_18695,N_18992);
nor U19240 (N_19240,N_18885,N_18907);
nor U19241 (N_19241,N_18783,N_18957);
nand U19242 (N_19242,N_18856,N_18930);
xnor U19243 (N_19243,N_18645,N_18943);
nand U19244 (N_19244,N_18711,N_18583);
and U19245 (N_19245,N_18593,N_18553);
nand U19246 (N_19246,N_18831,N_18805);
xnor U19247 (N_19247,N_18604,N_18991);
and U19248 (N_19248,N_18745,N_18777);
nand U19249 (N_19249,N_18639,N_18914);
nor U19250 (N_19250,N_18864,N_18704);
nor U19251 (N_19251,N_18999,N_18987);
nand U19252 (N_19252,N_18745,N_18583);
or U19253 (N_19253,N_18910,N_18745);
or U19254 (N_19254,N_18590,N_18922);
xor U19255 (N_19255,N_18627,N_18555);
and U19256 (N_19256,N_18581,N_18679);
or U19257 (N_19257,N_18975,N_18798);
xor U19258 (N_19258,N_18529,N_18725);
or U19259 (N_19259,N_18932,N_18622);
nor U19260 (N_19260,N_18836,N_18597);
xnor U19261 (N_19261,N_18904,N_18767);
and U19262 (N_19262,N_18595,N_18532);
or U19263 (N_19263,N_18765,N_18689);
and U19264 (N_19264,N_18901,N_18602);
or U19265 (N_19265,N_18545,N_18519);
nor U19266 (N_19266,N_18885,N_18541);
xor U19267 (N_19267,N_18975,N_18640);
or U19268 (N_19268,N_18859,N_18981);
or U19269 (N_19269,N_18850,N_18884);
nand U19270 (N_19270,N_18778,N_18725);
nand U19271 (N_19271,N_18691,N_18557);
nor U19272 (N_19272,N_18719,N_18805);
or U19273 (N_19273,N_18853,N_18670);
xor U19274 (N_19274,N_18831,N_18827);
xor U19275 (N_19275,N_18879,N_18674);
nor U19276 (N_19276,N_18780,N_18857);
nor U19277 (N_19277,N_18937,N_18901);
xnor U19278 (N_19278,N_18588,N_18626);
and U19279 (N_19279,N_18551,N_18969);
or U19280 (N_19280,N_18941,N_18989);
or U19281 (N_19281,N_18878,N_18912);
or U19282 (N_19282,N_18949,N_18922);
nor U19283 (N_19283,N_18952,N_18860);
nand U19284 (N_19284,N_18709,N_18571);
nor U19285 (N_19285,N_18845,N_18913);
xnor U19286 (N_19286,N_18947,N_18997);
and U19287 (N_19287,N_18662,N_18789);
and U19288 (N_19288,N_18534,N_18703);
nor U19289 (N_19289,N_18876,N_18933);
nand U19290 (N_19290,N_18523,N_18755);
or U19291 (N_19291,N_18506,N_18738);
nor U19292 (N_19292,N_18778,N_18667);
xnor U19293 (N_19293,N_18798,N_18567);
nand U19294 (N_19294,N_18969,N_18776);
xor U19295 (N_19295,N_18838,N_18752);
and U19296 (N_19296,N_18505,N_18832);
or U19297 (N_19297,N_18757,N_18582);
and U19298 (N_19298,N_18654,N_18879);
xor U19299 (N_19299,N_18813,N_18764);
xnor U19300 (N_19300,N_18621,N_18962);
nand U19301 (N_19301,N_18953,N_18535);
nand U19302 (N_19302,N_18675,N_18908);
or U19303 (N_19303,N_18951,N_18609);
or U19304 (N_19304,N_18550,N_18819);
nor U19305 (N_19305,N_18654,N_18931);
nand U19306 (N_19306,N_18793,N_18508);
nand U19307 (N_19307,N_18699,N_18507);
and U19308 (N_19308,N_18980,N_18724);
or U19309 (N_19309,N_18634,N_18991);
xor U19310 (N_19310,N_18578,N_18645);
nor U19311 (N_19311,N_18546,N_18613);
xnor U19312 (N_19312,N_18917,N_18842);
and U19313 (N_19313,N_18805,N_18541);
and U19314 (N_19314,N_18679,N_18566);
nor U19315 (N_19315,N_18663,N_18822);
and U19316 (N_19316,N_18693,N_18994);
nor U19317 (N_19317,N_18719,N_18705);
or U19318 (N_19318,N_18968,N_18811);
nand U19319 (N_19319,N_18940,N_18563);
nor U19320 (N_19320,N_18536,N_18564);
nand U19321 (N_19321,N_18806,N_18771);
xnor U19322 (N_19322,N_18971,N_18917);
or U19323 (N_19323,N_18899,N_18515);
or U19324 (N_19324,N_18560,N_18507);
xor U19325 (N_19325,N_18803,N_18805);
and U19326 (N_19326,N_18874,N_18884);
nand U19327 (N_19327,N_18532,N_18846);
nand U19328 (N_19328,N_18634,N_18917);
xor U19329 (N_19329,N_18573,N_18508);
nor U19330 (N_19330,N_18562,N_18553);
xnor U19331 (N_19331,N_18888,N_18571);
nor U19332 (N_19332,N_18718,N_18806);
nand U19333 (N_19333,N_18752,N_18902);
or U19334 (N_19334,N_18899,N_18590);
nand U19335 (N_19335,N_18565,N_18783);
nor U19336 (N_19336,N_18990,N_18719);
or U19337 (N_19337,N_18629,N_18568);
and U19338 (N_19338,N_18862,N_18528);
nor U19339 (N_19339,N_18894,N_18767);
xor U19340 (N_19340,N_18930,N_18827);
xor U19341 (N_19341,N_18759,N_18711);
nor U19342 (N_19342,N_18690,N_18702);
and U19343 (N_19343,N_18502,N_18623);
xnor U19344 (N_19344,N_18954,N_18553);
nand U19345 (N_19345,N_18943,N_18857);
xnor U19346 (N_19346,N_18949,N_18502);
nor U19347 (N_19347,N_18722,N_18932);
or U19348 (N_19348,N_18802,N_18572);
xor U19349 (N_19349,N_18832,N_18504);
nor U19350 (N_19350,N_18515,N_18807);
nand U19351 (N_19351,N_18529,N_18997);
nor U19352 (N_19352,N_18548,N_18576);
and U19353 (N_19353,N_18815,N_18609);
xnor U19354 (N_19354,N_18575,N_18842);
or U19355 (N_19355,N_18951,N_18996);
and U19356 (N_19356,N_18558,N_18744);
or U19357 (N_19357,N_18828,N_18705);
nand U19358 (N_19358,N_18848,N_18529);
nand U19359 (N_19359,N_18795,N_18882);
nand U19360 (N_19360,N_18522,N_18607);
or U19361 (N_19361,N_18613,N_18682);
or U19362 (N_19362,N_18728,N_18672);
nand U19363 (N_19363,N_18506,N_18502);
xor U19364 (N_19364,N_18999,N_18913);
and U19365 (N_19365,N_18567,N_18863);
xnor U19366 (N_19366,N_18706,N_18734);
or U19367 (N_19367,N_18726,N_18790);
nor U19368 (N_19368,N_18622,N_18756);
and U19369 (N_19369,N_18741,N_18835);
xor U19370 (N_19370,N_18597,N_18573);
nand U19371 (N_19371,N_18997,N_18989);
or U19372 (N_19372,N_18743,N_18944);
nor U19373 (N_19373,N_18986,N_18615);
xnor U19374 (N_19374,N_18792,N_18660);
xor U19375 (N_19375,N_18783,N_18714);
nand U19376 (N_19376,N_18935,N_18865);
nand U19377 (N_19377,N_18589,N_18833);
or U19378 (N_19378,N_18951,N_18979);
and U19379 (N_19379,N_18930,N_18853);
nand U19380 (N_19380,N_18774,N_18824);
xor U19381 (N_19381,N_18600,N_18518);
or U19382 (N_19382,N_18869,N_18904);
or U19383 (N_19383,N_18606,N_18651);
nand U19384 (N_19384,N_18876,N_18921);
xnor U19385 (N_19385,N_18798,N_18861);
nor U19386 (N_19386,N_18566,N_18620);
nor U19387 (N_19387,N_18637,N_18604);
or U19388 (N_19388,N_18620,N_18822);
nor U19389 (N_19389,N_18644,N_18737);
nand U19390 (N_19390,N_18667,N_18705);
xor U19391 (N_19391,N_18873,N_18785);
nor U19392 (N_19392,N_18938,N_18946);
and U19393 (N_19393,N_18915,N_18954);
nand U19394 (N_19394,N_18514,N_18575);
nand U19395 (N_19395,N_18914,N_18900);
or U19396 (N_19396,N_18694,N_18894);
and U19397 (N_19397,N_18602,N_18756);
xnor U19398 (N_19398,N_18940,N_18675);
and U19399 (N_19399,N_18700,N_18867);
nor U19400 (N_19400,N_18986,N_18913);
or U19401 (N_19401,N_18885,N_18795);
and U19402 (N_19402,N_18680,N_18675);
xnor U19403 (N_19403,N_18763,N_18823);
and U19404 (N_19404,N_18910,N_18605);
and U19405 (N_19405,N_18739,N_18843);
nand U19406 (N_19406,N_18807,N_18653);
and U19407 (N_19407,N_18638,N_18702);
xor U19408 (N_19408,N_18678,N_18959);
or U19409 (N_19409,N_18774,N_18873);
and U19410 (N_19410,N_18853,N_18675);
xnor U19411 (N_19411,N_18908,N_18508);
nand U19412 (N_19412,N_18564,N_18871);
xor U19413 (N_19413,N_18897,N_18743);
and U19414 (N_19414,N_18672,N_18569);
nand U19415 (N_19415,N_18844,N_18810);
xor U19416 (N_19416,N_18755,N_18792);
xnor U19417 (N_19417,N_18814,N_18693);
xnor U19418 (N_19418,N_18961,N_18671);
or U19419 (N_19419,N_18895,N_18626);
nand U19420 (N_19420,N_18510,N_18555);
or U19421 (N_19421,N_18545,N_18954);
nor U19422 (N_19422,N_18735,N_18536);
or U19423 (N_19423,N_18848,N_18844);
nand U19424 (N_19424,N_18849,N_18850);
xor U19425 (N_19425,N_18798,N_18754);
and U19426 (N_19426,N_18996,N_18911);
nor U19427 (N_19427,N_18843,N_18507);
or U19428 (N_19428,N_18769,N_18656);
and U19429 (N_19429,N_18553,N_18882);
xor U19430 (N_19430,N_18759,N_18726);
nand U19431 (N_19431,N_18624,N_18665);
xor U19432 (N_19432,N_18770,N_18528);
and U19433 (N_19433,N_18998,N_18641);
xnor U19434 (N_19434,N_18729,N_18837);
or U19435 (N_19435,N_18756,N_18941);
xnor U19436 (N_19436,N_18705,N_18607);
nand U19437 (N_19437,N_18801,N_18591);
nand U19438 (N_19438,N_18732,N_18713);
xnor U19439 (N_19439,N_18836,N_18512);
nor U19440 (N_19440,N_18914,N_18892);
nand U19441 (N_19441,N_18711,N_18835);
or U19442 (N_19442,N_18531,N_18677);
nor U19443 (N_19443,N_18929,N_18748);
xnor U19444 (N_19444,N_18798,N_18555);
xnor U19445 (N_19445,N_18954,N_18801);
or U19446 (N_19446,N_18752,N_18742);
nor U19447 (N_19447,N_18959,N_18722);
nand U19448 (N_19448,N_18883,N_18935);
and U19449 (N_19449,N_18769,N_18507);
nor U19450 (N_19450,N_18812,N_18793);
or U19451 (N_19451,N_18898,N_18605);
xnor U19452 (N_19452,N_18742,N_18642);
xor U19453 (N_19453,N_18886,N_18745);
and U19454 (N_19454,N_18821,N_18825);
and U19455 (N_19455,N_18846,N_18819);
nor U19456 (N_19456,N_18689,N_18503);
nor U19457 (N_19457,N_18747,N_18537);
xor U19458 (N_19458,N_18864,N_18696);
nand U19459 (N_19459,N_18642,N_18602);
and U19460 (N_19460,N_18950,N_18763);
nor U19461 (N_19461,N_18513,N_18525);
and U19462 (N_19462,N_18634,N_18890);
xor U19463 (N_19463,N_18980,N_18888);
or U19464 (N_19464,N_18780,N_18929);
nand U19465 (N_19465,N_18851,N_18812);
or U19466 (N_19466,N_18872,N_18898);
and U19467 (N_19467,N_18594,N_18724);
xnor U19468 (N_19468,N_18545,N_18814);
xor U19469 (N_19469,N_18884,N_18865);
nand U19470 (N_19470,N_18567,N_18945);
nor U19471 (N_19471,N_18737,N_18705);
and U19472 (N_19472,N_18682,N_18581);
or U19473 (N_19473,N_18760,N_18750);
xor U19474 (N_19474,N_18542,N_18669);
nor U19475 (N_19475,N_18553,N_18967);
nor U19476 (N_19476,N_18771,N_18707);
or U19477 (N_19477,N_18577,N_18769);
or U19478 (N_19478,N_18610,N_18830);
and U19479 (N_19479,N_18514,N_18807);
and U19480 (N_19480,N_18718,N_18898);
xnor U19481 (N_19481,N_18995,N_18559);
nand U19482 (N_19482,N_18828,N_18787);
and U19483 (N_19483,N_18684,N_18678);
xnor U19484 (N_19484,N_18840,N_18827);
or U19485 (N_19485,N_18866,N_18710);
nand U19486 (N_19486,N_18953,N_18759);
xnor U19487 (N_19487,N_18802,N_18840);
nor U19488 (N_19488,N_18656,N_18690);
xor U19489 (N_19489,N_18552,N_18866);
xor U19490 (N_19490,N_18646,N_18787);
nor U19491 (N_19491,N_18629,N_18640);
nor U19492 (N_19492,N_18612,N_18624);
or U19493 (N_19493,N_18733,N_18704);
xor U19494 (N_19494,N_18818,N_18573);
nand U19495 (N_19495,N_18593,N_18758);
nor U19496 (N_19496,N_18940,N_18736);
or U19497 (N_19497,N_18873,N_18545);
or U19498 (N_19498,N_18629,N_18545);
nand U19499 (N_19499,N_18981,N_18694);
and U19500 (N_19500,N_19225,N_19057);
xnor U19501 (N_19501,N_19453,N_19229);
or U19502 (N_19502,N_19422,N_19017);
and U19503 (N_19503,N_19353,N_19270);
nand U19504 (N_19504,N_19036,N_19288);
xnor U19505 (N_19505,N_19092,N_19321);
or U19506 (N_19506,N_19013,N_19255);
and U19507 (N_19507,N_19022,N_19393);
or U19508 (N_19508,N_19426,N_19074);
nor U19509 (N_19509,N_19146,N_19499);
xor U19510 (N_19510,N_19475,N_19459);
nor U19511 (N_19511,N_19480,N_19213);
nor U19512 (N_19512,N_19466,N_19169);
nand U19513 (N_19513,N_19091,N_19153);
nor U19514 (N_19514,N_19172,N_19341);
nand U19515 (N_19515,N_19399,N_19243);
xnor U19516 (N_19516,N_19355,N_19468);
nand U19517 (N_19517,N_19001,N_19107);
nand U19518 (N_19518,N_19100,N_19402);
or U19519 (N_19519,N_19285,N_19078);
nor U19520 (N_19520,N_19354,N_19224);
xor U19521 (N_19521,N_19377,N_19489);
or U19522 (N_19522,N_19164,N_19473);
nand U19523 (N_19523,N_19251,N_19240);
and U19524 (N_19524,N_19131,N_19405);
and U19525 (N_19525,N_19202,N_19315);
and U19526 (N_19526,N_19221,N_19051);
or U19527 (N_19527,N_19358,N_19147);
or U19528 (N_19528,N_19412,N_19299);
and U19529 (N_19529,N_19458,N_19332);
xnor U19530 (N_19530,N_19272,N_19083);
nand U19531 (N_19531,N_19351,N_19269);
and U19532 (N_19532,N_19309,N_19366);
or U19533 (N_19533,N_19382,N_19209);
nand U19534 (N_19534,N_19395,N_19201);
or U19535 (N_19535,N_19135,N_19231);
xnor U19536 (N_19536,N_19181,N_19049);
and U19537 (N_19537,N_19003,N_19494);
and U19538 (N_19538,N_19018,N_19449);
or U19539 (N_19539,N_19114,N_19227);
or U19540 (N_19540,N_19138,N_19342);
nor U19541 (N_19541,N_19418,N_19099);
and U19542 (N_19542,N_19215,N_19445);
nor U19543 (N_19543,N_19456,N_19126);
nand U19544 (N_19544,N_19308,N_19476);
or U19545 (N_19545,N_19190,N_19045);
and U19546 (N_19546,N_19248,N_19257);
or U19547 (N_19547,N_19180,N_19356);
or U19548 (N_19548,N_19261,N_19160);
or U19549 (N_19549,N_19496,N_19340);
and U19550 (N_19550,N_19154,N_19113);
or U19551 (N_19551,N_19441,N_19132);
nor U19552 (N_19552,N_19029,N_19439);
nand U19553 (N_19553,N_19168,N_19274);
xnor U19554 (N_19554,N_19219,N_19094);
nor U19555 (N_19555,N_19108,N_19266);
and U19556 (N_19556,N_19193,N_19088);
nor U19557 (N_19557,N_19007,N_19329);
and U19558 (N_19558,N_19203,N_19011);
or U19559 (N_19559,N_19484,N_19122);
nor U19560 (N_19560,N_19239,N_19296);
xnor U19561 (N_19561,N_19116,N_19322);
nor U19562 (N_19562,N_19333,N_19161);
nand U19563 (N_19563,N_19425,N_19157);
nand U19564 (N_19564,N_19348,N_19152);
or U19565 (N_19565,N_19046,N_19249);
or U19566 (N_19566,N_19256,N_19163);
and U19567 (N_19567,N_19442,N_19002);
nor U19568 (N_19568,N_19109,N_19428);
xor U19569 (N_19569,N_19452,N_19222);
nand U19570 (N_19570,N_19287,N_19121);
xnor U19571 (N_19571,N_19200,N_19063);
xor U19572 (N_19572,N_19303,N_19360);
or U19573 (N_19573,N_19214,N_19350);
nor U19574 (N_19574,N_19346,N_19433);
nor U19575 (N_19575,N_19183,N_19327);
xnor U19576 (N_19576,N_19103,N_19192);
or U19577 (N_19577,N_19175,N_19241);
xnor U19578 (N_19578,N_19483,N_19205);
nor U19579 (N_19579,N_19236,N_19349);
and U19580 (N_19580,N_19331,N_19050);
nand U19581 (N_19581,N_19386,N_19444);
xor U19582 (N_19582,N_19117,N_19362);
nor U19583 (N_19583,N_19254,N_19268);
nor U19584 (N_19584,N_19158,N_19167);
and U19585 (N_19585,N_19408,N_19486);
nand U19586 (N_19586,N_19010,N_19325);
xor U19587 (N_19587,N_19019,N_19199);
nor U19588 (N_19588,N_19477,N_19493);
or U19589 (N_19589,N_19195,N_19301);
nor U19590 (N_19590,N_19230,N_19436);
or U19591 (N_19591,N_19028,N_19435);
xor U19592 (N_19592,N_19216,N_19223);
nand U19593 (N_19593,N_19075,N_19335);
nor U19594 (N_19594,N_19027,N_19279);
or U19595 (N_19595,N_19352,N_19281);
or U19596 (N_19596,N_19463,N_19087);
nor U19597 (N_19597,N_19238,N_19413);
nor U19598 (N_19598,N_19271,N_19253);
and U19599 (N_19599,N_19390,N_19283);
or U19600 (N_19600,N_19485,N_19062);
and U19601 (N_19601,N_19015,N_19080);
nor U19602 (N_19602,N_19137,N_19110);
and U19603 (N_19603,N_19392,N_19026);
nor U19604 (N_19604,N_19089,N_19316);
nand U19605 (N_19605,N_19159,N_19124);
and U19606 (N_19606,N_19457,N_19318);
nand U19607 (N_19607,N_19372,N_19339);
nand U19608 (N_19608,N_19313,N_19375);
nand U19609 (N_19609,N_19077,N_19252);
or U19610 (N_19610,N_19284,N_19136);
and U19611 (N_19611,N_19166,N_19120);
and U19612 (N_19612,N_19307,N_19076);
xnor U19613 (N_19613,N_19064,N_19326);
nor U19614 (N_19614,N_19416,N_19177);
and U19615 (N_19615,N_19176,N_19041);
or U19616 (N_19616,N_19280,N_19492);
xor U19617 (N_19617,N_19361,N_19380);
nor U19618 (N_19618,N_19053,N_19328);
nand U19619 (N_19619,N_19278,N_19423);
or U19620 (N_19620,N_19171,N_19095);
or U19621 (N_19621,N_19208,N_19141);
and U19622 (N_19622,N_19298,N_19446);
nand U19623 (N_19623,N_19211,N_19042);
and U19624 (N_19624,N_19204,N_19273);
or U19625 (N_19625,N_19143,N_19388);
xor U19626 (N_19626,N_19367,N_19292);
xnor U19627 (N_19627,N_19082,N_19432);
and U19628 (N_19628,N_19337,N_19440);
xor U19629 (N_19629,N_19242,N_19497);
nor U19630 (N_19630,N_19282,N_19391);
or U19631 (N_19631,N_19093,N_19330);
or U19632 (N_19632,N_19039,N_19052);
nand U19633 (N_19633,N_19237,N_19396);
xor U19634 (N_19634,N_19068,N_19260);
nand U19635 (N_19635,N_19474,N_19244);
or U19636 (N_19636,N_19005,N_19374);
nor U19637 (N_19637,N_19004,N_19058);
or U19638 (N_19638,N_19196,N_19071);
or U19639 (N_19639,N_19482,N_19250);
nand U19640 (N_19640,N_19012,N_19479);
and U19641 (N_19641,N_19411,N_19319);
xnor U19642 (N_19642,N_19155,N_19228);
or U19643 (N_19643,N_19338,N_19376);
and U19644 (N_19644,N_19305,N_19185);
or U19645 (N_19645,N_19090,N_19119);
xnor U19646 (N_19646,N_19206,N_19182);
nand U19647 (N_19647,N_19455,N_19410);
nand U19648 (N_19648,N_19369,N_19096);
nand U19649 (N_19649,N_19234,N_19320);
and U19650 (N_19650,N_19291,N_19210);
nor U19651 (N_19651,N_19079,N_19072);
or U19652 (N_19652,N_19306,N_19020);
xor U19653 (N_19653,N_19347,N_19031);
nand U19654 (N_19654,N_19067,N_19462);
xor U19655 (N_19655,N_19295,N_19060);
nand U19656 (N_19656,N_19344,N_19187);
nor U19657 (N_19657,N_19478,N_19165);
nand U19658 (N_19658,N_19400,N_19371);
nand U19659 (N_19659,N_19490,N_19098);
nand U19660 (N_19660,N_19194,N_19140);
and U19661 (N_19661,N_19085,N_19414);
or U19662 (N_19662,N_19421,N_19084);
xor U19663 (N_19663,N_19434,N_19104);
nor U19664 (N_19664,N_19448,N_19186);
nand U19665 (N_19665,N_19389,N_19289);
or U19666 (N_19666,N_19430,N_19401);
nor U19667 (N_19667,N_19145,N_19179);
and U19668 (N_19668,N_19102,N_19324);
and U19669 (N_19669,N_19112,N_19404);
and U19670 (N_19670,N_19451,N_19118);
nand U19671 (N_19671,N_19212,N_19286);
and U19672 (N_19672,N_19304,N_19431);
nand U19673 (N_19673,N_19226,N_19334);
nor U19674 (N_19674,N_19394,N_19014);
xor U19675 (N_19675,N_19429,N_19105);
xor U19676 (N_19676,N_19488,N_19024);
nor U19677 (N_19677,N_19357,N_19220);
and U19678 (N_19678,N_19443,N_19297);
nand U19679 (N_19679,N_19368,N_19148);
nand U19680 (N_19680,N_19454,N_19021);
xor U19681 (N_19681,N_19232,N_19398);
and U19682 (N_19682,N_19464,N_19471);
nand U19683 (N_19683,N_19125,N_19427);
nand U19684 (N_19684,N_19262,N_19323);
nand U19685 (N_19685,N_19035,N_19008);
nand U19686 (N_19686,N_19056,N_19016);
and U19687 (N_19687,N_19073,N_19000);
xnor U19688 (N_19688,N_19363,N_19047);
nand U19689 (N_19689,N_19336,N_19415);
xor U19690 (N_19690,N_19263,N_19406);
or U19691 (N_19691,N_19198,N_19037);
or U19692 (N_19692,N_19156,N_19419);
and U19693 (N_19693,N_19397,N_19450);
and U19694 (N_19694,N_19173,N_19066);
or U19695 (N_19695,N_19150,N_19188);
and U19696 (N_19696,N_19461,N_19207);
or U19697 (N_19697,N_19481,N_19030);
or U19698 (N_19698,N_19314,N_19302);
and U19699 (N_19699,N_19417,N_19048);
or U19700 (N_19700,N_19069,N_19300);
and U19701 (N_19701,N_19364,N_19123);
nand U19702 (N_19702,N_19424,N_19277);
or U19703 (N_19703,N_19055,N_19365);
nand U19704 (N_19704,N_19312,N_19217);
nor U19705 (N_19705,N_19467,N_19469);
nor U19706 (N_19706,N_19460,N_19189);
nor U19707 (N_19707,N_19106,N_19127);
and U19708 (N_19708,N_19139,N_19097);
nor U19709 (N_19709,N_19383,N_19040);
nand U19710 (N_19710,N_19311,N_19149);
xor U19711 (N_19711,N_19465,N_19407);
nor U19712 (N_19712,N_19134,N_19033);
nor U19713 (N_19713,N_19130,N_19409);
or U19714 (N_19714,N_19174,N_19142);
nor U19715 (N_19715,N_19420,N_19385);
nand U19716 (N_19716,N_19317,N_19265);
and U19717 (N_19717,N_19370,N_19290);
nor U19718 (N_19718,N_19059,N_19191);
xnor U19719 (N_19719,N_19129,N_19043);
xnor U19720 (N_19720,N_19447,N_19259);
and U19721 (N_19721,N_19294,N_19111);
xnor U19722 (N_19722,N_19378,N_19498);
nand U19723 (N_19723,N_19006,N_19403);
nand U19724 (N_19724,N_19023,N_19144);
and U19725 (N_19725,N_19235,N_19054);
or U19726 (N_19726,N_19065,N_19310);
or U19727 (N_19727,N_19379,N_19267);
nand U19728 (N_19728,N_19151,N_19081);
and U19729 (N_19729,N_19491,N_19009);
or U19730 (N_19730,N_19246,N_19101);
nor U19731 (N_19731,N_19128,N_19133);
nand U19732 (N_19732,N_19343,N_19472);
or U19733 (N_19733,N_19373,N_19264);
nor U19734 (N_19734,N_19359,N_19197);
xnor U19735 (N_19735,N_19293,N_19470);
or U19736 (N_19736,N_19245,N_19070);
or U19737 (N_19737,N_19495,N_19275);
xor U19738 (N_19738,N_19086,N_19115);
nand U19739 (N_19739,N_19170,N_19034);
or U19740 (N_19740,N_19061,N_19162);
nor U19741 (N_19741,N_19438,N_19218);
nand U19742 (N_19742,N_19276,N_19437);
nor U19743 (N_19743,N_19233,N_19258);
xnor U19744 (N_19744,N_19384,N_19387);
nor U19745 (N_19745,N_19032,N_19038);
and U19746 (N_19746,N_19345,N_19178);
or U19747 (N_19747,N_19025,N_19381);
xor U19748 (N_19748,N_19184,N_19044);
xor U19749 (N_19749,N_19487,N_19247);
nand U19750 (N_19750,N_19118,N_19458);
or U19751 (N_19751,N_19107,N_19028);
or U19752 (N_19752,N_19135,N_19352);
nor U19753 (N_19753,N_19287,N_19259);
nor U19754 (N_19754,N_19282,N_19073);
nand U19755 (N_19755,N_19155,N_19070);
nor U19756 (N_19756,N_19445,N_19236);
xor U19757 (N_19757,N_19464,N_19215);
nand U19758 (N_19758,N_19445,N_19454);
nand U19759 (N_19759,N_19386,N_19482);
or U19760 (N_19760,N_19250,N_19338);
and U19761 (N_19761,N_19266,N_19457);
or U19762 (N_19762,N_19415,N_19352);
nor U19763 (N_19763,N_19352,N_19137);
xnor U19764 (N_19764,N_19226,N_19118);
or U19765 (N_19765,N_19413,N_19217);
nand U19766 (N_19766,N_19189,N_19478);
xor U19767 (N_19767,N_19370,N_19339);
nor U19768 (N_19768,N_19010,N_19450);
xor U19769 (N_19769,N_19368,N_19224);
or U19770 (N_19770,N_19490,N_19014);
and U19771 (N_19771,N_19012,N_19188);
or U19772 (N_19772,N_19268,N_19059);
xnor U19773 (N_19773,N_19253,N_19097);
nor U19774 (N_19774,N_19110,N_19341);
xnor U19775 (N_19775,N_19407,N_19295);
and U19776 (N_19776,N_19260,N_19025);
xnor U19777 (N_19777,N_19481,N_19210);
and U19778 (N_19778,N_19482,N_19426);
nor U19779 (N_19779,N_19048,N_19006);
xnor U19780 (N_19780,N_19342,N_19277);
nor U19781 (N_19781,N_19150,N_19402);
nand U19782 (N_19782,N_19113,N_19283);
nor U19783 (N_19783,N_19216,N_19008);
nor U19784 (N_19784,N_19016,N_19245);
xnor U19785 (N_19785,N_19084,N_19268);
or U19786 (N_19786,N_19146,N_19484);
and U19787 (N_19787,N_19436,N_19330);
and U19788 (N_19788,N_19265,N_19475);
or U19789 (N_19789,N_19027,N_19193);
xor U19790 (N_19790,N_19051,N_19123);
nand U19791 (N_19791,N_19188,N_19144);
or U19792 (N_19792,N_19255,N_19070);
xnor U19793 (N_19793,N_19301,N_19061);
nand U19794 (N_19794,N_19421,N_19438);
nand U19795 (N_19795,N_19198,N_19498);
and U19796 (N_19796,N_19276,N_19396);
nor U19797 (N_19797,N_19403,N_19313);
or U19798 (N_19798,N_19065,N_19499);
or U19799 (N_19799,N_19055,N_19312);
nand U19800 (N_19800,N_19188,N_19083);
nor U19801 (N_19801,N_19180,N_19488);
or U19802 (N_19802,N_19398,N_19291);
xnor U19803 (N_19803,N_19375,N_19130);
xor U19804 (N_19804,N_19058,N_19235);
or U19805 (N_19805,N_19209,N_19430);
and U19806 (N_19806,N_19162,N_19428);
and U19807 (N_19807,N_19497,N_19156);
xor U19808 (N_19808,N_19224,N_19428);
and U19809 (N_19809,N_19474,N_19415);
nor U19810 (N_19810,N_19400,N_19383);
nor U19811 (N_19811,N_19240,N_19156);
nor U19812 (N_19812,N_19063,N_19035);
nand U19813 (N_19813,N_19348,N_19115);
and U19814 (N_19814,N_19378,N_19240);
xnor U19815 (N_19815,N_19071,N_19427);
nor U19816 (N_19816,N_19047,N_19091);
xor U19817 (N_19817,N_19390,N_19327);
or U19818 (N_19818,N_19098,N_19152);
xor U19819 (N_19819,N_19061,N_19241);
nor U19820 (N_19820,N_19049,N_19426);
xnor U19821 (N_19821,N_19022,N_19435);
nand U19822 (N_19822,N_19181,N_19153);
or U19823 (N_19823,N_19124,N_19066);
nand U19824 (N_19824,N_19085,N_19399);
nand U19825 (N_19825,N_19145,N_19366);
nor U19826 (N_19826,N_19172,N_19256);
or U19827 (N_19827,N_19069,N_19484);
nand U19828 (N_19828,N_19471,N_19212);
nor U19829 (N_19829,N_19327,N_19060);
or U19830 (N_19830,N_19394,N_19375);
xnor U19831 (N_19831,N_19012,N_19306);
nand U19832 (N_19832,N_19478,N_19155);
or U19833 (N_19833,N_19370,N_19029);
nor U19834 (N_19834,N_19327,N_19230);
and U19835 (N_19835,N_19357,N_19133);
and U19836 (N_19836,N_19456,N_19039);
nand U19837 (N_19837,N_19241,N_19433);
xnor U19838 (N_19838,N_19264,N_19086);
nand U19839 (N_19839,N_19122,N_19120);
nand U19840 (N_19840,N_19151,N_19304);
xnor U19841 (N_19841,N_19089,N_19193);
or U19842 (N_19842,N_19490,N_19042);
nand U19843 (N_19843,N_19233,N_19207);
nor U19844 (N_19844,N_19019,N_19141);
or U19845 (N_19845,N_19466,N_19275);
or U19846 (N_19846,N_19029,N_19234);
or U19847 (N_19847,N_19438,N_19411);
nor U19848 (N_19848,N_19337,N_19400);
xor U19849 (N_19849,N_19157,N_19470);
nor U19850 (N_19850,N_19269,N_19477);
and U19851 (N_19851,N_19377,N_19062);
or U19852 (N_19852,N_19423,N_19265);
or U19853 (N_19853,N_19197,N_19345);
and U19854 (N_19854,N_19226,N_19459);
and U19855 (N_19855,N_19294,N_19194);
or U19856 (N_19856,N_19137,N_19115);
nand U19857 (N_19857,N_19449,N_19314);
nor U19858 (N_19858,N_19224,N_19497);
and U19859 (N_19859,N_19423,N_19460);
nor U19860 (N_19860,N_19199,N_19363);
nand U19861 (N_19861,N_19234,N_19190);
and U19862 (N_19862,N_19275,N_19452);
nand U19863 (N_19863,N_19341,N_19332);
or U19864 (N_19864,N_19243,N_19482);
nand U19865 (N_19865,N_19352,N_19410);
and U19866 (N_19866,N_19248,N_19486);
nor U19867 (N_19867,N_19276,N_19315);
xnor U19868 (N_19868,N_19333,N_19231);
and U19869 (N_19869,N_19056,N_19367);
or U19870 (N_19870,N_19189,N_19070);
and U19871 (N_19871,N_19015,N_19344);
xor U19872 (N_19872,N_19021,N_19053);
and U19873 (N_19873,N_19265,N_19236);
and U19874 (N_19874,N_19301,N_19259);
xnor U19875 (N_19875,N_19300,N_19472);
nor U19876 (N_19876,N_19079,N_19296);
and U19877 (N_19877,N_19426,N_19449);
nor U19878 (N_19878,N_19321,N_19449);
xnor U19879 (N_19879,N_19028,N_19282);
xnor U19880 (N_19880,N_19201,N_19369);
nor U19881 (N_19881,N_19125,N_19039);
xnor U19882 (N_19882,N_19065,N_19466);
xor U19883 (N_19883,N_19308,N_19047);
xor U19884 (N_19884,N_19237,N_19408);
nor U19885 (N_19885,N_19408,N_19293);
or U19886 (N_19886,N_19385,N_19459);
xnor U19887 (N_19887,N_19110,N_19446);
or U19888 (N_19888,N_19364,N_19212);
or U19889 (N_19889,N_19464,N_19129);
xnor U19890 (N_19890,N_19491,N_19136);
and U19891 (N_19891,N_19353,N_19272);
nor U19892 (N_19892,N_19334,N_19034);
nand U19893 (N_19893,N_19301,N_19043);
nor U19894 (N_19894,N_19213,N_19065);
and U19895 (N_19895,N_19428,N_19081);
nand U19896 (N_19896,N_19373,N_19299);
nand U19897 (N_19897,N_19298,N_19118);
or U19898 (N_19898,N_19475,N_19410);
nand U19899 (N_19899,N_19119,N_19497);
xor U19900 (N_19900,N_19286,N_19295);
nor U19901 (N_19901,N_19348,N_19430);
nor U19902 (N_19902,N_19271,N_19391);
and U19903 (N_19903,N_19325,N_19253);
or U19904 (N_19904,N_19093,N_19225);
and U19905 (N_19905,N_19389,N_19284);
nand U19906 (N_19906,N_19207,N_19379);
and U19907 (N_19907,N_19226,N_19120);
nand U19908 (N_19908,N_19053,N_19285);
or U19909 (N_19909,N_19014,N_19202);
and U19910 (N_19910,N_19155,N_19305);
and U19911 (N_19911,N_19149,N_19225);
xnor U19912 (N_19912,N_19020,N_19113);
nand U19913 (N_19913,N_19266,N_19171);
nand U19914 (N_19914,N_19331,N_19044);
nand U19915 (N_19915,N_19180,N_19449);
and U19916 (N_19916,N_19015,N_19021);
nand U19917 (N_19917,N_19019,N_19294);
xor U19918 (N_19918,N_19111,N_19407);
nor U19919 (N_19919,N_19326,N_19169);
nand U19920 (N_19920,N_19374,N_19154);
or U19921 (N_19921,N_19071,N_19209);
and U19922 (N_19922,N_19329,N_19367);
nor U19923 (N_19923,N_19040,N_19401);
nor U19924 (N_19924,N_19476,N_19281);
nand U19925 (N_19925,N_19416,N_19288);
nand U19926 (N_19926,N_19160,N_19224);
xnor U19927 (N_19927,N_19155,N_19338);
or U19928 (N_19928,N_19120,N_19220);
nand U19929 (N_19929,N_19143,N_19363);
xnor U19930 (N_19930,N_19005,N_19254);
nor U19931 (N_19931,N_19358,N_19418);
xor U19932 (N_19932,N_19115,N_19180);
or U19933 (N_19933,N_19411,N_19353);
nand U19934 (N_19934,N_19090,N_19483);
xnor U19935 (N_19935,N_19470,N_19388);
nand U19936 (N_19936,N_19485,N_19349);
nand U19937 (N_19937,N_19236,N_19234);
or U19938 (N_19938,N_19135,N_19396);
nor U19939 (N_19939,N_19475,N_19078);
xnor U19940 (N_19940,N_19033,N_19152);
or U19941 (N_19941,N_19277,N_19087);
xnor U19942 (N_19942,N_19144,N_19438);
nor U19943 (N_19943,N_19211,N_19062);
xnor U19944 (N_19944,N_19101,N_19167);
and U19945 (N_19945,N_19293,N_19248);
xnor U19946 (N_19946,N_19057,N_19415);
xnor U19947 (N_19947,N_19213,N_19047);
nor U19948 (N_19948,N_19422,N_19291);
or U19949 (N_19949,N_19179,N_19441);
or U19950 (N_19950,N_19210,N_19339);
nand U19951 (N_19951,N_19120,N_19420);
and U19952 (N_19952,N_19196,N_19029);
and U19953 (N_19953,N_19110,N_19074);
or U19954 (N_19954,N_19077,N_19216);
or U19955 (N_19955,N_19381,N_19464);
or U19956 (N_19956,N_19326,N_19032);
xnor U19957 (N_19957,N_19027,N_19493);
nand U19958 (N_19958,N_19028,N_19391);
nor U19959 (N_19959,N_19227,N_19242);
xnor U19960 (N_19960,N_19112,N_19030);
nand U19961 (N_19961,N_19377,N_19234);
or U19962 (N_19962,N_19277,N_19183);
nand U19963 (N_19963,N_19214,N_19411);
nand U19964 (N_19964,N_19275,N_19317);
or U19965 (N_19965,N_19166,N_19036);
and U19966 (N_19966,N_19015,N_19153);
and U19967 (N_19967,N_19443,N_19072);
and U19968 (N_19968,N_19354,N_19443);
nor U19969 (N_19969,N_19357,N_19014);
nor U19970 (N_19970,N_19390,N_19187);
nand U19971 (N_19971,N_19183,N_19374);
nand U19972 (N_19972,N_19412,N_19417);
xor U19973 (N_19973,N_19376,N_19246);
xnor U19974 (N_19974,N_19296,N_19058);
nand U19975 (N_19975,N_19094,N_19443);
or U19976 (N_19976,N_19132,N_19317);
nand U19977 (N_19977,N_19486,N_19351);
xnor U19978 (N_19978,N_19347,N_19123);
nor U19979 (N_19979,N_19069,N_19098);
nor U19980 (N_19980,N_19467,N_19160);
nor U19981 (N_19981,N_19183,N_19176);
nand U19982 (N_19982,N_19444,N_19490);
or U19983 (N_19983,N_19290,N_19255);
nand U19984 (N_19984,N_19168,N_19313);
and U19985 (N_19985,N_19287,N_19234);
nor U19986 (N_19986,N_19364,N_19221);
nor U19987 (N_19987,N_19450,N_19234);
and U19988 (N_19988,N_19335,N_19127);
or U19989 (N_19989,N_19493,N_19214);
xor U19990 (N_19990,N_19004,N_19064);
xnor U19991 (N_19991,N_19474,N_19419);
or U19992 (N_19992,N_19025,N_19394);
and U19993 (N_19993,N_19298,N_19432);
nand U19994 (N_19994,N_19375,N_19498);
nand U19995 (N_19995,N_19197,N_19198);
or U19996 (N_19996,N_19207,N_19467);
and U19997 (N_19997,N_19428,N_19078);
xnor U19998 (N_19998,N_19487,N_19428);
nand U19999 (N_19999,N_19466,N_19374);
nand UO_0 (O_0,N_19581,N_19865);
nor UO_1 (O_1,N_19744,N_19869);
nor UO_2 (O_2,N_19755,N_19781);
nor UO_3 (O_3,N_19709,N_19974);
nand UO_4 (O_4,N_19962,N_19702);
xor UO_5 (O_5,N_19897,N_19515);
and UO_6 (O_6,N_19589,N_19893);
or UO_7 (O_7,N_19970,N_19820);
and UO_8 (O_8,N_19513,N_19576);
and UO_9 (O_9,N_19705,N_19605);
nand UO_10 (O_10,N_19787,N_19566);
xnor UO_11 (O_11,N_19795,N_19935);
nor UO_12 (O_12,N_19915,N_19527);
nor UO_13 (O_13,N_19634,N_19908);
nand UO_14 (O_14,N_19983,N_19907);
nor UO_15 (O_15,N_19741,N_19789);
or UO_16 (O_16,N_19839,N_19534);
xnor UO_17 (O_17,N_19667,N_19827);
or UO_18 (O_18,N_19572,N_19958);
or UO_19 (O_19,N_19780,N_19875);
nor UO_20 (O_20,N_19852,N_19922);
and UO_21 (O_21,N_19841,N_19764);
nand UO_22 (O_22,N_19995,N_19866);
or UO_23 (O_23,N_19773,N_19782);
and UO_24 (O_24,N_19607,N_19919);
xnor UO_25 (O_25,N_19683,N_19536);
nor UO_26 (O_26,N_19956,N_19925);
nor UO_27 (O_27,N_19959,N_19554);
nor UO_28 (O_28,N_19552,N_19834);
xnor UO_29 (O_29,N_19950,N_19597);
nor UO_30 (O_30,N_19511,N_19853);
nor UO_31 (O_31,N_19717,N_19633);
nor UO_32 (O_32,N_19650,N_19553);
and UO_33 (O_33,N_19836,N_19507);
nor UO_34 (O_34,N_19750,N_19547);
and UO_35 (O_35,N_19766,N_19500);
or UO_36 (O_36,N_19942,N_19646);
xor UO_37 (O_37,N_19863,N_19535);
xnor UO_38 (O_38,N_19752,N_19695);
and UO_39 (O_39,N_19994,N_19842);
and UO_40 (O_40,N_19881,N_19867);
or UO_41 (O_41,N_19829,N_19545);
and UO_42 (O_42,N_19960,N_19616);
and UO_43 (O_43,N_19517,N_19903);
or UO_44 (O_44,N_19565,N_19564);
and UO_45 (O_45,N_19664,N_19877);
nor UO_46 (O_46,N_19886,N_19639);
and UO_47 (O_47,N_19889,N_19505);
nand UO_48 (O_48,N_19859,N_19518);
or UO_49 (O_49,N_19590,N_19767);
nand UO_50 (O_50,N_19934,N_19632);
nand UO_51 (O_51,N_19931,N_19508);
nand UO_52 (O_52,N_19519,N_19620);
nor UO_53 (O_53,N_19832,N_19879);
nand UO_54 (O_54,N_19777,N_19693);
nand UO_55 (O_55,N_19573,N_19596);
nand UO_56 (O_56,N_19567,N_19996);
xor UO_57 (O_57,N_19626,N_19591);
nand UO_58 (O_58,N_19860,N_19643);
nor UO_59 (O_59,N_19808,N_19711);
or UO_60 (O_60,N_19902,N_19801);
and UO_61 (O_61,N_19851,N_19720);
xor UO_62 (O_62,N_19965,N_19858);
nand UO_63 (O_63,N_19814,N_19817);
xnor UO_64 (O_64,N_19844,N_19622);
and UO_65 (O_65,N_19558,N_19964);
or UO_66 (O_66,N_19769,N_19855);
nor UO_67 (O_67,N_19598,N_19668);
and UO_68 (O_68,N_19543,N_19551);
nor UO_69 (O_69,N_19873,N_19775);
and UO_70 (O_70,N_19642,N_19503);
nor UO_71 (O_71,N_19763,N_19798);
xor UO_72 (O_72,N_19726,N_19888);
nor UO_73 (O_73,N_19712,N_19715);
nand UO_74 (O_74,N_19918,N_19625);
nor UO_75 (O_75,N_19945,N_19611);
xor UO_76 (O_76,N_19772,N_19629);
nand UO_77 (O_77,N_19927,N_19880);
xnor UO_78 (O_78,N_19791,N_19825);
nor UO_79 (O_79,N_19612,N_19778);
nor UO_80 (O_80,N_19774,N_19585);
and UO_81 (O_81,N_19949,N_19924);
and UO_82 (O_82,N_19848,N_19883);
or UO_83 (O_83,N_19753,N_19928);
or UO_84 (O_84,N_19525,N_19864);
xnor UO_85 (O_85,N_19516,N_19861);
or UO_86 (O_86,N_19916,N_19697);
or UO_87 (O_87,N_19509,N_19656);
and UO_88 (O_88,N_19735,N_19993);
or UO_89 (O_89,N_19833,N_19532);
or UO_90 (O_90,N_19951,N_19710);
xor UO_91 (O_91,N_19940,N_19846);
nor UO_92 (O_92,N_19665,N_19676);
xor UO_93 (O_93,N_19840,N_19784);
and UO_94 (O_94,N_19677,N_19701);
nor UO_95 (O_95,N_19990,N_19972);
or UO_96 (O_96,N_19723,N_19672);
and UO_97 (O_97,N_19561,N_19910);
and UO_98 (O_98,N_19706,N_19816);
and UO_99 (O_99,N_19673,N_19955);
nand UO_100 (O_100,N_19805,N_19930);
xor UO_101 (O_101,N_19725,N_19783);
and UO_102 (O_102,N_19968,N_19681);
or UO_103 (O_103,N_19608,N_19638);
nor UO_104 (O_104,N_19765,N_19937);
nand UO_105 (O_105,N_19943,N_19628);
and UO_106 (O_106,N_19898,N_19884);
nand UO_107 (O_107,N_19613,N_19653);
or UO_108 (O_108,N_19975,N_19533);
or UO_109 (O_109,N_19670,N_19980);
and UO_110 (O_110,N_19617,N_19663);
or UO_111 (O_111,N_19577,N_19818);
and UO_112 (O_112,N_19920,N_19809);
or UO_113 (O_113,N_19894,N_19522);
nand UO_114 (O_114,N_19731,N_19952);
and UO_115 (O_115,N_19571,N_19792);
nor UO_116 (O_116,N_19745,N_19954);
and UO_117 (O_117,N_19530,N_19679);
or UO_118 (O_118,N_19555,N_19810);
or UO_119 (O_119,N_19542,N_19714);
and UO_120 (O_120,N_19648,N_19803);
or UO_121 (O_121,N_19953,N_19799);
nand UO_122 (O_122,N_19982,N_19904);
xor UO_123 (O_123,N_19570,N_19574);
nand UO_124 (O_124,N_19872,N_19892);
nor UO_125 (O_125,N_19636,N_19826);
nand UO_126 (O_126,N_19979,N_19538);
or UO_127 (O_127,N_19973,N_19713);
or UO_128 (O_128,N_19797,N_19662);
xor UO_129 (O_129,N_19747,N_19946);
nand UO_130 (O_130,N_19978,N_19874);
or UO_131 (O_131,N_19926,N_19847);
xor UO_132 (O_132,N_19793,N_19976);
nor UO_133 (O_133,N_19691,N_19637);
nor UO_134 (O_134,N_19856,N_19708);
xor UO_135 (O_135,N_19660,N_19757);
nor UO_136 (O_136,N_19966,N_19680);
xnor UO_137 (O_137,N_19728,N_19540);
nand UO_138 (O_138,N_19619,N_19746);
or UO_139 (O_139,N_19690,N_19929);
nor UO_140 (O_140,N_19644,N_19748);
nand UO_141 (O_141,N_19546,N_19692);
nor UO_142 (O_142,N_19580,N_19578);
or UO_143 (O_143,N_19843,N_19901);
or UO_144 (O_144,N_19716,N_19602);
or UO_145 (O_145,N_19583,N_19742);
or UO_146 (O_146,N_19603,N_19604);
nor UO_147 (O_147,N_19609,N_19528);
nand UO_148 (O_148,N_19804,N_19624);
or UO_149 (O_149,N_19963,N_19790);
nor UO_150 (O_150,N_19722,N_19941);
nand UO_151 (O_151,N_19649,N_19734);
nor UO_152 (O_152,N_19600,N_19579);
nor UO_153 (O_153,N_19736,N_19694);
or UO_154 (O_154,N_19621,N_19759);
xor UO_155 (O_155,N_19770,N_19686);
nand UO_156 (O_156,N_19627,N_19685);
or UO_157 (O_157,N_19807,N_19917);
nor UO_158 (O_158,N_19896,N_19521);
nor UO_159 (O_159,N_19586,N_19997);
nand UO_160 (O_160,N_19991,N_19595);
xnor UO_161 (O_161,N_19761,N_19560);
nand UO_162 (O_162,N_19938,N_19549);
xnor UO_163 (O_163,N_19785,N_19615);
nand UO_164 (O_164,N_19849,N_19986);
nor UO_165 (O_165,N_19699,N_19882);
or UO_166 (O_166,N_19614,N_19788);
or UO_167 (O_167,N_19501,N_19806);
or UO_168 (O_168,N_19760,N_19878);
xor UO_169 (O_169,N_19811,N_19909);
xor UO_170 (O_170,N_19651,N_19640);
nand UO_171 (O_171,N_19923,N_19838);
nand UO_172 (O_172,N_19905,N_19599);
nand UO_173 (O_173,N_19740,N_19559);
or UO_174 (O_174,N_19666,N_19831);
nor UO_175 (O_175,N_19727,N_19835);
xnor UO_176 (O_176,N_19999,N_19821);
xnor UO_177 (O_177,N_19671,N_19661);
or UO_178 (O_178,N_19845,N_19912);
nor UO_179 (O_179,N_19900,N_19623);
and UO_180 (O_180,N_19678,N_19730);
nor UO_181 (O_181,N_19824,N_19606);
and UO_182 (O_182,N_19647,N_19768);
nand UO_183 (O_183,N_19718,N_19704);
xnor UO_184 (O_184,N_19652,N_19721);
xor UO_185 (O_185,N_19895,N_19890);
nand UO_186 (O_186,N_19674,N_19779);
and UO_187 (O_187,N_19911,N_19751);
or UO_188 (O_188,N_19887,N_19645);
nand UO_189 (O_189,N_19936,N_19684);
nand UO_190 (O_190,N_19985,N_19584);
and UO_191 (O_191,N_19815,N_19977);
or UO_192 (O_192,N_19512,N_19635);
xor UO_193 (O_193,N_19868,N_19987);
xnor UO_194 (O_194,N_19871,N_19506);
nand UO_195 (O_195,N_19669,N_19756);
xor UO_196 (O_196,N_19594,N_19906);
and UO_197 (O_197,N_19967,N_19689);
nand UO_198 (O_198,N_19531,N_19822);
or UO_199 (O_199,N_19688,N_19526);
nand UO_200 (O_200,N_19569,N_19575);
nor UO_201 (O_201,N_19556,N_19700);
or UO_202 (O_202,N_19998,N_19758);
and UO_203 (O_203,N_19539,N_19588);
or UO_204 (O_204,N_19502,N_19630);
or UO_205 (O_205,N_19969,N_19794);
or UO_206 (O_206,N_19984,N_19830);
nand UO_207 (O_207,N_19593,N_19550);
or UO_208 (O_208,N_19891,N_19682);
xnor UO_209 (O_209,N_19504,N_19514);
xor UO_210 (O_210,N_19557,N_19796);
nand UO_211 (O_211,N_19957,N_19738);
or UO_212 (O_212,N_19631,N_19562);
and UO_213 (O_213,N_19582,N_19563);
or UO_214 (O_214,N_19944,N_19762);
xor UO_215 (O_215,N_19641,N_19544);
nor UO_216 (O_216,N_19655,N_19659);
nor UO_217 (O_217,N_19548,N_19698);
nor UO_218 (O_218,N_19568,N_19971);
xor UO_219 (O_219,N_19828,N_19876);
nand UO_220 (O_220,N_19988,N_19813);
xnor UO_221 (O_221,N_19523,N_19654);
or UO_222 (O_222,N_19850,N_19947);
xnor UO_223 (O_223,N_19885,N_19771);
nor UO_224 (O_224,N_19592,N_19857);
and UO_225 (O_225,N_19754,N_19921);
or UO_226 (O_226,N_19913,N_19529);
xnor UO_227 (O_227,N_19939,N_19696);
nor UO_228 (O_228,N_19823,N_19862);
or UO_229 (O_229,N_19743,N_19687);
xor UO_230 (O_230,N_19739,N_19786);
nor UO_231 (O_231,N_19524,N_19719);
or UO_232 (O_232,N_19800,N_19675);
and UO_233 (O_233,N_19992,N_19854);
and UO_234 (O_234,N_19819,N_19541);
xor UO_235 (O_235,N_19776,N_19837);
nand UO_236 (O_236,N_19981,N_19729);
xor UO_237 (O_237,N_19658,N_19914);
or UO_238 (O_238,N_19733,N_19707);
nand UO_239 (O_239,N_19749,N_19989);
xnor UO_240 (O_240,N_19933,N_19510);
nor UO_241 (O_241,N_19899,N_19601);
or UO_242 (O_242,N_19703,N_19737);
nand UO_243 (O_243,N_19932,N_19657);
xor UO_244 (O_244,N_19610,N_19732);
nor UO_245 (O_245,N_19948,N_19802);
xor UO_246 (O_246,N_19961,N_19537);
and UO_247 (O_247,N_19724,N_19587);
xnor UO_248 (O_248,N_19520,N_19870);
or UO_249 (O_249,N_19618,N_19812);
xnor UO_250 (O_250,N_19852,N_19836);
nor UO_251 (O_251,N_19780,N_19816);
nand UO_252 (O_252,N_19786,N_19995);
xor UO_253 (O_253,N_19836,N_19795);
and UO_254 (O_254,N_19548,N_19696);
or UO_255 (O_255,N_19922,N_19869);
or UO_256 (O_256,N_19655,N_19922);
xor UO_257 (O_257,N_19991,N_19646);
and UO_258 (O_258,N_19979,N_19975);
or UO_259 (O_259,N_19924,N_19951);
nor UO_260 (O_260,N_19734,N_19518);
or UO_261 (O_261,N_19984,N_19589);
or UO_262 (O_262,N_19970,N_19883);
or UO_263 (O_263,N_19787,N_19851);
nand UO_264 (O_264,N_19601,N_19826);
nand UO_265 (O_265,N_19523,N_19711);
xor UO_266 (O_266,N_19712,N_19736);
xor UO_267 (O_267,N_19859,N_19708);
or UO_268 (O_268,N_19983,N_19951);
or UO_269 (O_269,N_19860,N_19830);
xnor UO_270 (O_270,N_19511,N_19742);
or UO_271 (O_271,N_19722,N_19533);
and UO_272 (O_272,N_19995,N_19778);
or UO_273 (O_273,N_19592,N_19676);
or UO_274 (O_274,N_19570,N_19692);
xor UO_275 (O_275,N_19758,N_19814);
and UO_276 (O_276,N_19999,N_19834);
and UO_277 (O_277,N_19859,N_19687);
xor UO_278 (O_278,N_19730,N_19966);
nand UO_279 (O_279,N_19597,N_19886);
and UO_280 (O_280,N_19882,N_19847);
and UO_281 (O_281,N_19773,N_19720);
xor UO_282 (O_282,N_19661,N_19925);
nand UO_283 (O_283,N_19651,N_19562);
or UO_284 (O_284,N_19854,N_19941);
xor UO_285 (O_285,N_19803,N_19635);
xor UO_286 (O_286,N_19966,N_19880);
xor UO_287 (O_287,N_19902,N_19916);
nand UO_288 (O_288,N_19905,N_19793);
nor UO_289 (O_289,N_19859,N_19938);
or UO_290 (O_290,N_19974,N_19578);
and UO_291 (O_291,N_19558,N_19842);
xnor UO_292 (O_292,N_19537,N_19784);
or UO_293 (O_293,N_19940,N_19578);
nand UO_294 (O_294,N_19936,N_19818);
nand UO_295 (O_295,N_19537,N_19983);
xnor UO_296 (O_296,N_19616,N_19561);
or UO_297 (O_297,N_19529,N_19818);
nand UO_298 (O_298,N_19992,N_19901);
xor UO_299 (O_299,N_19884,N_19715);
xnor UO_300 (O_300,N_19555,N_19917);
or UO_301 (O_301,N_19988,N_19707);
or UO_302 (O_302,N_19558,N_19830);
xor UO_303 (O_303,N_19905,N_19765);
nand UO_304 (O_304,N_19940,N_19877);
xor UO_305 (O_305,N_19883,N_19902);
or UO_306 (O_306,N_19975,N_19773);
nand UO_307 (O_307,N_19506,N_19516);
xor UO_308 (O_308,N_19890,N_19541);
nand UO_309 (O_309,N_19851,N_19651);
or UO_310 (O_310,N_19767,N_19528);
nand UO_311 (O_311,N_19862,N_19685);
nand UO_312 (O_312,N_19668,N_19536);
or UO_313 (O_313,N_19568,N_19804);
and UO_314 (O_314,N_19522,N_19897);
and UO_315 (O_315,N_19542,N_19698);
xor UO_316 (O_316,N_19970,N_19911);
xor UO_317 (O_317,N_19634,N_19780);
nor UO_318 (O_318,N_19653,N_19691);
and UO_319 (O_319,N_19931,N_19827);
nand UO_320 (O_320,N_19658,N_19950);
xor UO_321 (O_321,N_19555,N_19916);
nor UO_322 (O_322,N_19946,N_19963);
xor UO_323 (O_323,N_19606,N_19659);
nand UO_324 (O_324,N_19726,N_19936);
nor UO_325 (O_325,N_19760,N_19876);
nand UO_326 (O_326,N_19890,N_19915);
nand UO_327 (O_327,N_19652,N_19874);
or UO_328 (O_328,N_19781,N_19509);
or UO_329 (O_329,N_19934,N_19540);
and UO_330 (O_330,N_19712,N_19528);
and UO_331 (O_331,N_19934,N_19919);
xnor UO_332 (O_332,N_19896,N_19689);
and UO_333 (O_333,N_19622,N_19762);
and UO_334 (O_334,N_19622,N_19556);
xnor UO_335 (O_335,N_19942,N_19761);
nand UO_336 (O_336,N_19509,N_19542);
or UO_337 (O_337,N_19810,N_19503);
nor UO_338 (O_338,N_19607,N_19635);
nor UO_339 (O_339,N_19782,N_19858);
nor UO_340 (O_340,N_19782,N_19971);
or UO_341 (O_341,N_19753,N_19678);
and UO_342 (O_342,N_19964,N_19705);
and UO_343 (O_343,N_19982,N_19945);
xor UO_344 (O_344,N_19956,N_19943);
xor UO_345 (O_345,N_19775,N_19835);
nand UO_346 (O_346,N_19611,N_19859);
nand UO_347 (O_347,N_19652,N_19503);
or UO_348 (O_348,N_19690,N_19693);
and UO_349 (O_349,N_19780,N_19891);
and UO_350 (O_350,N_19841,N_19558);
nor UO_351 (O_351,N_19698,N_19774);
and UO_352 (O_352,N_19566,N_19589);
xnor UO_353 (O_353,N_19797,N_19693);
nand UO_354 (O_354,N_19985,N_19590);
or UO_355 (O_355,N_19531,N_19947);
nor UO_356 (O_356,N_19726,N_19581);
nand UO_357 (O_357,N_19603,N_19714);
xor UO_358 (O_358,N_19797,N_19624);
xnor UO_359 (O_359,N_19897,N_19715);
nand UO_360 (O_360,N_19736,N_19515);
nor UO_361 (O_361,N_19660,N_19817);
nor UO_362 (O_362,N_19891,N_19754);
and UO_363 (O_363,N_19935,N_19659);
or UO_364 (O_364,N_19654,N_19994);
xnor UO_365 (O_365,N_19859,N_19581);
nor UO_366 (O_366,N_19909,N_19551);
xor UO_367 (O_367,N_19959,N_19669);
xnor UO_368 (O_368,N_19722,N_19911);
and UO_369 (O_369,N_19595,N_19600);
and UO_370 (O_370,N_19982,N_19588);
or UO_371 (O_371,N_19824,N_19697);
xor UO_372 (O_372,N_19684,N_19850);
and UO_373 (O_373,N_19906,N_19802);
xor UO_374 (O_374,N_19814,N_19596);
nor UO_375 (O_375,N_19699,N_19750);
and UO_376 (O_376,N_19808,N_19850);
nor UO_377 (O_377,N_19673,N_19560);
nand UO_378 (O_378,N_19920,N_19835);
nor UO_379 (O_379,N_19917,N_19836);
nand UO_380 (O_380,N_19968,N_19967);
or UO_381 (O_381,N_19678,N_19543);
xnor UO_382 (O_382,N_19731,N_19610);
and UO_383 (O_383,N_19625,N_19532);
or UO_384 (O_384,N_19790,N_19972);
nand UO_385 (O_385,N_19507,N_19777);
and UO_386 (O_386,N_19951,N_19806);
or UO_387 (O_387,N_19736,N_19866);
nor UO_388 (O_388,N_19593,N_19949);
or UO_389 (O_389,N_19849,N_19711);
and UO_390 (O_390,N_19607,N_19862);
nor UO_391 (O_391,N_19874,N_19975);
and UO_392 (O_392,N_19811,N_19764);
nand UO_393 (O_393,N_19979,N_19528);
or UO_394 (O_394,N_19789,N_19846);
and UO_395 (O_395,N_19512,N_19907);
nand UO_396 (O_396,N_19913,N_19874);
nand UO_397 (O_397,N_19733,N_19627);
and UO_398 (O_398,N_19837,N_19894);
nor UO_399 (O_399,N_19753,N_19896);
and UO_400 (O_400,N_19812,N_19782);
nand UO_401 (O_401,N_19559,N_19612);
nor UO_402 (O_402,N_19949,N_19528);
nor UO_403 (O_403,N_19811,N_19819);
xnor UO_404 (O_404,N_19699,N_19980);
nor UO_405 (O_405,N_19854,N_19908);
and UO_406 (O_406,N_19914,N_19581);
xnor UO_407 (O_407,N_19717,N_19769);
or UO_408 (O_408,N_19709,N_19915);
nand UO_409 (O_409,N_19847,N_19592);
xor UO_410 (O_410,N_19700,N_19970);
xnor UO_411 (O_411,N_19519,N_19516);
xor UO_412 (O_412,N_19735,N_19786);
nand UO_413 (O_413,N_19754,N_19999);
or UO_414 (O_414,N_19934,N_19964);
and UO_415 (O_415,N_19600,N_19824);
or UO_416 (O_416,N_19631,N_19993);
xnor UO_417 (O_417,N_19620,N_19969);
xnor UO_418 (O_418,N_19652,N_19837);
xor UO_419 (O_419,N_19830,N_19809);
and UO_420 (O_420,N_19731,N_19539);
nand UO_421 (O_421,N_19570,N_19583);
nand UO_422 (O_422,N_19540,N_19702);
and UO_423 (O_423,N_19875,N_19835);
or UO_424 (O_424,N_19655,N_19900);
and UO_425 (O_425,N_19775,N_19535);
xor UO_426 (O_426,N_19578,N_19656);
nand UO_427 (O_427,N_19952,N_19818);
and UO_428 (O_428,N_19876,N_19692);
and UO_429 (O_429,N_19539,N_19814);
or UO_430 (O_430,N_19921,N_19611);
xor UO_431 (O_431,N_19844,N_19722);
nor UO_432 (O_432,N_19792,N_19515);
nand UO_433 (O_433,N_19771,N_19996);
xnor UO_434 (O_434,N_19992,N_19581);
nor UO_435 (O_435,N_19941,N_19674);
nand UO_436 (O_436,N_19531,N_19809);
xor UO_437 (O_437,N_19782,N_19882);
or UO_438 (O_438,N_19723,N_19569);
or UO_439 (O_439,N_19816,N_19731);
or UO_440 (O_440,N_19631,N_19679);
xnor UO_441 (O_441,N_19995,N_19991);
nand UO_442 (O_442,N_19654,N_19623);
or UO_443 (O_443,N_19692,N_19748);
xnor UO_444 (O_444,N_19686,N_19937);
and UO_445 (O_445,N_19631,N_19866);
xor UO_446 (O_446,N_19521,N_19916);
nor UO_447 (O_447,N_19873,N_19938);
and UO_448 (O_448,N_19723,N_19999);
nor UO_449 (O_449,N_19523,N_19941);
nand UO_450 (O_450,N_19584,N_19976);
and UO_451 (O_451,N_19942,N_19594);
or UO_452 (O_452,N_19639,N_19807);
nand UO_453 (O_453,N_19646,N_19895);
or UO_454 (O_454,N_19759,N_19780);
xor UO_455 (O_455,N_19595,N_19581);
xor UO_456 (O_456,N_19921,N_19664);
or UO_457 (O_457,N_19569,N_19990);
nand UO_458 (O_458,N_19767,N_19921);
nand UO_459 (O_459,N_19970,N_19830);
nor UO_460 (O_460,N_19836,N_19578);
or UO_461 (O_461,N_19707,N_19718);
and UO_462 (O_462,N_19829,N_19955);
nand UO_463 (O_463,N_19913,N_19637);
nor UO_464 (O_464,N_19964,N_19622);
and UO_465 (O_465,N_19677,N_19915);
and UO_466 (O_466,N_19555,N_19568);
and UO_467 (O_467,N_19707,N_19837);
or UO_468 (O_468,N_19810,N_19641);
nor UO_469 (O_469,N_19653,N_19774);
xor UO_470 (O_470,N_19979,N_19840);
nor UO_471 (O_471,N_19589,N_19892);
or UO_472 (O_472,N_19840,N_19586);
nand UO_473 (O_473,N_19611,N_19699);
and UO_474 (O_474,N_19706,N_19890);
xor UO_475 (O_475,N_19503,N_19539);
xor UO_476 (O_476,N_19505,N_19755);
nand UO_477 (O_477,N_19703,N_19914);
or UO_478 (O_478,N_19786,N_19628);
nand UO_479 (O_479,N_19646,N_19877);
nand UO_480 (O_480,N_19892,N_19957);
nand UO_481 (O_481,N_19646,N_19660);
and UO_482 (O_482,N_19558,N_19660);
nand UO_483 (O_483,N_19990,N_19736);
nand UO_484 (O_484,N_19926,N_19610);
nor UO_485 (O_485,N_19772,N_19759);
nand UO_486 (O_486,N_19985,N_19890);
or UO_487 (O_487,N_19672,N_19636);
nand UO_488 (O_488,N_19838,N_19871);
xnor UO_489 (O_489,N_19733,N_19939);
nor UO_490 (O_490,N_19630,N_19588);
nor UO_491 (O_491,N_19877,N_19601);
nor UO_492 (O_492,N_19820,N_19913);
nand UO_493 (O_493,N_19995,N_19823);
nand UO_494 (O_494,N_19751,N_19550);
or UO_495 (O_495,N_19579,N_19647);
and UO_496 (O_496,N_19959,N_19713);
xnor UO_497 (O_497,N_19922,N_19913);
or UO_498 (O_498,N_19693,N_19985);
nor UO_499 (O_499,N_19896,N_19831);
nor UO_500 (O_500,N_19911,N_19566);
or UO_501 (O_501,N_19618,N_19797);
or UO_502 (O_502,N_19934,N_19943);
nor UO_503 (O_503,N_19848,N_19658);
or UO_504 (O_504,N_19632,N_19778);
nand UO_505 (O_505,N_19996,N_19645);
and UO_506 (O_506,N_19603,N_19798);
xnor UO_507 (O_507,N_19852,N_19758);
nand UO_508 (O_508,N_19767,N_19699);
or UO_509 (O_509,N_19754,N_19910);
or UO_510 (O_510,N_19515,N_19770);
nor UO_511 (O_511,N_19976,N_19572);
and UO_512 (O_512,N_19747,N_19870);
xnor UO_513 (O_513,N_19743,N_19692);
nand UO_514 (O_514,N_19941,N_19839);
and UO_515 (O_515,N_19871,N_19666);
nand UO_516 (O_516,N_19593,N_19898);
xor UO_517 (O_517,N_19864,N_19758);
xnor UO_518 (O_518,N_19939,N_19935);
and UO_519 (O_519,N_19621,N_19726);
xor UO_520 (O_520,N_19889,N_19673);
nor UO_521 (O_521,N_19560,N_19762);
nand UO_522 (O_522,N_19855,N_19674);
or UO_523 (O_523,N_19614,N_19927);
xnor UO_524 (O_524,N_19994,N_19911);
nand UO_525 (O_525,N_19504,N_19745);
and UO_526 (O_526,N_19885,N_19639);
nand UO_527 (O_527,N_19949,N_19660);
nand UO_528 (O_528,N_19815,N_19627);
nand UO_529 (O_529,N_19979,N_19563);
nand UO_530 (O_530,N_19737,N_19844);
nand UO_531 (O_531,N_19813,N_19957);
and UO_532 (O_532,N_19991,N_19820);
nor UO_533 (O_533,N_19958,N_19646);
or UO_534 (O_534,N_19504,N_19673);
and UO_535 (O_535,N_19617,N_19524);
nand UO_536 (O_536,N_19619,N_19727);
xor UO_537 (O_537,N_19995,N_19581);
and UO_538 (O_538,N_19946,N_19809);
or UO_539 (O_539,N_19764,N_19585);
and UO_540 (O_540,N_19518,N_19515);
nor UO_541 (O_541,N_19737,N_19799);
nand UO_542 (O_542,N_19944,N_19542);
and UO_543 (O_543,N_19627,N_19979);
xor UO_544 (O_544,N_19927,N_19679);
nand UO_545 (O_545,N_19812,N_19805);
or UO_546 (O_546,N_19522,N_19678);
xnor UO_547 (O_547,N_19800,N_19510);
nand UO_548 (O_548,N_19811,N_19911);
nand UO_549 (O_549,N_19526,N_19800);
nand UO_550 (O_550,N_19531,N_19964);
and UO_551 (O_551,N_19525,N_19887);
and UO_552 (O_552,N_19628,N_19528);
nand UO_553 (O_553,N_19778,N_19592);
and UO_554 (O_554,N_19667,N_19877);
nor UO_555 (O_555,N_19921,N_19749);
or UO_556 (O_556,N_19902,N_19977);
xnor UO_557 (O_557,N_19922,N_19816);
nand UO_558 (O_558,N_19908,N_19650);
nor UO_559 (O_559,N_19833,N_19644);
nand UO_560 (O_560,N_19709,N_19503);
or UO_561 (O_561,N_19911,N_19716);
nand UO_562 (O_562,N_19831,N_19550);
nand UO_563 (O_563,N_19762,N_19634);
and UO_564 (O_564,N_19513,N_19571);
or UO_565 (O_565,N_19942,N_19713);
nand UO_566 (O_566,N_19526,N_19642);
or UO_567 (O_567,N_19970,N_19923);
nor UO_568 (O_568,N_19860,N_19726);
xor UO_569 (O_569,N_19885,N_19560);
xnor UO_570 (O_570,N_19653,N_19535);
and UO_571 (O_571,N_19762,N_19893);
or UO_572 (O_572,N_19876,N_19602);
nor UO_573 (O_573,N_19519,N_19736);
nor UO_574 (O_574,N_19737,N_19569);
and UO_575 (O_575,N_19652,N_19799);
nand UO_576 (O_576,N_19539,N_19626);
and UO_577 (O_577,N_19636,N_19802);
nand UO_578 (O_578,N_19893,N_19628);
xor UO_579 (O_579,N_19906,N_19967);
nand UO_580 (O_580,N_19867,N_19886);
and UO_581 (O_581,N_19785,N_19864);
nand UO_582 (O_582,N_19981,N_19547);
nand UO_583 (O_583,N_19900,N_19808);
nand UO_584 (O_584,N_19963,N_19913);
xnor UO_585 (O_585,N_19997,N_19742);
and UO_586 (O_586,N_19692,N_19696);
xor UO_587 (O_587,N_19685,N_19500);
and UO_588 (O_588,N_19875,N_19807);
nor UO_589 (O_589,N_19522,N_19717);
or UO_590 (O_590,N_19571,N_19949);
nor UO_591 (O_591,N_19843,N_19951);
nor UO_592 (O_592,N_19570,N_19884);
or UO_593 (O_593,N_19645,N_19927);
nand UO_594 (O_594,N_19553,N_19606);
nor UO_595 (O_595,N_19996,N_19653);
nand UO_596 (O_596,N_19759,N_19882);
nand UO_597 (O_597,N_19500,N_19807);
xor UO_598 (O_598,N_19670,N_19653);
xnor UO_599 (O_599,N_19754,N_19938);
or UO_600 (O_600,N_19584,N_19869);
xor UO_601 (O_601,N_19952,N_19975);
xor UO_602 (O_602,N_19959,N_19794);
xnor UO_603 (O_603,N_19973,N_19704);
nand UO_604 (O_604,N_19931,N_19994);
xor UO_605 (O_605,N_19575,N_19524);
or UO_606 (O_606,N_19759,N_19964);
nor UO_607 (O_607,N_19953,N_19589);
nand UO_608 (O_608,N_19914,N_19934);
nand UO_609 (O_609,N_19598,N_19834);
nor UO_610 (O_610,N_19561,N_19637);
xnor UO_611 (O_611,N_19737,N_19933);
nand UO_612 (O_612,N_19868,N_19759);
xnor UO_613 (O_613,N_19767,N_19764);
and UO_614 (O_614,N_19598,N_19944);
and UO_615 (O_615,N_19627,N_19870);
nor UO_616 (O_616,N_19804,N_19875);
nand UO_617 (O_617,N_19718,N_19591);
or UO_618 (O_618,N_19877,N_19924);
xnor UO_619 (O_619,N_19784,N_19745);
and UO_620 (O_620,N_19976,N_19872);
and UO_621 (O_621,N_19750,N_19586);
xor UO_622 (O_622,N_19960,N_19962);
xor UO_623 (O_623,N_19888,N_19972);
and UO_624 (O_624,N_19919,N_19614);
xor UO_625 (O_625,N_19871,N_19556);
xor UO_626 (O_626,N_19601,N_19533);
nand UO_627 (O_627,N_19717,N_19625);
and UO_628 (O_628,N_19914,N_19972);
nand UO_629 (O_629,N_19606,N_19578);
nor UO_630 (O_630,N_19765,N_19984);
or UO_631 (O_631,N_19818,N_19765);
or UO_632 (O_632,N_19509,N_19957);
and UO_633 (O_633,N_19654,N_19872);
nor UO_634 (O_634,N_19837,N_19509);
nor UO_635 (O_635,N_19740,N_19844);
or UO_636 (O_636,N_19911,N_19586);
xnor UO_637 (O_637,N_19768,N_19623);
nand UO_638 (O_638,N_19785,N_19789);
nor UO_639 (O_639,N_19937,N_19608);
xor UO_640 (O_640,N_19788,N_19936);
nand UO_641 (O_641,N_19696,N_19876);
nor UO_642 (O_642,N_19509,N_19673);
nand UO_643 (O_643,N_19641,N_19907);
or UO_644 (O_644,N_19743,N_19817);
xnor UO_645 (O_645,N_19554,N_19707);
and UO_646 (O_646,N_19660,N_19639);
nor UO_647 (O_647,N_19644,N_19664);
or UO_648 (O_648,N_19572,N_19556);
xnor UO_649 (O_649,N_19704,N_19791);
nand UO_650 (O_650,N_19517,N_19842);
nand UO_651 (O_651,N_19600,N_19625);
and UO_652 (O_652,N_19953,N_19870);
and UO_653 (O_653,N_19907,N_19852);
xor UO_654 (O_654,N_19527,N_19546);
xnor UO_655 (O_655,N_19945,N_19557);
or UO_656 (O_656,N_19500,N_19814);
xor UO_657 (O_657,N_19754,N_19721);
nor UO_658 (O_658,N_19598,N_19880);
xor UO_659 (O_659,N_19564,N_19940);
xor UO_660 (O_660,N_19521,N_19901);
xnor UO_661 (O_661,N_19861,N_19935);
xor UO_662 (O_662,N_19520,N_19979);
nand UO_663 (O_663,N_19587,N_19908);
or UO_664 (O_664,N_19536,N_19507);
xor UO_665 (O_665,N_19599,N_19640);
and UO_666 (O_666,N_19996,N_19591);
and UO_667 (O_667,N_19798,N_19679);
xor UO_668 (O_668,N_19509,N_19989);
xnor UO_669 (O_669,N_19545,N_19941);
and UO_670 (O_670,N_19945,N_19998);
nor UO_671 (O_671,N_19911,N_19662);
xnor UO_672 (O_672,N_19913,N_19846);
nand UO_673 (O_673,N_19702,N_19845);
nand UO_674 (O_674,N_19750,N_19853);
or UO_675 (O_675,N_19964,N_19658);
xnor UO_676 (O_676,N_19558,N_19682);
nand UO_677 (O_677,N_19569,N_19761);
nand UO_678 (O_678,N_19729,N_19915);
nand UO_679 (O_679,N_19719,N_19808);
nor UO_680 (O_680,N_19552,N_19776);
and UO_681 (O_681,N_19501,N_19786);
nand UO_682 (O_682,N_19581,N_19611);
nor UO_683 (O_683,N_19580,N_19501);
or UO_684 (O_684,N_19858,N_19791);
or UO_685 (O_685,N_19767,N_19772);
and UO_686 (O_686,N_19757,N_19597);
or UO_687 (O_687,N_19578,N_19603);
nor UO_688 (O_688,N_19883,N_19715);
and UO_689 (O_689,N_19699,N_19815);
or UO_690 (O_690,N_19850,N_19545);
nand UO_691 (O_691,N_19718,N_19721);
nor UO_692 (O_692,N_19544,N_19751);
nand UO_693 (O_693,N_19598,N_19932);
nand UO_694 (O_694,N_19681,N_19627);
nand UO_695 (O_695,N_19556,N_19911);
nor UO_696 (O_696,N_19558,N_19957);
xor UO_697 (O_697,N_19556,N_19694);
nand UO_698 (O_698,N_19646,N_19679);
nand UO_699 (O_699,N_19980,N_19798);
nor UO_700 (O_700,N_19744,N_19651);
nand UO_701 (O_701,N_19596,N_19761);
nor UO_702 (O_702,N_19528,N_19650);
nor UO_703 (O_703,N_19595,N_19657);
nor UO_704 (O_704,N_19982,N_19766);
and UO_705 (O_705,N_19965,N_19794);
and UO_706 (O_706,N_19928,N_19862);
nor UO_707 (O_707,N_19740,N_19640);
and UO_708 (O_708,N_19795,N_19528);
nand UO_709 (O_709,N_19778,N_19639);
xnor UO_710 (O_710,N_19653,N_19940);
nand UO_711 (O_711,N_19653,N_19927);
or UO_712 (O_712,N_19885,N_19950);
or UO_713 (O_713,N_19797,N_19750);
nor UO_714 (O_714,N_19759,N_19558);
or UO_715 (O_715,N_19730,N_19771);
and UO_716 (O_716,N_19775,N_19837);
and UO_717 (O_717,N_19593,N_19708);
nor UO_718 (O_718,N_19922,N_19981);
nand UO_719 (O_719,N_19945,N_19685);
nand UO_720 (O_720,N_19886,N_19767);
xor UO_721 (O_721,N_19686,N_19928);
nor UO_722 (O_722,N_19759,N_19997);
xor UO_723 (O_723,N_19852,N_19896);
and UO_724 (O_724,N_19831,N_19850);
or UO_725 (O_725,N_19581,N_19641);
nor UO_726 (O_726,N_19604,N_19584);
and UO_727 (O_727,N_19647,N_19548);
nand UO_728 (O_728,N_19996,N_19590);
nor UO_729 (O_729,N_19975,N_19630);
nor UO_730 (O_730,N_19932,N_19905);
nor UO_731 (O_731,N_19568,N_19875);
nor UO_732 (O_732,N_19917,N_19684);
xnor UO_733 (O_733,N_19973,N_19696);
nor UO_734 (O_734,N_19940,N_19835);
nor UO_735 (O_735,N_19670,N_19819);
xor UO_736 (O_736,N_19939,N_19734);
nand UO_737 (O_737,N_19571,N_19682);
nand UO_738 (O_738,N_19539,N_19894);
nor UO_739 (O_739,N_19812,N_19701);
xnor UO_740 (O_740,N_19644,N_19655);
xor UO_741 (O_741,N_19918,N_19882);
nor UO_742 (O_742,N_19752,N_19771);
nor UO_743 (O_743,N_19522,N_19514);
nand UO_744 (O_744,N_19955,N_19851);
xnor UO_745 (O_745,N_19777,N_19557);
and UO_746 (O_746,N_19683,N_19810);
xor UO_747 (O_747,N_19558,N_19828);
nand UO_748 (O_748,N_19535,N_19678);
xnor UO_749 (O_749,N_19898,N_19637);
and UO_750 (O_750,N_19630,N_19642);
xor UO_751 (O_751,N_19968,N_19784);
xor UO_752 (O_752,N_19564,N_19678);
and UO_753 (O_753,N_19963,N_19923);
nor UO_754 (O_754,N_19512,N_19918);
nor UO_755 (O_755,N_19797,N_19594);
nand UO_756 (O_756,N_19835,N_19850);
or UO_757 (O_757,N_19916,N_19825);
nand UO_758 (O_758,N_19736,N_19902);
and UO_759 (O_759,N_19780,N_19698);
nor UO_760 (O_760,N_19630,N_19584);
nor UO_761 (O_761,N_19945,N_19660);
nor UO_762 (O_762,N_19539,N_19727);
nor UO_763 (O_763,N_19524,N_19576);
xnor UO_764 (O_764,N_19759,N_19914);
nor UO_765 (O_765,N_19627,N_19989);
or UO_766 (O_766,N_19817,N_19616);
and UO_767 (O_767,N_19729,N_19636);
nor UO_768 (O_768,N_19655,N_19951);
nor UO_769 (O_769,N_19632,N_19843);
xor UO_770 (O_770,N_19651,N_19901);
nand UO_771 (O_771,N_19846,N_19942);
xnor UO_772 (O_772,N_19580,N_19656);
nor UO_773 (O_773,N_19607,N_19516);
and UO_774 (O_774,N_19830,N_19604);
and UO_775 (O_775,N_19821,N_19991);
xor UO_776 (O_776,N_19924,N_19969);
and UO_777 (O_777,N_19579,N_19713);
or UO_778 (O_778,N_19965,N_19940);
and UO_779 (O_779,N_19739,N_19575);
nor UO_780 (O_780,N_19680,N_19920);
xnor UO_781 (O_781,N_19928,N_19939);
xor UO_782 (O_782,N_19861,N_19690);
xor UO_783 (O_783,N_19617,N_19771);
nand UO_784 (O_784,N_19571,N_19989);
nor UO_785 (O_785,N_19556,N_19760);
nand UO_786 (O_786,N_19676,N_19581);
and UO_787 (O_787,N_19949,N_19882);
nor UO_788 (O_788,N_19532,N_19895);
and UO_789 (O_789,N_19733,N_19898);
xor UO_790 (O_790,N_19899,N_19928);
and UO_791 (O_791,N_19750,N_19643);
or UO_792 (O_792,N_19555,N_19746);
xnor UO_793 (O_793,N_19611,N_19564);
or UO_794 (O_794,N_19688,N_19987);
and UO_795 (O_795,N_19898,N_19854);
and UO_796 (O_796,N_19966,N_19702);
nand UO_797 (O_797,N_19854,N_19584);
and UO_798 (O_798,N_19977,N_19638);
nand UO_799 (O_799,N_19965,N_19787);
or UO_800 (O_800,N_19651,N_19821);
and UO_801 (O_801,N_19562,N_19589);
nand UO_802 (O_802,N_19962,N_19941);
nor UO_803 (O_803,N_19575,N_19521);
nor UO_804 (O_804,N_19927,N_19674);
xor UO_805 (O_805,N_19650,N_19939);
nor UO_806 (O_806,N_19620,N_19613);
and UO_807 (O_807,N_19887,N_19501);
nor UO_808 (O_808,N_19697,N_19571);
nor UO_809 (O_809,N_19652,N_19511);
nor UO_810 (O_810,N_19813,N_19972);
nor UO_811 (O_811,N_19841,N_19793);
and UO_812 (O_812,N_19977,N_19533);
and UO_813 (O_813,N_19626,N_19887);
and UO_814 (O_814,N_19560,N_19869);
nand UO_815 (O_815,N_19894,N_19712);
nor UO_816 (O_816,N_19805,N_19576);
or UO_817 (O_817,N_19548,N_19503);
xor UO_818 (O_818,N_19651,N_19770);
nand UO_819 (O_819,N_19597,N_19715);
xnor UO_820 (O_820,N_19650,N_19929);
xnor UO_821 (O_821,N_19829,N_19685);
nor UO_822 (O_822,N_19687,N_19839);
nand UO_823 (O_823,N_19616,N_19747);
nand UO_824 (O_824,N_19740,N_19614);
or UO_825 (O_825,N_19506,N_19938);
nor UO_826 (O_826,N_19690,N_19538);
or UO_827 (O_827,N_19718,N_19633);
or UO_828 (O_828,N_19902,N_19615);
or UO_829 (O_829,N_19596,N_19619);
or UO_830 (O_830,N_19808,N_19735);
nand UO_831 (O_831,N_19865,N_19989);
and UO_832 (O_832,N_19923,N_19712);
or UO_833 (O_833,N_19896,N_19804);
nor UO_834 (O_834,N_19906,N_19558);
nor UO_835 (O_835,N_19535,N_19868);
or UO_836 (O_836,N_19539,N_19823);
and UO_837 (O_837,N_19754,N_19755);
nor UO_838 (O_838,N_19603,N_19608);
and UO_839 (O_839,N_19928,N_19837);
xor UO_840 (O_840,N_19725,N_19959);
and UO_841 (O_841,N_19608,N_19944);
or UO_842 (O_842,N_19933,N_19981);
nor UO_843 (O_843,N_19710,N_19892);
nand UO_844 (O_844,N_19942,N_19522);
xnor UO_845 (O_845,N_19654,N_19554);
or UO_846 (O_846,N_19947,N_19752);
nor UO_847 (O_847,N_19760,N_19715);
nand UO_848 (O_848,N_19717,N_19718);
and UO_849 (O_849,N_19955,N_19528);
and UO_850 (O_850,N_19535,N_19641);
or UO_851 (O_851,N_19795,N_19516);
and UO_852 (O_852,N_19825,N_19692);
nand UO_853 (O_853,N_19698,N_19551);
nand UO_854 (O_854,N_19996,N_19857);
nand UO_855 (O_855,N_19593,N_19983);
and UO_856 (O_856,N_19511,N_19916);
nor UO_857 (O_857,N_19998,N_19780);
or UO_858 (O_858,N_19524,N_19628);
or UO_859 (O_859,N_19889,N_19508);
nor UO_860 (O_860,N_19687,N_19777);
and UO_861 (O_861,N_19674,N_19999);
and UO_862 (O_862,N_19578,N_19570);
or UO_863 (O_863,N_19734,N_19539);
or UO_864 (O_864,N_19858,N_19623);
xor UO_865 (O_865,N_19890,N_19546);
or UO_866 (O_866,N_19905,N_19839);
or UO_867 (O_867,N_19846,N_19733);
nand UO_868 (O_868,N_19958,N_19680);
or UO_869 (O_869,N_19862,N_19645);
nor UO_870 (O_870,N_19751,N_19703);
nand UO_871 (O_871,N_19646,N_19569);
xnor UO_872 (O_872,N_19796,N_19664);
or UO_873 (O_873,N_19864,N_19790);
and UO_874 (O_874,N_19802,N_19803);
nand UO_875 (O_875,N_19997,N_19907);
and UO_876 (O_876,N_19557,N_19728);
and UO_877 (O_877,N_19564,N_19682);
and UO_878 (O_878,N_19958,N_19608);
xnor UO_879 (O_879,N_19881,N_19732);
and UO_880 (O_880,N_19657,N_19504);
or UO_881 (O_881,N_19615,N_19911);
and UO_882 (O_882,N_19580,N_19935);
xor UO_883 (O_883,N_19596,N_19847);
nor UO_884 (O_884,N_19789,N_19925);
and UO_885 (O_885,N_19632,N_19961);
and UO_886 (O_886,N_19605,N_19972);
nor UO_887 (O_887,N_19678,N_19743);
xnor UO_888 (O_888,N_19567,N_19832);
nand UO_889 (O_889,N_19701,N_19570);
nor UO_890 (O_890,N_19926,N_19579);
xnor UO_891 (O_891,N_19837,N_19714);
nand UO_892 (O_892,N_19740,N_19968);
nor UO_893 (O_893,N_19806,N_19814);
nand UO_894 (O_894,N_19753,N_19780);
nor UO_895 (O_895,N_19612,N_19701);
nor UO_896 (O_896,N_19576,N_19628);
nand UO_897 (O_897,N_19827,N_19953);
or UO_898 (O_898,N_19874,N_19831);
xnor UO_899 (O_899,N_19935,N_19952);
nand UO_900 (O_900,N_19802,N_19628);
and UO_901 (O_901,N_19821,N_19586);
or UO_902 (O_902,N_19800,N_19585);
nand UO_903 (O_903,N_19694,N_19644);
and UO_904 (O_904,N_19716,N_19999);
or UO_905 (O_905,N_19705,N_19701);
nor UO_906 (O_906,N_19798,N_19772);
xnor UO_907 (O_907,N_19999,N_19788);
or UO_908 (O_908,N_19600,N_19745);
nand UO_909 (O_909,N_19738,N_19518);
nand UO_910 (O_910,N_19554,N_19708);
xor UO_911 (O_911,N_19749,N_19976);
xor UO_912 (O_912,N_19506,N_19866);
xnor UO_913 (O_913,N_19896,N_19817);
and UO_914 (O_914,N_19728,N_19967);
nor UO_915 (O_915,N_19912,N_19948);
nor UO_916 (O_916,N_19657,N_19827);
and UO_917 (O_917,N_19920,N_19776);
xnor UO_918 (O_918,N_19546,N_19588);
xnor UO_919 (O_919,N_19887,N_19943);
or UO_920 (O_920,N_19730,N_19578);
or UO_921 (O_921,N_19859,N_19614);
nand UO_922 (O_922,N_19856,N_19866);
nor UO_923 (O_923,N_19679,N_19723);
or UO_924 (O_924,N_19564,N_19881);
nand UO_925 (O_925,N_19663,N_19685);
xnor UO_926 (O_926,N_19869,N_19756);
and UO_927 (O_927,N_19571,N_19921);
nor UO_928 (O_928,N_19625,N_19546);
xor UO_929 (O_929,N_19698,N_19809);
nor UO_930 (O_930,N_19537,N_19590);
and UO_931 (O_931,N_19863,N_19973);
nor UO_932 (O_932,N_19881,N_19865);
xnor UO_933 (O_933,N_19746,N_19846);
or UO_934 (O_934,N_19930,N_19980);
nor UO_935 (O_935,N_19534,N_19833);
nand UO_936 (O_936,N_19724,N_19617);
xnor UO_937 (O_937,N_19883,N_19967);
nor UO_938 (O_938,N_19759,N_19870);
nor UO_939 (O_939,N_19846,N_19917);
or UO_940 (O_940,N_19759,N_19999);
and UO_941 (O_941,N_19911,N_19550);
nor UO_942 (O_942,N_19856,N_19742);
and UO_943 (O_943,N_19959,N_19884);
nand UO_944 (O_944,N_19927,N_19595);
nand UO_945 (O_945,N_19700,N_19716);
nor UO_946 (O_946,N_19846,N_19560);
nand UO_947 (O_947,N_19602,N_19717);
xor UO_948 (O_948,N_19834,N_19518);
nand UO_949 (O_949,N_19941,N_19665);
nand UO_950 (O_950,N_19760,N_19973);
xnor UO_951 (O_951,N_19629,N_19576);
nor UO_952 (O_952,N_19817,N_19579);
nand UO_953 (O_953,N_19739,N_19751);
xor UO_954 (O_954,N_19877,N_19893);
xnor UO_955 (O_955,N_19802,N_19855);
nand UO_956 (O_956,N_19725,N_19789);
xor UO_957 (O_957,N_19588,N_19580);
nand UO_958 (O_958,N_19698,N_19743);
and UO_959 (O_959,N_19571,N_19994);
xor UO_960 (O_960,N_19543,N_19564);
and UO_961 (O_961,N_19670,N_19638);
nor UO_962 (O_962,N_19639,N_19898);
xnor UO_963 (O_963,N_19661,N_19940);
nor UO_964 (O_964,N_19861,N_19937);
xnor UO_965 (O_965,N_19995,N_19652);
xnor UO_966 (O_966,N_19754,N_19594);
nand UO_967 (O_967,N_19991,N_19908);
nand UO_968 (O_968,N_19665,N_19849);
and UO_969 (O_969,N_19980,N_19595);
xnor UO_970 (O_970,N_19569,N_19573);
nand UO_971 (O_971,N_19888,N_19854);
xor UO_972 (O_972,N_19790,N_19622);
xor UO_973 (O_973,N_19565,N_19953);
nor UO_974 (O_974,N_19686,N_19763);
xnor UO_975 (O_975,N_19765,N_19523);
nand UO_976 (O_976,N_19524,N_19565);
and UO_977 (O_977,N_19557,N_19862);
xnor UO_978 (O_978,N_19768,N_19631);
or UO_979 (O_979,N_19863,N_19761);
or UO_980 (O_980,N_19823,N_19955);
nand UO_981 (O_981,N_19712,N_19566);
or UO_982 (O_982,N_19566,N_19725);
or UO_983 (O_983,N_19984,N_19704);
nor UO_984 (O_984,N_19756,N_19735);
xor UO_985 (O_985,N_19941,N_19850);
and UO_986 (O_986,N_19840,N_19731);
xor UO_987 (O_987,N_19993,N_19900);
and UO_988 (O_988,N_19876,N_19750);
xnor UO_989 (O_989,N_19967,N_19713);
nor UO_990 (O_990,N_19547,N_19728);
nor UO_991 (O_991,N_19883,N_19717);
nor UO_992 (O_992,N_19946,N_19671);
and UO_993 (O_993,N_19567,N_19743);
and UO_994 (O_994,N_19663,N_19592);
xnor UO_995 (O_995,N_19574,N_19988);
nand UO_996 (O_996,N_19810,N_19509);
nand UO_997 (O_997,N_19986,N_19896);
or UO_998 (O_998,N_19583,N_19538);
xnor UO_999 (O_999,N_19623,N_19715);
nand UO_1000 (O_1000,N_19559,N_19536);
nand UO_1001 (O_1001,N_19501,N_19999);
xor UO_1002 (O_1002,N_19791,N_19687);
or UO_1003 (O_1003,N_19664,N_19524);
or UO_1004 (O_1004,N_19834,N_19661);
nor UO_1005 (O_1005,N_19925,N_19984);
nor UO_1006 (O_1006,N_19776,N_19926);
nor UO_1007 (O_1007,N_19795,N_19897);
and UO_1008 (O_1008,N_19548,N_19650);
nand UO_1009 (O_1009,N_19996,N_19875);
or UO_1010 (O_1010,N_19657,N_19587);
nand UO_1011 (O_1011,N_19681,N_19557);
and UO_1012 (O_1012,N_19996,N_19777);
xor UO_1013 (O_1013,N_19728,N_19756);
nand UO_1014 (O_1014,N_19680,N_19799);
or UO_1015 (O_1015,N_19847,N_19570);
nor UO_1016 (O_1016,N_19560,N_19875);
nand UO_1017 (O_1017,N_19604,N_19976);
and UO_1018 (O_1018,N_19641,N_19533);
or UO_1019 (O_1019,N_19804,N_19756);
nand UO_1020 (O_1020,N_19683,N_19601);
nor UO_1021 (O_1021,N_19879,N_19576);
nand UO_1022 (O_1022,N_19728,N_19609);
nor UO_1023 (O_1023,N_19795,N_19895);
and UO_1024 (O_1024,N_19628,N_19619);
nor UO_1025 (O_1025,N_19561,N_19770);
or UO_1026 (O_1026,N_19855,N_19871);
nand UO_1027 (O_1027,N_19718,N_19625);
nand UO_1028 (O_1028,N_19571,N_19705);
nand UO_1029 (O_1029,N_19542,N_19855);
nand UO_1030 (O_1030,N_19896,N_19643);
nor UO_1031 (O_1031,N_19987,N_19682);
nor UO_1032 (O_1032,N_19721,N_19676);
nand UO_1033 (O_1033,N_19524,N_19569);
xor UO_1034 (O_1034,N_19871,N_19607);
and UO_1035 (O_1035,N_19585,N_19934);
nand UO_1036 (O_1036,N_19716,N_19846);
nor UO_1037 (O_1037,N_19649,N_19585);
and UO_1038 (O_1038,N_19995,N_19787);
nand UO_1039 (O_1039,N_19517,N_19847);
and UO_1040 (O_1040,N_19943,N_19687);
nand UO_1041 (O_1041,N_19843,N_19993);
and UO_1042 (O_1042,N_19978,N_19857);
nand UO_1043 (O_1043,N_19781,N_19580);
xor UO_1044 (O_1044,N_19546,N_19715);
xor UO_1045 (O_1045,N_19760,N_19865);
xnor UO_1046 (O_1046,N_19869,N_19592);
or UO_1047 (O_1047,N_19501,N_19948);
or UO_1048 (O_1048,N_19625,N_19954);
or UO_1049 (O_1049,N_19882,N_19896);
xor UO_1050 (O_1050,N_19990,N_19642);
nor UO_1051 (O_1051,N_19935,N_19613);
and UO_1052 (O_1052,N_19797,N_19890);
or UO_1053 (O_1053,N_19600,N_19776);
and UO_1054 (O_1054,N_19853,N_19857);
or UO_1055 (O_1055,N_19795,N_19505);
or UO_1056 (O_1056,N_19807,N_19696);
xnor UO_1057 (O_1057,N_19739,N_19641);
nand UO_1058 (O_1058,N_19927,N_19710);
or UO_1059 (O_1059,N_19947,N_19608);
nor UO_1060 (O_1060,N_19689,N_19996);
nand UO_1061 (O_1061,N_19625,N_19529);
xor UO_1062 (O_1062,N_19811,N_19867);
nor UO_1063 (O_1063,N_19862,N_19777);
or UO_1064 (O_1064,N_19674,N_19951);
xnor UO_1065 (O_1065,N_19952,N_19987);
or UO_1066 (O_1066,N_19668,N_19613);
nor UO_1067 (O_1067,N_19786,N_19561);
xor UO_1068 (O_1068,N_19745,N_19693);
xor UO_1069 (O_1069,N_19767,N_19879);
or UO_1070 (O_1070,N_19879,N_19702);
and UO_1071 (O_1071,N_19531,N_19735);
xor UO_1072 (O_1072,N_19602,N_19535);
xor UO_1073 (O_1073,N_19567,N_19784);
nand UO_1074 (O_1074,N_19935,N_19940);
xnor UO_1075 (O_1075,N_19824,N_19653);
and UO_1076 (O_1076,N_19576,N_19940);
nand UO_1077 (O_1077,N_19698,N_19903);
nor UO_1078 (O_1078,N_19930,N_19820);
nand UO_1079 (O_1079,N_19807,N_19608);
or UO_1080 (O_1080,N_19722,N_19535);
nand UO_1081 (O_1081,N_19935,N_19511);
xor UO_1082 (O_1082,N_19794,N_19964);
nand UO_1083 (O_1083,N_19640,N_19526);
nand UO_1084 (O_1084,N_19869,N_19515);
nor UO_1085 (O_1085,N_19680,N_19515);
and UO_1086 (O_1086,N_19654,N_19620);
and UO_1087 (O_1087,N_19853,N_19765);
and UO_1088 (O_1088,N_19653,N_19830);
nand UO_1089 (O_1089,N_19524,N_19997);
nand UO_1090 (O_1090,N_19986,N_19551);
and UO_1091 (O_1091,N_19768,N_19930);
nand UO_1092 (O_1092,N_19783,N_19941);
xor UO_1093 (O_1093,N_19997,N_19786);
and UO_1094 (O_1094,N_19539,N_19627);
nor UO_1095 (O_1095,N_19981,N_19769);
or UO_1096 (O_1096,N_19825,N_19713);
and UO_1097 (O_1097,N_19531,N_19600);
or UO_1098 (O_1098,N_19901,N_19570);
or UO_1099 (O_1099,N_19733,N_19995);
nor UO_1100 (O_1100,N_19596,N_19765);
nand UO_1101 (O_1101,N_19908,N_19681);
and UO_1102 (O_1102,N_19588,N_19578);
xor UO_1103 (O_1103,N_19615,N_19546);
nor UO_1104 (O_1104,N_19862,N_19932);
nand UO_1105 (O_1105,N_19744,N_19676);
nor UO_1106 (O_1106,N_19926,N_19980);
or UO_1107 (O_1107,N_19857,N_19536);
or UO_1108 (O_1108,N_19594,N_19728);
xnor UO_1109 (O_1109,N_19630,N_19957);
xor UO_1110 (O_1110,N_19663,N_19770);
nand UO_1111 (O_1111,N_19769,N_19509);
or UO_1112 (O_1112,N_19732,N_19702);
xor UO_1113 (O_1113,N_19517,N_19581);
or UO_1114 (O_1114,N_19504,N_19726);
nand UO_1115 (O_1115,N_19591,N_19531);
and UO_1116 (O_1116,N_19831,N_19512);
and UO_1117 (O_1117,N_19862,N_19735);
xor UO_1118 (O_1118,N_19927,N_19901);
nand UO_1119 (O_1119,N_19519,N_19857);
nor UO_1120 (O_1120,N_19980,N_19717);
xnor UO_1121 (O_1121,N_19826,N_19668);
nand UO_1122 (O_1122,N_19792,N_19526);
xnor UO_1123 (O_1123,N_19934,N_19536);
nor UO_1124 (O_1124,N_19961,N_19642);
nor UO_1125 (O_1125,N_19693,N_19503);
nor UO_1126 (O_1126,N_19802,N_19701);
or UO_1127 (O_1127,N_19931,N_19713);
and UO_1128 (O_1128,N_19701,N_19805);
and UO_1129 (O_1129,N_19688,N_19729);
xnor UO_1130 (O_1130,N_19939,N_19512);
xor UO_1131 (O_1131,N_19540,N_19592);
xor UO_1132 (O_1132,N_19725,N_19612);
nand UO_1133 (O_1133,N_19995,N_19785);
nor UO_1134 (O_1134,N_19900,N_19878);
nand UO_1135 (O_1135,N_19825,N_19712);
or UO_1136 (O_1136,N_19615,N_19935);
and UO_1137 (O_1137,N_19723,N_19859);
and UO_1138 (O_1138,N_19710,N_19708);
xnor UO_1139 (O_1139,N_19533,N_19611);
nand UO_1140 (O_1140,N_19533,N_19750);
nor UO_1141 (O_1141,N_19713,N_19960);
nor UO_1142 (O_1142,N_19956,N_19819);
and UO_1143 (O_1143,N_19850,N_19898);
and UO_1144 (O_1144,N_19718,N_19615);
xnor UO_1145 (O_1145,N_19932,N_19762);
nor UO_1146 (O_1146,N_19773,N_19658);
xor UO_1147 (O_1147,N_19891,N_19687);
xnor UO_1148 (O_1148,N_19693,N_19769);
nand UO_1149 (O_1149,N_19871,N_19549);
and UO_1150 (O_1150,N_19945,N_19645);
xnor UO_1151 (O_1151,N_19964,N_19525);
nor UO_1152 (O_1152,N_19794,N_19567);
or UO_1153 (O_1153,N_19663,N_19581);
nand UO_1154 (O_1154,N_19627,N_19716);
or UO_1155 (O_1155,N_19558,N_19907);
nor UO_1156 (O_1156,N_19939,N_19652);
nor UO_1157 (O_1157,N_19941,N_19972);
and UO_1158 (O_1158,N_19895,N_19555);
and UO_1159 (O_1159,N_19857,N_19665);
nor UO_1160 (O_1160,N_19629,N_19897);
xor UO_1161 (O_1161,N_19761,N_19877);
nand UO_1162 (O_1162,N_19583,N_19852);
nand UO_1163 (O_1163,N_19902,N_19986);
nand UO_1164 (O_1164,N_19873,N_19503);
and UO_1165 (O_1165,N_19896,N_19574);
or UO_1166 (O_1166,N_19665,N_19595);
nor UO_1167 (O_1167,N_19994,N_19613);
and UO_1168 (O_1168,N_19547,N_19568);
or UO_1169 (O_1169,N_19627,N_19506);
xor UO_1170 (O_1170,N_19732,N_19898);
xor UO_1171 (O_1171,N_19628,N_19980);
nor UO_1172 (O_1172,N_19644,N_19829);
or UO_1173 (O_1173,N_19858,N_19551);
or UO_1174 (O_1174,N_19568,N_19958);
or UO_1175 (O_1175,N_19643,N_19987);
and UO_1176 (O_1176,N_19871,N_19777);
nand UO_1177 (O_1177,N_19545,N_19665);
and UO_1178 (O_1178,N_19855,N_19800);
nor UO_1179 (O_1179,N_19861,N_19648);
xor UO_1180 (O_1180,N_19536,N_19986);
nor UO_1181 (O_1181,N_19636,N_19921);
or UO_1182 (O_1182,N_19665,N_19940);
and UO_1183 (O_1183,N_19512,N_19707);
nor UO_1184 (O_1184,N_19543,N_19672);
xor UO_1185 (O_1185,N_19887,N_19730);
xnor UO_1186 (O_1186,N_19764,N_19541);
nor UO_1187 (O_1187,N_19649,N_19555);
nor UO_1188 (O_1188,N_19699,N_19628);
or UO_1189 (O_1189,N_19904,N_19875);
and UO_1190 (O_1190,N_19536,N_19690);
nand UO_1191 (O_1191,N_19666,N_19796);
or UO_1192 (O_1192,N_19621,N_19583);
or UO_1193 (O_1193,N_19972,N_19772);
nor UO_1194 (O_1194,N_19751,N_19715);
xnor UO_1195 (O_1195,N_19726,N_19878);
and UO_1196 (O_1196,N_19641,N_19631);
or UO_1197 (O_1197,N_19860,N_19574);
nor UO_1198 (O_1198,N_19680,N_19948);
xnor UO_1199 (O_1199,N_19738,N_19843);
or UO_1200 (O_1200,N_19904,N_19570);
nand UO_1201 (O_1201,N_19744,N_19557);
xor UO_1202 (O_1202,N_19578,N_19502);
nand UO_1203 (O_1203,N_19508,N_19639);
nor UO_1204 (O_1204,N_19512,N_19740);
nand UO_1205 (O_1205,N_19668,N_19749);
xnor UO_1206 (O_1206,N_19686,N_19508);
xor UO_1207 (O_1207,N_19542,N_19646);
and UO_1208 (O_1208,N_19615,N_19891);
xor UO_1209 (O_1209,N_19707,N_19681);
xnor UO_1210 (O_1210,N_19809,N_19758);
nand UO_1211 (O_1211,N_19705,N_19579);
nand UO_1212 (O_1212,N_19755,N_19665);
or UO_1213 (O_1213,N_19550,N_19545);
nor UO_1214 (O_1214,N_19774,N_19518);
or UO_1215 (O_1215,N_19694,N_19964);
nand UO_1216 (O_1216,N_19702,N_19794);
or UO_1217 (O_1217,N_19761,N_19571);
or UO_1218 (O_1218,N_19574,N_19752);
nor UO_1219 (O_1219,N_19781,N_19923);
and UO_1220 (O_1220,N_19762,N_19990);
and UO_1221 (O_1221,N_19964,N_19889);
or UO_1222 (O_1222,N_19949,N_19938);
nand UO_1223 (O_1223,N_19583,N_19916);
xor UO_1224 (O_1224,N_19803,N_19513);
nor UO_1225 (O_1225,N_19932,N_19675);
nor UO_1226 (O_1226,N_19819,N_19737);
nand UO_1227 (O_1227,N_19754,N_19625);
xor UO_1228 (O_1228,N_19678,N_19783);
xor UO_1229 (O_1229,N_19947,N_19783);
nand UO_1230 (O_1230,N_19693,N_19927);
xnor UO_1231 (O_1231,N_19660,N_19746);
xor UO_1232 (O_1232,N_19505,N_19671);
and UO_1233 (O_1233,N_19605,N_19627);
xor UO_1234 (O_1234,N_19953,N_19625);
xnor UO_1235 (O_1235,N_19661,N_19612);
nor UO_1236 (O_1236,N_19776,N_19716);
or UO_1237 (O_1237,N_19538,N_19917);
xor UO_1238 (O_1238,N_19708,N_19946);
xor UO_1239 (O_1239,N_19561,N_19640);
or UO_1240 (O_1240,N_19787,N_19690);
and UO_1241 (O_1241,N_19912,N_19570);
nand UO_1242 (O_1242,N_19807,N_19601);
and UO_1243 (O_1243,N_19938,N_19609);
nor UO_1244 (O_1244,N_19866,N_19749);
xor UO_1245 (O_1245,N_19881,N_19502);
nor UO_1246 (O_1246,N_19606,N_19947);
nor UO_1247 (O_1247,N_19527,N_19508);
or UO_1248 (O_1248,N_19884,N_19523);
and UO_1249 (O_1249,N_19624,N_19558);
nand UO_1250 (O_1250,N_19906,N_19604);
nand UO_1251 (O_1251,N_19561,N_19760);
and UO_1252 (O_1252,N_19699,N_19825);
xnor UO_1253 (O_1253,N_19595,N_19633);
nor UO_1254 (O_1254,N_19733,N_19674);
xor UO_1255 (O_1255,N_19876,N_19607);
and UO_1256 (O_1256,N_19993,N_19635);
nand UO_1257 (O_1257,N_19524,N_19665);
nand UO_1258 (O_1258,N_19714,N_19512);
or UO_1259 (O_1259,N_19581,N_19667);
xnor UO_1260 (O_1260,N_19515,N_19604);
xor UO_1261 (O_1261,N_19791,N_19707);
nand UO_1262 (O_1262,N_19516,N_19708);
and UO_1263 (O_1263,N_19705,N_19700);
nor UO_1264 (O_1264,N_19765,N_19972);
nand UO_1265 (O_1265,N_19583,N_19834);
and UO_1266 (O_1266,N_19773,N_19685);
nor UO_1267 (O_1267,N_19830,N_19541);
nand UO_1268 (O_1268,N_19587,N_19763);
xnor UO_1269 (O_1269,N_19939,N_19851);
xnor UO_1270 (O_1270,N_19815,N_19611);
and UO_1271 (O_1271,N_19665,N_19910);
and UO_1272 (O_1272,N_19970,N_19843);
or UO_1273 (O_1273,N_19659,N_19814);
nor UO_1274 (O_1274,N_19526,N_19752);
or UO_1275 (O_1275,N_19826,N_19991);
nor UO_1276 (O_1276,N_19689,N_19551);
or UO_1277 (O_1277,N_19627,N_19662);
and UO_1278 (O_1278,N_19560,N_19897);
xor UO_1279 (O_1279,N_19868,N_19702);
or UO_1280 (O_1280,N_19700,N_19656);
nand UO_1281 (O_1281,N_19525,N_19743);
xnor UO_1282 (O_1282,N_19953,N_19797);
and UO_1283 (O_1283,N_19577,N_19977);
nand UO_1284 (O_1284,N_19814,N_19548);
and UO_1285 (O_1285,N_19920,N_19527);
xnor UO_1286 (O_1286,N_19944,N_19994);
or UO_1287 (O_1287,N_19611,N_19860);
nand UO_1288 (O_1288,N_19712,N_19585);
or UO_1289 (O_1289,N_19540,N_19912);
xor UO_1290 (O_1290,N_19821,N_19632);
nor UO_1291 (O_1291,N_19710,N_19678);
and UO_1292 (O_1292,N_19792,N_19842);
and UO_1293 (O_1293,N_19937,N_19577);
or UO_1294 (O_1294,N_19665,N_19763);
and UO_1295 (O_1295,N_19538,N_19716);
nand UO_1296 (O_1296,N_19730,N_19675);
nor UO_1297 (O_1297,N_19797,N_19786);
nand UO_1298 (O_1298,N_19869,N_19918);
nand UO_1299 (O_1299,N_19824,N_19599);
nor UO_1300 (O_1300,N_19981,N_19992);
and UO_1301 (O_1301,N_19737,N_19554);
nand UO_1302 (O_1302,N_19874,N_19519);
or UO_1303 (O_1303,N_19965,N_19963);
and UO_1304 (O_1304,N_19524,N_19901);
nand UO_1305 (O_1305,N_19575,N_19842);
nor UO_1306 (O_1306,N_19724,N_19733);
xnor UO_1307 (O_1307,N_19516,N_19995);
nand UO_1308 (O_1308,N_19614,N_19580);
or UO_1309 (O_1309,N_19920,N_19868);
or UO_1310 (O_1310,N_19926,N_19583);
and UO_1311 (O_1311,N_19690,N_19767);
xnor UO_1312 (O_1312,N_19565,N_19964);
xnor UO_1313 (O_1313,N_19509,N_19852);
nor UO_1314 (O_1314,N_19567,N_19936);
xnor UO_1315 (O_1315,N_19917,N_19803);
and UO_1316 (O_1316,N_19726,N_19855);
nor UO_1317 (O_1317,N_19745,N_19630);
nor UO_1318 (O_1318,N_19955,N_19653);
nor UO_1319 (O_1319,N_19876,N_19768);
or UO_1320 (O_1320,N_19517,N_19923);
and UO_1321 (O_1321,N_19825,N_19798);
nand UO_1322 (O_1322,N_19953,N_19902);
and UO_1323 (O_1323,N_19588,N_19674);
or UO_1324 (O_1324,N_19730,N_19935);
or UO_1325 (O_1325,N_19516,N_19855);
nand UO_1326 (O_1326,N_19621,N_19551);
xor UO_1327 (O_1327,N_19780,N_19723);
and UO_1328 (O_1328,N_19949,N_19718);
nor UO_1329 (O_1329,N_19624,N_19562);
and UO_1330 (O_1330,N_19535,N_19544);
or UO_1331 (O_1331,N_19988,N_19975);
nor UO_1332 (O_1332,N_19953,N_19828);
and UO_1333 (O_1333,N_19924,N_19886);
nand UO_1334 (O_1334,N_19500,N_19669);
and UO_1335 (O_1335,N_19679,N_19512);
xor UO_1336 (O_1336,N_19878,N_19980);
and UO_1337 (O_1337,N_19514,N_19572);
nand UO_1338 (O_1338,N_19529,N_19994);
nor UO_1339 (O_1339,N_19757,N_19603);
or UO_1340 (O_1340,N_19824,N_19737);
or UO_1341 (O_1341,N_19966,N_19862);
or UO_1342 (O_1342,N_19772,N_19990);
xor UO_1343 (O_1343,N_19890,N_19650);
xnor UO_1344 (O_1344,N_19836,N_19587);
nor UO_1345 (O_1345,N_19527,N_19793);
xnor UO_1346 (O_1346,N_19522,N_19575);
nor UO_1347 (O_1347,N_19580,N_19987);
nor UO_1348 (O_1348,N_19891,N_19974);
and UO_1349 (O_1349,N_19623,N_19619);
nand UO_1350 (O_1350,N_19702,N_19723);
nand UO_1351 (O_1351,N_19725,N_19510);
or UO_1352 (O_1352,N_19651,N_19937);
nand UO_1353 (O_1353,N_19978,N_19502);
and UO_1354 (O_1354,N_19529,N_19876);
and UO_1355 (O_1355,N_19774,N_19788);
nand UO_1356 (O_1356,N_19784,N_19503);
and UO_1357 (O_1357,N_19978,N_19616);
nand UO_1358 (O_1358,N_19793,N_19748);
or UO_1359 (O_1359,N_19644,N_19632);
nand UO_1360 (O_1360,N_19874,N_19666);
and UO_1361 (O_1361,N_19849,N_19608);
nand UO_1362 (O_1362,N_19582,N_19610);
xnor UO_1363 (O_1363,N_19530,N_19964);
nor UO_1364 (O_1364,N_19566,N_19971);
nor UO_1365 (O_1365,N_19893,N_19785);
nand UO_1366 (O_1366,N_19776,N_19581);
and UO_1367 (O_1367,N_19770,N_19777);
xor UO_1368 (O_1368,N_19991,N_19667);
and UO_1369 (O_1369,N_19550,N_19599);
nor UO_1370 (O_1370,N_19522,N_19919);
and UO_1371 (O_1371,N_19793,N_19510);
xor UO_1372 (O_1372,N_19932,N_19720);
xor UO_1373 (O_1373,N_19958,N_19640);
or UO_1374 (O_1374,N_19981,N_19540);
nor UO_1375 (O_1375,N_19713,N_19789);
xnor UO_1376 (O_1376,N_19580,N_19761);
nor UO_1377 (O_1377,N_19775,N_19878);
nor UO_1378 (O_1378,N_19534,N_19576);
nor UO_1379 (O_1379,N_19605,N_19950);
nor UO_1380 (O_1380,N_19989,N_19741);
nand UO_1381 (O_1381,N_19837,N_19575);
or UO_1382 (O_1382,N_19933,N_19785);
nand UO_1383 (O_1383,N_19653,N_19626);
nor UO_1384 (O_1384,N_19667,N_19803);
or UO_1385 (O_1385,N_19730,N_19932);
or UO_1386 (O_1386,N_19776,N_19784);
xnor UO_1387 (O_1387,N_19512,N_19618);
nand UO_1388 (O_1388,N_19661,N_19861);
xnor UO_1389 (O_1389,N_19673,N_19608);
or UO_1390 (O_1390,N_19798,N_19987);
or UO_1391 (O_1391,N_19876,N_19515);
or UO_1392 (O_1392,N_19607,N_19714);
nand UO_1393 (O_1393,N_19806,N_19641);
nand UO_1394 (O_1394,N_19988,N_19677);
xnor UO_1395 (O_1395,N_19613,N_19857);
or UO_1396 (O_1396,N_19757,N_19721);
xor UO_1397 (O_1397,N_19647,N_19988);
or UO_1398 (O_1398,N_19579,N_19559);
nor UO_1399 (O_1399,N_19748,N_19533);
nand UO_1400 (O_1400,N_19650,N_19719);
or UO_1401 (O_1401,N_19516,N_19859);
and UO_1402 (O_1402,N_19697,N_19775);
xor UO_1403 (O_1403,N_19724,N_19964);
or UO_1404 (O_1404,N_19976,N_19991);
and UO_1405 (O_1405,N_19889,N_19559);
xnor UO_1406 (O_1406,N_19728,N_19514);
or UO_1407 (O_1407,N_19702,N_19840);
and UO_1408 (O_1408,N_19906,N_19783);
or UO_1409 (O_1409,N_19736,N_19873);
nor UO_1410 (O_1410,N_19779,N_19706);
nand UO_1411 (O_1411,N_19988,N_19818);
nand UO_1412 (O_1412,N_19526,N_19890);
or UO_1413 (O_1413,N_19823,N_19681);
nor UO_1414 (O_1414,N_19896,N_19616);
xnor UO_1415 (O_1415,N_19518,N_19804);
or UO_1416 (O_1416,N_19690,N_19991);
or UO_1417 (O_1417,N_19877,N_19594);
or UO_1418 (O_1418,N_19925,N_19948);
or UO_1419 (O_1419,N_19634,N_19645);
nand UO_1420 (O_1420,N_19518,N_19782);
and UO_1421 (O_1421,N_19831,N_19638);
and UO_1422 (O_1422,N_19728,N_19711);
and UO_1423 (O_1423,N_19621,N_19859);
or UO_1424 (O_1424,N_19947,N_19610);
nor UO_1425 (O_1425,N_19787,N_19988);
and UO_1426 (O_1426,N_19827,N_19887);
xor UO_1427 (O_1427,N_19977,N_19881);
xnor UO_1428 (O_1428,N_19752,N_19710);
and UO_1429 (O_1429,N_19857,N_19925);
xor UO_1430 (O_1430,N_19772,N_19775);
xnor UO_1431 (O_1431,N_19668,N_19533);
nor UO_1432 (O_1432,N_19582,N_19985);
nor UO_1433 (O_1433,N_19689,N_19694);
or UO_1434 (O_1434,N_19602,N_19579);
and UO_1435 (O_1435,N_19817,N_19508);
and UO_1436 (O_1436,N_19538,N_19830);
and UO_1437 (O_1437,N_19539,N_19600);
nor UO_1438 (O_1438,N_19587,N_19906);
or UO_1439 (O_1439,N_19514,N_19636);
nand UO_1440 (O_1440,N_19809,N_19609);
nand UO_1441 (O_1441,N_19700,N_19512);
xnor UO_1442 (O_1442,N_19682,N_19920);
nor UO_1443 (O_1443,N_19859,N_19552);
nand UO_1444 (O_1444,N_19713,N_19700);
nand UO_1445 (O_1445,N_19647,N_19933);
or UO_1446 (O_1446,N_19869,N_19715);
or UO_1447 (O_1447,N_19854,N_19935);
and UO_1448 (O_1448,N_19858,N_19865);
nor UO_1449 (O_1449,N_19575,N_19743);
xor UO_1450 (O_1450,N_19933,N_19844);
and UO_1451 (O_1451,N_19894,N_19560);
or UO_1452 (O_1452,N_19599,N_19844);
or UO_1453 (O_1453,N_19880,N_19734);
and UO_1454 (O_1454,N_19553,N_19739);
nor UO_1455 (O_1455,N_19517,N_19883);
or UO_1456 (O_1456,N_19538,N_19580);
nand UO_1457 (O_1457,N_19964,N_19756);
nor UO_1458 (O_1458,N_19787,N_19968);
nor UO_1459 (O_1459,N_19587,N_19674);
xor UO_1460 (O_1460,N_19566,N_19705);
nor UO_1461 (O_1461,N_19702,N_19538);
nand UO_1462 (O_1462,N_19639,N_19802);
xor UO_1463 (O_1463,N_19593,N_19814);
and UO_1464 (O_1464,N_19670,N_19626);
nor UO_1465 (O_1465,N_19714,N_19533);
nand UO_1466 (O_1466,N_19727,N_19550);
and UO_1467 (O_1467,N_19980,N_19767);
or UO_1468 (O_1468,N_19592,N_19634);
or UO_1469 (O_1469,N_19910,N_19883);
nor UO_1470 (O_1470,N_19830,N_19684);
and UO_1471 (O_1471,N_19843,N_19798);
or UO_1472 (O_1472,N_19707,N_19658);
nor UO_1473 (O_1473,N_19951,N_19653);
nand UO_1474 (O_1474,N_19575,N_19633);
xor UO_1475 (O_1475,N_19756,N_19507);
nor UO_1476 (O_1476,N_19629,N_19683);
or UO_1477 (O_1477,N_19741,N_19749);
or UO_1478 (O_1478,N_19546,N_19898);
and UO_1479 (O_1479,N_19729,N_19819);
and UO_1480 (O_1480,N_19584,N_19636);
and UO_1481 (O_1481,N_19633,N_19740);
or UO_1482 (O_1482,N_19715,N_19855);
xnor UO_1483 (O_1483,N_19892,N_19739);
nand UO_1484 (O_1484,N_19981,N_19742);
xor UO_1485 (O_1485,N_19654,N_19726);
nand UO_1486 (O_1486,N_19573,N_19964);
xnor UO_1487 (O_1487,N_19929,N_19775);
xnor UO_1488 (O_1488,N_19693,N_19725);
or UO_1489 (O_1489,N_19571,N_19732);
xnor UO_1490 (O_1490,N_19950,N_19863);
xor UO_1491 (O_1491,N_19707,N_19981);
and UO_1492 (O_1492,N_19826,N_19650);
and UO_1493 (O_1493,N_19952,N_19914);
nand UO_1494 (O_1494,N_19895,N_19853);
nand UO_1495 (O_1495,N_19837,N_19952);
or UO_1496 (O_1496,N_19845,N_19800);
nor UO_1497 (O_1497,N_19777,N_19546);
and UO_1498 (O_1498,N_19765,N_19549);
and UO_1499 (O_1499,N_19803,N_19861);
nor UO_1500 (O_1500,N_19918,N_19790);
nand UO_1501 (O_1501,N_19767,N_19613);
nor UO_1502 (O_1502,N_19712,N_19921);
and UO_1503 (O_1503,N_19570,N_19878);
and UO_1504 (O_1504,N_19508,N_19590);
nor UO_1505 (O_1505,N_19970,N_19664);
nor UO_1506 (O_1506,N_19734,N_19971);
nand UO_1507 (O_1507,N_19801,N_19921);
nor UO_1508 (O_1508,N_19651,N_19951);
nand UO_1509 (O_1509,N_19973,N_19908);
nand UO_1510 (O_1510,N_19921,N_19550);
and UO_1511 (O_1511,N_19763,N_19793);
or UO_1512 (O_1512,N_19709,N_19951);
nand UO_1513 (O_1513,N_19532,N_19742);
nor UO_1514 (O_1514,N_19856,N_19895);
and UO_1515 (O_1515,N_19545,N_19570);
xor UO_1516 (O_1516,N_19978,N_19805);
or UO_1517 (O_1517,N_19759,N_19824);
nor UO_1518 (O_1518,N_19583,N_19640);
nor UO_1519 (O_1519,N_19776,N_19587);
xnor UO_1520 (O_1520,N_19932,N_19839);
nor UO_1521 (O_1521,N_19627,N_19754);
nor UO_1522 (O_1522,N_19788,N_19992);
and UO_1523 (O_1523,N_19575,N_19863);
or UO_1524 (O_1524,N_19807,N_19887);
nor UO_1525 (O_1525,N_19586,N_19677);
and UO_1526 (O_1526,N_19614,N_19726);
nand UO_1527 (O_1527,N_19514,N_19632);
and UO_1528 (O_1528,N_19758,N_19770);
or UO_1529 (O_1529,N_19688,N_19628);
or UO_1530 (O_1530,N_19997,N_19960);
and UO_1531 (O_1531,N_19766,N_19961);
nand UO_1532 (O_1532,N_19512,N_19537);
nor UO_1533 (O_1533,N_19824,N_19694);
nand UO_1534 (O_1534,N_19574,N_19976);
nand UO_1535 (O_1535,N_19503,N_19664);
and UO_1536 (O_1536,N_19936,N_19690);
and UO_1537 (O_1537,N_19662,N_19704);
nor UO_1538 (O_1538,N_19680,N_19648);
nand UO_1539 (O_1539,N_19892,N_19888);
nand UO_1540 (O_1540,N_19639,N_19587);
xnor UO_1541 (O_1541,N_19956,N_19815);
xnor UO_1542 (O_1542,N_19624,N_19693);
or UO_1543 (O_1543,N_19814,N_19730);
and UO_1544 (O_1544,N_19783,N_19670);
xnor UO_1545 (O_1545,N_19566,N_19599);
nand UO_1546 (O_1546,N_19799,N_19625);
or UO_1547 (O_1547,N_19515,N_19763);
or UO_1548 (O_1548,N_19678,N_19823);
and UO_1549 (O_1549,N_19766,N_19910);
nor UO_1550 (O_1550,N_19903,N_19536);
nand UO_1551 (O_1551,N_19535,N_19942);
nor UO_1552 (O_1552,N_19508,N_19607);
nand UO_1553 (O_1553,N_19853,N_19745);
nor UO_1554 (O_1554,N_19727,N_19522);
nor UO_1555 (O_1555,N_19831,N_19543);
nor UO_1556 (O_1556,N_19759,N_19777);
and UO_1557 (O_1557,N_19917,N_19891);
or UO_1558 (O_1558,N_19773,N_19617);
nor UO_1559 (O_1559,N_19899,N_19990);
or UO_1560 (O_1560,N_19960,N_19850);
or UO_1561 (O_1561,N_19516,N_19579);
nand UO_1562 (O_1562,N_19707,N_19854);
and UO_1563 (O_1563,N_19697,N_19519);
xor UO_1564 (O_1564,N_19862,N_19733);
nor UO_1565 (O_1565,N_19508,N_19636);
and UO_1566 (O_1566,N_19643,N_19950);
xnor UO_1567 (O_1567,N_19905,N_19734);
xor UO_1568 (O_1568,N_19534,N_19926);
xor UO_1569 (O_1569,N_19776,N_19991);
or UO_1570 (O_1570,N_19962,N_19696);
nor UO_1571 (O_1571,N_19806,N_19736);
xor UO_1572 (O_1572,N_19505,N_19605);
nand UO_1573 (O_1573,N_19865,N_19558);
or UO_1574 (O_1574,N_19728,N_19912);
nor UO_1575 (O_1575,N_19700,N_19886);
xor UO_1576 (O_1576,N_19680,N_19641);
or UO_1577 (O_1577,N_19570,N_19879);
or UO_1578 (O_1578,N_19959,N_19676);
or UO_1579 (O_1579,N_19950,N_19955);
nor UO_1580 (O_1580,N_19519,N_19893);
nand UO_1581 (O_1581,N_19956,N_19612);
nand UO_1582 (O_1582,N_19869,N_19780);
nor UO_1583 (O_1583,N_19939,N_19700);
and UO_1584 (O_1584,N_19635,N_19671);
nor UO_1585 (O_1585,N_19827,N_19704);
and UO_1586 (O_1586,N_19951,N_19990);
or UO_1587 (O_1587,N_19822,N_19631);
or UO_1588 (O_1588,N_19835,N_19637);
nand UO_1589 (O_1589,N_19533,N_19874);
and UO_1590 (O_1590,N_19878,N_19927);
nand UO_1591 (O_1591,N_19853,N_19986);
nand UO_1592 (O_1592,N_19608,N_19573);
nor UO_1593 (O_1593,N_19940,N_19726);
nand UO_1594 (O_1594,N_19600,N_19973);
nand UO_1595 (O_1595,N_19985,N_19948);
nand UO_1596 (O_1596,N_19631,N_19861);
nor UO_1597 (O_1597,N_19747,N_19963);
or UO_1598 (O_1598,N_19545,N_19757);
nor UO_1599 (O_1599,N_19648,N_19898);
nor UO_1600 (O_1600,N_19586,N_19657);
and UO_1601 (O_1601,N_19908,N_19507);
and UO_1602 (O_1602,N_19944,N_19736);
and UO_1603 (O_1603,N_19899,N_19818);
xnor UO_1604 (O_1604,N_19752,N_19589);
nand UO_1605 (O_1605,N_19816,N_19855);
nand UO_1606 (O_1606,N_19664,N_19768);
nand UO_1607 (O_1607,N_19687,N_19948);
or UO_1608 (O_1608,N_19776,N_19691);
or UO_1609 (O_1609,N_19587,N_19765);
or UO_1610 (O_1610,N_19545,N_19895);
nor UO_1611 (O_1611,N_19983,N_19716);
xnor UO_1612 (O_1612,N_19631,N_19831);
nor UO_1613 (O_1613,N_19768,N_19836);
xor UO_1614 (O_1614,N_19800,N_19754);
nor UO_1615 (O_1615,N_19778,N_19954);
or UO_1616 (O_1616,N_19557,N_19684);
and UO_1617 (O_1617,N_19965,N_19577);
xor UO_1618 (O_1618,N_19563,N_19997);
nor UO_1619 (O_1619,N_19754,N_19676);
and UO_1620 (O_1620,N_19512,N_19711);
xor UO_1621 (O_1621,N_19864,N_19868);
and UO_1622 (O_1622,N_19930,N_19920);
or UO_1623 (O_1623,N_19554,N_19760);
xor UO_1624 (O_1624,N_19707,N_19754);
or UO_1625 (O_1625,N_19659,N_19967);
nor UO_1626 (O_1626,N_19505,N_19536);
and UO_1627 (O_1627,N_19931,N_19733);
nor UO_1628 (O_1628,N_19516,N_19846);
and UO_1629 (O_1629,N_19744,N_19607);
nor UO_1630 (O_1630,N_19990,N_19756);
and UO_1631 (O_1631,N_19558,N_19739);
nand UO_1632 (O_1632,N_19526,N_19523);
nor UO_1633 (O_1633,N_19545,N_19775);
nor UO_1634 (O_1634,N_19717,N_19600);
nor UO_1635 (O_1635,N_19859,N_19925);
nor UO_1636 (O_1636,N_19696,N_19730);
xnor UO_1637 (O_1637,N_19621,N_19765);
nand UO_1638 (O_1638,N_19622,N_19678);
or UO_1639 (O_1639,N_19540,N_19717);
nor UO_1640 (O_1640,N_19574,N_19682);
nor UO_1641 (O_1641,N_19672,N_19959);
or UO_1642 (O_1642,N_19848,N_19706);
xnor UO_1643 (O_1643,N_19719,N_19995);
and UO_1644 (O_1644,N_19590,N_19709);
or UO_1645 (O_1645,N_19836,N_19799);
xor UO_1646 (O_1646,N_19790,N_19677);
nand UO_1647 (O_1647,N_19569,N_19589);
nand UO_1648 (O_1648,N_19584,N_19531);
or UO_1649 (O_1649,N_19722,N_19978);
xor UO_1650 (O_1650,N_19808,N_19829);
and UO_1651 (O_1651,N_19906,N_19975);
or UO_1652 (O_1652,N_19500,N_19802);
nor UO_1653 (O_1653,N_19715,N_19975);
or UO_1654 (O_1654,N_19664,N_19733);
xnor UO_1655 (O_1655,N_19591,N_19974);
nand UO_1656 (O_1656,N_19717,N_19840);
and UO_1657 (O_1657,N_19630,N_19987);
xor UO_1658 (O_1658,N_19574,N_19877);
or UO_1659 (O_1659,N_19932,N_19617);
xnor UO_1660 (O_1660,N_19534,N_19578);
nand UO_1661 (O_1661,N_19706,N_19815);
or UO_1662 (O_1662,N_19636,N_19590);
xnor UO_1663 (O_1663,N_19555,N_19853);
or UO_1664 (O_1664,N_19598,N_19558);
nor UO_1665 (O_1665,N_19796,N_19886);
nand UO_1666 (O_1666,N_19520,N_19584);
xnor UO_1667 (O_1667,N_19763,N_19706);
nor UO_1668 (O_1668,N_19557,N_19956);
nand UO_1669 (O_1669,N_19755,N_19822);
nand UO_1670 (O_1670,N_19771,N_19954);
nand UO_1671 (O_1671,N_19665,N_19506);
xor UO_1672 (O_1672,N_19807,N_19701);
xnor UO_1673 (O_1673,N_19580,N_19502);
xor UO_1674 (O_1674,N_19600,N_19819);
nand UO_1675 (O_1675,N_19826,N_19913);
and UO_1676 (O_1676,N_19885,N_19989);
xnor UO_1677 (O_1677,N_19524,N_19634);
xor UO_1678 (O_1678,N_19702,N_19905);
and UO_1679 (O_1679,N_19844,N_19806);
xor UO_1680 (O_1680,N_19582,N_19720);
or UO_1681 (O_1681,N_19692,N_19776);
nor UO_1682 (O_1682,N_19976,N_19828);
xor UO_1683 (O_1683,N_19758,N_19731);
xor UO_1684 (O_1684,N_19799,N_19715);
and UO_1685 (O_1685,N_19819,N_19854);
xor UO_1686 (O_1686,N_19594,N_19563);
nor UO_1687 (O_1687,N_19808,N_19562);
and UO_1688 (O_1688,N_19696,N_19905);
or UO_1689 (O_1689,N_19621,N_19782);
nand UO_1690 (O_1690,N_19809,N_19820);
xor UO_1691 (O_1691,N_19548,N_19699);
xnor UO_1692 (O_1692,N_19774,N_19717);
or UO_1693 (O_1693,N_19749,N_19717);
and UO_1694 (O_1694,N_19769,N_19768);
and UO_1695 (O_1695,N_19957,N_19963);
or UO_1696 (O_1696,N_19748,N_19579);
nand UO_1697 (O_1697,N_19838,N_19650);
or UO_1698 (O_1698,N_19664,N_19720);
or UO_1699 (O_1699,N_19637,N_19635);
and UO_1700 (O_1700,N_19782,N_19868);
nor UO_1701 (O_1701,N_19814,N_19602);
xnor UO_1702 (O_1702,N_19819,N_19731);
nand UO_1703 (O_1703,N_19807,N_19937);
or UO_1704 (O_1704,N_19974,N_19812);
nor UO_1705 (O_1705,N_19790,N_19710);
and UO_1706 (O_1706,N_19912,N_19904);
xor UO_1707 (O_1707,N_19598,N_19524);
nand UO_1708 (O_1708,N_19939,N_19943);
nand UO_1709 (O_1709,N_19564,N_19697);
and UO_1710 (O_1710,N_19986,N_19744);
nand UO_1711 (O_1711,N_19546,N_19706);
nand UO_1712 (O_1712,N_19542,N_19607);
or UO_1713 (O_1713,N_19540,N_19803);
or UO_1714 (O_1714,N_19744,N_19669);
or UO_1715 (O_1715,N_19516,N_19960);
nand UO_1716 (O_1716,N_19743,N_19938);
nand UO_1717 (O_1717,N_19873,N_19852);
nand UO_1718 (O_1718,N_19867,N_19769);
nand UO_1719 (O_1719,N_19718,N_19537);
and UO_1720 (O_1720,N_19710,N_19762);
nand UO_1721 (O_1721,N_19871,N_19722);
or UO_1722 (O_1722,N_19664,N_19771);
nand UO_1723 (O_1723,N_19611,N_19867);
xor UO_1724 (O_1724,N_19985,N_19837);
or UO_1725 (O_1725,N_19682,N_19536);
xor UO_1726 (O_1726,N_19897,N_19597);
nand UO_1727 (O_1727,N_19868,N_19743);
xor UO_1728 (O_1728,N_19696,N_19603);
nand UO_1729 (O_1729,N_19644,N_19704);
or UO_1730 (O_1730,N_19678,N_19744);
or UO_1731 (O_1731,N_19857,N_19553);
xor UO_1732 (O_1732,N_19684,N_19852);
xnor UO_1733 (O_1733,N_19859,N_19584);
or UO_1734 (O_1734,N_19617,N_19752);
nand UO_1735 (O_1735,N_19935,N_19905);
xnor UO_1736 (O_1736,N_19696,N_19901);
xnor UO_1737 (O_1737,N_19862,N_19946);
xnor UO_1738 (O_1738,N_19784,N_19618);
xnor UO_1739 (O_1739,N_19818,N_19624);
xnor UO_1740 (O_1740,N_19738,N_19573);
or UO_1741 (O_1741,N_19636,N_19930);
or UO_1742 (O_1742,N_19607,N_19749);
nor UO_1743 (O_1743,N_19629,N_19813);
nand UO_1744 (O_1744,N_19782,N_19988);
and UO_1745 (O_1745,N_19789,N_19933);
xor UO_1746 (O_1746,N_19990,N_19604);
or UO_1747 (O_1747,N_19933,N_19937);
or UO_1748 (O_1748,N_19697,N_19688);
and UO_1749 (O_1749,N_19591,N_19548);
nand UO_1750 (O_1750,N_19723,N_19626);
nor UO_1751 (O_1751,N_19919,N_19769);
and UO_1752 (O_1752,N_19760,N_19607);
xor UO_1753 (O_1753,N_19509,N_19633);
and UO_1754 (O_1754,N_19910,N_19793);
xnor UO_1755 (O_1755,N_19924,N_19917);
nor UO_1756 (O_1756,N_19809,N_19695);
nor UO_1757 (O_1757,N_19791,N_19958);
nand UO_1758 (O_1758,N_19803,N_19728);
nor UO_1759 (O_1759,N_19926,N_19820);
xor UO_1760 (O_1760,N_19785,N_19689);
xor UO_1761 (O_1761,N_19841,N_19893);
and UO_1762 (O_1762,N_19570,N_19989);
xnor UO_1763 (O_1763,N_19514,N_19553);
nor UO_1764 (O_1764,N_19775,N_19744);
xor UO_1765 (O_1765,N_19916,N_19831);
nor UO_1766 (O_1766,N_19774,N_19881);
or UO_1767 (O_1767,N_19716,N_19732);
nand UO_1768 (O_1768,N_19561,N_19711);
nor UO_1769 (O_1769,N_19731,N_19849);
nand UO_1770 (O_1770,N_19533,N_19536);
and UO_1771 (O_1771,N_19681,N_19523);
nor UO_1772 (O_1772,N_19970,N_19509);
and UO_1773 (O_1773,N_19720,N_19569);
nor UO_1774 (O_1774,N_19996,N_19538);
xnor UO_1775 (O_1775,N_19578,N_19669);
nor UO_1776 (O_1776,N_19729,N_19781);
nor UO_1777 (O_1777,N_19927,N_19649);
nor UO_1778 (O_1778,N_19573,N_19778);
nor UO_1779 (O_1779,N_19961,N_19610);
or UO_1780 (O_1780,N_19748,N_19886);
nand UO_1781 (O_1781,N_19541,N_19546);
nor UO_1782 (O_1782,N_19554,N_19685);
nand UO_1783 (O_1783,N_19904,N_19797);
nor UO_1784 (O_1784,N_19885,N_19658);
and UO_1785 (O_1785,N_19840,N_19869);
xnor UO_1786 (O_1786,N_19952,N_19745);
and UO_1787 (O_1787,N_19638,N_19631);
xnor UO_1788 (O_1788,N_19755,N_19975);
or UO_1789 (O_1789,N_19874,N_19725);
and UO_1790 (O_1790,N_19957,N_19722);
nor UO_1791 (O_1791,N_19821,N_19566);
nor UO_1792 (O_1792,N_19659,N_19968);
nor UO_1793 (O_1793,N_19818,N_19501);
nor UO_1794 (O_1794,N_19672,N_19516);
or UO_1795 (O_1795,N_19733,N_19698);
nor UO_1796 (O_1796,N_19666,N_19942);
nor UO_1797 (O_1797,N_19769,N_19621);
nand UO_1798 (O_1798,N_19815,N_19821);
xnor UO_1799 (O_1799,N_19841,N_19687);
nor UO_1800 (O_1800,N_19588,N_19728);
or UO_1801 (O_1801,N_19681,N_19997);
nand UO_1802 (O_1802,N_19760,N_19676);
nor UO_1803 (O_1803,N_19865,N_19819);
or UO_1804 (O_1804,N_19774,N_19791);
xor UO_1805 (O_1805,N_19850,N_19615);
and UO_1806 (O_1806,N_19607,N_19608);
nor UO_1807 (O_1807,N_19683,N_19509);
nand UO_1808 (O_1808,N_19796,N_19558);
nor UO_1809 (O_1809,N_19905,N_19821);
and UO_1810 (O_1810,N_19950,N_19788);
xnor UO_1811 (O_1811,N_19895,N_19668);
nand UO_1812 (O_1812,N_19886,N_19896);
nor UO_1813 (O_1813,N_19934,N_19713);
and UO_1814 (O_1814,N_19759,N_19724);
and UO_1815 (O_1815,N_19619,N_19888);
nand UO_1816 (O_1816,N_19543,N_19746);
and UO_1817 (O_1817,N_19598,N_19754);
nand UO_1818 (O_1818,N_19578,N_19787);
nand UO_1819 (O_1819,N_19728,N_19814);
nor UO_1820 (O_1820,N_19525,N_19997);
and UO_1821 (O_1821,N_19539,N_19816);
xnor UO_1822 (O_1822,N_19747,N_19569);
xor UO_1823 (O_1823,N_19599,N_19652);
xnor UO_1824 (O_1824,N_19746,N_19741);
nand UO_1825 (O_1825,N_19911,N_19596);
xor UO_1826 (O_1826,N_19739,N_19655);
nand UO_1827 (O_1827,N_19595,N_19576);
nand UO_1828 (O_1828,N_19737,N_19585);
xor UO_1829 (O_1829,N_19970,N_19671);
nand UO_1830 (O_1830,N_19544,N_19506);
nand UO_1831 (O_1831,N_19960,N_19852);
or UO_1832 (O_1832,N_19899,N_19814);
nor UO_1833 (O_1833,N_19571,N_19734);
nor UO_1834 (O_1834,N_19927,N_19791);
nand UO_1835 (O_1835,N_19651,N_19845);
or UO_1836 (O_1836,N_19694,N_19835);
or UO_1837 (O_1837,N_19847,N_19927);
and UO_1838 (O_1838,N_19800,N_19642);
and UO_1839 (O_1839,N_19885,N_19964);
and UO_1840 (O_1840,N_19676,N_19843);
or UO_1841 (O_1841,N_19600,N_19758);
xor UO_1842 (O_1842,N_19905,N_19794);
or UO_1843 (O_1843,N_19654,N_19714);
xnor UO_1844 (O_1844,N_19952,N_19695);
nand UO_1845 (O_1845,N_19698,N_19578);
xnor UO_1846 (O_1846,N_19797,N_19672);
xnor UO_1847 (O_1847,N_19919,N_19713);
or UO_1848 (O_1848,N_19789,N_19777);
xor UO_1849 (O_1849,N_19603,N_19980);
or UO_1850 (O_1850,N_19623,N_19662);
nand UO_1851 (O_1851,N_19883,N_19774);
nand UO_1852 (O_1852,N_19513,N_19761);
nand UO_1853 (O_1853,N_19957,N_19546);
nand UO_1854 (O_1854,N_19884,N_19611);
and UO_1855 (O_1855,N_19996,N_19503);
nand UO_1856 (O_1856,N_19731,N_19716);
xnor UO_1857 (O_1857,N_19694,N_19950);
xnor UO_1858 (O_1858,N_19925,N_19749);
xor UO_1859 (O_1859,N_19556,N_19914);
nor UO_1860 (O_1860,N_19621,N_19604);
nand UO_1861 (O_1861,N_19751,N_19893);
or UO_1862 (O_1862,N_19911,N_19824);
xor UO_1863 (O_1863,N_19811,N_19771);
and UO_1864 (O_1864,N_19793,N_19918);
or UO_1865 (O_1865,N_19911,N_19948);
xor UO_1866 (O_1866,N_19669,N_19822);
nor UO_1867 (O_1867,N_19702,N_19815);
nand UO_1868 (O_1868,N_19838,N_19774);
xor UO_1869 (O_1869,N_19620,N_19537);
nor UO_1870 (O_1870,N_19754,N_19515);
or UO_1871 (O_1871,N_19613,N_19539);
and UO_1872 (O_1872,N_19722,N_19789);
or UO_1873 (O_1873,N_19505,N_19598);
nand UO_1874 (O_1874,N_19939,N_19642);
xnor UO_1875 (O_1875,N_19553,N_19908);
and UO_1876 (O_1876,N_19512,N_19504);
and UO_1877 (O_1877,N_19918,N_19699);
and UO_1878 (O_1878,N_19934,N_19640);
nand UO_1879 (O_1879,N_19822,N_19689);
nor UO_1880 (O_1880,N_19918,N_19709);
nor UO_1881 (O_1881,N_19805,N_19730);
and UO_1882 (O_1882,N_19917,N_19546);
nand UO_1883 (O_1883,N_19582,N_19687);
nand UO_1884 (O_1884,N_19665,N_19743);
xor UO_1885 (O_1885,N_19623,N_19943);
nand UO_1886 (O_1886,N_19752,N_19624);
nor UO_1887 (O_1887,N_19663,N_19810);
nor UO_1888 (O_1888,N_19595,N_19854);
xnor UO_1889 (O_1889,N_19532,N_19835);
nor UO_1890 (O_1890,N_19887,N_19837);
xor UO_1891 (O_1891,N_19943,N_19626);
nor UO_1892 (O_1892,N_19769,N_19771);
or UO_1893 (O_1893,N_19766,N_19818);
xor UO_1894 (O_1894,N_19533,N_19839);
nor UO_1895 (O_1895,N_19871,N_19821);
and UO_1896 (O_1896,N_19753,N_19844);
and UO_1897 (O_1897,N_19702,N_19994);
nor UO_1898 (O_1898,N_19616,N_19506);
and UO_1899 (O_1899,N_19703,N_19536);
and UO_1900 (O_1900,N_19619,N_19527);
nor UO_1901 (O_1901,N_19715,N_19570);
and UO_1902 (O_1902,N_19544,N_19679);
nor UO_1903 (O_1903,N_19519,N_19948);
xnor UO_1904 (O_1904,N_19905,N_19668);
and UO_1905 (O_1905,N_19696,N_19524);
and UO_1906 (O_1906,N_19789,N_19910);
and UO_1907 (O_1907,N_19977,N_19505);
nor UO_1908 (O_1908,N_19875,N_19642);
nand UO_1909 (O_1909,N_19858,N_19919);
and UO_1910 (O_1910,N_19942,N_19880);
nand UO_1911 (O_1911,N_19755,N_19612);
or UO_1912 (O_1912,N_19512,N_19500);
nand UO_1913 (O_1913,N_19729,N_19909);
nor UO_1914 (O_1914,N_19572,N_19729);
nor UO_1915 (O_1915,N_19811,N_19561);
and UO_1916 (O_1916,N_19560,N_19995);
nor UO_1917 (O_1917,N_19617,N_19989);
xnor UO_1918 (O_1918,N_19675,N_19882);
nor UO_1919 (O_1919,N_19695,N_19938);
and UO_1920 (O_1920,N_19735,N_19803);
or UO_1921 (O_1921,N_19655,N_19615);
nand UO_1922 (O_1922,N_19524,N_19731);
nor UO_1923 (O_1923,N_19746,N_19613);
and UO_1924 (O_1924,N_19981,N_19557);
or UO_1925 (O_1925,N_19540,N_19657);
nor UO_1926 (O_1926,N_19849,N_19884);
or UO_1927 (O_1927,N_19549,N_19914);
xnor UO_1928 (O_1928,N_19915,N_19664);
nor UO_1929 (O_1929,N_19734,N_19792);
and UO_1930 (O_1930,N_19610,N_19727);
nor UO_1931 (O_1931,N_19778,N_19557);
xnor UO_1932 (O_1932,N_19681,N_19906);
and UO_1933 (O_1933,N_19782,N_19947);
xnor UO_1934 (O_1934,N_19503,N_19711);
or UO_1935 (O_1935,N_19701,N_19849);
xor UO_1936 (O_1936,N_19752,N_19891);
and UO_1937 (O_1937,N_19968,N_19799);
or UO_1938 (O_1938,N_19730,N_19599);
xor UO_1939 (O_1939,N_19553,N_19895);
xor UO_1940 (O_1940,N_19992,N_19799);
or UO_1941 (O_1941,N_19914,N_19522);
nand UO_1942 (O_1942,N_19973,N_19744);
and UO_1943 (O_1943,N_19853,N_19673);
xnor UO_1944 (O_1944,N_19524,N_19670);
and UO_1945 (O_1945,N_19924,N_19626);
nor UO_1946 (O_1946,N_19656,N_19988);
nor UO_1947 (O_1947,N_19923,N_19723);
xnor UO_1948 (O_1948,N_19855,N_19616);
xnor UO_1949 (O_1949,N_19605,N_19853);
and UO_1950 (O_1950,N_19503,N_19538);
or UO_1951 (O_1951,N_19744,N_19592);
and UO_1952 (O_1952,N_19762,N_19792);
xor UO_1953 (O_1953,N_19883,N_19726);
or UO_1954 (O_1954,N_19717,N_19953);
or UO_1955 (O_1955,N_19772,N_19577);
nand UO_1956 (O_1956,N_19544,N_19973);
xor UO_1957 (O_1957,N_19712,N_19768);
nor UO_1958 (O_1958,N_19775,N_19896);
or UO_1959 (O_1959,N_19659,N_19754);
nand UO_1960 (O_1960,N_19542,N_19667);
or UO_1961 (O_1961,N_19578,N_19586);
nand UO_1962 (O_1962,N_19908,N_19699);
or UO_1963 (O_1963,N_19918,N_19964);
nand UO_1964 (O_1964,N_19868,N_19862);
or UO_1965 (O_1965,N_19691,N_19668);
or UO_1966 (O_1966,N_19863,N_19693);
nor UO_1967 (O_1967,N_19863,N_19874);
nand UO_1968 (O_1968,N_19516,N_19919);
and UO_1969 (O_1969,N_19824,N_19703);
nand UO_1970 (O_1970,N_19613,N_19685);
nand UO_1971 (O_1971,N_19801,N_19670);
or UO_1972 (O_1972,N_19619,N_19748);
nand UO_1973 (O_1973,N_19853,N_19727);
nor UO_1974 (O_1974,N_19659,N_19555);
or UO_1975 (O_1975,N_19720,N_19904);
and UO_1976 (O_1976,N_19598,N_19984);
or UO_1977 (O_1977,N_19952,N_19684);
or UO_1978 (O_1978,N_19508,N_19815);
or UO_1979 (O_1979,N_19811,N_19759);
xor UO_1980 (O_1980,N_19589,N_19861);
xnor UO_1981 (O_1981,N_19949,N_19802);
xnor UO_1982 (O_1982,N_19511,N_19832);
nor UO_1983 (O_1983,N_19802,N_19890);
or UO_1984 (O_1984,N_19579,N_19807);
or UO_1985 (O_1985,N_19840,N_19891);
nand UO_1986 (O_1986,N_19855,N_19748);
or UO_1987 (O_1987,N_19903,N_19861);
or UO_1988 (O_1988,N_19916,N_19890);
nand UO_1989 (O_1989,N_19507,N_19625);
or UO_1990 (O_1990,N_19559,N_19735);
xor UO_1991 (O_1991,N_19872,N_19864);
nand UO_1992 (O_1992,N_19949,N_19799);
nor UO_1993 (O_1993,N_19859,N_19758);
nor UO_1994 (O_1994,N_19646,N_19730);
nand UO_1995 (O_1995,N_19519,N_19521);
xor UO_1996 (O_1996,N_19897,N_19917);
nor UO_1997 (O_1997,N_19563,N_19916);
nor UO_1998 (O_1998,N_19680,N_19767);
or UO_1999 (O_1999,N_19924,N_19989);
xnor UO_2000 (O_2000,N_19729,N_19993);
xnor UO_2001 (O_2001,N_19575,N_19802);
or UO_2002 (O_2002,N_19716,N_19778);
and UO_2003 (O_2003,N_19620,N_19558);
xor UO_2004 (O_2004,N_19820,N_19759);
or UO_2005 (O_2005,N_19921,N_19680);
nand UO_2006 (O_2006,N_19510,N_19705);
xnor UO_2007 (O_2007,N_19818,N_19581);
and UO_2008 (O_2008,N_19821,N_19509);
nand UO_2009 (O_2009,N_19622,N_19639);
and UO_2010 (O_2010,N_19918,N_19707);
or UO_2011 (O_2011,N_19857,N_19856);
and UO_2012 (O_2012,N_19638,N_19519);
xor UO_2013 (O_2013,N_19977,N_19949);
xor UO_2014 (O_2014,N_19812,N_19894);
or UO_2015 (O_2015,N_19807,N_19963);
nor UO_2016 (O_2016,N_19569,N_19907);
or UO_2017 (O_2017,N_19559,N_19540);
nor UO_2018 (O_2018,N_19866,N_19596);
nand UO_2019 (O_2019,N_19880,N_19782);
xnor UO_2020 (O_2020,N_19790,N_19660);
or UO_2021 (O_2021,N_19521,N_19977);
nor UO_2022 (O_2022,N_19834,N_19686);
and UO_2023 (O_2023,N_19570,N_19830);
or UO_2024 (O_2024,N_19896,N_19825);
or UO_2025 (O_2025,N_19693,N_19516);
and UO_2026 (O_2026,N_19716,N_19623);
or UO_2027 (O_2027,N_19982,N_19967);
and UO_2028 (O_2028,N_19914,N_19873);
xnor UO_2029 (O_2029,N_19565,N_19990);
and UO_2030 (O_2030,N_19878,N_19961);
and UO_2031 (O_2031,N_19543,N_19976);
xor UO_2032 (O_2032,N_19814,N_19504);
or UO_2033 (O_2033,N_19865,N_19671);
nand UO_2034 (O_2034,N_19682,N_19673);
xor UO_2035 (O_2035,N_19575,N_19572);
and UO_2036 (O_2036,N_19667,N_19974);
nor UO_2037 (O_2037,N_19963,N_19578);
and UO_2038 (O_2038,N_19824,N_19778);
nor UO_2039 (O_2039,N_19916,N_19851);
and UO_2040 (O_2040,N_19572,N_19542);
or UO_2041 (O_2041,N_19839,N_19639);
xor UO_2042 (O_2042,N_19608,N_19752);
xnor UO_2043 (O_2043,N_19835,N_19699);
nand UO_2044 (O_2044,N_19620,N_19720);
xor UO_2045 (O_2045,N_19899,N_19730);
nor UO_2046 (O_2046,N_19692,N_19840);
xnor UO_2047 (O_2047,N_19628,N_19797);
and UO_2048 (O_2048,N_19593,N_19884);
nor UO_2049 (O_2049,N_19841,N_19738);
and UO_2050 (O_2050,N_19978,N_19656);
or UO_2051 (O_2051,N_19913,N_19773);
and UO_2052 (O_2052,N_19764,N_19831);
and UO_2053 (O_2053,N_19866,N_19700);
nor UO_2054 (O_2054,N_19932,N_19969);
nand UO_2055 (O_2055,N_19951,N_19643);
or UO_2056 (O_2056,N_19671,N_19524);
xor UO_2057 (O_2057,N_19843,N_19621);
nor UO_2058 (O_2058,N_19796,N_19673);
xnor UO_2059 (O_2059,N_19778,N_19506);
or UO_2060 (O_2060,N_19764,N_19816);
or UO_2061 (O_2061,N_19995,N_19569);
or UO_2062 (O_2062,N_19617,N_19741);
nor UO_2063 (O_2063,N_19884,N_19823);
or UO_2064 (O_2064,N_19733,N_19746);
or UO_2065 (O_2065,N_19852,N_19665);
or UO_2066 (O_2066,N_19993,N_19848);
nand UO_2067 (O_2067,N_19580,N_19797);
and UO_2068 (O_2068,N_19862,N_19996);
xnor UO_2069 (O_2069,N_19837,N_19927);
and UO_2070 (O_2070,N_19524,N_19718);
or UO_2071 (O_2071,N_19982,N_19927);
xnor UO_2072 (O_2072,N_19800,N_19665);
nand UO_2073 (O_2073,N_19691,N_19575);
and UO_2074 (O_2074,N_19779,N_19679);
or UO_2075 (O_2075,N_19940,N_19691);
nand UO_2076 (O_2076,N_19748,N_19985);
nor UO_2077 (O_2077,N_19911,N_19549);
or UO_2078 (O_2078,N_19651,N_19580);
xnor UO_2079 (O_2079,N_19609,N_19642);
nand UO_2080 (O_2080,N_19621,N_19725);
or UO_2081 (O_2081,N_19826,N_19569);
xor UO_2082 (O_2082,N_19961,N_19806);
and UO_2083 (O_2083,N_19943,N_19851);
nand UO_2084 (O_2084,N_19794,N_19729);
xnor UO_2085 (O_2085,N_19979,N_19848);
or UO_2086 (O_2086,N_19837,N_19948);
nor UO_2087 (O_2087,N_19610,N_19546);
nand UO_2088 (O_2088,N_19570,N_19918);
nor UO_2089 (O_2089,N_19561,N_19813);
nor UO_2090 (O_2090,N_19997,N_19642);
nor UO_2091 (O_2091,N_19581,N_19784);
and UO_2092 (O_2092,N_19805,N_19696);
or UO_2093 (O_2093,N_19851,N_19560);
xnor UO_2094 (O_2094,N_19658,N_19576);
nand UO_2095 (O_2095,N_19694,N_19787);
and UO_2096 (O_2096,N_19641,N_19876);
xor UO_2097 (O_2097,N_19911,N_19790);
and UO_2098 (O_2098,N_19653,N_19814);
or UO_2099 (O_2099,N_19839,N_19766);
and UO_2100 (O_2100,N_19711,N_19895);
xor UO_2101 (O_2101,N_19993,N_19865);
and UO_2102 (O_2102,N_19853,N_19910);
nor UO_2103 (O_2103,N_19910,N_19724);
and UO_2104 (O_2104,N_19722,N_19744);
nand UO_2105 (O_2105,N_19672,N_19661);
or UO_2106 (O_2106,N_19929,N_19694);
xnor UO_2107 (O_2107,N_19686,N_19982);
or UO_2108 (O_2108,N_19740,N_19678);
or UO_2109 (O_2109,N_19830,N_19583);
or UO_2110 (O_2110,N_19553,N_19551);
nand UO_2111 (O_2111,N_19752,N_19705);
or UO_2112 (O_2112,N_19623,N_19905);
xor UO_2113 (O_2113,N_19712,N_19607);
or UO_2114 (O_2114,N_19919,N_19936);
and UO_2115 (O_2115,N_19934,N_19721);
xor UO_2116 (O_2116,N_19715,N_19943);
nand UO_2117 (O_2117,N_19684,N_19556);
xnor UO_2118 (O_2118,N_19539,N_19783);
nand UO_2119 (O_2119,N_19951,N_19872);
xor UO_2120 (O_2120,N_19828,N_19881);
or UO_2121 (O_2121,N_19643,N_19536);
nor UO_2122 (O_2122,N_19660,N_19704);
nand UO_2123 (O_2123,N_19721,N_19675);
nand UO_2124 (O_2124,N_19727,N_19983);
nand UO_2125 (O_2125,N_19924,N_19972);
and UO_2126 (O_2126,N_19881,N_19898);
nand UO_2127 (O_2127,N_19835,N_19944);
and UO_2128 (O_2128,N_19954,N_19836);
nand UO_2129 (O_2129,N_19701,N_19510);
xnor UO_2130 (O_2130,N_19977,N_19942);
and UO_2131 (O_2131,N_19710,N_19828);
or UO_2132 (O_2132,N_19731,N_19709);
nand UO_2133 (O_2133,N_19527,N_19607);
xor UO_2134 (O_2134,N_19541,N_19842);
or UO_2135 (O_2135,N_19722,N_19583);
xnor UO_2136 (O_2136,N_19766,N_19668);
and UO_2137 (O_2137,N_19903,N_19510);
and UO_2138 (O_2138,N_19836,N_19912);
nand UO_2139 (O_2139,N_19899,N_19540);
or UO_2140 (O_2140,N_19974,N_19626);
nor UO_2141 (O_2141,N_19757,N_19817);
xor UO_2142 (O_2142,N_19945,N_19720);
nor UO_2143 (O_2143,N_19575,N_19895);
nor UO_2144 (O_2144,N_19736,N_19611);
nor UO_2145 (O_2145,N_19836,N_19926);
xnor UO_2146 (O_2146,N_19560,N_19555);
nand UO_2147 (O_2147,N_19649,N_19639);
xor UO_2148 (O_2148,N_19546,N_19974);
xnor UO_2149 (O_2149,N_19844,N_19700);
nor UO_2150 (O_2150,N_19807,N_19894);
xnor UO_2151 (O_2151,N_19710,N_19645);
or UO_2152 (O_2152,N_19755,N_19785);
xor UO_2153 (O_2153,N_19862,N_19979);
and UO_2154 (O_2154,N_19762,N_19639);
or UO_2155 (O_2155,N_19628,N_19651);
nor UO_2156 (O_2156,N_19656,N_19579);
and UO_2157 (O_2157,N_19691,N_19564);
xnor UO_2158 (O_2158,N_19677,N_19711);
nor UO_2159 (O_2159,N_19513,N_19601);
or UO_2160 (O_2160,N_19954,N_19968);
nand UO_2161 (O_2161,N_19692,N_19588);
or UO_2162 (O_2162,N_19864,N_19632);
or UO_2163 (O_2163,N_19623,N_19626);
nor UO_2164 (O_2164,N_19762,N_19918);
nand UO_2165 (O_2165,N_19759,N_19511);
nand UO_2166 (O_2166,N_19599,N_19968);
nor UO_2167 (O_2167,N_19915,N_19582);
and UO_2168 (O_2168,N_19750,N_19507);
nand UO_2169 (O_2169,N_19831,N_19699);
xnor UO_2170 (O_2170,N_19720,N_19897);
and UO_2171 (O_2171,N_19919,N_19737);
xor UO_2172 (O_2172,N_19889,N_19690);
nand UO_2173 (O_2173,N_19556,N_19825);
and UO_2174 (O_2174,N_19841,N_19860);
nand UO_2175 (O_2175,N_19540,N_19729);
nor UO_2176 (O_2176,N_19934,N_19843);
nand UO_2177 (O_2177,N_19769,N_19923);
nand UO_2178 (O_2178,N_19741,N_19592);
or UO_2179 (O_2179,N_19831,N_19585);
nand UO_2180 (O_2180,N_19778,N_19965);
and UO_2181 (O_2181,N_19780,N_19793);
or UO_2182 (O_2182,N_19950,N_19887);
nand UO_2183 (O_2183,N_19932,N_19822);
xor UO_2184 (O_2184,N_19866,N_19767);
nor UO_2185 (O_2185,N_19975,N_19812);
xnor UO_2186 (O_2186,N_19791,N_19627);
nand UO_2187 (O_2187,N_19593,N_19824);
xnor UO_2188 (O_2188,N_19517,N_19586);
nand UO_2189 (O_2189,N_19829,N_19567);
nor UO_2190 (O_2190,N_19587,N_19567);
xnor UO_2191 (O_2191,N_19964,N_19834);
or UO_2192 (O_2192,N_19592,N_19894);
nor UO_2193 (O_2193,N_19612,N_19838);
xnor UO_2194 (O_2194,N_19874,N_19891);
and UO_2195 (O_2195,N_19909,N_19740);
nand UO_2196 (O_2196,N_19810,N_19966);
and UO_2197 (O_2197,N_19801,N_19789);
nand UO_2198 (O_2198,N_19949,N_19752);
xor UO_2199 (O_2199,N_19623,N_19565);
nor UO_2200 (O_2200,N_19581,N_19808);
xnor UO_2201 (O_2201,N_19526,N_19622);
or UO_2202 (O_2202,N_19516,N_19796);
or UO_2203 (O_2203,N_19708,N_19543);
nor UO_2204 (O_2204,N_19913,N_19970);
nor UO_2205 (O_2205,N_19822,N_19687);
or UO_2206 (O_2206,N_19519,N_19764);
or UO_2207 (O_2207,N_19539,N_19557);
and UO_2208 (O_2208,N_19651,N_19880);
and UO_2209 (O_2209,N_19518,N_19773);
nor UO_2210 (O_2210,N_19869,N_19598);
and UO_2211 (O_2211,N_19854,N_19549);
nand UO_2212 (O_2212,N_19676,N_19537);
xnor UO_2213 (O_2213,N_19872,N_19807);
and UO_2214 (O_2214,N_19676,N_19700);
and UO_2215 (O_2215,N_19558,N_19824);
nor UO_2216 (O_2216,N_19619,N_19696);
xor UO_2217 (O_2217,N_19593,N_19746);
nor UO_2218 (O_2218,N_19725,N_19931);
nor UO_2219 (O_2219,N_19549,N_19658);
xor UO_2220 (O_2220,N_19740,N_19808);
nand UO_2221 (O_2221,N_19869,N_19921);
or UO_2222 (O_2222,N_19640,N_19983);
xnor UO_2223 (O_2223,N_19880,N_19503);
or UO_2224 (O_2224,N_19612,N_19761);
and UO_2225 (O_2225,N_19696,N_19852);
xor UO_2226 (O_2226,N_19540,N_19949);
xor UO_2227 (O_2227,N_19544,N_19669);
nor UO_2228 (O_2228,N_19729,N_19637);
or UO_2229 (O_2229,N_19553,N_19905);
and UO_2230 (O_2230,N_19970,N_19973);
or UO_2231 (O_2231,N_19835,N_19622);
nor UO_2232 (O_2232,N_19784,N_19809);
or UO_2233 (O_2233,N_19571,N_19910);
nand UO_2234 (O_2234,N_19583,N_19749);
nand UO_2235 (O_2235,N_19903,N_19599);
or UO_2236 (O_2236,N_19522,N_19706);
xor UO_2237 (O_2237,N_19529,N_19974);
nor UO_2238 (O_2238,N_19743,N_19697);
nand UO_2239 (O_2239,N_19517,N_19527);
and UO_2240 (O_2240,N_19745,N_19978);
nor UO_2241 (O_2241,N_19698,N_19606);
xnor UO_2242 (O_2242,N_19737,N_19986);
or UO_2243 (O_2243,N_19567,N_19622);
and UO_2244 (O_2244,N_19888,N_19890);
nor UO_2245 (O_2245,N_19583,N_19891);
xnor UO_2246 (O_2246,N_19532,N_19735);
nand UO_2247 (O_2247,N_19891,N_19977);
nand UO_2248 (O_2248,N_19931,N_19888);
and UO_2249 (O_2249,N_19827,N_19967);
nand UO_2250 (O_2250,N_19933,N_19614);
nand UO_2251 (O_2251,N_19926,N_19684);
nor UO_2252 (O_2252,N_19605,N_19990);
nand UO_2253 (O_2253,N_19728,N_19616);
and UO_2254 (O_2254,N_19831,N_19687);
and UO_2255 (O_2255,N_19675,N_19566);
and UO_2256 (O_2256,N_19976,N_19686);
and UO_2257 (O_2257,N_19945,N_19564);
nand UO_2258 (O_2258,N_19831,N_19677);
and UO_2259 (O_2259,N_19954,N_19666);
and UO_2260 (O_2260,N_19866,N_19560);
nand UO_2261 (O_2261,N_19933,N_19958);
nor UO_2262 (O_2262,N_19953,N_19754);
nand UO_2263 (O_2263,N_19894,N_19972);
and UO_2264 (O_2264,N_19859,N_19844);
or UO_2265 (O_2265,N_19860,N_19605);
nand UO_2266 (O_2266,N_19525,N_19740);
and UO_2267 (O_2267,N_19827,N_19542);
nand UO_2268 (O_2268,N_19805,N_19628);
and UO_2269 (O_2269,N_19684,N_19633);
xnor UO_2270 (O_2270,N_19664,N_19967);
nor UO_2271 (O_2271,N_19685,N_19960);
and UO_2272 (O_2272,N_19680,N_19545);
xnor UO_2273 (O_2273,N_19897,N_19851);
nand UO_2274 (O_2274,N_19954,N_19608);
and UO_2275 (O_2275,N_19865,N_19639);
and UO_2276 (O_2276,N_19550,N_19877);
and UO_2277 (O_2277,N_19911,N_19739);
nand UO_2278 (O_2278,N_19926,N_19557);
nand UO_2279 (O_2279,N_19997,N_19717);
nand UO_2280 (O_2280,N_19857,N_19564);
nor UO_2281 (O_2281,N_19948,N_19758);
nand UO_2282 (O_2282,N_19625,N_19803);
or UO_2283 (O_2283,N_19646,N_19709);
nand UO_2284 (O_2284,N_19979,N_19774);
nand UO_2285 (O_2285,N_19544,N_19730);
and UO_2286 (O_2286,N_19633,N_19617);
nand UO_2287 (O_2287,N_19728,N_19565);
or UO_2288 (O_2288,N_19852,N_19904);
nor UO_2289 (O_2289,N_19796,N_19820);
xnor UO_2290 (O_2290,N_19965,N_19966);
nand UO_2291 (O_2291,N_19728,N_19880);
nor UO_2292 (O_2292,N_19534,N_19567);
xnor UO_2293 (O_2293,N_19806,N_19866);
or UO_2294 (O_2294,N_19664,N_19841);
and UO_2295 (O_2295,N_19583,N_19693);
and UO_2296 (O_2296,N_19903,N_19612);
or UO_2297 (O_2297,N_19577,N_19521);
xnor UO_2298 (O_2298,N_19859,N_19589);
nand UO_2299 (O_2299,N_19800,N_19854);
nor UO_2300 (O_2300,N_19575,N_19852);
nand UO_2301 (O_2301,N_19820,N_19652);
xnor UO_2302 (O_2302,N_19609,N_19546);
xnor UO_2303 (O_2303,N_19898,N_19622);
and UO_2304 (O_2304,N_19935,N_19608);
or UO_2305 (O_2305,N_19992,N_19714);
nor UO_2306 (O_2306,N_19557,N_19823);
xnor UO_2307 (O_2307,N_19848,N_19696);
nor UO_2308 (O_2308,N_19683,N_19804);
and UO_2309 (O_2309,N_19852,N_19972);
xnor UO_2310 (O_2310,N_19932,N_19883);
nor UO_2311 (O_2311,N_19848,N_19892);
and UO_2312 (O_2312,N_19578,N_19863);
xor UO_2313 (O_2313,N_19579,N_19724);
and UO_2314 (O_2314,N_19923,N_19666);
nand UO_2315 (O_2315,N_19983,N_19504);
xor UO_2316 (O_2316,N_19970,N_19723);
or UO_2317 (O_2317,N_19638,N_19704);
or UO_2318 (O_2318,N_19933,N_19818);
or UO_2319 (O_2319,N_19979,N_19530);
or UO_2320 (O_2320,N_19794,N_19514);
nor UO_2321 (O_2321,N_19543,N_19667);
or UO_2322 (O_2322,N_19858,N_19547);
nor UO_2323 (O_2323,N_19704,N_19587);
nor UO_2324 (O_2324,N_19820,N_19595);
nor UO_2325 (O_2325,N_19919,N_19665);
and UO_2326 (O_2326,N_19675,N_19548);
or UO_2327 (O_2327,N_19696,N_19889);
nand UO_2328 (O_2328,N_19639,N_19559);
and UO_2329 (O_2329,N_19866,N_19692);
nand UO_2330 (O_2330,N_19657,N_19879);
nand UO_2331 (O_2331,N_19502,N_19860);
xor UO_2332 (O_2332,N_19657,N_19714);
and UO_2333 (O_2333,N_19720,N_19668);
and UO_2334 (O_2334,N_19792,N_19775);
xor UO_2335 (O_2335,N_19526,N_19992);
nor UO_2336 (O_2336,N_19759,N_19786);
or UO_2337 (O_2337,N_19754,N_19821);
nand UO_2338 (O_2338,N_19608,N_19611);
xnor UO_2339 (O_2339,N_19761,N_19878);
nand UO_2340 (O_2340,N_19669,N_19943);
and UO_2341 (O_2341,N_19563,N_19881);
nand UO_2342 (O_2342,N_19609,N_19778);
nor UO_2343 (O_2343,N_19880,N_19913);
nand UO_2344 (O_2344,N_19829,N_19852);
xnor UO_2345 (O_2345,N_19530,N_19994);
and UO_2346 (O_2346,N_19789,N_19797);
xor UO_2347 (O_2347,N_19989,N_19999);
nand UO_2348 (O_2348,N_19525,N_19530);
xor UO_2349 (O_2349,N_19689,N_19668);
nand UO_2350 (O_2350,N_19764,N_19807);
nor UO_2351 (O_2351,N_19971,N_19827);
and UO_2352 (O_2352,N_19869,N_19833);
xor UO_2353 (O_2353,N_19574,N_19517);
or UO_2354 (O_2354,N_19735,N_19855);
nor UO_2355 (O_2355,N_19823,N_19922);
or UO_2356 (O_2356,N_19668,N_19773);
nand UO_2357 (O_2357,N_19826,N_19581);
or UO_2358 (O_2358,N_19526,N_19977);
xor UO_2359 (O_2359,N_19916,N_19940);
and UO_2360 (O_2360,N_19848,N_19606);
and UO_2361 (O_2361,N_19808,N_19522);
nand UO_2362 (O_2362,N_19675,N_19594);
nand UO_2363 (O_2363,N_19734,N_19778);
and UO_2364 (O_2364,N_19725,N_19967);
xnor UO_2365 (O_2365,N_19516,N_19807);
nor UO_2366 (O_2366,N_19710,N_19534);
nand UO_2367 (O_2367,N_19611,N_19542);
nand UO_2368 (O_2368,N_19587,N_19806);
and UO_2369 (O_2369,N_19641,N_19932);
nand UO_2370 (O_2370,N_19610,N_19617);
or UO_2371 (O_2371,N_19781,N_19787);
nor UO_2372 (O_2372,N_19971,N_19866);
or UO_2373 (O_2373,N_19890,N_19733);
nor UO_2374 (O_2374,N_19534,N_19753);
or UO_2375 (O_2375,N_19589,N_19836);
xnor UO_2376 (O_2376,N_19944,N_19776);
nand UO_2377 (O_2377,N_19745,N_19726);
nor UO_2378 (O_2378,N_19570,N_19883);
and UO_2379 (O_2379,N_19708,N_19798);
xnor UO_2380 (O_2380,N_19679,N_19840);
nor UO_2381 (O_2381,N_19976,N_19767);
nor UO_2382 (O_2382,N_19924,N_19942);
and UO_2383 (O_2383,N_19553,N_19533);
nand UO_2384 (O_2384,N_19834,N_19976);
nand UO_2385 (O_2385,N_19510,N_19966);
or UO_2386 (O_2386,N_19887,N_19589);
or UO_2387 (O_2387,N_19637,N_19888);
nand UO_2388 (O_2388,N_19624,N_19758);
and UO_2389 (O_2389,N_19580,N_19836);
and UO_2390 (O_2390,N_19844,N_19595);
xnor UO_2391 (O_2391,N_19644,N_19937);
nand UO_2392 (O_2392,N_19933,N_19819);
and UO_2393 (O_2393,N_19667,N_19606);
and UO_2394 (O_2394,N_19960,N_19638);
xor UO_2395 (O_2395,N_19884,N_19974);
nor UO_2396 (O_2396,N_19511,N_19807);
nand UO_2397 (O_2397,N_19879,N_19585);
nand UO_2398 (O_2398,N_19548,N_19993);
nor UO_2399 (O_2399,N_19617,N_19955);
and UO_2400 (O_2400,N_19705,N_19627);
nand UO_2401 (O_2401,N_19894,N_19779);
nor UO_2402 (O_2402,N_19726,N_19811);
xor UO_2403 (O_2403,N_19766,N_19911);
nand UO_2404 (O_2404,N_19512,N_19913);
or UO_2405 (O_2405,N_19693,N_19991);
nand UO_2406 (O_2406,N_19735,N_19980);
or UO_2407 (O_2407,N_19549,N_19645);
or UO_2408 (O_2408,N_19982,N_19558);
and UO_2409 (O_2409,N_19643,N_19674);
xor UO_2410 (O_2410,N_19592,N_19526);
and UO_2411 (O_2411,N_19763,N_19622);
nor UO_2412 (O_2412,N_19766,N_19894);
or UO_2413 (O_2413,N_19904,N_19587);
or UO_2414 (O_2414,N_19942,N_19712);
nor UO_2415 (O_2415,N_19798,N_19596);
xor UO_2416 (O_2416,N_19693,N_19711);
and UO_2417 (O_2417,N_19942,N_19543);
xnor UO_2418 (O_2418,N_19524,N_19582);
nor UO_2419 (O_2419,N_19741,N_19768);
nand UO_2420 (O_2420,N_19988,N_19699);
xor UO_2421 (O_2421,N_19754,N_19737);
or UO_2422 (O_2422,N_19599,N_19572);
and UO_2423 (O_2423,N_19874,N_19974);
nand UO_2424 (O_2424,N_19869,N_19754);
nor UO_2425 (O_2425,N_19864,N_19906);
and UO_2426 (O_2426,N_19517,N_19910);
or UO_2427 (O_2427,N_19536,N_19537);
and UO_2428 (O_2428,N_19800,N_19504);
nor UO_2429 (O_2429,N_19788,N_19553);
nor UO_2430 (O_2430,N_19729,N_19820);
and UO_2431 (O_2431,N_19544,N_19960);
nand UO_2432 (O_2432,N_19756,N_19782);
and UO_2433 (O_2433,N_19695,N_19846);
or UO_2434 (O_2434,N_19717,N_19748);
nand UO_2435 (O_2435,N_19651,N_19650);
and UO_2436 (O_2436,N_19814,N_19524);
and UO_2437 (O_2437,N_19972,N_19962);
and UO_2438 (O_2438,N_19964,N_19648);
or UO_2439 (O_2439,N_19976,N_19597);
nor UO_2440 (O_2440,N_19570,N_19650);
and UO_2441 (O_2441,N_19898,N_19895);
xnor UO_2442 (O_2442,N_19602,N_19599);
xnor UO_2443 (O_2443,N_19508,N_19893);
xor UO_2444 (O_2444,N_19537,N_19955);
xor UO_2445 (O_2445,N_19707,N_19888);
nand UO_2446 (O_2446,N_19690,N_19797);
or UO_2447 (O_2447,N_19784,N_19594);
nor UO_2448 (O_2448,N_19753,N_19665);
xnor UO_2449 (O_2449,N_19568,N_19777);
xor UO_2450 (O_2450,N_19829,N_19588);
nor UO_2451 (O_2451,N_19881,N_19709);
xor UO_2452 (O_2452,N_19878,N_19546);
nor UO_2453 (O_2453,N_19539,N_19705);
nor UO_2454 (O_2454,N_19570,N_19530);
nand UO_2455 (O_2455,N_19719,N_19561);
and UO_2456 (O_2456,N_19813,N_19857);
and UO_2457 (O_2457,N_19617,N_19996);
xnor UO_2458 (O_2458,N_19860,N_19573);
xor UO_2459 (O_2459,N_19703,N_19933);
nor UO_2460 (O_2460,N_19898,N_19738);
and UO_2461 (O_2461,N_19532,N_19724);
and UO_2462 (O_2462,N_19925,N_19668);
and UO_2463 (O_2463,N_19703,N_19520);
or UO_2464 (O_2464,N_19863,N_19669);
and UO_2465 (O_2465,N_19622,N_19599);
xnor UO_2466 (O_2466,N_19936,N_19609);
xnor UO_2467 (O_2467,N_19516,N_19839);
nor UO_2468 (O_2468,N_19775,N_19862);
and UO_2469 (O_2469,N_19881,N_19967);
or UO_2470 (O_2470,N_19564,N_19748);
nor UO_2471 (O_2471,N_19979,N_19918);
and UO_2472 (O_2472,N_19682,N_19665);
nor UO_2473 (O_2473,N_19777,N_19724);
xnor UO_2474 (O_2474,N_19888,N_19964);
or UO_2475 (O_2475,N_19594,N_19805);
xnor UO_2476 (O_2476,N_19617,N_19831);
nand UO_2477 (O_2477,N_19762,N_19729);
xor UO_2478 (O_2478,N_19995,N_19724);
and UO_2479 (O_2479,N_19859,N_19725);
and UO_2480 (O_2480,N_19831,N_19822);
or UO_2481 (O_2481,N_19787,N_19684);
nor UO_2482 (O_2482,N_19574,N_19765);
xor UO_2483 (O_2483,N_19948,N_19515);
and UO_2484 (O_2484,N_19895,N_19516);
and UO_2485 (O_2485,N_19715,N_19990);
nor UO_2486 (O_2486,N_19678,N_19565);
or UO_2487 (O_2487,N_19870,N_19576);
or UO_2488 (O_2488,N_19652,N_19738);
or UO_2489 (O_2489,N_19620,N_19825);
nor UO_2490 (O_2490,N_19948,N_19999);
nor UO_2491 (O_2491,N_19982,N_19827);
xor UO_2492 (O_2492,N_19549,N_19598);
nor UO_2493 (O_2493,N_19692,N_19935);
and UO_2494 (O_2494,N_19639,N_19573);
nand UO_2495 (O_2495,N_19580,N_19765);
xor UO_2496 (O_2496,N_19627,N_19823);
nor UO_2497 (O_2497,N_19601,N_19809);
nand UO_2498 (O_2498,N_19902,N_19729);
and UO_2499 (O_2499,N_19980,N_19608);
endmodule