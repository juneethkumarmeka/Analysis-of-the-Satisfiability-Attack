module basic_1500_15000_2000_15_levels_5xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nor U0 (N_0,In_734,In_432);
nor U1 (N_1,In_1169,In_879);
and U2 (N_2,In_990,In_860);
or U3 (N_3,In_1304,In_788);
nor U4 (N_4,In_1147,In_719);
nor U5 (N_5,In_1356,In_870);
xor U6 (N_6,In_1486,In_657);
nand U7 (N_7,In_101,In_1242);
nor U8 (N_8,In_341,In_762);
or U9 (N_9,In_1440,In_1129);
xnor U10 (N_10,In_371,In_764);
nor U11 (N_11,In_79,In_1205);
and U12 (N_12,In_752,In_1291);
or U13 (N_13,In_7,In_34);
nand U14 (N_14,In_386,In_1327);
and U15 (N_15,In_785,In_115);
xnor U16 (N_16,In_219,In_759);
xor U17 (N_17,In_302,In_1365);
nor U18 (N_18,In_464,In_1095);
nand U19 (N_19,In_201,In_1379);
or U20 (N_20,In_1284,In_455);
or U21 (N_21,In_425,In_512);
nor U22 (N_22,In_218,In_861);
nor U23 (N_23,In_520,In_1010);
xnor U24 (N_24,In_1191,In_1167);
nand U25 (N_25,In_1093,In_619);
nor U26 (N_26,In_924,In_296);
nand U27 (N_27,In_1250,In_775);
or U28 (N_28,In_210,In_435);
nor U29 (N_29,In_595,In_1405);
nand U30 (N_30,In_1233,In_1056);
nor U31 (N_31,In_636,In_1197);
or U32 (N_32,In_703,In_150);
or U33 (N_33,In_780,In_103);
or U34 (N_34,In_633,In_888);
and U35 (N_35,In_1319,In_890);
and U36 (N_36,In_1177,In_846);
or U37 (N_37,In_1376,In_1252);
or U38 (N_38,In_1413,In_173);
nor U39 (N_39,In_365,In_814);
and U40 (N_40,In_1288,In_1316);
xnor U41 (N_41,In_285,In_1151);
nor U42 (N_42,In_1354,In_1052);
nor U43 (N_43,In_1420,In_666);
nand U44 (N_44,In_1270,In_1450);
nand U45 (N_45,In_739,In_274);
nand U46 (N_46,In_549,In_100);
and U47 (N_47,In_899,In_1339);
and U48 (N_48,In_1078,In_504);
or U49 (N_49,In_248,In_68);
and U50 (N_50,In_685,In_1298);
or U51 (N_51,In_278,In_109);
and U52 (N_52,In_1211,In_774);
nor U53 (N_53,In_1436,In_1200);
or U54 (N_54,In_1439,In_337);
and U55 (N_55,In_1331,In_1328);
or U56 (N_56,In_1258,In_1320);
and U57 (N_57,In_1466,In_111);
or U58 (N_58,In_909,In_1255);
nor U59 (N_59,In_1238,In_208);
nand U60 (N_60,In_715,In_1481);
or U61 (N_61,In_184,In_1144);
nor U62 (N_62,In_1276,In_1231);
nand U63 (N_63,In_187,In_185);
nand U64 (N_64,In_997,In_445);
nand U65 (N_65,In_798,In_689);
nor U66 (N_66,In_982,In_236);
and U67 (N_67,In_1220,In_475);
and U68 (N_68,In_1476,In_229);
and U69 (N_69,In_427,In_704);
or U70 (N_70,In_713,In_894);
nor U71 (N_71,In_473,In_20);
xnor U72 (N_72,In_1090,In_367);
nand U73 (N_73,In_233,In_1071);
nor U74 (N_74,In_1047,In_695);
or U75 (N_75,In_63,In_148);
xor U76 (N_76,In_1221,In_1077);
nand U77 (N_77,In_738,In_571);
and U78 (N_78,In_1215,In_1092);
nor U79 (N_79,In_777,In_1337);
nor U80 (N_80,In_787,In_1059);
or U81 (N_81,In_126,In_378);
nand U82 (N_82,In_1117,In_947);
and U83 (N_83,In_1487,In_712);
or U84 (N_84,In_1108,In_1229);
nand U85 (N_85,In_950,In_962);
nor U86 (N_86,In_1335,In_1391);
or U87 (N_87,In_487,In_154);
or U88 (N_88,In_923,In_559);
xnor U89 (N_89,In_1037,In_1243);
nor U90 (N_90,In_615,In_272);
nor U91 (N_91,In_1332,In_585);
or U92 (N_92,In_682,In_1027);
nor U93 (N_93,In_1441,In_1290);
nor U94 (N_94,In_882,In_8);
xnor U95 (N_95,In_802,In_1397);
or U96 (N_96,In_576,In_749);
nor U97 (N_97,In_1455,In_1380);
and U98 (N_98,In_656,In_744);
nor U99 (N_99,In_467,In_1271);
xor U100 (N_100,In_1067,In_887);
nor U101 (N_101,In_963,In_240);
nor U102 (N_102,In_211,In_683);
nor U103 (N_103,In_1457,In_188);
xor U104 (N_104,In_472,In_304);
nor U105 (N_105,In_756,In_391);
nand U106 (N_106,In_1493,In_136);
nand U107 (N_107,In_1359,In_996);
nor U108 (N_108,In_877,In_723);
nand U109 (N_109,In_1370,In_1360);
xnor U110 (N_110,In_1425,In_90);
xnor U111 (N_111,In_80,In_515);
nor U112 (N_112,In_911,In_938);
and U113 (N_113,In_1187,In_493);
or U114 (N_114,In_1065,In_415);
nand U115 (N_115,In_369,In_1105);
nand U116 (N_116,In_1002,In_419);
nand U117 (N_117,In_99,In_740);
nand U118 (N_118,In_1015,In_376);
nor U119 (N_119,In_338,In_1388);
nor U120 (N_120,In_1449,In_399);
or U121 (N_121,In_1334,In_937);
nor U122 (N_122,In_755,In_70);
and U123 (N_123,In_36,In_157);
and U124 (N_124,In_776,In_38);
nand U125 (N_125,In_838,In_805);
and U126 (N_126,In_466,In_1196);
or U127 (N_127,In_929,In_773);
nor U128 (N_128,In_231,In_255);
nor U129 (N_129,In_339,In_429);
or U130 (N_130,In_541,In_1340);
nand U131 (N_131,In_1404,In_1333);
or U132 (N_132,In_352,In_1305);
or U133 (N_133,In_885,In_468);
nand U134 (N_134,In_209,In_1091);
or U135 (N_135,In_1463,In_556);
and U136 (N_136,In_494,In_514);
nand U137 (N_137,In_266,In_624);
and U138 (N_138,In_58,In_1294);
xor U139 (N_139,In_1350,In_907);
or U140 (N_140,In_1412,In_867);
and U141 (N_141,In_1377,In_1495);
and U142 (N_142,In_603,In_1249);
nor U143 (N_143,In_364,In_293);
nor U144 (N_144,In_292,In_344);
or U145 (N_145,In_360,In_460);
and U146 (N_146,In_592,In_193);
and U147 (N_147,In_1175,In_315);
nand U148 (N_148,In_1366,In_1207);
xor U149 (N_149,In_841,In_134);
nor U150 (N_150,In_417,In_324);
nand U151 (N_151,In_1223,In_1313);
xnor U152 (N_152,In_416,In_599);
nor U153 (N_153,In_1121,In_359);
nor U154 (N_154,In_954,In_825);
nor U155 (N_155,In_469,In_1087);
nand U156 (N_156,In_1003,In_202);
and U157 (N_157,In_1153,In_1448);
nor U158 (N_158,In_1145,In_574);
or U159 (N_159,In_530,In_396);
or U160 (N_160,In_17,In_1409);
or U161 (N_161,In_10,In_325);
nand U162 (N_162,In_641,In_44);
xnor U163 (N_163,In_54,In_1073);
and U164 (N_164,In_1491,In_659);
xnor U165 (N_165,In_518,In_323);
xor U166 (N_166,In_1011,In_1384);
nor U167 (N_167,In_639,In_1259);
or U168 (N_168,In_562,In_731);
xor U169 (N_169,In_198,In_390);
or U170 (N_170,In_1085,In_610);
nor U171 (N_171,In_829,In_1429);
or U172 (N_172,In_1364,In_801);
or U173 (N_173,In_497,In_392);
xor U174 (N_174,In_637,In_1396);
nand U175 (N_175,In_884,In_13);
or U176 (N_176,In_981,In_856);
nand U177 (N_177,In_459,In_1499);
and U178 (N_178,In_161,In_539);
xnor U179 (N_179,In_830,In_797);
and U180 (N_180,In_783,In_151);
nor U181 (N_181,In_946,In_1034);
xnor U182 (N_182,In_290,In_1451);
and U183 (N_183,In_89,In_751);
nor U184 (N_184,In_977,In_71);
nand U185 (N_185,In_1393,In_1201);
nand U186 (N_186,In_537,In_186);
nand U187 (N_187,In_1104,In_673);
or U188 (N_188,In_872,In_1082);
and U189 (N_189,In_1355,In_930);
and U190 (N_190,In_140,In_15);
nand U191 (N_191,In_1143,In_265);
or U192 (N_192,In_1120,In_22);
and U193 (N_193,In_532,In_928);
or U194 (N_194,In_893,In_69);
xor U195 (N_195,In_736,In_1212);
nand U196 (N_196,In_326,In_267);
or U197 (N_197,In_564,In_1431);
or U198 (N_198,In_1410,In_1444);
nand U199 (N_199,In_11,In_1421);
nand U200 (N_200,In_1484,In_1127);
or U201 (N_201,In_1023,In_1239);
nand U202 (N_202,In_1186,In_874);
or U203 (N_203,In_1454,In_816);
and U204 (N_204,In_1054,In_672);
and U205 (N_205,In_1106,In_627);
and U206 (N_206,In_550,In_1088);
nand U207 (N_207,In_892,In_531);
nor U208 (N_208,In_1443,In_936);
nor U209 (N_209,In_771,In_349);
and U210 (N_210,In_398,In_1283);
nor U211 (N_211,In_602,In_516);
nand U212 (N_212,In_457,In_1357);
nand U213 (N_213,In_920,In_1174);
or U214 (N_214,In_589,In_1209);
or U215 (N_215,In_1324,In_1447);
or U216 (N_216,In_1134,In_1321);
nand U217 (N_217,In_165,In_223);
xor U218 (N_218,In_1038,In_289);
and U219 (N_219,In_60,In_544);
or U220 (N_220,In_593,In_48);
and U221 (N_221,In_594,In_401);
or U222 (N_222,In_350,In_995);
or U223 (N_223,In_1061,In_1066);
nor U224 (N_224,In_1162,In_96);
nand U225 (N_225,In_845,In_903);
or U226 (N_226,In_540,In_1032);
nand U227 (N_227,In_507,In_264);
nand U228 (N_228,In_1490,In_242);
and U229 (N_229,In_728,In_567);
nand U230 (N_230,In_688,In_1107);
xnor U231 (N_231,In_998,In_474);
nor U232 (N_232,In_1394,In_854);
nand U233 (N_233,In_869,In_971);
and U234 (N_234,In_94,In_908);
xor U235 (N_235,In_575,In_384);
nor U236 (N_236,In_217,In_840);
nand U237 (N_237,In_1230,In_456);
nand U238 (N_238,In_1202,In_1247);
nand U239 (N_239,In_87,In_696);
nor U240 (N_240,In_3,In_1057);
nor U241 (N_241,In_614,In_73);
nand U242 (N_242,In_31,In_978);
nor U243 (N_243,In_137,In_334);
and U244 (N_244,In_1020,In_499);
and U245 (N_245,In_972,In_479);
and U246 (N_246,In_440,In_561);
nor U247 (N_247,In_833,In_1184);
or U248 (N_248,In_1138,In_421);
nand U249 (N_249,In_1055,In_183);
and U250 (N_250,In_170,In_1374);
or U251 (N_251,In_678,In_975);
xor U252 (N_252,In_934,In_484);
and U253 (N_253,In_1253,In_298);
nand U254 (N_254,In_477,In_608);
or U255 (N_255,In_118,In_129);
or U256 (N_256,In_1341,In_192);
or U257 (N_257,In_1387,In_1123);
and U258 (N_258,In_72,In_1286);
xor U259 (N_259,In_271,In_895);
nand U260 (N_260,In_1089,In_1217);
or U261 (N_261,In_317,In_47);
nand U262 (N_262,In_1392,In_340);
xnor U263 (N_263,In_1475,In_1301);
nor U264 (N_264,In_426,In_307);
and U265 (N_265,In_1483,In_708);
nor U266 (N_266,In_230,In_407);
xnor U267 (N_267,In_85,In_393);
nand U268 (N_268,In_199,In_301);
and U269 (N_269,In_647,In_716);
or U270 (N_270,In_281,In_563);
or U271 (N_271,In_842,In_650);
nand U272 (N_272,In_1157,In_701);
nor U273 (N_273,In_1009,In_1028);
or U274 (N_274,In_1140,In_1264);
and U275 (N_275,In_1307,In_758);
nor U276 (N_276,In_1228,In_698);
or U277 (N_277,In_1399,In_273);
xnor U278 (N_278,In_297,In_117);
nor U279 (N_279,In_784,In_143);
or U280 (N_280,In_256,In_965);
or U281 (N_281,In_1173,In_1470);
or U282 (N_282,In_761,In_116);
nor U283 (N_283,In_1437,In_374);
or U284 (N_284,In_1137,In_649);
xnor U285 (N_285,In_448,In_824);
or U286 (N_286,In_1048,In_142);
nor U287 (N_287,In_1345,In_692);
nand U288 (N_288,In_387,In_560);
xor U289 (N_289,In_742,In_700);
nor U290 (N_290,In_991,In_110);
xnor U291 (N_291,In_902,In_1445);
xnor U292 (N_292,In_1411,In_1241);
or U293 (N_293,In_164,In_1194);
and U294 (N_294,In_1171,In_163);
nand U295 (N_295,In_912,In_394);
nand U296 (N_296,In_623,In_1007);
and U297 (N_297,In_1383,In_159);
nand U298 (N_298,In_182,In_1214);
xor U299 (N_299,In_826,In_855);
and U300 (N_300,In_1362,In_737);
and U301 (N_301,In_631,In_35);
or U302 (N_302,In_97,In_463);
or U303 (N_303,In_252,In_1489);
nand U304 (N_304,In_1244,In_1072);
xor U305 (N_305,In_1203,In_1348);
nand U306 (N_306,In_27,In_629);
nor U307 (N_307,In_1183,In_699);
and U308 (N_308,In_1060,In_707);
nor U309 (N_309,In_1235,In_961);
nor U310 (N_310,In_449,In_662);
nor U311 (N_311,In_625,In_521);
or U312 (N_312,In_886,In_722);
nand U313 (N_313,In_1323,In_1232);
nand U314 (N_314,In_400,In_1478);
nor U315 (N_315,In_667,In_511);
xor U316 (N_316,In_1155,In_1043);
xnor U317 (N_317,In_1414,In_406);
nand U318 (N_318,In_19,In_146);
nand U319 (N_319,In_612,In_132);
nor U320 (N_320,In_727,In_1198);
nand U321 (N_321,In_106,In_1017);
or U322 (N_322,In_1180,In_1389);
nor U323 (N_323,In_1152,In_820);
or U324 (N_324,In_300,In_1423);
or U325 (N_325,In_1395,In_613);
and U326 (N_326,In_1016,In_462);
nor U327 (N_327,In_653,In_320);
and U328 (N_328,In_442,In_587);
nand U329 (N_329,In_385,In_1018);
or U330 (N_330,In_221,In_772);
or U331 (N_331,In_939,In_628);
and U332 (N_332,In_420,In_1062);
nor U333 (N_333,In_546,In_212);
and U334 (N_334,In_941,In_717);
nor U335 (N_335,In_482,In_312);
nor U336 (N_336,In_5,In_1302);
and U337 (N_337,In_850,In_853);
nor U338 (N_338,In_983,In_489);
and U339 (N_339,In_1135,In_724);
or U340 (N_340,In_1130,In_55);
nand U341 (N_341,In_1219,In_24);
nor U342 (N_342,In_1468,In_496);
xor U343 (N_343,In_1372,In_646);
nor U344 (N_344,In_213,In_257);
nor U345 (N_345,In_1049,In_569);
nor U346 (N_346,In_598,In_710);
and U347 (N_347,In_1245,In_336);
and U348 (N_348,In_1248,In_451);
nor U349 (N_349,In_1459,In_1480);
or U350 (N_350,In_711,In_26);
nand U351 (N_351,In_174,In_1081);
nor U352 (N_352,In_232,In_554);
nor U353 (N_353,In_513,In_864);
nand U354 (N_354,In_83,In_697);
and U355 (N_355,In_66,In_402);
xor U356 (N_356,In_1080,In_921);
and U357 (N_357,In_0,In_122);
nor U358 (N_358,In_373,In_268);
and U359 (N_359,In_1257,In_176);
xor U360 (N_360,In_1118,In_851);
nor U361 (N_361,In_935,In_640);
nand U362 (N_362,In_75,In_1382);
nand U363 (N_363,In_1110,In_450);
nand U364 (N_364,In_347,In_1);
and U365 (N_365,In_876,In_490);
nor U366 (N_366,In_1021,In_294);
nand U367 (N_367,In_478,In_966);
and U368 (N_368,In_718,In_93);
or U369 (N_369,In_506,In_1343);
or U370 (N_370,In_979,In_1042);
nor U371 (N_371,In_355,In_486);
nand U372 (N_372,In_942,In_1299);
nor U373 (N_373,In_725,In_366);
and U374 (N_374,In_1352,In_1456);
nand U375 (N_375,In_873,In_234);
nand U376 (N_376,In_957,In_606);
nand U377 (N_377,In_992,In_434);
nor U378 (N_378,In_967,In_1013);
nand U379 (N_379,In_588,In_1315);
nor U380 (N_380,In_280,In_4);
and U381 (N_381,In_388,In_1116);
nor U382 (N_382,In_1461,In_1096);
nor U383 (N_383,In_726,In_1190);
nand U384 (N_384,In_1240,In_1251);
nand U385 (N_385,In_1216,In_308);
nor U386 (N_386,In_1398,In_831);
and U387 (N_387,In_803,In_735);
nor U388 (N_388,In_327,In_1426);
nor U389 (N_389,In_162,In_1044);
or U390 (N_390,In_1179,In_153);
and U391 (N_391,In_408,In_621);
nand U392 (N_392,In_331,In_1465);
nand U393 (N_393,In_253,In_536);
and U394 (N_394,In_249,In_1136);
nand U395 (N_395,In_1064,In_1422);
nand U396 (N_396,In_1070,In_433);
xor U397 (N_397,In_679,In_88);
or U398 (N_398,In_1285,In_880);
or U399 (N_399,In_730,In_956);
nor U400 (N_400,In_220,In_524);
and U401 (N_401,In_823,In_127);
or U402 (N_402,In_346,In_225);
and U403 (N_403,In_691,In_9);
nor U404 (N_404,In_1417,In_102);
and U405 (N_405,In_1008,In_131);
and U406 (N_406,In_834,In_411);
nand U407 (N_407,In_1369,In_693);
or U408 (N_408,In_871,In_1317);
or U409 (N_409,In_32,In_702);
nand U410 (N_410,In_25,In_1150);
and U411 (N_411,In_568,In_945);
and U412 (N_412,In_342,In_1074);
and U413 (N_413,In_596,In_37);
and U414 (N_414,In_241,In_668);
nor U415 (N_415,In_172,In_1260);
and U416 (N_416,In_453,In_332);
nor U417 (N_417,In_284,In_262);
nor U418 (N_418,In_694,In_953);
and U419 (N_419,In_1040,In_809);
or U420 (N_420,In_1373,In_769);
nor U421 (N_421,In_1462,In_1192);
and U422 (N_422,In_1261,In_77);
and U423 (N_423,In_1029,In_1496);
nor U424 (N_424,In_428,In_1000);
or U425 (N_425,In_847,In_1166);
or U426 (N_426,In_61,In_149);
nor U427 (N_427,In_1300,In_709);
nor U428 (N_428,In_306,In_465);
nand U429 (N_429,In_1269,In_583);
nor U430 (N_430,In_618,In_1236);
nand U431 (N_431,In_189,In_286);
nor U432 (N_432,In_124,In_686);
xor U433 (N_433,In_1122,In_669);
nor U434 (N_434,In_1224,In_205);
nand U435 (N_435,In_681,In_1272);
nor U436 (N_436,In_1094,In_254);
or U437 (N_437,In_1322,In_1309);
and U438 (N_438,In_635,In_1099);
nand U439 (N_439,In_1477,In_1292);
or U440 (N_440,In_330,In_1326);
and U441 (N_441,In_969,In_120);
nand U442 (N_442,In_922,In_1342);
and U443 (N_443,In_321,In_889);
nor U444 (N_444,In_1111,In_191);
or U445 (N_445,In_1275,In_988);
xor U446 (N_446,In_553,In_1051);
nand U447 (N_447,In_354,In_955);
nor U448 (N_448,In_875,In_781);
nand U449 (N_449,In_1101,In_1378);
nor U450 (N_450,In_914,In_1103);
nor U451 (N_451,In_1402,In_259);
nor U452 (N_452,In_1109,In_1329);
nor U453 (N_453,In_779,In_1119);
nand U454 (N_454,In_793,In_207);
nand U455 (N_455,In_770,In_1277);
or U456 (N_456,In_105,In_1353);
and U457 (N_457,In_796,In_1428);
xor U458 (N_458,In_1154,In_1368);
nand U459 (N_459,In_852,In_476);
nand U460 (N_460,In_970,In_351);
nand U461 (N_461,In_543,In_310);
and U462 (N_462,In_177,In_1318);
nor U463 (N_463,In_380,In_818);
and U464 (N_464,In_896,In_1164);
nand U465 (N_465,In_1498,In_245);
nor U466 (N_466,In_430,In_309);
and U467 (N_467,In_368,In_1160);
nand U468 (N_468,In_12,In_1408);
and U469 (N_469,In_169,In_243);
and U470 (N_470,In_152,In_444);
or U471 (N_471,In_237,In_333);
or U472 (N_472,In_626,In_1142);
or U473 (N_473,In_1296,In_817);
nand U474 (N_474,In_1131,In_480);
xor U475 (N_475,In_295,In_488);
and U476 (N_476,In_765,In_362);
nand U477 (N_477,In_1053,In_651);
or U478 (N_478,In_750,In_418);
or U479 (N_479,In_206,In_913);
nor U480 (N_480,In_441,In_1165);
and U481 (N_481,In_807,In_1218);
xor U482 (N_482,In_525,In_655);
nor U483 (N_483,In_714,In_753);
nand U484 (N_484,In_1246,In_548);
nand U485 (N_485,In_50,In_1039);
nand U486 (N_486,In_591,In_314);
and U487 (N_487,In_144,In_318);
or U488 (N_488,In_181,In_891);
or U489 (N_489,In_973,In_760);
and U490 (N_490,In_436,In_439);
and U491 (N_491,In_458,In_1189);
nand U492 (N_492,In_878,In_690);
or U493 (N_493,In_795,In_1452);
nor U494 (N_494,In_1159,In_422);
or U495 (N_495,In_1325,In_200);
and U496 (N_496,In_108,In_78);
or U497 (N_497,In_508,In_1156);
or U498 (N_498,In_813,In_1293);
nor U499 (N_499,In_835,In_86);
and U500 (N_500,In_452,In_674);
nor U501 (N_501,In_46,In_810);
nand U502 (N_502,In_1100,In_1204);
nor U503 (N_503,In_389,In_282);
or U504 (N_504,In_578,In_1280);
nor U505 (N_505,In_168,In_1458);
or U506 (N_506,In_985,In_1041);
or U507 (N_507,In_30,In_1227);
or U508 (N_508,In_470,In_812);
xor U509 (N_509,In_461,In_82);
or U510 (N_510,In_98,In_343);
and U511 (N_511,In_501,In_502);
and U512 (N_512,In_1281,In_958);
or U513 (N_513,In_989,In_405);
and U514 (N_514,In_721,In_258);
xnor U515 (N_515,In_745,In_250);
and U516 (N_516,In_1349,In_190);
nor U517 (N_517,In_1430,In_933);
nand U518 (N_518,In_763,In_1086);
and U519 (N_519,In_789,In_95);
and U520 (N_520,In_1406,In_277);
nor U521 (N_521,In_658,In_766);
and U522 (N_522,In_720,In_1006);
and U523 (N_523,In_1344,In_1022);
and U524 (N_524,In_580,In_584);
or U525 (N_525,In_733,In_1226);
or U526 (N_526,In_431,In_832);
and U527 (N_527,In_1188,In_804);
and U528 (N_528,In_125,In_791);
or U529 (N_529,In_897,In_1193);
nor U530 (N_530,In_1442,In_1185);
nand U531 (N_531,In_863,In_557);
and U532 (N_532,In_214,In_1222);
or U533 (N_533,In_361,In_1063);
and U534 (N_534,In_203,In_1208);
nand U535 (N_535,In_906,In_1482);
nand U536 (N_536,In_741,In_1195);
xnor U537 (N_537,In_1033,In_21);
nor U538 (N_538,In_363,In_483);
nand U539 (N_539,In_677,In_849);
nor U540 (N_540,In_519,In_792);
nand U541 (N_541,In_883,In_815);
and U542 (N_542,In_862,In_447);
xnor U543 (N_543,In_660,In_51);
nand U544 (N_544,In_1225,In_28);
or U545 (N_545,In_551,In_1390);
nand U546 (N_546,In_56,In_263);
nand U547 (N_547,In_1297,In_1381);
nand U548 (N_548,In_53,In_987);
nor U549 (N_549,In_33,In_1416);
or U550 (N_550,In_403,In_632);
or U551 (N_551,In_276,In_1266);
nor U552 (N_552,In_216,In_808);
xor U553 (N_553,In_527,In_664);
or U554 (N_554,In_1076,In_1035);
nand U555 (N_555,In_1464,In_1149);
nor U556 (N_556,In_194,In_944);
and U557 (N_557,In_287,In_1400);
nand U558 (N_558,In_729,In_948);
or U559 (N_559,In_915,In_1312);
nand U560 (N_560,In_305,In_247);
nand U561 (N_561,In_1336,In_1004);
or U562 (N_562,In_121,In_844);
nor U563 (N_563,In_622,In_1069);
nor U564 (N_564,In_1433,In_597);
xor U565 (N_565,In_607,In_353);
or U566 (N_566,In_133,In_328);
and U567 (N_567,In_239,In_114);
or U568 (N_568,In_705,In_1098);
nor U569 (N_569,In_375,In_329);
nor U570 (N_570,In_1068,In_819);
xor U571 (N_571,In_348,In_155);
or U572 (N_572,In_481,In_238);
nor U573 (N_573,In_976,In_684);
nand U574 (N_574,In_919,In_952);
or U575 (N_575,In_1361,In_1282);
or U576 (N_576,In_372,In_107);
and U577 (N_577,In_768,In_904);
and U578 (N_578,In_1265,In_43);
nand U579 (N_579,In_535,In_16);
nor U580 (N_580,In_1289,In_1182);
and U581 (N_581,In_1295,In_45);
nand U582 (N_582,In_1479,In_1446);
nor U583 (N_583,In_523,In_382);
and U584 (N_584,In_757,In_377);
nand U585 (N_585,In_1432,In_529);
or U586 (N_586,In_570,In_1424);
nor U587 (N_587,In_1358,In_542);
nor U588 (N_588,In_748,In_1058);
or U589 (N_589,In_64,In_1128);
and U590 (N_590,In_865,In_454);
and U591 (N_591,In_251,In_1001);
nor U592 (N_592,In_404,In_74);
or U593 (N_593,In_113,In_687);
nand U594 (N_594,In_663,In_676);
and U595 (N_595,In_671,In_316);
nand U596 (N_596,In_345,In_141);
nand U597 (N_597,In_837,In_1267);
xor U598 (N_598,In_600,In_313);
nand U599 (N_599,In_881,In_1310);
nand U600 (N_600,In_918,In_14);
and U601 (N_601,In_1163,In_800);
nor U602 (N_602,In_582,In_604);
and U603 (N_603,In_522,In_1132);
and U604 (N_604,In_1386,In_943);
or U605 (N_605,In_379,In_746);
nor U606 (N_606,In_423,In_654);
xor U607 (N_607,In_579,In_552);
and U608 (N_608,In_577,In_1178);
or U609 (N_609,In_898,In_437);
nor U610 (N_610,In_652,In_558);
nand U611 (N_611,In_1453,In_839);
and U612 (N_612,In_926,In_1139);
or U613 (N_613,In_555,In_41);
or U614 (N_614,In_538,In_917);
or U615 (N_615,In_959,In_59);
nor U616 (N_616,In_171,In_23);
and U617 (N_617,In_1206,In_492);
xnor U618 (N_618,In_799,In_1172);
xnor U619 (N_619,In_224,In_446);
nor U620 (N_620,In_1401,In_1427);
nand U621 (N_621,In_868,In_510);
nor U622 (N_622,In_1494,In_859);
or U623 (N_623,In_397,In_1351);
and U624 (N_624,In_1367,In_980);
or U625 (N_625,In_1308,In_179);
or U626 (N_626,In_130,In_1114);
or U627 (N_627,In_1438,In_128);
nor U628 (N_628,In_438,In_1031);
or U629 (N_629,In_644,In_547);
nor U630 (N_630,In_634,In_29);
xor U631 (N_631,In_605,In_828);
nor U632 (N_632,In_498,In_1474);
and U633 (N_633,In_1403,In_670);
and U634 (N_634,In_1419,In_1254);
nand U635 (N_635,In_616,In_786);
nor U636 (N_636,In_1330,In_545);
nor U637 (N_637,In_1084,In_1314);
and U638 (N_638,In_1210,In_932);
and U639 (N_639,In_573,In_1046);
xor U640 (N_640,In_566,In_178);
or U641 (N_641,In_848,In_222);
or U642 (N_642,In_166,In_601);
and U643 (N_643,In_1311,In_1471);
nand U644 (N_644,In_1050,In_1472);
and U645 (N_645,In_509,In_123);
or U646 (N_646,In_565,In_767);
nand U647 (N_647,In_1262,In_528);
and U648 (N_648,In_158,In_1287);
and U649 (N_649,In_1181,In_383);
or U650 (N_650,In_260,In_858);
or U651 (N_651,In_999,In_1102);
xor U652 (N_652,In_269,In_414);
nand U653 (N_653,In_235,In_743);
nand U654 (N_654,In_1492,In_1170);
and U655 (N_655,In_244,In_1019);
and U656 (N_656,In_806,In_279);
and U657 (N_657,In_1278,In_609);
nand U658 (N_658,In_960,In_1306);
xor U659 (N_659,In_1036,In_747);
and U660 (N_660,In_288,In_500);
nor U661 (N_661,In_638,In_1346);
nor U662 (N_662,In_620,In_381);
and U663 (N_663,In_84,In_1237);
xor U664 (N_664,In_526,In_1075);
and U665 (N_665,In_1030,In_62);
nand U666 (N_666,In_1263,In_413);
nor U667 (N_667,In_196,In_993);
or U668 (N_668,In_586,In_794);
nor U669 (N_669,In_335,In_485);
nand U670 (N_670,In_590,In_39);
xor U671 (N_671,In_925,In_581);
nor U672 (N_672,In_1014,In_283);
nand U673 (N_673,In_572,In_901);
xnor U674 (N_674,In_65,In_505);
or U675 (N_675,In_1045,In_994);
xor U676 (N_676,In_927,In_139);
xnor U677 (N_677,In_949,In_180);
and U678 (N_678,In_790,In_1141);
nand U679 (N_679,In_1012,In_52);
nor U680 (N_680,In_910,In_665);
nand U681 (N_681,In_517,In_67);
and U682 (N_682,In_1133,In_471);
nor U683 (N_683,In_18,In_357);
nand U684 (N_684,In_1005,In_495);
nor U685 (N_685,In_195,In_104);
xnor U686 (N_686,In_931,In_1435);
and U687 (N_687,In_1274,In_900);
nor U688 (N_688,In_358,In_732);
and U689 (N_689,In_630,In_754);
nor U690 (N_690,In_1146,In_275);
xor U691 (N_691,In_76,In_42);
nor U692 (N_692,In_951,In_778);
nand U693 (N_693,In_156,In_1415);
nor U694 (N_694,In_1168,In_1434);
nor U695 (N_695,In_215,In_167);
nor U696 (N_696,In_91,In_303);
or U697 (N_697,In_1158,In_135);
nor U698 (N_698,In_410,In_534);
and U699 (N_699,In_986,In_1097);
or U700 (N_700,In_1371,In_1024);
xnor U701 (N_701,In_291,In_197);
or U702 (N_702,In_1126,In_138);
xnor U703 (N_703,In_1488,In_160);
and U704 (N_704,In_356,In_6);
and U705 (N_705,In_311,In_643);
nor U706 (N_706,In_57,In_175);
or U707 (N_707,In_1418,In_866);
nor U708 (N_708,In_1025,In_1083);
nor U709 (N_709,In_822,In_40);
nand U710 (N_710,In_964,In_1363);
nor U711 (N_711,In_503,In_843);
nor U712 (N_712,In_968,In_226);
and U713 (N_713,In_1125,In_1234);
and U714 (N_714,In_49,In_811);
and U715 (N_715,In_1338,In_119);
xor U716 (N_716,In_1303,In_533);
or U717 (N_717,In_246,In_261);
nand U718 (N_718,In_491,In_322);
xnor U719 (N_719,In_1256,In_1115);
and U720 (N_720,In_2,In_827);
nand U721 (N_721,In_1375,In_1460);
and U722 (N_722,In_1148,In_1347);
xnor U723 (N_723,In_112,In_227);
or U724 (N_724,In_145,In_940);
or U725 (N_725,In_147,In_1112);
or U726 (N_726,In_1473,In_645);
xnor U727 (N_727,In_675,In_661);
or U728 (N_728,In_1199,In_1079);
or U729 (N_729,In_1176,In_81);
or U730 (N_730,In_1407,In_611);
nand U731 (N_731,In_395,In_905);
and U732 (N_732,In_1279,In_617);
nand U733 (N_733,In_1467,In_642);
nand U734 (N_734,In_270,In_821);
and U735 (N_735,In_1213,In_974);
nand U736 (N_736,In_1161,In_680);
and U737 (N_737,In_1385,In_1113);
and U738 (N_738,In_706,In_1124);
nand U739 (N_739,In_648,In_1268);
nand U740 (N_740,In_412,In_984);
or U741 (N_741,In_92,In_1273);
nand U742 (N_742,In_299,In_409);
nor U743 (N_743,In_1026,In_1469);
nor U744 (N_744,In_782,In_443);
and U745 (N_745,In_836,In_1497);
or U746 (N_746,In_424,In_916);
and U747 (N_747,In_319,In_1485);
and U748 (N_748,In_370,In_204);
nor U749 (N_749,In_857,In_228);
or U750 (N_750,In_1304,In_91);
nor U751 (N_751,In_1263,In_1244);
nor U752 (N_752,In_1065,In_96);
nand U753 (N_753,In_1376,In_1455);
nand U754 (N_754,In_1250,In_1020);
nand U755 (N_755,In_88,In_312);
and U756 (N_756,In_615,In_301);
nand U757 (N_757,In_638,In_1355);
nand U758 (N_758,In_286,In_673);
nor U759 (N_759,In_332,In_28);
or U760 (N_760,In_953,In_1118);
nand U761 (N_761,In_1151,In_14);
nand U762 (N_762,In_1286,In_77);
and U763 (N_763,In_1263,In_727);
and U764 (N_764,In_654,In_576);
nand U765 (N_765,In_493,In_837);
nand U766 (N_766,In_36,In_238);
and U767 (N_767,In_289,In_687);
nand U768 (N_768,In_1101,In_801);
nand U769 (N_769,In_1381,In_893);
or U770 (N_770,In_1391,In_515);
nand U771 (N_771,In_1498,In_3);
nand U772 (N_772,In_102,In_1237);
and U773 (N_773,In_925,In_635);
nand U774 (N_774,In_955,In_274);
nor U775 (N_775,In_652,In_1442);
and U776 (N_776,In_1226,In_74);
nand U777 (N_777,In_384,In_282);
xnor U778 (N_778,In_96,In_62);
or U779 (N_779,In_531,In_1052);
and U780 (N_780,In_1421,In_430);
or U781 (N_781,In_703,In_567);
or U782 (N_782,In_1270,In_1207);
nand U783 (N_783,In_62,In_1236);
nor U784 (N_784,In_1304,In_885);
or U785 (N_785,In_259,In_1416);
and U786 (N_786,In_1215,In_844);
nand U787 (N_787,In_700,In_1362);
nand U788 (N_788,In_331,In_989);
and U789 (N_789,In_962,In_1249);
or U790 (N_790,In_952,In_1305);
and U791 (N_791,In_957,In_1286);
nor U792 (N_792,In_729,In_428);
nand U793 (N_793,In_1065,In_318);
nor U794 (N_794,In_1006,In_1204);
nand U795 (N_795,In_339,In_1031);
nor U796 (N_796,In_879,In_545);
nand U797 (N_797,In_1471,In_46);
nand U798 (N_798,In_553,In_867);
nor U799 (N_799,In_1406,In_1103);
xnor U800 (N_800,In_429,In_134);
nand U801 (N_801,In_4,In_538);
and U802 (N_802,In_463,In_532);
nor U803 (N_803,In_849,In_1169);
nand U804 (N_804,In_79,In_433);
nand U805 (N_805,In_924,In_250);
and U806 (N_806,In_783,In_1329);
nand U807 (N_807,In_1031,In_1046);
and U808 (N_808,In_1380,In_951);
nor U809 (N_809,In_1070,In_705);
nand U810 (N_810,In_1444,In_306);
nor U811 (N_811,In_958,In_448);
or U812 (N_812,In_142,In_1446);
xnor U813 (N_813,In_619,In_1224);
or U814 (N_814,In_541,In_312);
xor U815 (N_815,In_157,In_61);
nor U816 (N_816,In_500,In_344);
nand U817 (N_817,In_1380,In_1150);
or U818 (N_818,In_1397,In_1297);
xor U819 (N_819,In_994,In_123);
nand U820 (N_820,In_1015,In_1456);
and U821 (N_821,In_1138,In_715);
nand U822 (N_822,In_1321,In_1413);
nand U823 (N_823,In_873,In_1068);
nor U824 (N_824,In_123,In_524);
nand U825 (N_825,In_407,In_764);
and U826 (N_826,In_45,In_484);
nor U827 (N_827,In_1239,In_1421);
nand U828 (N_828,In_1163,In_953);
nand U829 (N_829,In_1387,In_955);
nor U830 (N_830,In_66,In_1304);
and U831 (N_831,In_1274,In_796);
or U832 (N_832,In_267,In_864);
and U833 (N_833,In_417,In_845);
or U834 (N_834,In_787,In_1259);
and U835 (N_835,In_1109,In_1312);
and U836 (N_836,In_980,In_269);
nand U837 (N_837,In_410,In_564);
nor U838 (N_838,In_897,In_816);
nor U839 (N_839,In_895,In_120);
and U840 (N_840,In_472,In_758);
nor U841 (N_841,In_738,In_1022);
and U842 (N_842,In_857,In_1399);
nor U843 (N_843,In_1228,In_138);
nand U844 (N_844,In_870,In_483);
or U845 (N_845,In_1275,In_8);
nor U846 (N_846,In_393,In_178);
and U847 (N_847,In_411,In_51);
or U848 (N_848,In_399,In_329);
nor U849 (N_849,In_625,In_721);
xor U850 (N_850,In_782,In_1445);
nand U851 (N_851,In_443,In_348);
or U852 (N_852,In_1335,In_1465);
nand U853 (N_853,In_1079,In_301);
nand U854 (N_854,In_1372,In_7);
or U855 (N_855,In_719,In_658);
nand U856 (N_856,In_709,In_710);
or U857 (N_857,In_905,In_900);
or U858 (N_858,In_1152,In_902);
or U859 (N_859,In_737,In_793);
and U860 (N_860,In_1297,In_206);
or U861 (N_861,In_1234,In_359);
nand U862 (N_862,In_136,In_437);
nand U863 (N_863,In_1159,In_1233);
nand U864 (N_864,In_1274,In_165);
nand U865 (N_865,In_1276,In_1243);
nand U866 (N_866,In_353,In_394);
nor U867 (N_867,In_479,In_115);
or U868 (N_868,In_1314,In_350);
or U869 (N_869,In_637,In_1426);
and U870 (N_870,In_976,In_554);
nor U871 (N_871,In_1432,In_1000);
nand U872 (N_872,In_311,In_1028);
or U873 (N_873,In_79,In_821);
nor U874 (N_874,In_416,In_830);
or U875 (N_875,In_1179,In_876);
and U876 (N_876,In_1169,In_544);
or U877 (N_877,In_159,In_976);
and U878 (N_878,In_594,In_528);
nand U879 (N_879,In_712,In_758);
or U880 (N_880,In_390,In_1384);
xnor U881 (N_881,In_526,In_517);
and U882 (N_882,In_889,In_457);
nand U883 (N_883,In_528,In_870);
xor U884 (N_884,In_732,In_1412);
or U885 (N_885,In_236,In_1125);
nor U886 (N_886,In_1089,In_31);
nand U887 (N_887,In_390,In_861);
nand U888 (N_888,In_384,In_638);
xor U889 (N_889,In_209,In_101);
xnor U890 (N_890,In_1227,In_1397);
or U891 (N_891,In_1167,In_803);
nand U892 (N_892,In_1356,In_1422);
or U893 (N_893,In_1422,In_362);
nor U894 (N_894,In_391,In_773);
or U895 (N_895,In_246,In_563);
and U896 (N_896,In_475,In_747);
xnor U897 (N_897,In_1232,In_450);
nand U898 (N_898,In_1028,In_1353);
or U899 (N_899,In_961,In_584);
nor U900 (N_900,In_741,In_866);
or U901 (N_901,In_19,In_366);
nand U902 (N_902,In_1153,In_772);
nand U903 (N_903,In_48,In_388);
xor U904 (N_904,In_315,In_1281);
nand U905 (N_905,In_948,In_1301);
and U906 (N_906,In_633,In_552);
nor U907 (N_907,In_1143,In_1024);
or U908 (N_908,In_272,In_903);
nor U909 (N_909,In_1366,In_39);
nor U910 (N_910,In_475,In_1238);
nor U911 (N_911,In_101,In_1402);
nand U912 (N_912,In_1437,In_238);
or U913 (N_913,In_1201,In_766);
and U914 (N_914,In_593,In_79);
and U915 (N_915,In_740,In_801);
nand U916 (N_916,In_107,In_627);
nor U917 (N_917,In_806,In_712);
nor U918 (N_918,In_1058,In_1403);
nand U919 (N_919,In_670,In_630);
nand U920 (N_920,In_434,In_1271);
nor U921 (N_921,In_31,In_514);
and U922 (N_922,In_1414,In_1308);
and U923 (N_923,In_1001,In_274);
nor U924 (N_924,In_65,In_863);
or U925 (N_925,In_354,In_1333);
or U926 (N_926,In_1487,In_1386);
or U927 (N_927,In_1166,In_1221);
and U928 (N_928,In_653,In_599);
xnor U929 (N_929,In_361,In_419);
or U930 (N_930,In_828,In_929);
nor U931 (N_931,In_1046,In_1383);
nor U932 (N_932,In_989,In_551);
nor U933 (N_933,In_216,In_910);
or U934 (N_934,In_1389,In_1145);
and U935 (N_935,In_658,In_519);
or U936 (N_936,In_291,In_88);
or U937 (N_937,In_1073,In_1313);
or U938 (N_938,In_1066,In_618);
and U939 (N_939,In_651,In_997);
and U940 (N_940,In_175,In_223);
and U941 (N_941,In_60,In_365);
nor U942 (N_942,In_259,In_114);
nand U943 (N_943,In_1001,In_433);
nor U944 (N_944,In_1044,In_52);
nand U945 (N_945,In_739,In_1380);
xnor U946 (N_946,In_942,In_254);
or U947 (N_947,In_875,In_601);
nand U948 (N_948,In_1370,In_1170);
or U949 (N_949,In_1273,In_791);
or U950 (N_950,In_920,In_798);
and U951 (N_951,In_415,In_230);
nand U952 (N_952,In_270,In_1375);
or U953 (N_953,In_986,In_1022);
nand U954 (N_954,In_276,In_1423);
and U955 (N_955,In_212,In_588);
or U956 (N_956,In_531,In_176);
nor U957 (N_957,In_152,In_313);
or U958 (N_958,In_1275,In_563);
xnor U959 (N_959,In_853,In_788);
nand U960 (N_960,In_292,In_212);
and U961 (N_961,In_906,In_150);
nor U962 (N_962,In_1105,In_47);
or U963 (N_963,In_589,In_453);
nand U964 (N_964,In_637,In_1401);
nor U965 (N_965,In_30,In_932);
or U966 (N_966,In_382,In_432);
and U967 (N_967,In_1156,In_702);
nand U968 (N_968,In_259,In_460);
nor U969 (N_969,In_385,In_1241);
and U970 (N_970,In_804,In_1163);
nor U971 (N_971,In_1378,In_518);
and U972 (N_972,In_622,In_847);
xnor U973 (N_973,In_182,In_1161);
nor U974 (N_974,In_415,In_354);
xor U975 (N_975,In_61,In_209);
and U976 (N_976,In_440,In_1123);
and U977 (N_977,In_1380,In_711);
nor U978 (N_978,In_782,In_675);
nor U979 (N_979,In_188,In_203);
nand U980 (N_980,In_1039,In_756);
nor U981 (N_981,In_493,In_1349);
nand U982 (N_982,In_935,In_738);
nor U983 (N_983,In_777,In_232);
nand U984 (N_984,In_768,In_278);
nor U985 (N_985,In_1417,In_1122);
nor U986 (N_986,In_437,In_846);
nor U987 (N_987,In_1224,In_1187);
nor U988 (N_988,In_72,In_1342);
or U989 (N_989,In_326,In_1469);
or U990 (N_990,In_1409,In_1247);
nor U991 (N_991,In_788,In_320);
or U992 (N_992,In_264,In_1283);
or U993 (N_993,In_930,In_56);
nand U994 (N_994,In_1050,In_1222);
or U995 (N_995,In_240,In_1154);
xnor U996 (N_996,In_321,In_598);
xnor U997 (N_997,In_235,In_877);
nor U998 (N_998,In_752,In_1051);
nor U999 (N_999,In_405,In_623);
or U1000 (N_1000,N_634,N_727);
or U1001 (N_1001,N_230,N_126);
or U1002 (N_1002,N_325,N_939);
xor U1003 (N_1003,N_602,N_938);
or U1004 (N_1004,N_879,N_814);
nand U1005 (N_1005,N_416,N_599);
and U1006 (N_1006,N_391,N_684);
nor U1007 (N_1007,N_921,N_151);
xor U1008 (N_1008,N_401,N_72);
nand U1009 (N_1009,N_421,N_918);
or U1010 (N_1010,N_486,N_20);
nand U1011 (N_1011,N_514,N_121);
or U1012 (N_1012,N_440,N_790);
or U1013 (N_1013,N_503,N_975);
and U1014 (N_1014,N_622,N_469);
nand U1015 (N_1015,N_701,N_323);
nor U1016 (N_1016,N_800,N_772);
and U1017 (N_1017,N_659,N_76);
and U1018 (N_1018,N_821,N_474);
xnor U1019 (N_1019,N_653,N_519);
xor U1020 (N_1020,N_53,N_499);
nor U1021 (N_1021,N_862,N_604);
or U1022 (N_1022,N_806,N_644);
or U1023 (N_1023,N_1,N_471);
or U1024 (N_1024,N_402,N_115);
or U1025 (N_1025,N_32,N_992);
and U1026 (N_1026,N_920,N_985);
and U1027 (N_1027,N_84,N_465);
xor U1028 (N_1028,N_216,N_118);
nand U1029 (N_1029,N_298,N_615);
nand U1030 (N_1030,N_613,N_949);
nor U1031 (N_1031,N_271,N_28);
nor U1032 (N_1032,N_864,N_40);
nor U1033 (N_1033,N_650,N_691);
xor U1034 (N_1034,N_572,N_453);
nand U1035 (N_1035,N_686,N_587);
and U1036 (N_1036,N_224,N_117);
xnor U1037 (N_1037,N_415,N_770);
or U1038 (N_1038,N_193,N_746);
or U1039 (N_1039,N_427,N_501);
nand U1040 (N_1040,N_529,N_609);
and U1041 (N_1041,N_630,N_595);
nor U1042 (N_1042,N_768,N_124);
nor U1043 (N_1043,N_422,N_694);
nand U1044 (N_1044,N_158,N_867);
nor U1045 (N_1045,N_467,N_850);
nor U1046 (N_1046,N_911,N_747);
or U1047 (N_1047,N_835,N_637);
and U1048 (N_1048,N_581,N_181);
or U1049 (N_1049,N_400,N_853);
nor U1050 (N_1050,N_733,N_530);
xor U1051 (N_1051,N_66,N_69);
or U1052 (N_1052,N_131,N_108);
nand U1053 (N_1053,N_885,N_424);
nand U1054 (N_1054,N_33,N_668);
nor U1055 (N_1055,N_218,N_771);
nor U1056 (N_1056,N_948,N_296);
nor U1057 (N_1057,N_342,N_950);
nor U1058 (N_1058,N_783,N_873);
and U1059 (N_1059,N_497,N_669);
nand U1060 (N_1060,N_278,N_163);
nand U1061 (N_1061,N_246,N_157);
nor U1062 (N_1062,N_756,N_833);
nor U1063 (N_1063,N_951,N_575);
xnor U1064 (N_1064,N_740,N_174);
nand U1065 (N_1065,N_364,N_194);
nand U1066 (N_1066,N_754,N_886);
or U1067 (N_1067,N_801,N_103);
nand U1068 (N_1068,N_683,N_468);
and U1069 (N_1069,N_914,N_852);
and U1070 (N_1070,N_138,N_444);
and U1071 (N_1071,N_973,N_39);
and U1072 (N_1072,N_347,N_667);
or U1073 (N_1073,N_95,N_372);
and U1074 (N_1074,N_751,N_954);
xnor U1075 (N_1075,N_607,N_127);
nand U1076 (N_1076,N_627,N_989);
nand U1077 (N_1077,N_155,N_113);
nand U1078 (N_1078,N_829,N_591);
or U1079 (N_1079,N_169,N_997);
and U1080 (N_1080,N_847,N_438);
nand U1081 (N_1081,N_696,N_279);
or U1082 (N_1082,N_681,N_226);
nor U1083 (N_1083,N_904,N_393);
or U1084 (N_1084,N_930,N_809);
nor U1085 (N_1085,N_620,N_721);
nor U1086 (N_1086,N_414,N_319);
nor U1087 (N_1087,N_349,N_924);
nor U1088 (N_1088,N_354,N_260);
or U1089 (N_1089,N_326,N_91);
xor U1090 (N_1090,N_542,N_909);
nand U1091 (N_1091,N_826,N_880);
nor U1092 (N_1092,N_242,N_656);
or U1093 (N_1093,N_738,N_173);
nor U1094 (N_1094,N_359,N_310);
nand U1095 (N_1095,N_420,N_692);
nand U1096 (N_1096,N_726,N_413);
or U1097 (N_1097,N_365,N_578);
or U1098 (N_1098,N_146,N_883);
or U1099 (N_1099,N_858,N_657);
nand U1100 (N_1100,N_875,N_429);
and U1101 (N_1101,N_535,N_189);
and U1102 (N_1102,N_273,N_720);
and U1103 (N_1103,N_957,N_967);
or U1104 (N_1104,N_605,N_635);
and U1105 (N_1105,N_133,N_380);
or U1106 (N_1106,N_254,N_943);
and U1107 (N_1107,N_177,N_141);
or U1108 (N_1108,N_191,N_869);
or U1109 (N_1109,N_19,N_144);
nor U1110 (N_1110,N_616,N_63);
or U1111 (N_1111,N_648,N_176);
nand U1112 (N_1112,N_68,N_636);
or U1113 (N_1113,N_742,N_27);
nand U1114 (N_1114,N_80,N_901);
or U1115 (N_1115,N_43,N_825);
or U1116 (N_1116,N_752,N_94);
or U1117 (N_1117,N_167,N_135);
and U1118 (N_1118,N_456,N_820);
and U1119 (N_1119,N_944,N_446);
and U1120 (N_1120,N_228,N_837);
or U1121 (N_1121,N_990,N_284);
nor U1122 (N_1122,N_494,N_30);
nand U1123 (N_1123,N_512,N_705);
and U1124 (N_1124,N_162,N_23);
and U1125 (N_1125,N_328,N_580);
nor U1126 (N_1126,N_351,N_455);
nand U1127 (N_1127,N_817,N_376);
nor U1128 (N_1128,N_286,N_898);
nand U1129 (N_1129,N_788,N_2);
nand U1130 (N_1130,N_406,N_164);
nand U1131 (N_1131,N_331,N_903);
xnor U1132 (N_1132,N_798,N_891);
and U1133 (N_1133,N_227,N_498);
xnor U1134 (N_1134,N_900,N_571);
xnor U1135 (N_1135,N_588,N_831);
nor U1136 (N_1136,N_240,N_116);
xor U1137 (N_1137,N_263,N_965);
nor U1138 (N_1138,N_827,N_905);
or U1139 (N_1139,N_513,N_120);
nand U1140 (N_1140,N_466,N_407);
nand U1141 (N_1141,N_638,N_457);
nor U1142 (N_1142,N_172,N_600);
or U1143 (N_1143,N_92,N_309);
and U1144 (N_1144,N_225,N_878);
and U1145 (N_1145,N_674,N_972);
and U1146 (N_1146,N_596,N_360);
or U1147 (N_1147,N_672,N_171);
and U1148 (N_1148,N_504,N_710);
and U1149 (N_1149,N_44,N_663);
and U1150 (N_1150,N_371,N_366);
nor U1151 (N_1151,N_197,N_662);
nand U1152 (N_1152,N_507,N_941);
nor U1153 (N_1153,N_262,N_538);
and U1154 (N_1154,N_554,N_524);
nand U1155 (N_1155,N_160,N_122);
and U1156 (N_1156,N_527,N_166);
and U1157 (N_1157,N_755,N_714);
and U1158 (N_1158,N_409,N_687);
nor U1159 (N_1159,N_9,N_848);
nor U1160 (N_1160,N_841,N_540);
or U1161 (N_1161,N_132,N_556);
nand U1162 (N_1162,N_428,N_633);
or U1163 (N_1163,N_435,N_38);
and U1164 (N_1164,N_37,N_153);
or U1165 (N_1165,N_509,N_815);
nor U1166 (N_1166,N_358,N_758);
or U1167 (N_1167,N_79,N_589);
and U1168 (N_1168,N_405,N_152);
or U1169 (N_1169,N_487,N_114);
or U1170 (N_1170,N_699,N_55);
and U1171 (N_1171,N_386,N_688);
and U1172 (N_1172,N_411,N_250);
and U1173 (N_1173,N_221,N_110);
nor U1174 (N_1174,N_215,N_492);
nand U1175 (N_1175,N_547,N_551);
xnor U1176 (N_1176,N_399,N_212);
nor U1177 (N_1177,N_234,N_346);
and U1178 (N_1178,N_59,N_410);
nand U1179 (N_1179,N_846,N_179);
or U1180 (N_1180,N_676,N_645);
nor U1181 (N_1181,N_332,N_628);
or U1182 (N_1182,N_22,N_16);
nor U1183 (N_1183,N_933,N_643);
nor U1184 (N_1184,N_24,N_956);
nand U1185 (N_1185,N_489,N_287);
nand U1186 (N_1186,N_805,N_830);
nand U1187 (N_1187,N_460,N_966);
or U1188 (N_1188,N_31,N_881);
and U1189 (N_1189,N_362,N_205);
and U1190 (N_1190,N_111,N_813);
nand U1191 (N_1191,N_397,N_838);
nor U1192 (N_1192,N_266,N_808);
or U1193 (N_1193,N_586,N_836);
nand U1194 (N_1194,N_545,N_889);
or U1195 (N_1195,N_490,N_969);
or U1196 (N_1196,N_77,N_180);
or U1197 (N_1197,N_539,N_477);
nand U1198 (N_1198,N_762,N_106);
nor U1199 (N_1199,N_308,N_65);
and U1200 (N_1200,N_876,N_626);
or U1201 (N_1201,N_573,N_741);
nand U1202 (N_1202,N_553,N_811);
nand U1203 (N_1203,N_321,N_845);
nor U1204 (N_1204,N_819,N_47);
nor U1205 (N_1205,N_353,N_685);
or U1206 (N_1206,N_670,N_139);
nor U1207 (N_1207,N_217,N_15);
nand U1208 (N_1208,N_147,N_717);
xor U1209 (N_1209,N_960,N_984);
or U1210 (N_1210,N_666,N_612);
nand U1211 (N_1211,N_508,N_196);
nor U1212 (N_1212,N_912,N_919);
nor U1213 (N_1213,N_282,N_640);
xor U1214 (N_1214,N_404,N_90);
or U1215 (N_1215,N_269,N_175);
xnor U1216 (N_1216,N_462,N_201);
nor U1217 (N_1217,N_373,N_293);
and U1218 (N_1218,N_865,N_274);
or U1219 (N_1219,N_963,N_202);
or U1220 (N_1220,N_988,N_849);
xor U1221 (N_1221,N_96,N_673);
and U1222 (N_1222,N_934,N_98);
nor U1223 (N_1223,N_646,N_974);
or U1224 (N_1224,N_178,N_515);
nand U1225 (N_1225,N_761,N_412);
nor U1226 (N_1226,N_536,N_148);
or U1227 (N_1227,N_582,N_842);
or U1228 (N_1228,N_102,N_767);
nand U1229 (N_1229,N_464,N_60);
nor U1230 (N_1230,N_704,N_355);
or U1231 (N_1231,N_680,N_11);
nand U1232 (N_1232,N_82,N_970);
and U1233 (N_1233,N_57,N_394);
nand U1234 (N_1234,N_629,N_367);
nand U1235 (N_1235,N_526,N_500);
and U1236 (N_1236,N_606,N_5);
or U1237 (N_1237,N_495,N_384);
and U1238 (N_1238,N_781,N_759);
and U1239 (N_1239,N_61,N_285);
or U1240 (N_1240,N_736,N_136);
or U1241 (N_1241,N_395,N_327);
or U1242 (N_1242,N_214,N_339);
and U1243 (N_1243,N_249,N_565);
nor U1244 (N_1244,N_42,N_485);
or U1245 (N_1245,N_952,N_834);
or U1246 (N_1246,N_961,N_665);
nor U1247 (N_1247,N_336,N_443);
and U1248 (N_1248,N_947,N_923);
nand U1249 (N_1249,N_543,N_516);
xor U1250 (N_1250,N_312,N_142);
or U1251 (N_1251,N_773,N_190);
and U1252 (N_1252,N_804,N_213);
and U1253 (N_1253,N_154,N_978);
xnor U1254 (N_1254,N_344,N_678);
nand U1255 (N_1255,N_238,N_283);
and U1256 (N_1256,N_50,N_598);
nor U1257 (N_1257,N_859,N_549);
and U1258 (N_1258,N_706,N_567);
and U1259 (N_1259,N_46,N_112);
nor U1260 (N_1260,N_480,N_807);
nor U1261 (N_1261,N_780,N_302);
nor U1262 (N_1262,N_318,N_7);
nor U1263 (N_1263,N_658,N_281);
xor U1264 (N_1264,N_942,N_786);
and U1265 (N_1265,N_425,N_335);
xnor U1266 (N_1266,N_430,N_334);
nor U1267 (N_1267,N_265,N_451);
xor U1268 (N_1268,N_906,N_145);
nor U1269 (N_1269,N_583,N_590);
nand U1270 (N_1270,N_245,N_233);
and U1271 (N_1271,N_315,N_361);
nand U1272 (N_1272,N_832,N_744);
or U1273 (N_1273,N_313,N_532);
and U1274 (N_1274,N_971,N_481);
xor U1275 (N_1275,N_895,N_743);
and U1276 (N_1276,N_324,N_140);
nand U1277 (N_1277,N_470,N_763);
or U1278 (N_1278,N_774,N_936);
or U1279 (N_1279,N_463,N_436);
or U1280 (N_1280,N_908,N_893);
and U1281 (N_1281,N_541,N_198);
nand U1282 (N_1282,N_610,N_439);
nor U1283 (N_1283,N_623,N_803);
nor U1284 (N_1284,N_937,N_925);
nor U1285 (N_1285,N_21,N_458);
nand U1286 (N_1286,N_484,N_161);
or U1287 (N_1287,N_252,N_247);
and U1288 (N_1288,N_712,N_654);
nor U1289 (N_1289,N_700,N_356);
and U1290 (N_1290,N_619,N_75);
or U1291 (N_1291,N_100,N_964);
or U1292 (N_1292,N_702,N_856);
and U1293 (N_1293,N_861,N_304);
xnor U1294 (N_1294,N_894,N_769);
and U1295 (N_1295,N_4,N_632);
and U1296 (N_1296,N_206,N_698);
nor U1297 (N_1297,N_54,N_259);
or U1298 (N_1298,N_624,N_417);
nor U1299 (N_1299,N_728,N_560);
and U1300 (N_1300,N_475,N_268);
nand U1301 (N_1301,N_868,N_383);
nor U1302 (N_1302,N_204,N_253);
nor U1303 (N_1303,N_182,N_426);
nand U1304 (N_1304,N_995,N_311);
and U1305 (N_1305,N_718,N_41);
nor U1306 (N_1306,N_896,N_557);
or U1307 (N_1307,N_917,N_922);
nand U1308 (N_1308,N_614,N_377);
and U1309 (N_1309,N_730,N_398);
and U1310 (N_1310,N_523,N_306);
xor U1311 (N_1311,N_340,N_199);
nand U1312 (N_1312,N_818,N_611);
nor U1313 (N_1313,N_101,N_945);
xor U1314 (N_1314,N_872,N_352);
and U1315 (N_1315,N_729,N_592);
and U1316 (N_1316,N_928,N_996);
nor U1317 (N_1317,N_454,N_796);
nand U1318 (N_1318,N_337,N_220);
or U1319 (N_1319,N_946,N_418);
nand U1320 (N_1320,N_6,N_631);
or U1321 (N_1321,N_493,N_647);
or U1322 (N_1322,N_49,N_459);
xnor U1323 (N_1323,N_472,N_107);
xor U1324 (N_1324,N_156,N_83);
nor U1325 (N_1325,N_338,N_528);
and U1326 (N_1326,N_791,N_45);
or U1327 (N_1327,N_231,N_675);
and U1328 (N_1328,N_816,N_58);
or U1329 (N_1329,N_552,N_305);
or U1330 (N_1330,N_211,N_387);
and U1331 (N_1331,N_345,N_929);
nand U1332 (N_1332,N_195,N_320);
or U1333 (N_1333,N_874,N_732);
nand U1334 (N_1334,N_374,N_34);
or U1335 (N_1335,N_276,N_379);
or U1336 (N_1336,N_745,N_130);
xnor U1337 (N_1337,N_291,N_731);
or U1338 (N_1338,N_150,N_660);
nand U1339 (N_1339,N_300,N_13);
nor U1340 (N_1340,N_749,N_866);
or U1341 (N_1341,N_73,N_993);
and U1342 (N_1342,N_51,N_200);
nand U1343 (N_1343,N_257,N_682);
or U1344 (N_1344,N_986,N_843);
nor U1345 (N_1345,N_275,N_317);
or U1346 (N_1346,N_299,N_608);
xor U1347 (N_1347,N_777,N_902);
nor U1348 (N_1348,N_86,N_870);
nor U1349 (N_1349,N_982,N_277);
and U1350 (N_1350,N_649,N_403);
and U1351 (N_1351,N_735,N_863);
nor U1352 (N_1352,N_85,N_375);
nor U1353 (N_1353,N_188,N_776);
nand U1354 (N_1354,N_787,N_258);
or U1355 (N_1355,N_959,N_860);
and U1356 (N_1356,N_29,N_857);
nand U1357 (N_1357,N_237,N_236);
and U1358 (N_1358,N_795,N_105);
or U1359 (N_1359,N_184,N_792);
nor U1360 (N_1360,N_569,N_778);
xnor U1361 (N_1361,N_496,N_149);
or U1362 (N_1362,N_168,N_882);
nor U1363 (N_1363,N_550,N_561);
nor U1364 (N_1364,N_170,N_267);
xor U1365 (N_1365,N_981,N_664);
nand U1366 (N_1366,N_737,N_478);
and U1367 (N_1367,N_913,N_264);
xnor U1368 (N_1368,N_899,N_953);
or U1369 (N_1369,N_433,N_958);
xnor U1370 (N_1370,N_562,N_725);
or U1371 (N_1371,N_408,N_87);
nor U1372 (N_1372,N_764,N_382);
nand U1373 (N_1373,N_935,N_396);
nor U1374 (N_1374,N_434,N_350);
or U1375 (N_1375,N_128,N_518);
and U1376 (N_1376,N_52,N_256);
xnor U1377 (N_1377,N_307,N_143);
nor U1378 (N_1378,N_574,N_679);
and U1379 (N_1379,N_564,N_99);
nor U1380 (N_1380,N_348,N_280);
nor U1381 (N_1381,N_887,N_566);
or U1382 (N_1382,N_799,N_854);
and U1383 (N_1383,N_525,N_448);
nand U1384 (N_1384,N_292,N_36);
nor U1385 (N_1385,N_521,N_594);
nor U1386 (N_1386,N_229,N_210);
or U1387 (N_1387,N_748,N_915);
nand U1388 (N_1388,N_449,N_357);
nor U1389 (N_1389,N_389,N_476);
or U1390 (N_1390,N_134,N_782);
nor U1391 (N_1391,N_555,N_482);
nor U1392 (N_1392,N_423,N_597);
or U1393 (N_1393,N_812,N_71);
or U1394 (N_1394,N_232,N_81);
and U1395 (N_1395,N_890,N_968);
nor U1396 (N_1396,N_187,N_689);
nand U1397 (N_1397,N_388,N_109);
nand U1398 (N_1398,N_766,N_239);
nand U1399 (N_1399,N_159,N_822);
nand U1400 (N_1400,N_534,N_724);
nor U1401 (N_1401,N_442,N_385);
nand U1402 (N_1402,N_558,N_381);
and U1403 (N_1403,N_35,N_505);
or U1404 (N_1404,N_74,N_980);
and U1405 (N_1405,N_431,N_78);
and U1406 (N_1406,N_3,N_690);
or U1407 (N_1407,N_88,N_765);
nand U1408 (N_1408,N_707,N_301);
nor U1409 (N_1409,N_955,N_926);
or U1410 (N_1410,N_368,N_17);
nor U1411 (N_1411,N_185,N_844);
or U1412 (N_1412,N_165,N_506);
nand U1413 (N_1413,N_784,N_390);
or U1414 (N_1414,N_760,N_241);
xnor U1415 (N_1415,N_502,N_12);
nor U1416 (N_1416,N_962,N_641);
nor U1417 (N_1417,N_445,N_927);
and U1418 (N_1418,N_137,N_884);
or U1419 (N_1419,N_897,N_93);
or U1420 (N_1420,N_243,N_288);
xor U1421 (N_1421,N_708,N_651);
nor U1422 (N_1422,N_999,N_125);
or U1423 (N_1423,N_983,N_601);
nor U1424 (N_1424,N_719,N_824);
nand U1425 (N_1425,N_26,N_270);
or U1426 (N_1426,N_652,N_25);
nor U1427 (N_1427,N_709,N_907);
or U1428 (N_1428,N_998,N_56);
and U1429 (N_1429,N_207,N_810);
and U1430 (N_1430,N_931,N_779);
nand U1431 (N_1431,N_419,N_579);
nor U1432 (N_1432,N_655,N_793);
nand U1433 (N_1433,N_208,N_703);
or U1434 (N_1434,N_452,N_203);
or U1435 (N_1435,N_695,N_251);
nand U1436 (N_1436,N_473,N_785);
nor U1437 (N_1437,N_479,N_70);
and U1438 (N_1438,N_261,N_584);
nor U1439 (N_1439,N_522,N_244);
nor U1440 (N_1440,N_104,N_723);
and U1441 (N_1441,N_129,N_341);
xnor U1442 (N_1442,N_693,N_855);
nor U1443 (N_1443,N_290,N_888);
or U1444 (N_1444,N_333,N_932);
or U1445 (N_1445,N_533,N_750);
and U1446 (N_1446,N_544,N_910);
and U1447 (N_1447,N_517,N_10);
xor U1448 (N_1448,N_510,N_8);
and U1449 (N_1449,N_235,N_219);
xnor U1450 (N_1450,N_491,N_223);
xnor U1451 (N_1451,N_330,N_209);
or U1452 (N_1452,N_322,N_314);
nand U1453 (N_1453,N_940,N_64);
and U1454 (N_1454,N_297,N_775);
and U1455 (N_1455,N_186,N_97);
or U1456 (N_1456,N_828,N_531);
nand U1457 (N_1457,N_289,N_840);
or U1458 (N_1458,N_295,N_369);
or U1459 (N_1459,N_67,N_839);
nand U1460 (N_1460,N_851,N_991);
and U1461 (N_1461,N_976,N_447);
or U1462 (N_1462,N_639,N_450);
or U1463 (N_1463,N_89,N_48);
xor U1464 (N_1464,N_979,N_255);
and U1465 (N_1465,N_294,N_713);
and U1466 (N_1466,N_789,N_593);
nand U1467 (N_1467,N_18,N_222);
nor U1468 (N_1468,N_753,N_794);
or U1469 (N_1469,N_316,N_363);
and U1470 (N_1470,N_697,N_441);
nor U1471 (N_1471,N_671,N_272);
nand U1472 (N_1472,N_123,N_548);
or U1473 (N_1473,N_461,N_546);
or U1474 (N_1474,N_378,N_488);
and U1475 (N_1475,N_392,N_568);
or U1476 (N_1476,N_559,N_303);
or U1477 (N_1477,N_62,N_625);
and U1478 (N_1478,N_585,N_432);
nor U1479 (N_1479,N_877,N_994);
nor U1480 (N_1480,N_618,N_563);
nor U1481 (N_1481,N_892,N_183);
xor U1482 (N_1482,N_642,N_192);
xor U1483 (N_1483,N_823,N_916);
or U1484 (N_1484,N_711,N_437);
nor U1485 (N_1485,N_119,N_343);
nand U1486 (N_1486,N_520,N_577);
nor U1487 (N_1487,N_715,N_248);
nand U1488 (N_1488,N_739,N_757);
nand U1489 (N_1489,N_734,N_716);
nor U1490 (N_1490,N_370,N_802);
and U1491 (N_1491,N_621,N_576);
or U1492 (N_1492,N_661,N_0);
or U1493 (N_1493,N_14,N_871);
nand U1494 (N_1494,N_570,N_329);
nor U1495 (N_1495,N_722,N_511);
xor U1496 (N_1496,N_537,N_977);
or U1497 (N_1497,N_617,N_677);
nand U1498 (N_1498,N_603,N_797);
nand U1499 (N_1499,N_483,N_987);
and U1500 (N_1500,N_963,N_224);
nand U1501 (N_1501,N_580,N_810);
xnor U1502 (N_1502,N_326,N_87);
and U1503 (N_1503,N_925,N_928);
nand U1504 (N_1504,N_455,N_20);
and U1505 (N_1505,N_572,N_781);
and U1506 (N_1506,N_95,N_364);
xnor U1507 (N_1507,N_376,N_885);
nor U1508 (N_1508,N_951,N_854);
or U1509 (N_1509,N_29,N_677);
and U1510 (N_1510,N_748,N_269);
and U1511 (N_1511,N_784,N_794);
and U1512 (N_1512,N_326,N_167);
or U1513 (N_1513,N_351,N_405);
and U1514 (N_1514,N_413,N_157);
nor U1515 (N_1515,N_191,N_927);
nand U1516 (N_1516,N_93,N_791);
xor U1517 (N_1517,N_518,N_467);
nand U1518 (N_1518,N_673,N_1);
nor U1519 (N_1519,N_953,N_82);
or U1520 (N_1520,N_194,N_259);
nor U1521 (N_1521,N_615,N_944);
nor U1522 (N_1522,N_917,N_975);
nor U1523 (N_1523,N_240,N_482);
nand U1524 (N_1524,N_525,N_897);
xnor U1525 (N_1525,N_391,N_697);
and U1526 (N_1526,N_564,N_572);
nand U1527 (N_1527,N_810,N_138);
nor U1528 (N_1528,N_505,N_479);
nor U1529 (N_1529,N_655,N_70);
xor U1530 (N_1530,N_362,N_874);
nor U1531 (N_1531,N_540,N_664);
or U1532 (N_1532,N_44,N_479);
nand U1533 (N_1533,N_238,N_10);
xor U1534 (N_1534,N_713,N_912);
nor U1535 (N_1535,N_887,N_49);
and U1536 (N_1536,N_758,N_299);
nor U1537 (N_1537,N_818,N_474);
nor U1538 (N_1538,N_131,N_361);
nand U1539 (N_1539,N_946,N_185);
or U1540 (N_1540,N_382,N_994);
nor U1541 (N_1541,N_884,N_359);
nor U1542 (N_1542,N_846,N_989);
and U1543 (N_1543,N_35,N_413);
nand U1544 (N_1544,N_255,N_555);
xor U1545 (N_1545,N_614,N_736);
or U1546 (N_1546,N_890,N_412);
or U1547 (N_1547,N_141,N_692);
and U1548 (N_1548,N_113,N_134);
and U1549 (N_1549,N_207,N_556);
and U1550 (N_1550,N_202,N_979);
nand U1551 (N_1551,N_395,N_992);
or U1552 (N_1552,N_117,N_764);
or U1553 (N_1553,N_553,N_540);
and U1554 (N_1554,N_897,N_418);
and U1555 (N_1555,N_42,N_904);
or U1556 (N_1556,N_683,N_930);
and U1557 (N_1557,N_452,N_573);
nor U1558 (N_1558,N_493,N_187);
xnor U1559 (N_1559,N_595,N_785);
and U1560 (N_1560,N_581,N_867);
and U1561 (N_1561,N_803,N_833);
or U1562 (N_1562,N_309,N_90);
and U1563 (N_1563,N_822,N_969);
and U1564 (N_1564,N_245,N_243);
and U1565 (N_1565,N_281,N_47);
or U1566 (N_1566,N_86,N_651);
nand U1567 (N_1567,N_259,N_653);
nor U1568 (N_1568,N_658,N_25);
nand U1569 (N_1569,N_757,N_700);
and U1570 (N_1570,N_330,N_909);
xnor U1571 (N_1571,N_567,N_683);
nand U1572 (N_1572,N_100,N_673);
nor U1573 (N_1573,N_643,N_736);
nor U1574 (N_1574,N_545,N_810);
nor U1575 (N_1575,N_742,N_392);
or U1576 (N_1576,N_95,N_46);
nand U1577 (N_1577,N_211,N_386);
nor U1578 (N_1578,N_215,N_705);
and U1579 (N_1579,N_84,N_949);
or U1580 (N_1580,N_664,N_120);
or U1581 (N_1581,N_871,N_917);
nor U1582 (N_1582,N_755,N_699);
nor U1583 (N_1583,N_737,N_73);
nand U1584 (N_1584,N_346,N_916);
or U1585 (N_1585,N_205,N_43);
or U1586 (N_1586,N_961,N_443);
or U1587 (N_1587,N_690,N_322);
or U1588 (N_1588,N_702,N_87);
nand U1589 (N_1589,N_781,N_504);
nor U1590 (N_1590,N_127,N_208);
nand U1591 (N_1591,N_813,N_723);
and U1592 (N_1592,N_155,N_311);
and U1593 (N_1593,N_627,N_34);
nor U1594 (N_1594,N_617,N_354);
nand U1595 (N_1595,N_87,N_823);
or U1596 (N_1596,N_845,N_240);
xnor U1597 (N_1597,N_751,N_486);
nand U1598 (N_1598,N_613,N_98);
nand U1599 (N_1599,N_631,N_82);
or U1600 (N_1600,N_613,N_802);
and U1601 (N_1601,N_943,N_702);
or U1602 (N_1602,N_830,N_564);
nor U1603 (N_1603,N_748,N_830);
xor U1604 (N_1604,N_891,N_367);
and U1605 (N_1605,N_884,N_911);
xor U1606 (N_1606,N_427,N_717);
nor U1607 (N_1607,N_170,N_181);
or U1608 (N_1608,N_501,N_962);
or U1609 (N_1609,N_267,N_79);
nand U1610 (N_1610,N_74,N_955);
nor U1611 (N_1611,N_865,N_137);
and U1612 (N_1612,N_493,N_946);
xor U1613 (N_1613,N_53,N_738);
nand U1614 (N_1614,N_769,N_332);
xnor U1615 (N_1615,N_91,N_302);
nand U1616 (N_1616,N_899,N_999);
and U1617 (N_1617,N_211,N_107);
nand U1618 (N_1618,N_600,N_145);
and U1619 (N_1619,N_25,N_276);
and U1620 (N_1620,N_78,N_692);
nor U1621 (N_1621,N_553,N_614);
or U1622 (N_1622,N_173,N_495);
or U1623 (N_1623,N_404,N_202);
xnor U1624 (N_1624,N_411,N_255);
nand U1625 (N_1625,N_544,N_130);
or U1626 (N_1626,N_274,N_66);
nor U1627 (N_1627,N_821,N_705);
xor U1628 (N_1628,N_604,N_736);
or U1629 (N_1629,N_336,N_453);
nor U1630 (N_1630,N_854,N_722);
and U1631 (N_1631,N_638,N_662);
xnor U1632 (N_1632,N_586,N_118);
or U1633 (N_1633,N_266,N_197);
and U1634 (N_1634,N_709,N_62);
or U1635 (N_1635,N_286,N_838);
nand U1636 (N_1636,N_52,N_331);
and U1637 (N_1637,N_751,N_359);
nor U1638 (N_1638,N_164,N_574);
and U1639 (N_1639,N_827,N_286);
and U1640 (N_1640,N_569,N_179);
or U1641 (N_1641,N_156,N_577);
nor U1642 (N_1642,N_837,N_202);
nor U1643 (N_1643,N_227,N_305);
xnor U1644 (N_1644,N_187,N_313);
nor U1645 (N_1645,N_844,N_339);
nor U1646 (N_1646,N_452,N_249);
and U1647 (N_1647,N_137,N_890);
nor U1648 (N_1648,N_510,N_563);
nand U1649 (N_1649,N_688,N_323);
nor U1650 (N_1650,N_926,N_653);
or U1651 (N_1651,N_260,N_47);
and U1652 (N_1652,N_58,N_0);
nand U1653 (N_1653,N_123,N_676);
nor U1654 (N_1654,N_282,N_431);
nand U1655 (N_1655,N_87,N_539);
nand U1656 (N_1656,N_333,N_353);
or U1657 (N_1657,N_594,N_951);
nand U1658 (N_1658,N_290,N_921);
xnor U1659 (N_1659,N_481,N_865);
or U1660 (N_1660,N_229,N_942);
or U1661 (N_1661,N_138,N_908);
nor U1662 (N_1662,N_957,N_685);
nor U1663 (N_1663,N_790,N_220);
nor U1664 (N_1664,N_560,N_710);
nand U1665 (N_1665,N_994,N_506);
or U1666 (N_1666,N_429,N_300);
and U1667 (N_1667,N_368,N_869);
and U1668 (N_1668,N_268,N_114);
and U1669 (N_1669,N_462,N_86);
and U1670 (N_1670,N_288,N_902);
and U1671 (N_1671,N_48,N_894);
or U1672 (N_1672,N_704,N_684);
nand U1673 (N_1673,N_982,N_155);
nor U1674 (N_1674,N_965,N_738);
and U1675 (N_1675,N_652,N_342);
xnor U1676 (N_1676,N_529,N_595);
nor U1677 (N_1677,N_329,N_711);
or U1678 (N_1678,N_334,N_576);
nor U1679 (N_1679,N_576,N_865);
nor U1680 (N_1680,N_51,N_177);
and U1681 (N_1681,N_671,N_778);
and U1682 (N_1682,N_412,N_446);
or U1683 (N_1683,N_215,N_104);
or U1684 (N_1684,N_524,N_71);
or U1685 (N_1685,N_294,N_783);
or U1686 (N_1686,N_986,N_534);
xor U1687 (N_1687,N_644,N_20);
or U1688 (N_1688,N_949,N_547);
nor U1689 (N_1689,N_666,N_351);
or U1690 (N_1690,N_839,N_813);
and U1691 (N_1691,N_771,N_49);
nor U1692 (N_1692,N_892,N_130);
or U1693 (N_1693,N_110,N_52);
nor U1694 (N_1694,N_573,N_42);
nand U1695 (N_1695,N_314,N_941);
and U1696 (N_1696,N_960,N_625);
and U1697 (N_1697,N_4,N_286);
nand U1698 (N_1698,N_305,N_646);
nor U1699 (N_1699,N_479,N_888);
nand U1700 (N_1700,N_669,N_496);
nor U1701 (N_1701,N_780,N_48);
and U1702 (N_1702,N_838,N_407);
and U1703 (N_1703,N_441,N_181);
nor U1704 (N_1704,N_704,N_798);
nor U1705 (N_1705,N_669,N_482);
and U1706 (N_1706,N_203,N_937);
or U1707 (N_1707,N_457,N_546);
and U1708 (N_1708,N_163,N_911);
or U1709 (N_1709,N_152,N_2);
or U1710 (N_1710,N_56,N_376);
nand U1711 (N_1711,N_144,N_195);
or U1712 (N_1712,N_832,N_331);
nor U1713 (N_1713,N_59,N_671);
nor U1714 (N_1714,N_939,N_408);
nand U1715 (N_1715,N_968,N_683);
xnor U1716 (N_1716,N_785,N_555);
nand U1717 (N_1717,N_543,N_904);
and U1718 (N_1718,N_844,N_216);
and U1719 (N_1719,N_223,N_850);
nand U1720 (N_1720,N_974,N_736);
nor U1721 (N_1721,N_424,N_201);
nor U1722 (N_1722,N_815,N_966);
xnor U1723 (N_1723,N_838,N_453);
nand U1724 (N_1724,N_209,N_399);
or U1725 (N_1725,N_16,N_237);
and U1726 (N_1726,N_314,N_86);
or U1727 (N_1727,N_374,N_681);
or U1728 (N_1728,N_70,N_150);
nor U1729 (N_1729,N_689,N_769);
or U1730 (N_1730,N_757,N_248);
or U1731 (N_1731,N_380,N_732);
or U1732 (N_1732,N_72,N_402);
nor U1733 (N_1733,N_454,N_777);
and U1734 (N_1734,N_688,N_757);
nand U1735 (N_1735,N_684,N_99);
nor U1736 (N_1736,N_698,N_912);
or U1737 (N_1737,N_383,N_105);
nand U1738 (N_1738,N_165,N_220);
nor U1739 (N_1739,N_353,N_570);
or U1740 (N_1740,N_18,N_66);
and U1741 (N_1741,N_202,N_165);
or U1742 (N_1742,N_981,N_154);
and U1743 (N_1743,N_749,N_487);
or U1744 (N_1744,N_455,N_686);
and U1745 (N_1745,N_855,N_471);
and U1746 (N_1746,N_765,N_326);
or U1747 (N_1747,N_176,N_740);
nor U1748 (N_1748,N_145,N_200);
or U1749 (N_1749,N_677,N_307);
xnor U1750 (N_1750,N_74,N_620);
and U1751 (N_1751,N_461,N_566);
or U1752 (N_1752,N_453,N_517);
xnor U1753 (N_1753,N_126,N_322);
nand U1754 (N_1754,N_639,N_250);
nand U1755 (N_1755,N_898,N_385);
nand U1756 (N_1756,N_397,N_40);
and U1757 (N_1757,N_935,N_173);
and U1758 (N_1758,N_104,N_529);
or U1759 (N_1759,N_745,N_220);
and U1760 (N_1760,N_766,N_172);
or U1761 (N_1761,N_588,N_569);
and U1762 (N_1762,N_300,N_223);
nor U1763 (N_1763,N_65,N_600);
and U1764 (N_1764,N_657,N_183);
nor U1765 (N_1765,N_32,N_854);
xor U1766 (N_1766,N_415,N_511);
or U1767 (N_1767,N_320,N_191);
or U1768 (N_1768,N_242,N_360);
or U1769 (N_1769,N_316,N_159);
xnor U1770 (N_1770,N_235,N_160);
nand U1771 (N_1771,N_459,N_40);
nand U1772 (N_1772,N_281,N_691);
nor U1773 (N_1773,N_235,N_715);
and U1774 (N_1774,N_622,N_361);
nor U1775 (N_1775,N_118,N_266);
nor U1776 (N_1776,N_925,N_667);
and U1777 (N_1777,N_34,N_508);
nor U1778 (N_1778,N_892,N_312);
xor U1779 (N_1779,N_123,N_784);
or U1780 (N_1780,N_115,N_971);
xor U1781 (N_1781,N_284,N_824);
or U1782 (N_1782,N_194,N_121);
or U1783 (N_1783,N_911,N_172);
or U1784 (N_1784,N_846,N_616);
or U1785 (N_1785,N_675,N_404);
or U1786 (N_1786,N_609,N_601);
or U1787 (N_1787,N_973,N_659);
or U1788 (N_1788,N_176,N_615);
xnor U1789 (N_1789,N_402,N_532);
nor U1790 (N_1790,N_675,N_447);
or U1791 (N_1791,N_217,N_743);
and U1792 (N_1792,N_322,N_591);
nor U1793 (N_1793,N_968,N_762);
nand U1794 (N_1794,N_703,N_576);
nand U1795 (N_1795,N_923,N_697);
nor U1796 (N_1796,N_738,N_371);
nand U1797 (N_1797,N_39,N_465);
nand U1798 (N_1798,N_573,N_694);
xnor U1799 (N_1799,N_993,N_709);
or U1800 (N_1800,N_246,N_203);
nor U1801 (N_1801,N_797,N_708);
xnor U1802 (N_1802,N_573,N_91);
and U1803 (N_1803,N_360,N_127);
and U1804 (N_1804,N_431,N_581);
and U1805 (N_1805,N_425,N_223);
or U1806 (N_1806,N_926,N_634);
nand U1807 (N_1807,N_216,N_960);
and U1808 (N_1808,N_794,N_20);
xor U1809 (N_1809,N_449,N_599);
or U1810 (N_1810,N_464,N_514);
or U1811 (N_1811,N_325,N_954);
nand U1812 (N_1812,N_936,N_413);
xnor U1813 (N_1813,N_755,N_632);
and U1814 (N_1814,N_353,N_253);
nor U1815 (N_1815,N_178,N_666);
xnor U1816 (N_1816,N_905,N_73);
nor U1817 (N_1817,N_308,N_957);
xnor U1818 (N_1818,N_498,N_3);
nand U1819 (N_1819,N_813,N_371);
or U1820 (N_1820,N_600,N_685);
nand U1821 (N_1821,N_474,N_488);
or U1822 (N_1822,N_876,N_773);
xnor U1823 (N_1823,N_263,N_705);
nor U1824 (N_1824,N_480,N_801);
xnor U1825 (N_1825,N_386,N_438);
nand U1826 (N_1826,N_738,N_8);
nand U1827 (N_1827,N_946,N_813);
and U1828 (N_1828,N_769,N_567);
or U1829 (N_1829,N_8,N_595);
xnor U1830 (N_1830,N_232,N_124);
and U1831 (N_1831,N_434,N_432);
and U1832 (N_1832,N_878,N_765);
or U1833 (N_1833,N_950,N_809);
nand U1834 (N_1834,N_654,N_400);
or U1835 (N_1835,N_732,N_968);
xnor U1836 (N_1836,N_898,N_853);
nor U1837 (N_1837,N_809,N_129);
xor U1838 (N_1838,N_579,N_517);
and U1839 (N_1839,N_662,N_126);
or U1840 (N_1840,N_395,N_874);
or U1841 (N_1841,N_933,N_824);
nand U1842 (N_1842,N_297,N_29);
or U1843 (N_1843,N_248,N_549);
xor U1844 (N_1844,N_940,N_948);
xnor U1845 (N_1845,N_433,N_274);
or U1846 (N_1846,N_641,N_404);
nand U1847 (N_1847,N_68,N_544);
nor U1848 (N_1848,N_447,N_181);
and U1849 (N_1849,N_675,N_553);
or U1850 (N_1850,N_728,N_627);
nand U1851 (N_1851,N_759,N_551);
nor U1852 (N_1852,N_438,N_421);
nand U1853 (N_1853,N_793,N_104);
nor U1854 (N_1854,N_777,N_549);
and U1855 (N_1855,N_736,N_407);
and U1856 (N_1856,N_977,N_688);
xor U1857 (N_1857,N_806,N_285);
nor U1858 (N_1858,N_683,N_195);
and U1859 (N_1859,N_106,N_165);
and U1860 (N_1860,N_72,N_389);
nand U1861 (N_1861,N_214,N_763);
or U1862 (N_1862,N_117,N_453);
xor U1863 (N_1863,N_558,N_527);
nand U1864 (N_1864,N_784,N_228);
and U1865 (N_1865,N_140,N_968);
and U1866 (N_1866,N_85,N_238);
or U1867 (N_1867,N_383,N_785);
and U1868 (N_1868,N_82,N_635);
nand U1869 (N_1869,N_90,N_882);
or U1870 (N_1870,N_178,N_319);
xor U1871 (N_1871,N_231,N_393);
and U1872 (N_1872,N_3,N_382);
and U1873 (N_1873,N_232,N_489);
and U1874 (N_1874,N_634,N_180);
or U1875 (N_1875,N_545,N_77);
or U1876 (N_1876,N_293,N_483);
nor U1877 (N_1877,N_63,N_786);
and U1878 (N_1878,N_71,N_854);
and U1879 (N_1879,N_915,N_881);
nand U1880 (N_1880,N_345,N_825);
and U1881 (N_1881,N_780,N_86);
xor U1882 (N_1882,N_150,N_709);
nor U1883 (N_1883,N_392,N_755);
nand U1884 (N_1884,N_241,N_952);
and U1885 (N_1885,N_572,N_443);
xnor U1886 (N_1886,N_781,N_384);
and U1887 (N_1887,N_312,N_722);
xnor U1888 (N_1888,N_494,N_245);
nand U1889 (N_1889,N_743,N_998);
nor U1890 (N_1890,N_463,N_154);
xor U1891 (N_1891,N_922,N_64);
and U1892 (N_1892,N_717,N_412);
xor U1893 (N_1893,N_0,N_21);
and U1894 (N_1894,N_686,N_121);
or U1895 (N_1895,N_338,N_112);
or U1896 (N_1896,N_140,N_39);
nor U1897 (N_1897,N_525,N_602);
and U1898 (N_1898,N_804,N_305);
or U1899 (N_1899,N_340,N_198);
or U1900 (N_1900,N_92,N_429);
and U1901 (N_1901,N_346,N_334);
xor U1902 (N_1902,N_43,N_865);
and U1903 (N_1903,N_876,N_772);
nor U1904 (N_1904,N_239,N_740);
nand U1905 (N_1905,N_928,N_922);
and U1906 (N_1906,N_180,N_384);
or U1907 (N_1907,N_723,N_637);
or U1908 (N_1908,N_719,N_942);
nand U1909 (N_1909,N_199,N_428);
or U1910 (N_1910,N_353,N_290);
nand U1911 (N_1911,N_575,N_778);
or U1912 (N_1912,N_578,N_264);
nand U1913 (N_1913,N_875,N_606);
and U1914 (N_1914,N_389,N_285);
nand U1915 (N_1915,N_483,N_856);
xor U1916 (N_1916,N_96,N_169);
nor U1917 (N_1917,N_524,N_552);
nor U1918 (N_1918,N_999,N_897);
nand U1919 (N_1919,N_644,N_483);
xor U1920 (N_1920,N_507,N_67);
or U1921 (N_1921,N_242,N_478);
or U1922 (N_1922,N_151,N_518);
nand U1923 (N_1923,N_325,N_213);
or U1924 (N_1924,N_6,N_869);
and U1925 (N_1925,N_833,N_595);
or U1926 (N_1926,N_336,N_953);
xnor U1927 (N_1927,N_716,N_992);
nor U1928 (N_1928,N_68,N_218);
xnor U1929 (N_1929,N_220,N_15);
or U1930 (N_1930,N_631,N_339);
and U1931 (N_1931,N_234,N_723);
nand U1932 (N_1932,N_222,N_565);
and U1933 (N_1933,N_437,N_664);
nand U1934 (N_1934,N_588,N_877);
or U1935 (N_1935,N_887,N_64);
and U1936 (N_1936,N_638,N_461);
and U1937 (N_1937,N_472,N_668);
and U1938 (N_1938,N_953,N_340);
xnor U1939 (N_1939,N_807,N_176);
nand U1940 (N_1940,N_264,N_226);
nor U1941 (N_1941,N_790,N_170);
nor U1942 (N_1942,N_613,N_896);
nand U1943 (N_1943,N_16,N_931);
and U1944 (N_1944,N_542,N_88);
nand U1945 (N_1945,N_238,N_264);
xor U1946 (N_1946,N_103,N_656);
nor U1947 (N_1947,N_612,N_550);
nor U1948 (N_1948,N_111,N_215);
or U1949 (N_1949,N_174,N_135);
nor U1950 (N_1950,N_138,N_84);
nor U1951 (N_1951,N_919,N_446);
and U1952 (N_1952,N_818,N_865);
or U1953 (N_1953,N_783,N_727);
and U1954 (N_1954,N_247,N_756);
nand U1955 (N_1955,N_307,N_279);
and U1956 (N_1956,N_698,N_490);
or U1957 (N_1957,N_594,N_586);
xor U1958 (N_1958,N_383,N_700);
nand U1959 (N_1959,N_228,N_188);
nor U1960 (N_1960,N_151,N_801);
and U1961 (N_1961,N_201,N_104);
and U1962 (N_1962,N_898,N_716);
or U1963 (N_1963,N_139,N_227);
or U1964 (N_1964,N_727,N_140);
or U1965 (N_1965,N_969,N_794);
and U1966 (N_1966,N_730,N_381);
nor U1967 (N_1967,N_980,N_855);
nand U1968 (N_1968,N_405,N_33);
nand U1969 (N_1969,N_59,N_740);
and U1970 (N_1970,N_251,N_907);
xnor U1971 (N_1971,N_528,N_979);
nand U1972 (N_1972,N_180,N_356);
and U1973 (N_1973,N_556,N_153);
nand U1974 (N_1974,N_850,N_750);
nand U1975 (N_1975,N_684,N_573);
or U1976 (N_1976,N_350,N_59);
or U1977 (N_1977,N_180,N_550);
nand U1978 (N_1978,N_881,N_585);
or U1979 (N_1979,N_246,N_670);
or U1980 (N_1980,N_625,N_243);
nor U1981 (N_1981,N_293,N_806);
xnor U1982 (N_1982,N_613,N_314);
xor U1983 (N_1983,N_744,N_295);
xnor U1984 (N_1984,N_215,N_742);
and U1985 (N_1985,N_22,N_754);
and U1986 (N_1986,N_429,N_487);
or U1987 (N_1987,N_423,N_871);
xor U1988 (N_1988,N_428,N_835);
or U1989 (N_1989,N_442,N_957);
nor U1990 (N_1990,N_574,N_654);
xnor U1991 (N_1991,N_452,N_407);
xor U1992 (N_1992,N_203,N_144);
nor U1993 (N_1993,N_771,N_328);
nand U1994 (N_1994,N_758,N_389);
nor U1995 (N_1995,N_745,N_809);
and U1996 (N_1996,N_412,N_4);
or U1997 (N_1997,N_114,N_555);
and U1998 (N_1998,N_884,N_243);
or U1999 (N_1999,N_738,N_84);
nor U2000 (N_2000,N_1071,N_1237);
nand U2001 (N_2001,N_1040,N_1406);
xnor U2002 (N_2002,N_1060,N_1990);
nor U2003 (N_2003,N_1612,N_1076);
or U2004 (N_2004,N_1368,N_1678);
nor U2005 (N_2005,N_1572,N_1426);
xor U2006 (N_2006,N_1552,N_1641);
nand U2007 (N_2007,N_1998,N_1831);
and U2008 (N_2008,N_1110,N_1282);
xor U2009 (N_2009,N_1954,N_1232);
nor U2010 (N_2010,N_1058,N_1116);
nor U2011 (N_2011,N_1720,N_1752);
and U2012 (N_2012,N_1979,N_1953);
nand U2013 (N_2013,N_1545,N_1035);
and U2014 (N_2014,N_1689,N_1947);
and U2015 (N_2015,N_1622,N_1288);
nor U2016 (N_2016,N_1492,N_1475);
and U2017 (N_2017,N_1878,N_1699);
or U2018 (N_2018,N_1049,N_1790);
nor U2019 (N_2019,N_1412,N_1117);
and U2020 (N_2020,N_1774,N_1201);
or U2021 (N_2021,N_1263,N_1649);
nand U2022 (N_2022,N_1149,N_1765);
nand U2023 (N_2023,N_1322,N_1051);
or U2024 (N_2024,N_1369,N_1984);
nor U2025 (N_2025,N_1348,N_1888);
nor U2026 (N_2026,N_1815,N_1440);
nor U2027 (N_2027,N_1850,N_1827);
nor U2028 (N_2028,N_1949,N_1208);
or U2029 (N_2029,N_1745,N_1472);
xor U2030 (N_2030,N_1046,N_1707);
and U2031 (N_2031,N_1402,N_1166);
or U2032 (N_2032,N_1659,N_1638);
or U2033 (N_2033,N_1764,N_1628);
nor U2034 (N_2034,N_1653,N_1303);
and U2035 (N_2035,N_1000,N_1889);
nand U2036 (N_2036,N_1528,N_1523);
nor U2037 (N_2037,N_1977,N_1449);
nor U2038 (N_2038,N_1045,N_1775);
nor U2039 (N_2039,N_1967,N_1608);
or U2040 (N_2040,N_1724,N_1456);
nand U2041 (N_2041,N_1769,N_1909);
or U2042 (N_2042,N_1531,N_1139);
nor U2043 (N_2043,N_1511,N_1673);
and U2044 (N_2044,N_1065,N_1665);
nand U2045 (N_2045,N_1395,N_1399);
or U2046 (N_2046,N_1454,N_1924);
nand U2047 (N_2047,N_1107,N_1778);
nor U2048 (N_2048,N_1017,N_1494);
nor U2049 (N_2049,N_1258,N_1372);
nand U2050 (N_2050,N_1508,N_1662);
and U2051 (N_2051,N_1078,N_1739);
nand U2052 (N_2052,N_1112,N_1548);
nor U2053 (N_2053,N_1129,N_1427);
or U2054 (N_2054,N_1629,N_1123);
nor U2055 (N_2055,N_1347,N_1230);
nor U2056 (N_2056,N_1184,N_1124);
nor U2057 (N_2057,N_1316,N_1679);
and U2058 (N_2058,N_1816,N_1398);
xor U2059 (N_2059,N_1863,N_1580);
or U2060 (N_2060,N_1565,N_1926);
nand U2061 (N_2061,N_1175,N_1377);
or U2062 (N_2062,N_1593,N_1259);
nand U2063 (N_2063,N_1703,N_1605);
or U2064 (N_2064,N_1906,N_1877);
or U2065 (N_2065,N_1595,N_1599);
nor U2066 (N_2066,N_1932,N_1442);
and U2067 (N_2067,N_1274,N_1709);
and U2068 (N_2068,N_1457,N_1003);
nor U2069 (N_2069,N_1293,N_1776);
nand U2070 (N_2070,N_1610,N_1483);
xnor U2071 (N_2071,N_1140,N_1178);
nor U2072 (N_2072,N_1247,N_1225);
and U2073 (N_2073,N_1052,N_1213);
nand U2074 (N_2074,N_1180,N_1591);
or U2075 (N_2075,N_1154,N_1798);
or U2076 (N_2076,N_1200,N_1023);
or U2077 (N_2077,N_1019,N_1471);
xor U2078 (N_2078,N_1872,N_1385);
nor U2079 (N_2079,N_1683,N_1105);
nor U2080 (N_2080,N_1787,N_1537);
nor U2081 (N_2081,N_1323,N_1777);
nand U2082 (N_2082,N_1391,N_1711);
nor U2083 (N_2083,N_1940,N_1148);
xnor U2084 (N_2084,N_1246,N_1820);
nor U2085 (N_2085,N_1946,N_1310);
and U2086 (N_2086,N_1205,N_1186);
and U2087 (N_2087,N_1069,N_1054);
nor U2088 (N_2088,N_1895,N_1285);
nor U2089 (N_2089,N_1617,N_1841);
nor U2090 (N_2090,N_1750,N_1064);
or U2091 (N_2091,N_1788,N_1174);
or U2092 (N_2092,N_1725,N_1055);
or U2093 (N_2093,N_1738,N_1497);
and U2094 (N_2094,N_1854,N_1858);
xnor U2095 (N_2095,N_1267,N_1829);
and U2096 (N_2096,N_1417,N_1448);
and U2097 (N_2097,N_1428,N_1957);
or U2098 (N_2098,N_1460,N_1084);
nor U2099 (N_2099,N_1606,N_1630);
xnor U2100 (N_2100,N_1340,N_1011);
nor U2101 (N_2101,N_1163,N_1309);
or U2102 (N_2102,N_1283,N_1128);
nand U2103 (N_2103,N_1644,N_1042);
nor U2104 (N_2104,N_1009,N_1740);
or U2105 (N_2105,N_1190,N_1435);
nor U2106 (N_2106,N_1031,N_1748);
and U2107 (N_2107,N_1873,N_1639);
nand U2108 (N_2108,N_1362,N_1592);
and U2109 (N_2109,N_1164,N_1618);
or U2110 (N_2110,N_1900,N_1389);
nand U2111 (N_2111,N_1634,N_1539);
or U2112 (N_2112,N_1423,N_1091);
xor U2113 (N_2113,N_1027,N_1640);
or U2114 (N_2114,N_1373,N_1999);
nand U2115 (N_2115,N_1083,N_1532);
or U2116 (N_2116,N_1431,N_1991);
or U2117 (N_2117,N_1575,N_1536);
and U2118 (N_2118,N_1062,N_1546);
nand U2119 (N_2119,N_1498,N_1302);
nand U2120 (N_2120,N_1378,N_1603);
and U2121 (N_2121,N_1944,N_1367);
and U2122 (N_2122,N_1292,N_1446);
nand U2123 (N_2123,N_1419,N_1624);
nor U2124 (N_2124,N_1966,N_1680);
nand U2125 (N_2125,N_1196,N_1059);
or U2126 (N_2126,N_1266,N_1847);
and U2127 (N_2127,N_1884,N_1681);
nor U2128 (N_2128,N_1008,N_1929);
xor U2129 (N_2129,N_1490,N_1988);
nand U2130 (N_2130,N_1682,N_1613);
and U2131 (N_2131,N_1321,N_1963);
and U2132 (N_2132,N_1094,N_1138);
nand U2133 (N_2133,N_1611,N_1692);
nor U2134 (N_2134,N_1474,N_1666);
xor U2135 (N_2135,N_1482,N_1082);
and U2136 (N_2136,N_1239,N_1095);
nand U2137 (N_2137,N_1501,N_1315);
nand U2138 (N_2138,N_1969,N_1115);
or U2139 (N_2139,N_1080,N_1466);
and U2140 (N_2140,N_1325,N_1358);
xnor U2141 (N_2141,N_1330,N_1899);
nand U2142 (N_2142,N_1824,N_1789);
nor U2143 (N_2143,N_1210,N_1403);
xor U2144 (N_2144,N_1708,N_1136);
nand U2145 (N_2145,N_1228,N_1014);
xor U2146 (N_2146,N_1207,N_1874);
or U2147 (N_2147,N_1422,N_1041);
and U2148 (N_2148,N_1652,N_1749);
nand U2149 (N_2149,N_1733,N_1307);
xnor U2150 (N_2150,N_1028,N_1951);
or U2151 (N_2151,N_1212,N_1254);
nand U2152 (N_2152,N_1390,N_1029);
nand U2153 (N_2153,N_1279,N_1505);
and U2154 (N_2154,N_1549,N_1530);
nor U2155 (N_2155,N_1182,N_1919);
or U2156 (N_2156,N_1560,N_1363);
and U2157 (N_2157,N_1300,N_1382);
and U2158 (N_2158,N_1981,N_1381);
or U2159 (N_2159,N_1489,N_1890);
and U2160 (N_2160,N_1291,N_1146);
nand U2161 (N_2161,N_1849,N_1360);
nand U2162 (N_2162,N_1231,N_1693);
nor U2163 (N_2163,N_1277,N_1500);
nor U2164 (N_2164,N_1394,N_1936);
and U2165 (N_2165,N_1879,N_1473);
or U2166 (N_2166,N_1928,N_1913);
nand U2167 (N_2167,N_1920,N_1584);
nand U2168 (N_2168,N_1862,N_1719);
or U2169 (N_2169,N_1766,N_1507);
or U2170 (N_2170,N_1102,N_1783);
xnor U2171 (N_2171,N_1521,N_1865);
nand U2172 (N_2172,N_1660,N_1432);
xnor U2173 (N_2173,N_1597,N_1669);
or U2174 (N_2174,N_1127,N_1677);
and U2175 (N_2175,N_1939,N_1852);
or U2176 (N_2176,N_1965,N_1415);
and U2177 (N_2177,N_1686,N_1836);
and U2178 (N_2178,N_1077,N_1098);
nand U2179 (N_2179,N_1276,N_1491);
xor U2180 (N_2180,N_1173,N_1756);
xor U2181 (N_2181,N_1903,N_1700);
and U2182 (N_2182,N_1192,N_1336);
and U2183 (N_2183,N_1509,N_1063);
nand U2184 (N_2184,N_1219,N_1941);
nor U2185 (N_2185,N_1972,N_1897);
nor U2186 (N_2186,N_1244,N_1452);
and U2187 (N_2187,N_1499,N_1418);
nor U2188 (N_2188,N_1637,N_1758);
nor U2189 (N_2189,N_1633,N_1604);
or U2190 (N_2190,N_1021,N_1191);
nor U2191 (N_2191,N_1642,N_1131);
nor U2192 (N_2192,N_1943,N_1596);
nand U2193 (N_2193,N_1864,N_1444);
and U2194 (N_2194,N_1187,N_1251);
nand U2195 (N_2195,N_1664,N_1761);
nand U2196 (N_2196,N_1918,N_1762);
nand U2197 (N_2197,N_1488,N_1631);
nor U2198 (N_2198,N_1656,N_1355);
nand U2199 (N_2199,N_1807,N_1317);
and U2200 (N_2200,N_1671,N_1024);
or U2201 (N_2201,N_1731,N_1741);
or U2202 (N_2202,N_1632,N_1968);
nand U2203 (N_2203,N_1512,N_1645);
nor U2204 (N_2204,N_1695,N_1485);
nand U2205 (N_2205,N_1691,N_1085);
and U2206 (N_2206,N_1704,N_1496);
nor U2207 (N_2207,N_1275,N_1722);
and U2208 (N_2208,N_1272,N_1875);
nand U2209 (N_2209,N_1757,N_1713);
and U2210 (N_2210,N_1238,N_1882);
nand U2211 (N_2211,N_1171,N_1694);
nor U2212 (N_2212,N_1667,N_1141);
nor U2213 (N_2213,N_1464,N_1945);
or U2214 (N_2214,N_1948,N_1760);
or U2215 (N_2215,N_1635,N_1338);
xnor U2216 (N_2216,N_1763,N_1142);
and U2217 (N_2217,N_1737,N_1516);
xnor U2218 (N_2218,N_1675,N_1155);
or U2219 (N_2219,N_1144,N_1840);
nand U2220 (N_2220,N_1996,N_1157);
nor U2221 (N_2221,N_1623,N_1006);
xor U2222 (N_2222,N_1172,N_1281);
and U2223 (N_2223,N_1455,N_1411);
nor U2224 (N_2224,N_1795,N_1318);
and U2225 (N_2225,N_1688,N_1794);
or U2226 (N_2226,N_1755,N_1962);
and U2227 (N_2227,N_1843,N_1992);
or U2228 (N_2228,N_1135,N_1844);
or U2229 (N_2229,N_1329,N_1600);
nand U2230 (N_2230,N_1893,N_1493);
or U2231 (N_2231,N_1658,N_1320);
nor U2232 (N_2232,N_1197,N_1598);
nand U2233 (N_2233,N_1371,N_1621);
xor U2234 (N_2234,N_1925,N_1594);
nand U2235 (N_2235,N_1746,N_1562);
nor U2236 (N_2236,N_1100,N_1696);
nand U2237 (N_2237,N_1170,N_1535);
nor U2238 (N_2238,N_1480,N_1469);
nor U2239 (N_2239,N_1551,N_1033);
nor U2240 (N_2240,N_1721,N_1313);
or U2241 (N_2241,N_1066,N_1147);
nor U2242 (N_2242,N_1927,N_1993);
or U2243 (N_2243,N_1985,N_1802);
nand U2244 (N_2244,N_1384,N_1233);
or U2245 (N_2245,N_1034,N_1013);
or U2246 (N_2246,N_1159,N_1930);
nand U2247 (N_2247,N_1072,N_1352);
nand U2248 (N_2248,N_1183,N_1162);
nand U2249 (N_2249,N_1801,N_1436);
and U2250 (N_2250,N_1911,N_1216);
and U2251 (N_2251,N_1477,N_1445);
nor U2252 (N_2252,N_1269,N_1821);
and U2253 (N_2253,N_1533,N_1273);
nand U2254 (N_2254,N_1414,N_1383);
or U2255 (N_2255,N_1299,N_1010);
or U2256 (N_2256,N_1817,N_1767);
nand U2257 (N_2257,N_1994,N_1312);
and U2258 (N_2258,N_1204,N_1554);
nor U2259 (N_2259,N_1447,N_1294);
and U2260 (N_2260,N_1881,N_1375);
nand U2261 (N_2261,N_1169,N_1942);
nand U2262 (N_2262,N_1915,N_1038);
or U2263 (N_2263,N_1380,N_1161);
nand U2264 (N_2264,N_1995,N_1870);
or U2265 (N_2265,N_1729,N_1295);
and U2266 (N_2266,N_1518,N_1822);
nor U2267 (N_2267,N_1754,N_1253);
nand U2268 (N_2268,N_1438,N_1022);
or U2269 (N_2269,N_1120,N_1643);
nor U2270 (N_2270,N_1674,N_1855);
nor U2271 (N_2271,N_1566,N_1458);
and U2272 (N_2272,N_1811,N_1651);
xnor U2273 (N_2273,N_1654,N_1487);
and U2274 (N_2274,N_1958,N_1796);
nor U2275 (N_2275,N_1089,N_1647);
nand U2276 (N_2276,N_1346,N_1558);
xor U2277 (N_2277,N_1826,N_1068);
nand U2278 (N_2278,N_1564,N_1809);
or U2279 (N_2279,N_1194,N_1217);
nand U2280 (N_2280,N_1308,N_1079);
and U2281 (N_2281,N_1868,N_1479);
nand U2282 (N_2282,N_1590,N_1048);
nor U2283 (N_2283,N_1751,N_1910);
nor U2284 (N_2284,N_1241,N_1938);
and U2285 (N_2285,N_1718,N_1914);
and U2286 (N_2286,N_1952,N_1387);
or U2287 (N_2287,N_1086,N_1289);
or U2288 (N_2288,N_1478,N_1133);
nor U2289 (N_2289,N_1090,N_1176);
and U2290 (N_2290,N_1211,N_1986);
or U2291 (N_2291,N_1121,N_1401);
xnor U2292 (N_2292,N_1736,N_1887);
and U2293 (N_2293,N_1353,N_1290);
and U2294 (N_2294,N_1734,N_1366);
and U2295 (N_2295,N_1328,N_1556);
nor U2296 (N_2296,N_1715,N_1252);
or U2297 (N_2297,N_1262,N_1143);
and U2298 (N_2298,N_1744,N_1810);
and U2299 (N_2299,N_1278,N_1931);
and U2300 (N_2300,N_1583,N_1341);
and U2301 (N_2301,N_1015,N_1203);
nor U2302 (N_2302,N_1574,N_1800);
xor U2303 (N_2303,N_1607,N_1663);
or U2304 (N_2304,N_1894,N_1343);
xnor U2305 (N_2305,N_1921,N_1588);
or U2306 (N_2306,N_1030,N_1805);
nor U2307 (N_2307,N_1209,N_1134);
xor U2308 (N_2308,N_1514,N_1037);
xor U2309 (N_2309,N_1502,N_1772);
and U2310 (N_2310,N_1917,N_1356);
and U2311 (N_2311,N_1495,N_1793);
nand U2312 (N_2312,N_1421,N_1032);
or U2313 (N_2313,N_1185,N_1525);
xor U2314 (N_2314,N_1544,N_1297);
nor U2315 (N_2315,N_1886,N_1818);
nand U2316 (N_2316,N_1132,N_1450);
and U2317 (N_2317,N_1109,N_1687);
xor U2318 (N_2318,N_1576,N_1020);
nor U2319 (N_2319,N_1335,N_1898);
nand U2320 (N_2320,N_1425,N_1825);
and U2321 (N_2321,N_1408,N_1710);
and U2322 (N_2322,N_1304,N_1959);
or U2323 (N_2323,N_1370,N_1056);
and U2324 (N_2324,N_1242,N_1908);
and U2325 (N_2325,N_1214,N_1803);
nor U2326 (N_2326,N_1527,N_1036);
nor U2327 (N_2327,N_1467,N_1570);
and U2328 (N_2328,N_1424,N_1188);
nand U2329 (N_2329,N_1627,N_1301);
nor U2330 (N_2330,N_1812,N_1547);
or U2331 (N_2331,N_1202,N_1240);
and U2332 (N_2332,N_1326,N_1255);
nand U2333 (N_2333,N_1344,N_1983);
or U2334 (N_2334,N_1108,N_1506);
nor U2335 (N_2335,N_1218,N_1782);
or U2336 (N_2336,N_1626,N_1484);
nor U2337 (N_2337,N_1397,N_1876);
and U2338 (N_2338,N_1451,N_1937);
or U2339 (N_2339,N_1221,N_1961);
or U2340 (N_2340,N_1250,N_1950);
and U2341 (N_2341,N_1130,N_1561);
nand U2342 (N_2342,N_1337,N_1223);
nor U2343 (N_2343,N_1160,N_1256);
nor U2344 (N_2344,N_1759,N_1248);
and U2345 (N_2345,N_1327,N_1193);
nand U2346 (N_2346,N_1672,N_1785);
nand U2347 (N_2347,N_1851,N_1111);
and U2348 (N_2348,N_1268,N_1018);
nand U2349 (N_2349,N_1837,N_1571);
or U2350 (N_2350,N_1074,N_1177);
and U2351 (N_2351,N_1698,N_1061);
nor U2352 (N_2352,N_1792,N_1075);
or U2353 (N_2353,N_1122,N_1465);
and U2354 (N_2354,N_1092,N_1043);
and U2355 (N_2355,N_1270,N_1839);
nor U2356 (N_2356,N_1434,N_1459);
nor U2357 (N_2357,N_1860,N_1589);
nor U2358 (N_2358,N_1916,N_1025);
nor U2359 (N_2359,N_1206,N_1265);
nor U2360 (N_2360,N_1298,N_1980);
nor U2361 (N_2361,N_1376,N_1437);
and U2362 (N_2362,N_1838,N_1264);
xnor U2363 (N_2363,N_1819,N_1413);
nor U2364 (N_2364,N_1016,N_1386);
or U2365 (N_2365,N_1165,N_1705);
nand U2366 (N_2366,N_1339,N_1541);
xor U2367 (N_2367,N_1296,N_1396);
nor U2368 (N_2368,N_1728,N_1410);
or U2369 (N_2369,N_1797,N_1567);
nor U2370 (N_2370,N_1093,N_1004);
and U2371 (N_2371,N_1158,N_1892);
xor U2372 (N_2372,N_1405,N_1234);
nand U2373 (N_2373,N_1620,N_1880);
or U2374 (N_2374,N_1409,N_1615);
nand U2375 (N_2375,N_1732,N_1747);
xnor U2376 (N_2376,N_1706,N_1334);
or U2377 (N_2377,N_1463,N_1503);
nand U2378 (N_2378,N_1476,N_1830);
or U2379 (N_2379,N_1104,N_1646);
or U2380 (N_2380,N_1784,N_1902);
nand U2381 (N_2381,N_1717,N_1280);
nand U2382 (N_2382,N_1891,N_1319);
nor U2383 (N_2383,N_1271,N_1901);
and U2384 (N_2384,N_1520,N_1771);
nor U2385 (N_2385,N_1430,N_1354);
nand U2386 (N_2386,N_1388,N_1439);
or U2387 (N_2387,N_1702,N_1780);
and U2388 (N_2388,N_1859,N_1832);
nand U2389 (N_2389,N_1374,N_1861);
or U2390 (N_2390,N_1614,N_1668);
or U2391 (N_2391,N_1150,N_1249);
xor U2392 (N_2392,N_1260,N_1716);
nand U2393 (N_2393,N_1625,N_1103);
or U2394 (N_2394,N_1226,N_1168);
or U2395 (N_2395,N_1609,N_1619);
or U2396 (N_2396,N_1806,N_1753);
nand U2397 (N_2397,N_1845,N_1126);
and U2398 (N_2398,N_1462,N_1723);
nand U2399 (N_2399,N_1770,N_1578);
xnor U2400 (N_2400,N_1441,N_1684);
or U2401 (N_2401,N_1224,N_1311);
nand U2402 (N_2402,N_1714,N_1236);
or U2403 (N_2403,N_1586,N_1922);
xnor U2404 (N_2404,N_1935,N_1470);
nand U2405 (N_2405,N_1791,N_1198);
nor U2406 (N_2406,N_1151,N_1057);
nand U2407 (N_2407,N_1987,N_1834);
nand U2408 (N_2408,N_1510,N_1883);
nor U2409 (N_2409,N_1853,N_1542);
or U2410 (N_2410,N_1429,N_1529);
nand U2411 (N_2411,N_1885,N_1314);
and U2412 (N_2412,N_1114,N_1361);
or U2413 (N_2413,N_1676,N_1912);
or U2414 (N_2414,N_1960,N_1044);
and U2415 (N_2415,N_1357,N_1039);
and U2416 (N_2416,N_1235,N_1848);
or U2417 (N_2417,N_1543,N_1726);
or U2418 (N_2418,N_1522,N_1538);
or U2419 (N_2419,N_1661,N_1690);
or U2420 (N_2420,N_1743,N_1420);
nor U2421 (N_2421,N_1324,N_1828);
xnor U2422 (N_2422,N_1835,N_1181);
nor U2423 (N_2423,N_1359,N_1416);
nor U2424 (N_2424,N_1975,N_1125);
nor U2425 (N_2425,N_1342,N_1650);
and U2426 (N_2426,N_1768,N_1167);
xor U2427 (N_2427,N_1305,N_1005);
and U2428 (N_2428,N_1443,N_1730);
nor U2429 (N_2429,N_1101,N_1550);
nand U2430 (N_2430,N_1997,N_1814);
and U2431 (N_2431,N_1587,N_1517);
xor U2432 (N_2432,N_1284,N_1067);
nand U2433 (N_2433,N_1365,N_1735);
or U2434 (N_2434,N_1907,N_1227);
nand U2435 (N_2435,N_1199,N_1026);
or U2436 (N_2436,N_1976,N_1287);
nand U2437 (N_2437,N_1786,N_1779);
xnor U2438 (N_2438,N_1773,N_1113);
nand U2439 (N_2439,N_1559,N_1156);
and U2440 (N_2440,N_1616,N_1804);
and U2441 (N_2441,N_1012,N_1602);
xnor U2442 (N_2442,N_1842,N_1670);
and U2443 (N_2443,N_1364,N_1582);
nor U2444 (N_2444,N_1070,N_1867);
nand U2445 (N_2445,N_1229,N_1971);
or U2446 (N_2446,N_1195,N_1964);
and U2447 (N_2447,N_1153,N_1351);
nand U2448 (N_2448,N_1306,N_1978);
nor U2449 (N_2449,N_1515,N_1137);
and U2450 (N_2450,N_1220,N_1982);
nor U2451 (N_2451,N_1569,N_1392);
or U2452 (N_2452,N_1513,N_1823);
nor U2453 (N_2453,N_1856,N_1896);
xnor U2454 (N_2454,N_1697,N_1097);
nand U2455 (N_2455,N_1563,N_1453);
xnor U2456 (N_2456,N_1286,N_1257);
nand U2457 (N_2457,N_1002,N_1973);
or U2458 (N_2458,N_1433,N_1581);
and U2459 (N_2459,N_1379,N_1050);
xnor U2460 (N_2460,N_1519,N_1096);
or U2461 (N_2461,N_1648,N_1970);
or U2462 (N_2462,N_1577,N_1087);
nor U2463 (N_2463,N_1573,N_1557);
nand U2464 (N_2464,N_1243,N_1081);
xor U2465 (N_2465,N_1106,N_1261);
nor U2466 (N_2466,N_1869,N_1727);
xnor U2467 (N_2467,N_1486,N_1345);
and U2468 (N_2468,N_1904,N_1400);
xnor U2469 (N_2469,N_1701,N_1119);
nand U2470 (N_2470,N_1152,N_1657);
nand U2471 (N_2471,N_1332,N_1934);
and U2472 (N_2472,N_1866,N_1504);
nor U2473 (N_2473,N_1933,N_1407);
and U2474 (N_2474,N_1179,N_1685);
xnor U2475 (N_2475,N_1846,N_1601);
nor U2476 (N_2476,N_1540,N_1808);
or U2477 (N_2477,N_1579,N_1568);
nor U2478 (N_2478,N_1333,N_1461);
or U2479 (N_2479,N_1813,N_1923);
nand U2480 (N_2480,N_1534,N_1007);
nor U2481 (N_2481,N_1393,N_1955);
or U2482 (N_2482,N_1871,N_1245);
nor U2483 (N_2483,N_1553,N_1073);
and U2484 (N_2484,N_1118,N_1088);
nor U2485 (N_2485,N_1585,N_1742);
or U2486 (N_2486,N_1468,N_1145);
and U2487 (N_2487,N_1404,N_1555);
xor U2488 (N_2488,N_1857,N_1047);
and U2489 (N_2489,N_1781,N_1215);
nor U2490 (N_2490,N_1481,N_1974);
nand U2491 (N_2491,N_1524,N_1526);
or U2492 (N_2492,N_1099,N_1956);
nand U2493 (N_2493,N_1001,N_1833);
and U2494 (N_2494,N_1712,N_1636);
xor U2495 (N_2495,N_1189,N_1222);
or U2496 (N_2496,N_1350,N_1799);
nand U2497 (N_2497,N_1655,N_1989);
xor U2498 (N_2498,N_1905,N_1349);
nand U2499 (N_2499,N_1331,N_1053);
nand U2500 (N_2500,N_1752,N_1753);
nor U2501 (N_2501,N_1330,N_1870);
xor U2502 (N_2502,N_1991,N_1769);
and U2503 (N_2503,N_1278,N_1292);
and U2504 (N_2504,N_1763,N_1667);
nand U2505 (N_2505,N_1627,N_1537);
and U2506 (N_2506,N_1462,N_1550);
nand U2507 (N_2507,N_1566,N_1338);
nand U2508 (N_2508,N_1064,N_1027);
nand U2509 (N_2509,N_1893,N_1032);
xnor U2510 (N_2510,N_1730,N_1585);
or U2511 (N_2511,N_1950,N_1580);
nor U2512 (N_2512,N_1233,N_1153);
nor U2513 (N_2513,N_1901,N_1247);
nand U2514 (N_2514,N_1633,N_1037);
nand U2515 (N_2515,N_1794,N_1313);
or U2516 (N_2516,N_1966,N_1216);
nor U2517 (N_2517,N_1943,N_1231);
xor U2518 (N_2518,N_1693,N_1111);
and U2519 (N_2519,N_1345,N_1863);
nor U2520 (N_2520,N_1237,N_1772);
nand U2521 (N_2521,N_1801,N_1096);
nor U2522 (N_2522,N_1728,N_1061);
nor U2523 (N_2523,N_1750,N_1150);
nand U2524 (N_2524,N_1619,N_1383);
nand U2525 (N_2525,N_1104,N_1980);
xor U2526 (N_2526,N_1860,N_1380);
nor U2527 (N_2527,N_1470,N_1816);
xnor U2528 (N_2528,N_1187,N_1988);
nor U2529 (N_2529,N_1788,N_1333);
or U2530 (N_2530,N_1092,N_1882);
nand U2531 (N_2531,N_1606,N_1133);
and U2532 (N_2532,N_1948,N_1215);
nor U2533 (N_2533,N_1413,N_1671);
xor U2534 (N_2534,N_1756,N_1955);
or U2535 (N_2535,N_1926,N_1781);
xnor U2536 (N_2536,N_1742,N_1494);
or U2537 (N_2537,N_1331,N_1169);
nor U2538 (N_2538,N_1928,N_1580);
or U2539 (N_2539,N_1063,N_1779);
and U2540 (N_2540,N_1574,N_1609);
nor U2541 (N_2541,N_1862,N_1354);
nand U2542 (N_2542,N_1029,N_1523);
nand U2543 (N_2543,N_1050,N_1212);
or U2544 (N_2544,N_1831,N_1199);
nor U2545 (N_2545,N_1506,N_1888);
and U2546 (N_2546,N_1149,N_1321);
nand U2547 (N_2547,N_1588,N_1965);
and U2548 (N_2548,N_1758,N_1213);
or U2549 (N_2549,N_1358,N_1659);
nand U2550 (N_2550,N_1417,N_1581);
nand U2551 (N_2551,N_1360,N_1071);
and U2552 (N_2552,N_1680,N_1419);
and U2553 (N_2553,N_1325,N_1311);
and U2554 (N_2554,N_1973,N_1571);
or U2555 (N_2555,N_1261,N_1896);
xnor U2556 (N_2556,N_1772,N_1647);
or U2557 (N_2557,N_1360,N_1583);
nand U2558 (N_2558,N_1922,N_1246);
nor U2559 (N_2559,N_1273,N_1266);
and U2560 (N_2560,N_1524,N_1162);
and U2561 (N_2561,N_1429,N_1330);
or U2562 (N_2562,N_1561,N_1342);
or U2563 (N_2563,N_1426,N_1095);
or U2564 (N_2564,N_1726,N_1422);
or U2565 (N_2565,N_1283,N_1606);
and U2566 (N_2566,N_1575,N_1139);
nor U2567 (N_2567,N_1055,N_1317);
nand U2568 (N_2568,N_1893,N_1428);
or U2569 (N_2569,N_1417,N_1252);
nor U2570 (N_2570,N_1638,N_1794);
or U2571 (N_2571,N_1330,N_1554);
and U2572 (N_2572,N_1695,N_1238);
or U2573 (N_2573,N_1923,N_1031);
nor U2574 (N_2574,N_1485,N_1414);
nor U2575 (N_2575,N_1659,N_1651);
or U2576 (N_2576,N_1849,N_1229);
or U2577 (N_2577,N_1337,N_1816);
nor U2578 (N_2578,N_1572,N_1401);
nand U2579 (N_2579,N_1047,N_1159);
or U2580 (N_2580,N_1658,N_1826);
nor U2581 (N_2581,N_1333,N_1713);
nand U2582 (N_2582,N_1204,N_1469);
nor U2583 (N_2583,N_1093,N_1704);
nand U2584 (N_2584,N_1186,N_1992);
or U2585 (N_2585,N_1371,N_1613);
or U2586 (N_2586,N_1713,N_1246);
or U2587 (N_2587,N_1876,N_1501);
and U2588 (N_2588,N_1191,N_1510);
nand U2589 (N_2589,N_1406,N_1565);
and U2590 (N_2590,N_1380,N_1278);
xnor U2591 (N_2591,N_1047,N_1156);
nor U2592 (N_2592,N_1630,N_1807);
nand U2593 (N_2593,N_1427,N_1853);
nand U2594 (N_2594,N_1640,N_1469);
nand U2595 (N_2595,N_1847,N_1288);
nand U2596 (N_2596,N_1665,N_1491);
and U2597 (N_2597,N_1577,N_1013);
or U2598 (N_2598,N_1035,N_1633);
xnor U2599 (N_2599,N_1219,N_1446);
nor U2600 (N_2600,N_1353,N_1846);
nor U2601 (N_2601,N_1777,N_1834);
or U2602 (N_2602,N_1799,N_1359);
nand U2603 (N_2603,N_1869,N_1351);
nand U2604 (N_2604,N_1559,N_1071);
or U2605 (N_2605,N_1488,N_1753);
or U2606 (N_2606,N_1981,N_1081);
or U2607 (N_2607,N_1635,N_1515);
nor U2608 (N_2608,N_1690,N_1940);
nand U2609 (N_2609,N_1628,N_1856);
or U2610 (N_2610,N_1235,N_1076);
or U2611 (N_2611,N_1871,N_1800);
or U2612 (N_2612,N_1065,N_1037);
nor U2613 (N_2613,N_1069,N_1145);
nand U2614 (N_2614,N_1491,N_1971);
nand U2615 (N_2615,N_1589,N_1845);
nand U2616 (N_2616,N_1385,N_1750);
or U2617 (N_2617,N_1708,N_1654);
or U2618 (N_2618,N_1713,N_1197);
or U2619 (N_2619,N_1540,N_1112);
nor U2620 (N_2620,N_1439,N_1056);
nand U2621 (N_2621,N_1457,N_1973);
or U2622 (N_2622,N_1995,N_1920);
nor U2623 (N_2623,N_1122,N_1442);
and U2624 (N_2624,N_1647,N_1640);
and U2625 (N_2625,N_1899,N_1993);
and U2626 (N_2626,N_1546,N_1635);
nand U2627 (N_2627,N_1541,N_1283);
and U2628 (N_2628,N_1674,N_1376);
nand U2629 (N_2629,N_1694,N_1873);
nand U2630 (N_2630,N_1684,N_1794);
nand U2631 (N_2631,N_1144,N_1008);
nor U2632 (N_2632,N_1157,N_1685);
and U2633 (N_2633,N_1342,N_1219);
xnor U2634 (N_2634,N_1363,N_1964);
nand U2635 (N_2635,N_1728,N_1268);
or U2636 (N_2636,N_1376,N_1655);
and U2637 (N_2637,N_1768,N_1323);
or U2638 (N_2638,N_1533,N_1057);
xnor U2639 (N_2639,N_1145,N_1916);
nor U2640 (N_2640,N_1971,N_1711);
nand U2641 (N_2641,N_1142,N_1685);
or U2642 (N_2642,N_1205,N_1907);
nand U2643 (N_2643,N_1377,N_1360);
and U2644 (N_2644,N_1596,N_1683);
and U2645 (N_2645,N_1859,N_1996);
nor U2646 (N_2646,N_1304,N_1909);
nor U2647 (N_2647,N_1754,N_1888);
or U2648 (N_2648,N_1642,N_1974);
nand U2649 (N_2649,N_1784,N_1294);
nor U2650 (N_2650,N_1749,N_1943);
nor U2651 (N_2651,N_1070,N_1461);
and U2652 (N_2652,N_1783,N_1456);
and U2653 (N_2653,N_1326,N_1733);
nand U2654 (N_2654,N_1562,N_1401);
nand U2655 (N_2655,N_1540,N_1066);
nor U2656 (N_2656,N_1944,N_1286);
nor U2657 (N_2657,N_1330,N_1970);
and U2658 (N_2658,N_1816,N_1154);
nand U2659 (N_2659,N_1243,N_1955);
nor U2660 (N_2660,N_1786,N_1624);
nand U2661 (N_2661,N_1892,N_1600);
nor U2662 (N_2662,N_1815,N_1614);
nor U2663 (N_2663,N_1401,N_1319);
nand U2664 (N_2664,N_1903,N_1824);
or U2665 (N_2665,N_1237,N_1714);
xor U2666 (N_2666,N_1888,N_1163);
nand U2667 (N_2667,N_1855,N_1526);
nor U2668 (N_2668,N_1457,N_1639);
nor U2669 (N_2669,N_1737,N_1303);
xor U2670 (N_2670,N_1339,N_1881);
nor U2671 (N_2671,N_1080,N_1880);
nand U2672 (N_2672,N_1310,N_1608);
or U2673 (N_2673,N_1987,N_1517);
nand U2674 (N_2674,N_1862,N_1460);
and U2675 (N_2675,N_1656,N_1903);
nor U2676 (N_2676,N_1142,N_1490);
and U2677 (N_2677,N_1254,N_1008);
xnor U2678 (N_2678,N_1816,N_1952);
nand U2679 (N_2679,N_1601,N_1331);
or U2680 (N_2680,N_1084,N_1725);
or U2681 (N_2681,N_1023,N_1198);
or U2682 (N_2682,N_1341,N_1692);
and U2683 (N_2683,N_1044,N_1213);
nor U2684 (N_2684,N_1252,N_1677);
or U2685 (N_2685,N_1404,N_1077);
and U2686 (N_2686,N_1867,N_1576);
or U2687 (N_2687,N_1938,N_1993);
and U2688 (N_2688,N_1808,N_1603);
nor U2689 (N_2689,N_1963,N_1783);
nand U2690 (N_2690,N_1528,N_1107);
nor U2691 (N_2691,N_1426,N_1115);
nand U2692 (N_2692,N_1556,N_1479);
and U2693 (N_2693,N_1782,N_1813);
nand U2694 (N_2694,N_1839,N_1535);
xor U2695 (N_2695,N_1109,N_1841);
and U2696 (N_2696,N_1911,N_1403);
nand U2697 (N_2697,N_1610,N_1849);
and U2698 (N_2698,N_1418,N_1911);
xor U2699 (N_2699,N_1844,N_1377);
nand U2700 (N_2700,N_1445,N_1627);
nand U2701 (N_2701,N_1831,N_1219);
or U2702 (N_2702,N_1176,N_1981);
nor U2703 (N_2703,N_1911,N_1108);
or U2704 (N_2704,N_1772,N_1922);
nand U2705 (N_2705,N_1005,N_1659);
and U2706 (N_2706,N_1309,N_1027);
and U2707 (N_2707,N_1067,N_1101);
xor U2708 (N_2708,N_1747,N_1698);
xor U2709 (N_2709,N_1104,N_1042);
and U2710 (N_2710,N_1168,N_1374);
or U2711 (N_2711,N_1498,N_1977);
and U2712 (N_2712,N_1277,N_1118);
nor U2713 (N_2713,N_1408,N_1216);
nand U2714 (N_2714,N_1424,N_1507);
nor U2715 (N_2715,N_1215,N_1703);
and U2716 (N_2716,N_1636,N_1514);
or U2717 (N_2717,N_1388,N_1941);
nor U2718 (N_2718,N_1093,N_1967);
nand U2719 (N_2719,N_1324,N_1011);
or U2720 (N_2720,N_1834,N_1439);
xnor U2721 (N_2721,N_1212,N_1245);
nor U2722 (N_2722,N_1026,N_1753);
and U2723 (N_2723,N_1140,N_1598);
nand U2724 (N_2724,N_1000,N_1546);
or U2725 (N_2725,N_1110,N_1300);
or U2726 (N_2726,N_1395,N_1863);
nand U2727 (N_2727,N_1051,N_1220);
nor U2728 (N_2728,N_1242,N_1663);
nand U2729 (N_2729,N_1366,N_1685);
or U2730 (N_2730,N_1947,N_1855);
nor U2731 (N_2731,N_1580,N_1820);
and U2732 (N_2732,N_1740,N_1529);
nor U2733 (N_2733,N_1300,N_1330);
xor U2734 (N_2734,N_1544,N_1332);
and U2735 (N_2735,N_1475,N_1235);
or U2736 (N_2736,N_1223,N_1052);
xnor U2737 (N_2737,N_1445,N_1154);
or U2738 (N_2738,N_1021,N_1817);
and U2739 (N_2739,N_1800,N_1167);
nand U2740 (N_2740,N_1074,N_1917);
xnor U2741 (N_2741,N_1049,N_1434);
and U2742 (N_2742,N_1811,N_1884);
nand U2743 (N_2743,N_1206,N_1317);
or U2744 (N_2744,N_1438,N_1503);
nand U2745 (N_2745,N_1186,N_1166);
or U2746 (N_2746,N_1232,N_1941);
nor U2747 (N_2747,N_1440,N_1484);
and U2748 (N_2748,N_1895,N_1181);
or U2749 (N_2749,N_1114,N_1351);
nand U2750 (N_2750,N_1443,N_1733);
and U2751 (N_2751,N_1130,N_1424);
and U2752 (N_2752,N_1435,N_1622);
nor U2753 (N_2753,N_1420,N_1490);
or U2754 (N_2754,N_1237,N_1358);
xnor U2755 (N_2755,N_1860,N_1900);
nand U2756 (N_2756,N_1758,N_1650);
or U2757 (N_2757,N_1474,N_1067);
nor U2758 (N_2758,N_1789,N_1547);
or U2759 (N_2759,N_1509,N_1926);
nand U2760 (N_2760,N_1803,N_1315);
nor U2761 (N_2761,N_1806,N_1688);
nor U2762 (N_2762,N_1520,N_1258);
and U2763 (N_2763,N_1072,N_1857);
or U2764 (N_2764,N_1257,N_1647);
nand U2765 (N_2765,N_1437,N_1623);
xnor U2766 (N_2766,N_1455,N_1856);
or U2767 (N_2767,N_1206,N_1361);
nor U2768 (N_2768,N_1523,N_1042);
nand U2769 (N_2769,N_1836,N_1559);
and U2770 (N_2770,N_1412,N_1145);
nand U2771 (N_2771,N_1671,N_1718);
and U2772 (N_2772,N_1917,N_1994);
and U2773 (N_2773,N_1932,N_1290);
or U2774 (N_2774,N_1202,N_1107);
or U2775 (N_2775,N_1178,N_1756);
nor U2776 (N_2776,N_1863,N_1922);
nor U2777 (N_2777,N_1962,N_1431);
nor U2778 (N_2778,N_1028,N_1243);
or U2779 (N_2779,N_1346,N_1103);
or U2780 (N_2780,N_1837,N_1285);
or U2781 (N_2781,N_1446,N_1028);
or U2782 (N_2782,N_1320,N_1339);
or U2783 (N_2783,N_1844,N_1176);
or U2784 (N_2784,N_1741,N_1678);
xnor U2785 (N_2785,N_1725,N_1764);
or U2786 (N_2786,N_1671,N_1542);
nor U2787 (N_2787,N_1598,N_1154);
or U2788 (N_2788,N_1579,N_1379);
and U2789 (N_2789,N_1022,N_1044);
xor U2790 (N_2790,N_1455,N_1612);
nand U2791 (N_2791,N_1333,N_1108);
xor U2792 (N_2792,N_1507,N_1033);
and U2793 (N_2793,N_1932,N_1076);
or U2794 (N_2794,N_1204,N_1057);
and U2795 (N_2795,N_1463,N_1846);
nor U2796 (N_2796,N_1089,N_1065);
and U2797 (N_2797,N_1202,N_1382);
nor U2798 (N_2798,N_1996,N_1223);
nand U2799 (N_2799,N_1623,N_1567);
nand U2800 (N_2800,N_1456,N_1203);
or U2801 (N_2801,N_1293,N_1352);
or U2802 (N_2802,N_1195,N_1683);
nand U2803 (N_2803,N_1011,N_1976);
nand U2804 (N_2804,N_1824,N_1888);
nand U2805 (N_2805,N_1126,N_1536);
xnor U2806 (N_2806,N_1418,N_1529);
and U2807 (N_2807,N_1638,N_1872);
nor U2808 (N_2808,N_1467,N_1833);
nand U2809 (N_2809,N_1547,N_1729);
xnor U2810 (N_2810,N_1264,N_1358);
and U2811 (N_2811,N_1064,N_1817);
nor U2812 (N_2812,N_1755,N_1443);
or U2813 (N_2813,N_1966,N_1909);
or U2814 (N_2814,N_1920,N_1386);
nor U2815 (N_2815,N_1793,N_1108);
nor U2816 (N_2816,N_1326,N_1717);
xnor U2817 (N_2817,N_1021,N_1629);
xor U2818 (N_2818,N_1581,N_1601);
and U2819 (N_2819,N_1904,N_1734);
or U2820 (N_2820,N_1304,N_1095);
nor U2821 (N_2821,N_1689,N_1979);
nand U2822 (N_2822,N_1657,N_1662);
or U2823 (N_2823,N_1268,N_1058);
and U2824 (N_2824,N_1797,N_1961);
and U2825 (N_2825,N_1021,N_1099);
nand U2826 (N_2826,N_1109,N_1317);
or U2827 (N_2827,N_1118,N_1514);
and U2828 (N_2828,N_1524,N_1623);
nor U2829 (N_2829,N_1760,N_1819);
nand U2830 (N_2830,N_1262,N_1913);
nor U2831 (N_2831,N_1400,N_1635);
nand U2832 (N_2832,N_1694,N_1968);
and U2833 (N_2833,N_1878,N_1078);
and U2834 (N_2834,N_1299,N_1814);
nor U2835 (N_2835,N_1144,N_1101);
and U2836 (N_2836,N_1274,N_1074);
or U2837 (N_2837,N_1933,N_1967);
and U2838 (N_2838,N_1302,N_1802);
or U2839 (N_2839,N_1826,N_1274);
nand U2840 (N_2840,N_1843,N_1290);
nand U2841 (N_2841,N_1448,N_1687);
or U2842 (N_2842,N_1896,N_1912);
xor U2843 (N_2843,N_1807,N_1486);
nor U2844 (N_2844,N_1734,N_1389);
nor U2845 (N_2845,N_1812,N_1932);
nand U2846 (N_2846,N_1193,N_1736);
nand U2847 (N_2847,N_1984,N_1450);
and U2848 (N_2848,N_1375,N_1227);
xor U2849 (N_2849,N_1850,N_1414);
nand U2850 (N_2850,N_1164,N_1773);
or U2851 (N_2851,N_1125,N_1291);
and U2852 (N_2852,N_1850,N_1343);
nand U2853 (N_2853,N_1703,N_1347);
nand U2854 (N_2854,N_1653,N_1088);
and U2855 (N_2855,N_1432,N_1042);
nand U2856 (N_2856,N_1880,N_1284);
nor U2857 (N_2857,N_1910,N_1509);
nor U2858 (N_2858,N_1056,N_1975);
or U2859 (N_2859,N_1711,N_1665);
xnor U2860 (N_2860,N_1694,N_1055);
nand U2861 (N_2861,N_1736,N_1170);
and U2862 (N_2862,N_1191,N_1633);
or U2863 (N_2863,N_1574,N_1241);
nor U2864 (N_2864,N_1180,N_1366);
xor U2865 (N_2865,N_1781,N_1288);
or U2866 (N_2866,N_1611,N_1270);
nor U2867 (N_2867,N_1443,N_1619);
nor U2868 (N_2868,N_1361,N_1665);
xnor U2869 (N_2869,N_1297,N_1972);
nand U2870 (N_2870,N_1449,N_1516);
or U2871 (N_2871,N_1906,N_1163);
nor U2872 (N_2872,N_1393,N_1558);
nand U2873 (N_2873,N_1647,N_1592);
nor U2874 (N_2874,N_1111,N_1543);
nor U2875 (N_2875,N_1595,N_1301);
nand U2876 (N_2876,N_1635,N_1869);
and U2877 (N_2877,N_1297,N_1292);
or U2878 (N_2878,N_1138,N_1793);
nor U2879 (N_2879,N_1894,N_1159);
nor U2880 (N_2880,N_1277,N_1725);
nand U2881 (N_2881,N_1588,N_1990);
nand U2882 (N_2882,N_1160,N_1550);
nand U2883 (N_2883,N_1799,N_1687);
and U2884 (N_2884,N_1686,N_1799);
and U2885 (N_2885,N_1297,N_1763);
and U2886 (N_2886,N_1543,N_1976);
and U2887 (N_2887,N_1818,N_1177);
and U2888 (N_2888,N_1195,N_1748);
nor U2889 (N_2889,N_1001,N_1438);
nor U2890 (N_2890,N_1119,N_1814);
nor U2891 (N_2891,N_1380,N_1312);
and U2892 (N_2892,N_1514,N_1848);
and U2893 (N_2893,N_1864,N_1220);
or U2894 (N_2894,N_1259,N_1557);
nand U2895 (N_2895,N_1105,N_1387);
or U2896 (N_2896,N_1186,N_1201);
or U2897 (N_2897,N_1394,N_1012);
or U2898 (N_2898,N_1318,N_1451);
nor U2899 (N_2899,N_1662,N_1737);
nand U2900 (N_2900,N_1089,N_1699);
nor U2901 (N_2901,N_1690,N_1012);
and U2902 (N_2902,N_1476,N_1551);
or U2903 (N_2903,N_1797,N_1896);
or U2904 (N_2904,N_1124,N_1256);
nand U2905 (N_2905,N_1666,N_1536);
nor U2906 (N_2906,N_1242,N_1636);
nand U2907 (N_2907,N_1997,N_1198);
or U2908 (N_2908,N_1350,N_1265);
nand U2909 (N_2909,N_1649,N_1708);
nand U2910 (N_2910,N_1525,N_1490);
or U2911 (N_2911,N_1157,N_1817);
nand U2912 (N_2912,N_1143,N_1582);
nor U2913 (N_2913,N_1387,N_1438);
and U2914 (N_2914,N_1194,N_1966);
and U2915 (N_2915,N_1068,N_1844);
nand U2916 (N_2916,N_1569,N_1898);
or U2917 (N_2917,N_1048,N_1846);
and U2918 (N_2918,N_1798,N_1719);
and U2919 (N_2919,N_1187,N_1575);
nor U2920 (N_2920,N_1663,N_1059);
or U2921 (N_2921,N_1238,N_1972);
nand U2922 (N_2922,N_1312,N_1514);
nor U2923 (N_2923,N_1180,N_1923);
nor U2924 (N_2924,N_1118,N_1996);
nand U2925 (N_2925,N_1809,N_1387);
nand U2926 (N_2926,N_1188,N_1486);
nor U2927 (N_2927,N_1759,N_1740);
nand U2928 (N_2928,N_1983,N_1708);
or U2929 (N_2929,N_1916,N_1968);
nor U2930 (N_2930,N_1604,N_1829);
and U2931 (N_2931,N_1781,N_1454);
nand U2932 (N_2932,N_1057,N_1817);
nor U2933 (N_2933,N_1788,N_1254);
or U2934 (N_2934,N_1096,N_1964);
and U2935 (N_2935,N_1040,N_1086);
or U2936 (N_2936,N_1146,N_1175);
nand U2937 (N_2937,N_1457,N_1376);
nor U2938 (N_2938,N_1571,N_1807);
nand U2939 (N_2939,N_1191,N_1150);
nand U2940 (N_2940,N_1027,N_1720);
nor U2941 (N_2941,N_1495,N_1408);
nand U2942 (N_2942,N_1045,N_1937);
nand U2943 (N_2943,N_1107,N_1187);
nor U2944 (N_2944,N_1986,N_1009);
nand U2945 (N_2945,N_1090,N_1422);
or U2946 (N_2946,N_1338,N_1954);
and U2947 (N_2947,N_1398,N_1099);
and U2948 (N_2948,N_1833,N_1353);
nand U2949 (N_2949,N_1946,N_1740);
nand U2950 (N_2950,N_1345,N_1414);
nor U2951 (N_2951,N_1592,N_1897);
nor U2952 (N_2952,N_1214,N_1777);
nor U2953 (N_2953,N_1223,N_1815);
nand U2954 (N_2954,N_1205,N_1705);
nand U2955 (N_2955,N_1955,N_1520);
or U2956 (N_2956,N_1770,N_1626);
or U2957 (N_2957,N_1008,N_1979);
and U2958 (N_2958,N_1025,N_1262);
and U2959 (N_2959,N_1953,N_1651);
nand U2960 (N_2960,N_1257,N_1877);
and U2961 (N_2961,N_1678,N_1123);
or U2962 (N_2962,N_1787,N_1873);
xor U2963 (N_2963,N_1807,N_1505);
nand U2964 (N_2964,N_1349,N_1763);
nand U2965 (N_2965,N_1669,N_1588);
nand U2966 (N_2966,N_1076,N_1438);
nand U2967 (N_2967,N_1215,N_1950);
nand U2968 (N_2968,N_1181,N_1414);
nand U2969 (N_2969,N_1952,N_1770);
xnor U2970 (N_2970,N_1311,N_1182);
or U2971 (N_2971,N_1906,N_1980);
or U2972 (N_2972,N_1807,N_1260);
or U2973 (N_2973,N_1854,N_1184);
xor U2974 (N_2974,N_1613,N_1587);
nor U2975 (N_2975,N_1811,N_1432);
and U2976 (N_2976,N_1020,N_1532);
nand U2977 (N_2977,N_1661,N_1994);
or U2978 (N_2978,N_1184,N_1735);
or U2979 (N_2979,N_1617,N_1402);
or U2980 (N_2980,N_1353,N_1888);
and U2981 (N_2981,N_1514,N_1232);
xnor U2982 (N_2982,N_1918,N_1765);
or U2983 (N_2983,N_1075,N_1511);
or U2984 (N_2984,N_1340,N_1024);
nand U2985 (N_2985,N_1274,N_1385);
and U2986 (N_2986,N_1559,N_1263);
nand U2987 (N_2987,N_1805,N_1248);
or U2988 (N_2988,N_1414,N_1463);
and U2989 (N_2989,N_1913,N_1780);
nor U2990 (N_2990,N_1621,N_1656);
and U2991 (N_2991,N_1077,N_1326);
nand U2992 (N_2992,N_1066,N_1823);
nor U2993 (N_2993,N_1949,N_1897);
xor U2994 (N_2994,N_1788,N_1760);
and U2995 (N_2995,N_1555,N_1336);
and U2996 (N_2996,N_1441,N_1014);
or U2997 (N_2997,N_1732,N_1831);
nand U2998 (N_2998,N_1407,N_1684);
and U2999 (N_2999,N_1100,N_1760);
xor U3000 (N_3000,N_2828,N_2272);
nand U3001 (N_3001,N_2519,N_2479);
nor U3002 (N_3002,N_2124,N_2549);
nand U3003 (N_3003,N_2105,N_2924);
and U3004 (N_3004,N_2987,N_2862);
nand U3005 (N_3005,N_2192,N_2866);
or U3006 (N_3006,N_2205,N_2363);
nand U3007 (N_3007,N_2947,N_2850);
nand U3008 (N_3008,N_2029,N_2035);
nand U3009 (N_3009,N_2212,N_2431);
or U3010 (N_3010,N_2097,N_2079);
nor U3011 (N_3011,N_2166,N_2755);
nor U3012 (N_3012,N_2720,N_2422);
nor U3013 (N_3013,N_2238,N_2584);
nor U3014 (N_3014,N_2872,N_2989);
xor U3015 (N_3015,N_2896,N_2633);
or U3016 (N_3016,N_2067,N_2647);
and U3017 (N_3017,N_2476,N_2569);
or U3018 (N_3018,N_2425,N_2570);
and U3019 (N_3019,N_2714,N_2466);
xor U3020 (N_3020,N_2201,N_2426);
xnor U3021 (N_3021,N_2214,N_2120);
nand U3022 (N_3022,N_2344,N_2387);
nor U3023 (N_3023,N_2604,N_2080);
and U3024 (N_3024,N_2279,N_2348);
xor U3025 (N_3025,N_2565,N_2992);
nor U3026 (N_3026,N_2652,N_2318);
or U3027 (N_3027,N_2965,N_2028);
and U3028 (N_3028,N_2651,N_2036);
or U3029 (N_3029,N_2394,N_2677);
and U3030 (N_3030,N_2456,N_2768);
and U3031 (N_3031,N_2874,N_2958);
and U3032 (N_3032,N_2390,N_2611);
or U3033 (N_3033,N_2158,N_2188);
nand U3034 (N_3034,N_2870,N_2087);
nor U3035 (N_3035,N_2858,N_2421);
nand U3036 (N_3036,N_2146,N_2187);
or U3037 (N_3037,N_2017,N_2962);
nor U3038 (N_3038,N_2050,N_2985);
nor U3039 (N_3039,N_2278,N_2015);
or U3040 (N_3040,N_2857,N_2262);
nor U3041 (N_3041,N_2708,N_2402);
or U3042 (N_3042,N_2692,N_2073);
xnor U3043 (N_3043,N_2592,N_2027);
nand U3044 (N_3044,N_2655,N_2732);
or U3045 (N_3045,N_2518,N_2054);
nor U3046 (N_3046,N_2762,N_2718);
and U3047 (N_3047,N_2091,N_2354);
xnor U3048 (N_3048,N_2928,N_2014);
nand U3049 (N_3049,N_2753,N_2645);
nor U3050 (N_3050,N_2040,N_2642);
nor U3051 (N_3051,N_2399,N_2313);
nand U3052 (N_3052,N_2574,N_2690);
or U3053 (N_3053,N_2323,N_2957);
nor U3054 (N_3054,N_2922,N_2761);
nor U3055 (N_3055,N_2107,N_2436);
nand U3056 (N_3056,N_2328,N_2472);
nand U3057 (N_3057,N_2150,N_2917);
nand U3058 (N_3058,N_2268,N_2285);
and U3059 (N_3059,N_2034,N_2156);
and U3060 (N_3060,N_2243,N_2170);
nand U3061 (N_3061,N_2736,N_2974);
nor U3062 (N_3062,N_2134,N_2667);
or U3063 (N_3063,N_2599,N_2649);
and U3064 (N_3064,N_2137,N_2590);
or U3065 (N_3065,N_2779,N_2427);
nor U3066 (N_3066,N_2048,N_2159);
xor U3067 (N_3067,N_2101,N_2259);
nand U3068 (N_3068,N_2112,N_2345);
and U3069 (N_3069,N_2566,N_2787);
or U3070 (N_3070,N_2596,N_2455);
and U3071 (N_3071,N_2379,N_2774);
and U3072 (N_3072,N_2795,N_2705);
or U3073 (N_3073,N_2338,N_2993);
or U3074 (N_3074,N_2898,N_2614);
nand U3075 (N_3075,N_2509,N_2771);
or U3076 (N_3076,N_2904,N_2467);
nor U3077 (N_3077,N_2253,N_2304);
nand U3078 (N_3078,N_2620,N_2024);
and U3079 (N_3079,N_2481,N_2157);
or U3080 (N_3080,N_2788,N_2143);
nand U3081 (N_3081,N_2662,N_2103);
and U3082 (N_3082,N_2817,N_2092);
and U3083 (N_3083,N_2636,N_2486);
nand U3084 (N_3084,N_2218,N_2716);
nor U3085 (N_3085,N_2179,N_2556);
nor U3086 (N_3086,N_2007,N_2491);
nor U3087 (N_3087,N_2721,N_2452);
nor U3088 (N_3088,N_2406,N_2948);
and U3089 (N_3089,N_2229,N_2089);
nand U3090 (N_3090,N_2901,N_2859);
nor U3091 (N_3091,N_2333,N_2608);
nor U3092 (N_3092,N_2940,N_2109);
and U3093 (N_3093,N_2542,N_2543);
nor U3094 (N_3094,N_2084,N_2075);
or U3095 (N_3095,N_2117,N_2325);
nor U3096 (N_3096,N_2177,N_2265);
or U3097 (N_3097,N_2401,N_2060);
nand U3098 (N_3098,N_2942,N_2322);
or U3099 (N_3099,N_2497,N_2236);
or U3100 (N_3100,N_2640,N_2625);
and U3101 (N_3101,N_2767,N_2292);
or U3102 (N_3102,N_2280,N_2587);
nor U3103 (N_3103,N_2042,N_2807);
nor U3104 (N_3104,N_2415,N_2326);
and U3105 (N_3105,N_2598,N_2700);
and U3106 (N_3106,N_2384,N_2175);
nor U3107 (N_3107,N_2738,N_2725);
or U3108 (N_3108,N_2811,N_2658);
xor U3109 (N_3109,N_2271,N_2386);
nor U3110 (N_3110,N_2521,N_2737);
and U3111 (N_3111,N_2062,N_2722);
and U3112 (N_3112,N_2801,N_2059);
nand U3113 (N_3113,N_2849,N_2806);
or U3114 (N_3114,N_2506,N_2461);
and U3115 (N_3115,N_2507,N_2302);
nand U3116 (N_3116,N_2226,N_2835);
nand U3117 (N_3117,N_2227,N_2217);
or U3118 (N_3118,N_2680,N_2113);
nand U3119 (N_3119,N_2135,N_2471);
and U3120 (N_3120,N_2077,N_2726);
and U3121 (N_3121,N_2897,N_2578);
xor U3122 (N_3122,N_2263,N_2641);
and U3123 (N_3123,N_2398,N_2595);
xnor U3124 (N_3124,N_2536,N_2260);
nor U3125 (N_3125,N_2269,N_2020);
nand U3126 (N_3126,N_2485,N_2139);
nand U3127 (N_3127,N_2867,N_2520);
nand U3128 (N_3128,N_2167,N_2085);
xor U3129 (N_3129,N_2881,N_2295);
or U3130 (N_3130,N_2972,N_2750);
xor U3131 (N_3131,N_2508,N_2930);
xnor U3132 (N_3132,N_2256,N_2539);
and U3133 (N_3133,N_2529,N_2453);
nor U3134 (N_3134,N_2395,N_2316);
nand U3135 (N_3135,N_2887,N_2936);
or U3136 (N_3136,N_2448,N_2005);
xor U3137 (N_3137,N_2743,N_2963);
nand U3138 (N_3138,N_2678,N_2953);
or U3139 (N_3139,N_2289,N_2648);
or U3140 (N_3140,N_2697,N_2251);
nand U3141 (N_3141,N_2908,N_2824);
and U3142 (N_3142,N_2078,N_2357);
and U3143 (N_3143,N_2430,N_2882);
nand U3144 (N_3144,N_2548,N_2562);
or U3145 (N_3145,N_2002,N_2961);
xor U3146 (N_3146,N_2552,N_2951);
xor U3147 (N_3147,N_2791,N_2827);
or U3148 (N_3148,N_2952,N_2588);
nand U3149 (N_3149,N_2239,N_2559);
nor U3150 (N_3150,N_2628,N_2819);
or U3151 (N_3151,N_2712,N_2274);
nor U3152 (N_3152,N_2808,N_2056);
nand U3153 (N_3153,N_2912,N_2830);
nor U3154 (N_3154,N_2102,N_2638);
nand U3155 (N_3155,N_2222,N_2441);
nand U3156 (N_3156,N_2149,N_2997);
xnor U3157 (N_3157,N_2799,N_2407);
and U3158 (N_3158,N_2907,N_2138);
or U3159 (N_3159,N_2305,N_2173);
or U3160 (N_3160,N_2465,N_2707);
xnor U3161 (N_3161,N_2735,N_2586);
and U3162 (N_3162,N_2086,N_2082);
and U3163 (N_3163,N_2329,N_2511);
nor U3164 (N_3164,N_2478,N_2500);
and U3165 (N_3165,N_2684,N_2861);
or U3166 (N_3166,N_2290,N_2419);
and U3167 (N_3167,N_2053,N_2128);
and U3168 (N_3168,N_2475,N_2327);
and U3169 (N_3169,N_2848,N_2317);
and U3170 (N_3170,N_2999,N_2920);
or U3171 (N_3171,N_2840,N_2668);
and U3172 (N_3172,N_2624,N_2096);
nand U3173 (N_3173,N_2759,N_2110);
or U3174 (N_3174,N_2030,N_2216);
nor U3175 (N_3175,N_2568,N_2039);
nor U3176 (N_3176,N_2734,N_2293);
and U3177 (N_3177,N_2825,N_2046);
nand U3178 (N_3178,N_2763,N_2764);
xnor U3179 (N_3179,N_2148,N_2675);
nor U3180 (N_3180,N_2136,N_2739);
and U3181 (N_3181,N_2051,N_2489);
or U3182 (N_3182,N_2623,N_2267);
nor U3183 (N_3183,N_2356,N_2070);
or U3184 (N_3184,N_2551,N_2673);
nand U3185 (N_3185,N_2909,N_2129);
and U3186 (N_3186,N_2434,N_2286);
nor U3187 (N_3187,N_2303,N_2541);
and U3188 (N_3188,N_2903,N_2396);
or U3189 (N_3189,N_2656,N_2458);
and U3190 (N_3190,N_2281,N_2012);
nor U3191 (N_3191,N_2785,N_2603);
xnor U3192 (N_3192,N_2480,N_2186);
nor U3193 (N_3193,N_2927,N_2902);
and U3194 (N_3194,N_2932,N_2564);
or U3195 (N_3195,N_2976,N_2145);
and U3196 (N_3196,N_2609,N_2760);
nand U3197 (N_3197,N_2021,N_2695);
or U3198 (N_3198,N_2526,N_2470);
nor U3199 (N_3199,N_2810,N_2748);
and U3200 (N_3200,N_2729,N_2198);
and U3201 (N_3201,N_2831,N_2180);
nor U3202 (N_3202,N_2626,N_2772);
nor U3203 (N_3203,N_2044,N_2713);
or U3204 (N_3204,N_2378,N_2424);
xor U3205 (N_3205,N_2501,N_2443);
nor U3206 (N_3206,N_2423,N_2412);
nand U3207 (N_3207,N_2373,N_2127);
and U3208 (N_3208,N_2880,N_2343);
nand U3209 (N_3209,N_2189,N_2778);
nor U3210 (N_3210,N_2288,N_2408);
or U3211 (N_3211,N_2495,N_2594);
and U3212 (N_3212,N_2161,N_2445);
nor U3213 (N_3213,N_2747,N_2207);
xor U3214 (N_3214,N_2093,N_2884);
nand U3215 (N_3215,N_2754,N_2249);
or U3216 (N_3216,N_2661,N_2477);
nand U3217 (N_3217,N_2664,N_2533);
nand U3218 (N_3218,N_2194,N_2474);
or U3219 (N_3219,N_2525,N_2561);
nand U3220 (N_3220,N_2314,N_2210);
and U3221 (N_3221,N_2809,N_2644);
or U3222 (N_3222,N_2023,N_2273);
and U3223 (N_3223,N_2306,N_2581);
nand U3224 (N_3224,N_2499,N_2998);
or U3225 (N_3225,N_2659,N_2765);
and U3226 (N_3226,N_2248,N_2654);
or U3227 (N_3227,N_2504,N_2460);
nor U3228 (N_3228,N_2417,N_2710);
and U3229 (N_3229,N_2049,N_2769);
and U3230 (N_3230,N_2503,N_2488);
nand U3231 (N_3231,N_2100,N_2382);
and U3232 (N_3232,N_2597,N_2190);
xor U3233 (N_3233,N_2944,N_2493);
nand U3234 (N_3234,N_2823,N_2794);
nor U3235 (N_3235,N_2601,N_2914);
nand U3236 (N_3236,N_2943,N_2008);
nand U3237 (N_3237,N_2444,N_2671);
or U3238 (N_3238,N_2929,N_2964);
and U3239 (N_3239,N_2532,N_2950);
nand U3240 (N_3240,N_2114,N_2414);
nor U3241 (N_3241,N_2530,N_2704);
and U3242 (N_3242,N_2308,N_2528);
nand U3243 (N_3243,N_2287,N_2682);
nand U3244 (N_3244,N_2320,N_2487);
nand U3245 (N_3245,N_2437,N_2340);
or U3246 (N_3246,N_2111,N_2631);
nor U3247 (N_3247,N_2294,N_2839);
xnor U3248 (N_3248,N_2300,N_2283);
xnor U3249 (N_3249,N_2342,N_2815);
nor U3250 (N_3250,N_2063,N_2984);
xor U3251 (N_3251,N_2266,N_2757);
or U3252 (N_3252,N_2770,N_2978);
nor U3253 (N_3253,N_2330,N_2833);
nor U3254 (N_3254,N_2247,N_2983);
and U3255 (N_3255,N_2037,N_2245);
nand U3256 (N_3256,N_2234,N_2746);
and U3257 (N_3257,N_2153,N_2879);
xor U3258 (N_3258,N_2733,N_2935);
or U3259 (N_3259,N_2674,N_2646);
and U3260 (N_3260,N_2967,N_2719);
nand U3261 (N_3261,N_2841,N_2450);
xor U3262 (N_3262,N_2171,N_2061);
or U3263 (N_3263,N_2199,N_2593);
and U3264 (N_3264,N_2405,N_2178);
or U3265 (N_3265,N_2886,N_2132);
nor U3266 (N_3266,N_2168,N_2703);
or U3267 (N_3267,N_2851,N_2990);
nor U3268 (N_3268,N_2670,N_2900);
or U3269 (N_3269,N_2971,N_2986);
nand U3270 (N_3270,N_2071,N_2832);
nor U3271 (N_3271,N_2740,N_2540);
xnor U3272 (N_3272,N_2813,N_2955);
or U3273 (N_3273,N_2496,N_2038);
xnor U3274 (N_3274,N_2232,N_2041);
nor U3275 (N_3275,N_2505,N_2863);
nand U3276 (N_3276,N_2782,N_2428);
or U3277 (N_3277,N_2449,N_2918);
nor U3278 (N_3278,N_2200,N_2074);
and U3279 (N_3279,N_2792,N_2066);
nand U3280 (N_3280,N_2375,N_2181);
nand U3281 (N_3281,N_2282,N_2195);
or U3282 (N_3282,N_2013,N_2058);
nand U3283 (N_3283,N_2244,N_2147);
or U3284 (N_3284,N_2923,N_2650);
nand U3285 (N_3285,N_2968,N_2681);
or U3286 (N_3286,N_2573,N_2104);
or U3287 (N_3287,N_2583,N_2711);
nor U3288 (N_3288,N_2871,N_2018);
and U3289 (N_3289,N_2400,N_2358);
and U3290 (N_3290,N_2208,N_2404);
or U3291 (N_3291,N_2213,N_2355);
or U3292 (N_3292,N_2215,N_2558);
or U3293 (N_3293,N_2223,N_2687);
xnor U3294 (N_3294,N_2440,N_2197);
nor U3295 (N_3295,N_2446,N_2865);
and U3296 (N_3296,N_2435,N_2803);
nand U3297 (N_3297,N_2696,N_2176);
and U3298 (N_3298,N_2883,N_2557);
nand U3299 (N_3299,N_2727,N_2381);
nand U3300 (N_3300,N_2413,N_2174);
xor U3301 (N_3301,N_2099,N_2531);
xor U3302 (N_3302,N_2106,N_2892);
nand U3303 (N_3303,N_2960,N_2906);
and U3304 (N_3304,N_2522,N_2602);
and U3305 (N_3305,N_2837,N_2994);
xor U3306 (N_3306,N_2921,N_2545);
nand U3307 (N_3307,N_2309,N_2366);
or U3308 (N_3308,N_2630,N_2605);
or U3309 (N_3309,N_2933,N_2126);
or U3310 (N_3310,N_2022,N_2834);
nor U3311 (N_3311,N_2261,N_2691);
or U3312 (N_3312,N_2131,N_2349);
nor U3313 (N_3313,N_2484,N_2959);
xor U3314 (N_3314,N_2560,N_2125);
nand U3315 (N_3315,N_2370,N_2847);
nand U3316 (N_3316,N_2816,N_2116);
and U3317 (N_3317,N_2154,N_2321);
or U3318 (N_3318,N_2065,N_2347);
xor U3319 (N_3319,N_2606,N_2184);
nand U3320 (N_3320,N_2941,N_2784);
xnor U3321 (N_3321,N_2339,N_2169);
nand U3322 (N_3322,N_2016,N_2275);
and U3323 (N_3323,N_2246,N_2706);
and U3324 (N_3324,N_2621,N_2081);
nand U3325 (N_3325,N_2334,N_2982);
xor U3326 (N_3326,N_2009,N_2291);
and U3327 (N_3327,N_2916,N_2731);
xnor U3328 (N_3328,N_2397,N_2411);
and U3329 (N_3329,N_2473,N_2805);
nand U3330 (N_3330,N_2544,N_2307);
and U3331 (N_3331,N_2513,N_2252);
or U3332 (N_3332,N_2353,N_2004);
xnor U3333 (N_3333,N_2165,N_2514);
or U3334 (N_3334,N_2374,N_2255);
nor U3335 (N_3335,N_2890,N_2211);
nor U3336 (N_3336,N_2403,N_2362);
xor U3337 (N_3337,N_2889,N_2498);
nor U3338 (N_3338,N_2196,N_2172);
nand U3339 (N_3339,N_2350,N_2820);
nor U3340 (N_3340,N_2524,N_2796);
or U3341 (N_3341,N_2776,N_2814);
nand U3342 (N_3342,N_2970,N_2869);
xor U3343 (N_3343,N_2826,N_2264);
or U3344 (N_3344,N_2447,N_2140);
nand U3345 (N_3345,N_2003,N_2072);
nor U3346 (N_3346,N_2418,N_2873);
and U3347 (N_3347,N_2699,N_2224);
or U3348 (N_3348,N_2853,N_2310);
or U3349 (N_3349,N_2535,N_2821);
nor U3350 (N_3350,N_2749,N_2877);
nor U3351 (N_3351,N_2351,N_2416);
nor U3352 (N_3352,N_2838,N_2966);
and U3353 (N_3353,N_2547,N_2409);
xnor U3354 (N_3354,N_2221,N_2822);
nor U3355 (N_3355,N_2133,N_2006);
nor U3356 (N_3356,N_2991,N_2025);
nor U3357 (N_3357,N_2995,N_2676);
nand U3358 (N_3358,N_2368,N_2895);
nand U3359 (N_3359,N_2660,N_2463);
nor U3360 (N_3360,N_2800,N_2001);
nor U3361 (N_3361,N_2164,N_2257);
xor U3362 (N_3362,N_2119,N_2802);
and U3363 (N_3363,N_2155,N_2361);
and U3364 (N_3364,N_2876,N_2393);
nand U3365 (N_3365,N_2319,N_2332);
and U3366 (N_3366,N_2988,N_2141);
or U3367 (N_3367,N_2618,N_2752);
or U3368 (N_3368,N_2885,N_2534);
nand U3369 (N_3369,N_2019,N_2553);
nand U3370 (N_3370,N_2372,N_2000);
or U3371 (N_3371,N_2864,N_2756);
nand U3372 (N_3372,N_2385,N_2438);
or U3373 (N_3373,N_2582,N_2980);
xnor U3374 (N_3374,N_2121,N_2537);
or U3375 (N_3375,N_2206,N_2193);
and U3376 (N_3376,N_2804,N_2459);
and U3377 (N_3377,N_2931,N_2672);
and U3378 (N_3378,N_2380,N_2629);
or U3379 (N_3379,N_2299,N_2919);
and U3380 (N_3380,N_2494,N_2790);
nor U3381 (N_3381,N_2669,N_2377);
or U3382 (N_3382,N_2392,N_2634);
nand U3383 (N_3383,N_2312,N_2315);
nand U3384 (N_3384,N_2457,N_2546);
nor U3385 (N_3385,N_2679,N_2615);
xnor U3386 (N_3386,N_2946,N_2878);
and U3387 (N_3387,N_2846,N_2766);
nand U3388 (N_3388,N_2842,N_2185);
nor U3389 (N_3389,N_2237,N_2875);
nor U3390 (N_3390,N_2780,N_2975);
or U3391 (N_3391,N_2331,N_2225);
nand U3392 (N_3392,N_2938,N_2639);
or U3393 (N_3393,N_2758,N_2694);
nor U3394 (N_3394,N_2616,N_2433);
and U3395 (N_3395,N_2429,N_2773);
nand U3396 (N_3396,N_2538,N_2981);
nor U3397 (N_3397,N_2359,N_2612);
nand U3398 (N_3398,N_2492,N_2945);
xor U3399 (N_3399,N_2836,N_2969);
nor U3400 (N_3400,N_2554,N_2702);
nor U3401 (N_3401,N_2891,N_2632);
or U3402 (N_3402,N_2130,N_2610);
or U3403 (N_3403,N_2240,N_2899);
or U3404 (N_3404,N_2341,N_2915);
and U3405 (N_3405,N_2144,N_2956);
and U3406 (N_3406,N_2346,N_2793);
xor U3407 (N_3407,N_2183,N_2032);
or U3408 (N_3408,N_2576,N_2613);
or U3409 (N_3409,N_2868,N_2439);
nand U3410 (N_3410,N_2893,N_2163);
or U3411 (N_3411,N_2088,N_2230);
or U3412 (N_3412,N_2665,N_2219);
xor U3413 (N_3413,N_2517,N_2657);
or U3414 (N_3414,N_2977,N_2228);
or U3415 (N_3415,N_2555,N_2383);
or U3416 (N_3416,N_2115,N_2937);
and U3417 (N_3417,N_2777,N_2856);
nand U3418 (N_3418,N_2516,N_2242);
or U3419 (N_3419,N_2666,N_2360);
or U3420 (N_3420,N_2142,N_2203);
nand U3421 (N_3421,N_2202,N_2469);
nand U3422 (N_3422,N_2996,N_2254);
nand U3423 (N_3423,N_2052,N_2797);
xor U3424 (N_3424,N_2069,N_2741);
or U3425 (N_3425,N_2855,N_2798);
nand U3426 (N_3426,N_2160,N_2812);
and U3427 (N_3427,N_2627,N_2689);
or U3428 (N_3428,N_2490,N_2575);
and U3429 (N_3429,N_2462,N_2683);
and U3430 (N_3430,N_2235,N_2209);
or U3431 (N_3431,N_2420,N_2352);
nor U3432 (N_3432,N_2095,N_2055);
or U3433 (N_3433,N_2789,N_2860);
nor U3434 (N_3434,N_2949,N_2643);
xnor U3435 (N_3435,N_2335,N_2122);
nand U3436 (N_3436,N_2979,N_2745);
nor U3437 (N_3437,N_2090,N_2926);
nand U3438 (N_3438,N_2888,N_2512);
xor U3439 (N_3439,N_2277,N_2258);
or U3440 (N_3440,N_2934,N_2270);
or U3441 (N_3441,N_2033,N_2728);
nor U3442 (N_3442,N_2905,N_2910);
or U3443 (N_3443,N_2010,N_2123);
nor U3444 (N_3444,N_2527,N_2468);
nor U3445 (N_3445,N_2031,N_2693);
or U3446 (N_3446,N_2709,N_2064);
nor U3447 (N_3447,N_2567,N_2786);
nand U3448 (N_3448,N_2389,N_2685);
xor U3449 (N_3449,N_2571,N_2775);
or U3450 (N_3450,N_2451,N_2118);
or U3451 (N_3451,N_2744,N_2454);
or U3452 (N_3452,N_2502,N_2954);
nand U3453 (N_3453,N_2367,N_2730);
and U3454 (N_3454,N_2284,N_2043);
nor U3455 (N_3455,N_2076,N_2047);
or U3456 (N_3456,N_2098,N_2577);
nand U3457 (N_3457,N_2298,N_2619);
nand U3458 (N_3458,N_2410,N_2364);
nor U3459 (N_3459,N_2296,N_2845);
nand U3460 (N_3460,N_2483,N_2717);
nor U3461 (N_3461,N_2724,N_2607);
nor U3462 (N_3462,N_2723,N_2151);
or U3463 (N_3463,N_2152,N_2337);
and U3464 (N_3464,N_2688,N_2622);
or U3465 (N_3465,N_2220,N_2432);
or U3466 (N_3466,N_2482,N_2894);
xor U3467 (N_3467,N_2925,N_2742);
nor U3468 (N_3468,N_2510,N_2580);
xnor U3469 (N_3469,N_2715,N_2585);
nor U3470 (N_3470,N_2371,N_2068);
or U3471 (N_3471,N_2011,N_2913);
or U3472 (N_3472,N_2464,N_2241);
nand U3473 (N_3473,N_2191,N_2635);
or U3474 (N_3474,N_2108,N_2442);
xnor U3475 (N_3475,N_2301,N_2182);
or U3476 (N_3476,N_2045,N_2939);
and U3477 (N_3477,N_2783,N_2391);
nor U3478 (N_3478,N_2973,N_2818);
and U3479 (N_3479,N_2233,N_2852);
xor U3480 (N_3480,N_2515,N_2911);
nor U3481 (N_3481,N_2701,N_2324);
and U3482 (N_3482,N_2311,N_2550);
nand U3483 (N_3483,N_2204,N_2781);
or U3484 (N_3484,N_2523,N_2686);
nand U3485 (N_3485,N_2829,N_2843);
and U3486 (N_3486,N_2276,N_2591);
xor U3487 (N_3487,N_2388,N_2637);
nor U3488 (N_3488,N_2250,N_2376);
and U3489 (N_3489,N_2563,N_2162);
and U3490 (N_3490,N_2663,N_2083);
and U3491 (N_3491,N_2336,N_2231);
nor U3492 (N_3492,N_2579,N_2365);
and U3493 (N_3493,N_2589,N_2026);
and U3494 (N_3494,N_2698,N_2094);
nand U3495 (N_3495,N_2854,N_2369);
and U3496 (N_3496,N_2600,N_2297);
or U3497 (N_3497,N_2751,N_2617);
and U3498 (N_3498,N_2572,N_2844);
or U3499 (N_3499,N_2653,N_2057);
nand U3500 (N_3500,N_2967,N_2068);
nand U3501 (N_3501,N_2065,N_2697);
nand U3502 (N_3502,N_2409,N_2979);
nor U3503 (N_3503,N_2661,N_2533);
nor U3504 (N_3504,N_2128,N_2932);
nor U3505 (N_3505,N_2008,N_2101);
and U3506 (N_3506,N_2169,N_2239);
and U3507 (N_3507,N_2504,N_2089);
nand U3508 (N_3508,N_2612,N_2528);
nand U3509 (N_3509,N_2344,N_2709);
or U3510 (N_3510,N_2571,N_2591);
nor U3511 (N_3511,N_2746,N_2601);
or U3512 (N_3512,N_2858,N_2882);
nor U3513 (N_3513,N_2274,N_2046);
or U3514 (N_3514,N_2996,N_2497);
nor U3515 (N_3515,N_2963,N_2674);
and U3516 (N_3516,N_2060,N_2231);
nor U3517 (N_3517,N_2113,N_2723);
nor U3518 (N_3518,N_2020,N_2776);
nor U3519 (N_3519,N_2014,N_2176);
and U3520 (N_3520,N_2207,N_2678);
nor U3521 (N_3521,N_2934,N_2732);
and U3522 (N_3522,N_2810,N_2191);
and U3523 (N_3523,N_2520,N_2472);
nor U3524 (N_3524,N_2513,N_2878);
nor U3525 (N_3525,N_2624,N_2361);
or U3526 (N_3526,N_2505,N_2158);
or U3527 (N_3527,N_2178,N_2618);
nand U3528 (N_3528,N_2069,N_2888);
nor U3529 (N_3529,N_2198,N_2319);
nand U3530 (N_3530,N_2018,N_2483);
nand U3531 (N_3531,N_2875,N_2905);
and U3532 (N_3532,N_2821,N_2188);
nor U3533 (N_3533,N_2242,N_2858);
and U3534 (N_3534,N_2466,N_2248);
xor U3535 (N_3535,N_2874,N_2849);
nand U3536 (N_3536,N_2148,N_2917);
nor U3537 (N_3537,N_2000,N_2113);
xnor U3538 (N_3538,N_2687,N_2669);
nand U3539 (N_3539,N_2674,N_2817);
or U3540 (N_3540,N_2509,N_2356);
and U3541 (N_3541,N_2445,N_2016);
xor U3542 (N_3542,N_2715,N_2139);
or U3543 (N_3543,N_2743,N_2552);
or U3544 (N_3544,N_2921,N_2578);
xor U3545 (N_3545,N_2599,N_2600);
or U3546 (N_3546,N_2588,N_2899);
nor U3547 (N_3547,N_2278,N_2403);
and U3548 (N_3548,N_2002,N_2823);
xnor U3549 (N_3549,N_2181,N_2762);
nor U3550 (N_3550,N_2490,N_2176);
nand U3551 (N_3551,N_2136,N_2444);
or U3552 (N_3552,N_2898,N_2927);
nand U3553 (N_3553,N_2801,N_2527);
and U3554 (N_3554,N_2350,N_2577);
nor U3555 (N_3555,N_2249,N_2112);
xnor U3556 (N_3556,N_2895,N_2875);
and U3557 (N_3557,N_2002,N_2474);
nor U3558 (N_3558,N_2264,N_2254);
or U3559 (N_3559,N_2408,N_2051);
nand U3560 (N_3560,N_2102,N_2771);
nand U3561 (N_3561,N_2851,N_2365);
and U3562 (N_3562,N_2213,N_2476);
nor U3563 (N_3563,N_2190,N_2563);
nand U3564 (N_3564,N_2419,N_2495);
and U3565 (N_3565,N_2440,N_2666);
and U3566 (N_3566,N_2374,N_2475);
and U3567 (N_3567,N_2596,N_2276);
or U3568 (N_3568,N_2405,N_2906);
nand U3569 (N_3569,N_2959,N_2379);
nand U3570 (N_3570,N_2500,N_2238);
nand U3571 (N_3571,N_2929,N_2053);
and U3572 (N_3572,N_2066,N_2020);
nor U3573 (N_3573,N_2158,N_2053);
xnor U3574 (N_3574,N_2251,N_2703);
and U3575 (N_3575,N_2151,N_2076);
xor U3576 (N_3576,N_2795,N_2534);
nand U3577 (N_3577,N_2229,N_2061);
and U3578 (N_3578,N_2321,N_2750);
nor U3579 (N_3579,N_2458,N_2754);
or U3580 (N_3580,N_2145,N_2699);
nand U3581 (N_3581,N_2856,N_2088);
nor U3582 (N_3582,N_2198,N_2246);
or U3583 (N_3583,N_2251,N_2846);
xor U3584 (N_3584,N_2521,N_2752);
or U3585 (N_3585,N_2960,N_2719);
and U3586 (N_3586,N_2793,N_2396);
or U3587 (N_3587,N_2109,N_2790);
nand U3588 (N_3588,N_2207,N_2669);
xor U3589 (N_3589,N_2862,N_2408);
and U3590 (N_3590,N_2264,N_2150);
or U3591 (N_3591,N_2698,N_2121);
or U3592 (N_3592,N_2814,N_2684);
or U3593 (N_3593,N_2035,N_2130);
or U3594 (N_3594,N_2434,N_2833);
or U3595 (N_3595,N_2866,N_2474);
and U3596 (N_3596,N_2982,N_2020);
nand U3597 (N_3597,N_2666,N_2243);
xnor U3598 (N_3598,N_2468,N_2722);
or U3599 (N_3599,N_2157,N_2527);
xnor U3600 (N_3600,N_2642,N_2238);
or U3601 (N_3601,N_2754,N_2136);
xor U3602 (N_3602,N_2601,N_2602);
and U3603 (N_3603,N_2856,N_2125);
xnor U3604 (N_3604,N_2398,N_2034);
and U3605 (N_3605,N_2214,N_2384);
nand U3606 (N_3606,N_2857,N_2809);
nor U3607 (N_3607,N_2193,N_2596);
nand U3608 (N_3608,N_2229,N_2108);
xnor U3609 (N_3609,N_2581,N_2466);
nor U3610 (N_3610,N_2917,N_2141);
nand U3611 (N_3611,N_2055,N_2090);
and U3612 (N_3612,N_2127,N_2482);
or U3613 (N_3613,N_2787,N_2742);
or U3614 (N_3614,N_2632,N_2797);
xnor U3615 (N_3615,N_2121,N_2407);
nand U3616 (N_3616,N_2454,N_2308);
nand U3617 (N_3617,N_2239,N_2085);
and U3618 (N_3618,N_2967,N_2583);
nand U3619 (N_3619,N_2412,N_2210);
or U3620 (N_3620,N_2949,N_2683);
nand U3621 (N_3621,N_2451,N_2791);
and U3622 (N_3622,N_2359,N_2766);
nand U3623 (N_3623,N_2184,N_2712);
or U3624 (N_3624,N_2716,N_2360);
xnor U3625 (N_3625,N_2143,N_2556);
or U3626 (N_3626,N_2256,N_2774);
nor U3627 (N_3627,N_2311,N_2037);
and U3628 (N_3628,N_2295,N_2146);
nand U3629 (N_3629,N_2308,N_2274);
nor U3630 (N_3630,N_2386,N_2589);
nand U3631 (N_3631,N_2834,N_2950);
nand U3632 (N_3632,N_2437,N_2930);
nor U3633 (N_3633,N_2213,N_2652);
and U3634 (N_3634,N_2729,N_2455);
and U3635 (N_3635,N_2239,N_2123);
nor U3636 (N_3636,N_2181,N_2399);
nor U3637 (N_3637,N_2856,N_2846);
and U3638 (N_3638,N_2600,N_2162);
nand U3639 (N_3639,N_2545,N_2271);
xnor U3640 (N_3640,N_2913,N_2062);
and U3641 (N_3641,N_2264,N_2996);
or U3642 (N_3642,N_2317,N_2099);
and U3643 (N_3643,N_2754,N_2532);
nand U3644 (N_3644,N_2815,N_2895);
nor U3645 (N_3645,N_2315,N_2323);
nand U3646 (N_3646,N_2025,N_2020);
nand U3647 (N_3647,N_2224,N_2778);
and U3648 (N_3648,N_2179,N_2666);
nor U3649 (N_3649,N_2452,N_2587);
nor U3650 (N_3650,N_2004,N_2100);
and U3651 (N_3651,N_2492,N_2473);
and U3652 (N_3652,N_2379,N_2064);
and U3653 (N_3653,N_2617,N_2182);
nor U3654 (N_3654,N_2701,N_2844);
nor U3655 (N_3655,N_2501,N_2234);
nor U3656 (N_3656,N_2139,N_2561);
or U3657 (N_3657,N_2401,N_2752);
nor U3658 (N_3658,N_2490,N_2602);
or U3659 (N_3659,N_2873,N_2745);
and U3660 (N_3660,N_2579,N_2509);
nand U3661 (N_3661,N_2570,N_2673);
or U3662 (N_3662,N_2204,N_2106);
nand U3663 (N_3663,N_2412,N_2556);
xor U3664 (N_3664,N_2904,N_2677);
and U3665 (N_3665,N_2046,N_2346);
nor U3666 (N_3666,N_2887,N_2760);
nand U3667 (N_3667,N_2874,N_2075);
nor U3668 (N_3668,N_2806,N_2979);
or U3669 (N_3669,N_2373,N_2718);
nand U3670 (N_3670,N_2538,N_2783);
nand U3671 (N_3671,N_2116,N_2857);
nor U3672 (N_3672,N_2986,N_2303);
nor U3673 (N_3673,N_2810,N_2066);
or U3674 (N_3674,N_2988,N_2914);
and U3675 (N_3675,N_2202,N_2687);
or U3676 (N_3676,N_2366,N_2806);
nand U3677 (N_3677,N_2963,N_2487);
nand U3678 (N_3678,N_2631,N_2758);
or U3679 (N_3679,N_2238,N_2600);
nand U3680 (N_3680,N_2945,N_2791);
nand U3681 (N_3681,N_2263,N_2035);
or U3682 (N_3682,N_2027,N_2768);
nor U3683 (N_3683,N_2677,N_2690);
and U3684 (N_3684,N_2112,N_2076);
nand U3685 (N_3685,N_2971,N_2623);
xnor U3686 (N_3686,N_2296,N_2396);
and U3687 (N_3687,N_2192,N_2567);
xor U3688 (N_3688,N_2821,N_2602);
or U3689 (N_3689,N_2126,N_2568);
nor U3690 (N_3690,N_2963,N_2540);
or U3691 (N_3691,N_2116,N_2867);
nand U3692 (N_3692,N_2447,N_2608);
nor U3693 (N_3693,N_2187,N_2183);
nand U3694 (N_3694,N_2828,N_2681);
and U3695 (N_3695,N_2989,N_2901);
xor U3696 (N_3696,N_2649,N_2514);
or U3697 (N_3697,N_2813,N_2860);
nand U3698 (N_3698,N_2605,N_2703);
or U3699 (N_3699,N_2792,N_2794);
or U3700 (N_3700,N_2224,N_2937);
nor U3701 (N_3701,N_2656,N_2286);
nor U3702 (N_3702,N_2649,N_2484);
and U3703 (N_3703,N_2116,N_2660);
nand U3704 (N_3704,N_2804,N_2438);
nand U3705 (N_3705,N_2397,N_2799);
and U3706 (N_3706,N_2204,N_2619);
nand U3707 (N_3707,N_2576,N_2751);
nand U3708 (N_3708,N_2741,N_2477);
nand U3709 (N_3709,N_2471,N_2937);
nor U3710 (N_3710,N_2221,N_2283);
nand U3711 (N_3711,N_2759,N_2761);
nand U3712 (N_3712,N_2161,N_2695);
and U3713 (N_3713,N_2733,N_2787);
and U3714 (N_3714,N_2495,N_2124);
xor U3715 (N_3715,N_2137,N_2897);
or U3716 (N_3716,N_2604,N_2261);
nand U3717 (N_3717,N_2425,N_2622);
and U3718 (N_3718,N_2884,N_2721);
and U3719 (N_3719,N_2839,N_2032);
or U3720 (N_3720,N_2943,N_2856);
xor U3721 (N_3721,N_2347,N_2921);
nor U3722 (N_3722,N_2286,N_2894);
nand U3723 (N_3723,N_2556,N_2897);
nand U3724 (N_3724,N_2959,N_2299);
or U3725 (N_3725,N_2256,N_2684);
and U3726 (N_3726,N_2761,N_2252);
nand U3727 (N_3727,N_2161,N_2419);
nor U3728 (N_3728,N_2277,N_2434);
and U3729 (N_3729,N_2738,N_2019);
and U3730 (N_3730,N_2597,N_2010);
or U3731 (N_3731,N_2708,N_2909);
nor U3732 (N_3732,N_2855,N_2635);
nor U3733 (N_3733,N_2247,N_2636);
xnor U3734 (N_3734,N_2780,N_2906);
or U3735 (N_3735,N_2099,N_2820);
and U3736 (N_3736,N_2405,N_2593);
nand U3737 (N_3737,N_2925,N_2137);
and U3738 (N_3738,N_2406,N_2644);
nand U3739 (N_3739,N_2941,N_2659);
or U3740 (N_3740,N_2274,N_2418);
and U3741 (N_3741,N_2120,N_2045);
and U3742 (N_3742,N_2988,N_2812);
nor U3743 (N_3743,N_2359,N_2592);
and U3744 (N_3744,N_2845,N_2037);
nor U3745 (N_3745,N_2560,N_2944);
nor U3746 (N_3746,N_2248,N_2592);
and U3747 (N_3747,N_2528,N_2738);
and U3748 (N_3748,N_2283,N_2480);
or U3749 (N_3749,N_2915,N_2863);
and U3750 (N_3750,N_2180,N_2452);
or U3751 (N_3751,N_2912,N_2385);
or U3752 (N_3752,N_2475,N_2425);
xnor U3753 (N_3753,N_2702,N_2293);
xnor U3754 (N_3754,N_2013,N_2948);
and U3755 (N_3755,N_2026,N_2942);
or U3756 (N_3756,N_2435,N_2577);
and U3757 (N_3757,N_2456,N_2606);
xor U3758 (N_3758,N_2478,N_2349);
nand U3759 (N_3759,N_2076,N_2606);
nor U3760 (N_3760,N_2111,N_2045);
nor U3761 (N_3761,N_2259,N_2775);
or U3762 (N_3762,N_2262,N_2742);
xor U3763 (N_3763,N_2178,N_2282);
nand U3764 (N_3764,N_2459,N_2454);
or U3765 (N_3765,N_2908,N_2211);
nand U3766 (N_3766,N_2210,N_2639);
nor U3767 (N_3767,N_2552,N_2617);
nor U3768 (N_3768,N_2207,N_2133);
and U3769 (N_3769,N_2520,N_2852);
and U3770 (N_3770,N_2276,N_2409);
or U3771 (N_3771,N_2112,N_2425);
nor U3772 (N_3772,N_2185,N_2523);
and U3773 (N_3773,N_2887,N_2619);
or U3774 (N_3774,N_2887,N_2568);
or U3775 (N_3775,N_2077,N_2758);
or U3776 (N_3776,N_2481,N_2082);
nor U3777 (N_3777,N_2983,N_2073);
or U3778 (N_3778,N_2424,N_2348);
and U3779 (N_3779,N_2347,N_2748);
or U3780 (N_3780,N_2579,N_2480);
nor U3781 (N_3781,N_2698,N_2332);
xnor U3782 (N_3782,N_2795,N_2663);
and U3783 (N_3783,N_2132,N_2266);
nand U3784 (N_3784,N_2318,N_2439);
xor U3785 (N_3785,N_2273,N_2153);
nand U3786 (N_3786,N_2098,N_2745);
nor U3787 (N_3787,N_2723,N_2253);
nor U3788 (N_3788,N_2178,N_2276);
or U3789 (N_3789,N_2140,N_2024);
and U3790 (N_3790,N_2948,N_2492);
and U3791 (N_3791,N_2169,N_2825);
and U3792 (N_3792,N_2210,N_2973);
and U3793 (N_3793,N_2064,N_2435);
nand U3794 (N_3794,N_2155,N_2538);
nor U3795 (N_3795,N_2842,N_2126);
nand U3796 (N_3796,N_2134,N_2547);
nand U3797 (N_3797,N_2981,N_2911);
nand U3798 (N_3798,N_2444,N_2156);
nand U3799 (N_3799,N_2094,N_2413);
nand U3800 (N_3800,N_2316,N_2501);
nand U3801 (N_3801,N_2641,N_2159);
or U3802 (N_3802,N_2929,N_2286);
nand U3803 (N_3803,N_2762,N_2479);
nor U3804 (N_3804,N_2212,N_2153);
and U3805 (N_3805,N_2016,N_2082);
nand U3806 (N_3806,N_2791,N_2380);
nand U3807 (N_3807,N_2994,N_2234);
nor U3808 (N_3808,N_2175,N_2290);
nor U3809 (N_3809,N_2075,N_2273);
or U3810 (N_3810,N_2496,N_2528);
nor U3811 (N_3811,N_2776,N_2938);
and U3812 (N_3812,N_2585,N_2089);
xor U3813 (N_3813,N_2016,N_2337);
nor U3814 (N_3814,N_2232,N_2079);
and U3815 (N_3815,N_2378,N_2286);
or U3816 (N_3816,N_2058,N_2164);
xor U3817 (N_3817,N_2654,N_2604);
and U3818 (N_3818,N_2018,N_2549);
and U3819 (N_3819,N_2051,N_2218);
or U3820 (N_3820,N_2851,N_2666);
and U3821 (N_3821,N_2464,N_2307);
or U3822 (N_3822,N_2114,N_2491);
and U3823 (N_3823,N_2400,N_2290);
and U3824 (N_3824,N_2597,N_2237);
nand U3825 (N_3825,N_2362,N_2955);
nor U3826 (N_3826,N_2412,N_2673);
nor U3827 (N_3827,N_2534,N_2255);
xor U3828 (N_3828,N_2513,N_2394);
and U3829 (N_3829,N_2373,N_2692);
nor U3830 (N_3830,N_2445,N_2238);
xnor U3831 (N_3831,N_2379,N_2914);
and U3832 (N_3832,N_2452,N_2487);
or U3833 (N_3833,N_2185,N_2042);
nor U3834 (N_3834,N_2615,N_2526);
or U3835 (N_3835,N_2940,N_2672);
nor U3836 (N_3836,N_2212,N_2140);
or U3837 (N_3837,N_2922,N_2134);
nor U3838 (N_3838,N_2453,N_2548);
and U3839 (N_3839,N_2565,N_2328);
nand U3840 (N_3840,N_2059,N_2968);
nor U3841 (N_3841,N_2182,N_2479);
nor U3842 (N_3842,N_2318,N_2116);
or U3843 (N_3843,N_2530,N_2154);
or U3844 (N_3844,N_2228,N_2147);
nand U3845 (N_3845,N_2116,N_2359);
xnor U3846 (N_3846,N_2132,N_2908);
and U3847 (N_3847,N_2482,N_2556);
nor U3848 (N_3848,N_2447,N_2778);
xor U3849 (N_3849,N_2000,N_2076);
or U3850 (N_3850,N_2656,N_2394);
or U3851 (N_3851,N_2977,N_2279);
nor U3852 (N_3852,N_2408,N_2518);
nand U3853 (N_3853,N_2557,N_2234);
and U3854 (N_3854,N_2211,N_2478);
nor U3855 (N_3855,N_2710,N_2944);
or U3856 (N_3856,N_2213,N_2899);
or U3857 (N_3857,N_2566,N_2227);
or U3858 (N_3858,N_2450,N_2832);
xnor U3859 (N_3859,N_2334,N_2676);
nor U3860 (N_3860,N_2481,N_2208);
xnor U3861 (N_3861,N_2893,N_2667);
xnor U3862 (N_3862,N_2412,N_2835);
nand U3863 (N_3863,N_2316,N_2831);
and U3864 (N_3864,N_2371,N_2901);
or U3865 (N_3865,N_2425,N_2655);
nor U3866 (N_3866,N_2051,N_2369);
nand U3867 (N_3867,N_2515,N_2149);
or U3868 (N_3868,N_2449,N_2003);
and U3869 (N_3869,N_2603,N_2399);
nand U3870 (N_3870,N_2035,N_2171);
or U3871 (N_3871,N_2665,N_2680);
nand U3872 (N_3872,N_2572,N_2494);
xor U3873 (N_3873,N_2791,N_2173);
and U3874 (N_3874,N_2145,N_2759);
or U3875 (N_3875,N_2592,N_2105);
and U3876 (N_3876,N_2356,N_2819);
and U3877 (N_3877,N_2770,N_2330);
and U3878 (N_3878,N_2758,N_2996);
and U3879 (N_3879,N_2693,N_2549);
and U3880 (N_3880,N_2610,N_2358);
xor U3881 (N_3881,N_2728,N_2017);
xnor U3882 (N_3882,N_2083,N_2421);
nor U3883 (N_3883,N_2774,N_2817);
nand U3884 (N_3884,N_2845,N_2682);
xor U3885 (N_3885,N_2935,N_2680);
and U3886 (N_3886,N_2571,N_2243);
nor U3887 (N_3887,N_2807,N_2476);
nand U3888 (N_3888,N_2667,N_2344);
nor U3889 (N_3889,N_2797,N_2058);
xor U3890 (N_3890,N_2847,N_2017);
or U3891 (N_3891,N_2418,N_2606);
nand U3892 (N_3892,N_2526,N_2749);
or U3893 (N_3893,N_2586,N_2449);
nor U3894 (N_3894,N_2263,N_2775);
nand U3895 (N_3895,N_2324,N_2876);
and U3896 (N_3896,N_2677,N_2107);
and U3897 (N_3897,N_2185,N_2104);
nand U3898 (N_3898,N_2990,N_2975);
xor U3899 (N_3899,N_2889,N_2725);
or U3900 (N_3900,N_2046,N_2359);
nor U3901 (N_3901,N_2376,N_2464);
or U3902 (N_3902,N_2697,N_2016);
nor U3903 (N_3903,N_2166,N_2065);
and U3904 (N_3904,N_2979,N_2131);
nor U3905 (N_3905,N_2549,N_2482);
or U3906 (N_3906,N_2481,N_2584);
nor U3907 (N_3907,N_2893,N_2721);
nand U3908 (N_3908,N_2735,N_2550);
or U3909 (N_3909,N_2110,N_2150);
nor U3910 (N_3910,N_2189,N_2677);
nor U3911 (N_3911,N_2739,N_2338);
or U3912 (N_3912,N_2445,N_2243);
or U3913 (N_3913,N_2172,N_2493);
or U3914 (N_3914,N_2287,N_2083);
or U3915 (N_3915,N_2559,N_2882);
or U3916 (N_3916,N_2160,N_2374);
and U3917 (N_3917,N_2234,N_2083);
xnor U3918 (N_3918,N_2616,N_2294);
or U3919 (N_3919,N_2734,N_2708);
xor U3920 (N_3920,N_2865,N_2962);
and U3921 (N_3921,N_2377,N_2929);
or U3922 (N_3922,N_2355,N_2223);
nand U3923 (N_3923,N_2095,N_2937);
nand U3924 (N_3924,N_2430,N_2295);
nor U3925 (N_3925,N_2999,N_2251);
nand U3926 (N_3926,N_2294,N_2805);
or U3927 (N_3927,N_2201,N_2883);
or U3928 (N_3928,N_2781,N_2549);
or U3929 (N_3929,N_2796,N_2673);
nor U3930 (N_3930,N_2367,N_2930);
nand U3931 (N_3931,N_2805,N_2656);
nor U3932 (N_3932,N_2344,N_2310);
xor U3933 (N_3933,N_2154,N_2088);
nor U3934 (N_3934,N_2895,N_2606);
and U3935 (N_3935,N_2883,N_2154);
or U3936 (N_3936,N_2615,N_2603);
or U3937 (N_3937,N_2746,N_2101);
nor U3938 (N_3938,N_2360,N_2221);
or U3939 (N_3939,N_2842,N_2626);
nand U3940 (N_3940,N_2158,N_2021);
nor U3941 (N_3941,N_2017,N_2247);
and U3942 (N_3942,N_2909,N_2984);
or U3943 (N_3943,N_2326,N_2186);
nor U3944 (N_3944,N_2179,N_2288);
nor U3945 (N_3945,N_2808,N_2643);
and U3946 (N_3946,N_2952,N_2175);
or U3947 (N_3947,N_2755,N_2290);
nor U3948 (N_3948,N_2236,N_2652);
or U3949 (N_3949,N_2044,N_2581);
nor U3950 (N_3950,N_2389,N_2206);
or U3951 (N_3951,N_2574,N_2458);
nor U3952 (N_3952,N_2598,N_2008);
xnor U3953 (N_3953,N_2129,N_2210);
and U3954 (N_3954,N_2016,N_2670);
or U3955 (N_3955,N_2045,N_2833);
or U3956 (N_3956,N_2806,N_2974);
xnor U3957 (N_3957,N_2232,N_2419);
nand U3958 (N_3958,N_2639,N_2629);
nor U3959 (N_3959,N_2488,N_2960);
and U3960 (N_3960,N_2722,N_2794);
nor U3961 (N_3961,N_2638,N_2340);
and U3962 (N_3962,N_2120,N_2041);
nand U3963 (N_3963,N_2864,N_2389);
and U3964 (N_3964,N_2057,N_2119);
nor U3965 (N_3965,N_2983,N_2553);
nand U3966 (N_3966,N_2519,N_2883);
nand U3967 (N_3967,N_2759,N_2299);
xor U3968 (N_3968,N_2740,N_2744);
nor U3969 (N_3969,N_2435,N_2789);
or U3970 (N_3970,N_2783,N_2543);
and U3971 (N_3971,N_2853,N_2223);
xor U3972 (N_3972,N_2211,N_2325);
and U3973 (N_3973,N_2548,N_2420);
xnor U3974 (N_3974,N_2380,N_2389);
nand U3975 (N_3975,N_2056,N_2492);
and U3976 (N_3976,N_2233,N_2584);
or U3977 (N_3977,N_2764,N_2771);
nand U3978 (N_3978,N_2141,N_2794);
nand U3979 (N_3979,N_2973,N_2706);
nor U3980 (N_3980,N_2821,N_2019);
nor U3981 (N_3981,N_2186,N_2211);
nor U3982 (N_3982,N_2949,N_2096);
and U3983 (N_3983,N_2064,N_2723);
nand U3984 (N_3984,N_2412,N_2910);
nor U3985 (N_3985,N_2476,N_2959);
and U3986 (N_3986,N_2933,N_2341);
nand U3987 (N_3987,N_2328,N_2503);
nand U3988 (N_3988,N_2043,N_2267);
nor U3989 (N_3989,N_2324,N_2170);
and U3990 (N_3990,N_2415,N_2194);
nor U3991 (N_3991,N_2290,N_2452);
or U3992 (N_3992,N_2719,N_2907);
nand U3993 (N_3993,N_2197,N_2229);
and U3994 (N_3994,N_2973,N_2997);
and U3995 (N_3995,N_2407,N_2856);
xor U3996 (N_3996,N_2510,N_2082);
or U3997 (N_3997,N_2993,N_2841);
nand U3998 (N_3998,N_2783,N_2429);
nor U3999 (N_3999,N_2682,N_2400);
nand U4000 (N_4000,N_3183,N_3094);
or U4001 (N_4001,N_3068,N_3249);
or U4002 (N_4002,N_3607,N_3694);
nor U4003 (N_4003,N_3794,N_3987);
nand U4004 (N_4004,N_3863,N_3801);
and U4005 (N_4005,N_3588,N_3245);
xnor U4006 (N_4006,N_3495,N_3133);
nor U4007 (N_4007,N_3367,N_3505);
and U4008 (N_4008,N_3030,N_3115);
and U4009 (N_4009,N_3867,N_3540);
or U4010 (N_4010,N_3331,N_3691);
nor U4011 (N_4011,N_3004,N_3826);
and U4012 (N_4012,N_3810,N_3374);
xnor U4013 (N_4013,N_3017,N_3005);
or U4014 (N_4014,N_3101,N_3922);
and U4015 (N_4015,N_3015,N_3384);
nor U4016 (N_4016,N_3699,N_3668);
nor U4017 (N_4017,N_3656,N_3636);
or U4018 (N_4018,N_3104,N_3494);
nand U4019 (N_4019,N_3811,N_3338);
nor U4020 (N_4020,N_3585,N_3918);
nor U4021 (N_4021,N_3186,N_3665);
nor U4022 (N_4022,N_3560,N_3000);
or U4023 (N_4023,N_3066,N_3662);
and U4024 (N_4024,N_3731,N_3406);
or U4025 (N_4025,N_3012,N_3988);
nor U4026 (N_4026,N_3622,N_3532);
nand U4027 (N_4027,N_3110,N_3873);
and U4028 (N_4028,N_3837,N_3126);
xor U4029 (N_4029,N_3599,N_3284);
or U4030 (N_4030,N_3309,N_3677);
and U4031 (N_4031,N_3928,N_3483);
nor U4032 (N_4032,N_3380,N_3836);
or U4033 (N_4033,N_3805,N_3959);
nand U4034 (N_4034,N_3261,N_3725);
xor U4035 (N_4035,N_3717,N_3021);
or U4036 (N_4036,N_3514,N_3973);
or U4037 (N_4037,N_3264,N_3402);
and U4038 (N_4038,N_3070,N_3872);
xor U4039 (N_4039,N_3184,N_3020);
nor U4040 (N_4040,N_3536,N_3736);
nand U4041 (N_4041,N_3465,N_3033);
or U4042 (N_4042,N_3117,N_3137);
nor U4043 (N_4043,N_3630,N_3625);
and U4044 (N_4044,N_3577,N_3010);
nand U4045 (N_4045,N_3452,N_3541);
nor U4046 (N_4046,N_3831,N_3266);
and U4047 (N_4047,N_3940,N_3617);
and U4048 (N_4048,N_3300,N_3236);
and U4049 (N_4049,N_3008,N_3527);
and U4050 (N_4050,N_3597,N_3006);
nand U4051 (N_4051,N_3660,N_3459);
nand U4052 (N_4052,N_3220,N_3774);
nor U4053 (N_4053,N_3968,N_3571);
and U4054 (N_4054,N_3263,N_3210);
nand U4055 (N_4055,N_3082,N_3684);
and U4056 (N_4056,N_3568,N_3433);
and U4057 (N_4057,N_3390,N_3590);
nor U4058 (N_4058,N_3565,N_3637);
or U4059 (N_4059,N_3611,N_3854);
or U4060 (N_4060,N_3050,N_3596);
xor U4061 (N_4061,N_3173,N_3693);
nor U4062 (N_4062,N_3071,N_3517);
nor U4063 (N_4063,N_3790,N_3623);
nor U4064 (N_4064,N_3205,N_3286);
nand U4065 (N_4065,N_3127,N_3086);
and U4066 (N_4066,N_3169,N_3724);
or U4067 (N_4067,N_3681,N_3387);
or U4068 (N_4068,N_3105,N_3237);
and U4069 (N_4069,N_3009,N_3657);
nand U4070 (N_4070,N_3519,N_3889);
and U4071 (N_4071,N_3492,N_3217);
nand U4072 (N_4072,N_3703,N_3129);
nand U4073 (N_4073,N_3641,N_3412);
nand U4074 (N_4074,N_3933,N_3531);
or U4075 (N_4075,N_3160,N_3573);
or U4076 (N_4076,N_3156,N_3972);
and U4077 (N_4077,N_3464,N_3537);
nor U4078 (N_4078,N_3159,N_3243);
nor U4079 (N_4079,N_3706,N_3062);
nor U4080 (N_4080,N_3314,N_3513);
and U4081 (N_4081,N_3733,N_3784);
and U4082 (N_4082,N_3092,N_3842);
nand U4083 (N_4083,N_3153,N_3634);
xor U4084 (N_4084,N_3043,N_3089);
xor U4085 (N_4085,N_3757,N_3895);
nand U4086 (N_4086,N_3179,N_3077);
or U4087 (N_4087,N_3510,N_3342);
or U4088 (N_4088,N_3290,N_3440);
nor U4089 (N_4089,N_3269,N_3230);
and U4090 (N_4090,N_3157,N_3315);
and U4091 (N_4091,N_3177,N_3721);
nor U4092 (N_4092,N_3899,N_3116);
and U4093 (N_4093,N_3368,N_3675);
nor U4094 (N_4094,N_3956,N_3403);
and U4095 (N_4095,N_3888,N_3470);
or U4096 (N_4096,N_3938,N_3026);
or U4097 (N_4097,N_3651,N_3904);
nand U4098 (N_4098,N_3248,N_3851);
and U4099 (N_4099,N_3524,N_3576);
or U4100 (N_4100,N_3530,N_3818);
and U4101 (N_4101,N_3233,N_3754);
or U4102 (N_4102,N_3806,N_3913);
nand U4103 (N_4103,N_3287,N_3554);
nand U4104 (N_4104,N_3631,N_3934);
xnor U4105 (N_4105,N_3658,N_3544);
nor U4106 (N_4106,N_3609,N_3711);
nand U4107 (N_4107,N_3073,N_3923);
nand U4108 (N_4108,N_3164,N_3511);
and U4109 (N_4109,N_3983,N_3445);
or U4110 (N_4110,N_3078,N_3714);
or U4111 (N_4111,N_3798,N_3386);
and U4112 (N_4112,N_3874,N_3521);
nor U4113 (N_4113,N_3778,N_3962);
nand U4114 (N_4114,N_3466,N_3546);
or U4115 (N_4115,N_3697,N_3768);
nand U4116 (N_4116,N_3083,N_3683);
nor U4117 (N_4117,N_3362,N_3924);
and U4118 (N_4118,N_3946,N_3887);
nor U4119 (N_4119,N_3844,N_3392);
nand U4120 (N_4120,N_3726,N_3476);
or U4121 (N_4121,N_3399,N_3966);
nor U4122 (N_4122,N_3011,N_3321);
and U4123 (N_4123,N_3337,N_3219);
and U4124 (N_4124,N_3722,N_3646);
nor U4125 (N_4125,N_3860,N_3161);
nor U4126 (N_4126,N_3310,N_3743);
xor U4127 (N_4127,N_3339,N_3378);
or U4128 (N_4128,N_3639,N_3047);
nor U4129 (N_4129,N_3529,N_3620);
or U4130 (N_4130,N_3750,N_3328);
nor U4131 (N_4131,N_3642,N_3882);
nand U4132 (N_4132,N_3958,N_3980);
and U4133 (N_4133,N_3600,N_3563);
and U4134 (N_4134,N_3791,N_3324);
nor U4135 (N_4135,N_3203,N_3221);
nor U4136 (N_4136,N_3821,N_3520);
or U4137 (N_4137,N_3312,N_3682);
and U4138 (N_4138,N_3343,N_3190);
and U4139 (N_4139,N_3752,N_3740);
or U4140 (N_4140,N_3866,N_3032);
nor U4141 (N_4141,N_3674,N_3277);
and U4142 (N_4142,N_3274,N_3382);
nand U4143 (N_4143,N_3151,N_3451);
and U4144 (N_4144,N_3346,N_3100);
nor U4145 (N_4145,N_3467,N_3979);
nand U4146 (N_4146,N_3618,N_3167);
nor U4147 (N_4147,N_3120,N_3256);
and U4148 (N_4148,N_3292,N_3950);
nor U4149 (N_4149,N_3985,N_3253);
nor U4150 (N_4150,N_3175,N_3493);
and U4151 (N_4151,N_3431,N_3500);
xor U4152 (N_4152,N_3136,N_3921);
xnor U4153 (N_4153,N_3478,N_3356);
and U4154 (N_4154,N_3695,N_3689);
nor U4155 (N_4155,N_3425,N_3592);
or U4156 (N_4156,N_3508,N_3861);
and U4157 (N_4157,N_3297,N_3051);
xnor U4158 (N_4158,N_3046,N_3799);
or U4159 (N_4159,N_3215,N_3223);
and U4160 (N_4160,N_3834,N_3293);
nor U4161 (N_4161,N_3195,N_3145);
nand U4162 (N_4162,N_3262,N_3613);
nor U4163 (N_4163,N_3593,N_3316);
xor U4164 (N_4164,N_3629,N_3663);
nand U4165 (N_4165,N_3268,N_3458);
nand U4166 (N_4166,N_3871,N_3931);
nand U4167 (N_4167,N_3594,N_3163);
xor U4168 (N_4168,N_3589,N_3393);
or U4169 (N_4169,N_3640,N_3063);
nand U4170 (N_4170,N_3947,N_3974);
nor U4171 (N_4171,N_3422,N_3712);
nand U4172 (N_4172,N_3036,N_3745);
and U4173 (N_4173,N_3619,N_3612);
nor U4174 (N_4174,N_3401,N_3807);
and U4175 (N_4175,N_3949,N_3621);
nor U4176 (N_4176,N_3491,N_3567);
or U4177 (N_4177,N_3883,N_3761);
nor U4178 (N_4178,N_3969,N_3789);
nor U4179 (N_4179,N_3408,N_3448);
nor U4180 (N_4180,N_3014,N_3538);
or U4181 (N_4181,N_3042,N_3917);
nand U4182 (N_4182,N_3049,N_3438);
nand U4183 (N_4183,N_3064,N_3246);
or U4184 (N_4184,N_3606,N_3766);
and U4185 (N_4185,N_3961,N_3019);
or U4186 (N_4186,N_3603,N_3441);
nand U4187 (N_4187,N_3772,N_3518);
and U4188 (N_4188,N_3423,N_3664);
and U4189 (N_4189,N_3295,N_3583);
or U4190 (N_4190,N_3898,N_3472);
xnor U4191 (N_4191,N_3251,N_3890);
and U4192 (N_4192,N_3626,N_3855);
and U4193 (N_4193,N_3809,N_3782);
nand U4194 (N_4194,N_3345,N_3003);
or U4195 (N_4195,N_3424,N_3580);
and U4196 (N_4196,N_3052,N_3013);
xnor U4197 (N_4197,N_3391,N_3696);
nand U4198 (N_4198,N_3574,N_3479);
and U4199 (N_4199,N_3528,N_3841);
nand U4200 (N_4200,N_3022,N_3352);
nor U4201 (N_4201,N_3397,N_3498);
and U4202 (N_4202,N_3713,N_3832);
or U4203 (N_4203,N_3037,N_3932);
xor U4204 (N_4204,N_3558,N_3561);
and U4205 (N_4205,N_3085,N_3140);
and U4206 (N_4206,N_3031,N_3812);
nand U4207 (N_4207,N_3525,N_3614);
or U4208 (N_4208,N_3303,N_3208);
or U4209 (N_4209,N_3911,N_3690);
nand U4210 (N_4210,N_3542,N_3655);
or U4211 (N_4211,N_3096,N_3381);
nor U4212 (N_4212,N_3845,N_3672);
nor U4213 (N_4213,N_3212,N_3886);
nand U4214 (N_4214,N_3727,N_3948);
and U4215 (N_4215,N_3952,N_3490);
and U4216 (N_4216,N_3853,N_3201);
nand U4217 (N_4217,N_3322,N_3978);
and U4218 (N_4218,N_3435,N_3468);
or U4219 (N_4219,N_3856,N_3276);
or U4220 (N_4220,N_3900,N_3825);
nand U4221 (N_4221,N_3119,N_3076);
and U4222 (N_4222,N_3708,N_3123);
and U4223 (N_4223,N_3819,N_3124);
nor U4224 (N_4224,N_3881,N_3038);
nand U4225 (N_4225,N_3864,N_3715);
nor U4226 (N_4226,N_3474,N_3072);
nor U4227 (N_4227,N_3785,N_3209);
and U4228 (N_4228,N_3045,N_3552);
nor U4229 (N_4229,N_3769,N_3741);
or U4230 (N_4230,N_3704,N_3647);
nand U4231 (N_4231,N_3060,N_3484);
and U4232 (N_4232,N_3131,N_3598);
nand U4233 (N_4233,N_3383,N_3206);
and U4234 (N_4234,N_3462,N_3114);
nor U4235 (N_4235,N_3056,N_3473);
nand U4236 (N_4236,N_3787,N_3814);
or U4237 (N_4237,N_3087,N_3482);
or U4238 (N_4238,N_3896,N_3275);
nand U4239 (N_4239,N_3211,N_3349);
or U4240 (N_4240,N_3228,N_3875);
and U4241 (N_4241,N_3868,N_3143);
nand U4242 (N_4242,N_3041,N_3828);
xnor U4243 (N_4243,N_3318,N_3953);
or U4244 (N_4244,N_3502,N_3447);
or U4245 (N_4245,N_3936,N_3204);
nand U4246 (N_4246,N_3150,N_3199);
and U4247 (N_4247,N_3735,N_3415);
and U4248 (N_4248,N_3570,N_3564);
nand U4249 (N_4249,N_3624,N_3121);
or U4250 (N_4250,N_3709,N_3385);
xor U4251 (N_4251,N_3428,N_3394);
xor U4252 (N_4252,N_3549,N_3180);
and U4253 (N_4253,N_3515,N_3398);
or U4254 (N_4254,N_3756,N_3539);
and U4255 (N_4255,N_3838,N_3591);
and U4256 (N_4256,N_3363,N_3702);
nand U4257 (N_4257,N_3840,N_3319);
nor U4258 (N_4258,N_3059,N_3698);
and U4259 (N_4259,N_3943,N_3654);
nor U4260 (N_4260,N_3587,N_3701);
nand U4261 (N_4261,N_3800,N_3763);
or U4262 (N_4262,N_3281,N_3975);
xnor U4263 (N_4263,N_3165,N_3128);
or U4264 (N_4264,N_3377,N_3080);
nor U4265 (N_4265,N_3920,N_3941);
and U4266 (N_4266,N_3870,N_3644);
or U4267 (N_4267,N_3700,N_3369);
or U4268 (N_4268,N_3016,N_3793);
and U4269 (N_4269,N_3240,N_3154);
nand U4270 (N_4270,N_3301,N_3776);
or U4271 (N_4271,N_3065,N_3523);
nand U4272 (N_4272,N_3200,N_3797);
nor U4273 (N_4273,N_3430,N_3892);
nand U4274 (N_4274,N_3347,N_3294);
nand U4275 (N_4275,N_3299,N_3499);
xnor U4276 (N_4276,N_3437,N_3118);
or U4277 (N_4277,N_3993,N_3185);
or U4278 (N_4278,N_3601,N_3191);
nor U4279 (N_4279,N_3409,N_3048);
and U4280 (N_4280,N_3330,N_3350);
nor U4281 (N_4281,N_3351,N_3770);
and U4282 (N_4282,N_3850,N_3182);
and U4283 (N_4283,N_3497,N_3427);
nor U4284 (N_4284,N_3575,N_3334);
nor U4285 (N_4285,N_3891,N_3192);
or U4286 (N_4286,N_3088,N_3992);
nor U4287 (N_4287,N_3395,N_3361);
nor U4288 (N_4288,N_3915,N_3652);
or U4289 (N_4289,N_3313,N_3335);
nor U4290 (N_4290,N_3707,N_3566);
and U4291 (N_4291,N_3418,N_3141);
xnor U4292 (N_4292,N_3372,N_3976);
and U4293 (N_4293,N_3905,N_3218);
nand U4294 (N_4294,N_3375,N_3138);
or U4295 (N_4295,N_3097,N_3122);
or U4296 (N_4296,N_3091,N_3605);
nor U4297 (N_4297,N_3410,N_3442);
or U4298 (N_4298,N_3242,N_3130);
and U4299 (N_4299,N_3257,N_3053);
or U4300 (N_4300,N_3417,N_3547);
or U4301 (N_4301,N_3170,N_3001);
nor U4302 (N_4302,N_3912,N_3680);
and U4303 (N_4303,N_3916,N_3687);
xnor U4304 (N_4304,N_3653,N_3635);
nand U4305 (N_4305,N_3504,N_3885);
and U4306 (N_4306,N_3488,N_3710);
or U4307 (N_4307,N_3659,N_3827);
nand U4308 (N_4308,N_3308,N_3481);
nor U4309 (N_4309,N_3278,N_3282);
xnor U4310 (N_4310,N_3102,N_3325);
or U4311 (N_4311,N_3739,N_3443);
nand U4312 (N_4312,N_3461,N_3884);
and U4313 (N_4313,N_3945,N_3556);
xnor U4314 (N_4314,N_3229,N_3044);
nand U4315 (N_4315,N_3955,N_3507);
and U4316 (N_4316,N_3964,N_3288);
nor U4317 (N_4317,N_3880,N_3457);
and U4318 (N_4318,N_3688,N_3503);
or U4319 (N_4319,N_3551,N_3234);
nand U4320 (N_4320,N_3035,N_3633);
xnor U4321 (N_4321,N_3804,N_3628);
and U4322 (N_4322,N_3986,N_3166);
nand U4323 (N_4323,N_3099,N_3765);
nand U4324 (N_4324,N_3359,N_3152);
and U4325 (N_4325,N_3815,N_3742);
or U4326 (N_4326,N_3877,N_3796);
and U4327 (N_4327,N_3661,N_3930);
xor U4328 (N_4328,N_3779,N_3250);
nand U4329 (N_4329,N_3719,N_3550);
nor U4330 (N_4330,N_3802,N_3453);
xnor U4331 (N_4331,N_3732,N_3951);
or U4332 (N_4332,N_3232,N_3994);
nand U4333 (N_4333,N_3139,N_3388);
nor U4334 (N_4334,N_3759,N_3239);
nand U4335 (N_4335,N_3876,N_3981);
nor U4336 (N_4336,N_3579,N_3991);
and U4337 (N_4337,N_3595,N_3323);
or U4338 (N_4338,N_3216,N_3578);
nor U4339 (N_4339,N_3258,N_3207);
nand U4340 (N_4340,N_3908,N_3054);
nor U4341 (N_4341,N_3728,N_3280);
and U4342 (N_4342,N_3509,N_3291);
and U4343 (N_4343,N_3830,N_3196);
nand U4344 (N_4344,N_3751,N_3907);
or U4345 (N_4345,N_3977,N_3616);
nand U4346 (N_4346,N_3172,N_3103);
and U4347 (N_4347,N_3489,N_3061);
nor U4348 (N_4348,N_3632,N_3178);
and U4349 (N_4349,N_3265,N_3247);
xnor U4350 (N_4350,N_3501,N_3067);
and U4351 (N_4351,N_3029,N_3260);
nor U4352 (N_4352,N_3069,N_3762);
nor U4353 (N_4353,N_3764,N_3439);
and U4354 (N_4354,N_3999,N_3777);
nand U4355 (N_4355,N_3786,N_3718);
or U4356 (N_4356,N_3198,N_3255);
or U4357 (N_4357,N_3413,N_3231);
nor U4358 (N_4358,N_3332,N_3098);
nor U4359 (N_4359,N_3176,N_3989);
and U4360 (N_4360,N_3729,N_3317);
xor U4361 (N_4361,N_3553,N_3108);
xnor U4362 (N_4362,N_3079,N_3929);
and U4363 (N_4363,N_3839,N_3925);
or U4364 (N_4364,N_3516,N_3107);
or U4365 (N_4365,N_3093,N_3336);
nand U4366 (N_4366,N_3944,N_3865);
nand U4367 (N_4367,N_3997,N_3400);
nand U4368 (N_4368,N_3954,N_3716);
or U4369 (N_4369,N_3271,N_3436);
nand U4370 (N_4370,N_3957,N_3747);
nor U4371 (N_4371,N_3775,N_3364);
nand U4372 (N_4372,N_3469,N_3643);
and U4373 (N_4373,N_3548,N_3627);
nor U4374 (N_4374,N_3534,N_3817);
and U4375 (N_4375,N_3901,N_3746);
and U4376 (N_4376,N_3155,N_3648);
or U4377 (N_4377,N_3376,N_3894);
or U4378 (N_4378,N_3148,N_3327);
xor U4379 (N_4379,N_3584,N_3935);
nor U4380 (N_4380,N_3454,N_3002);
nor U4381 (N_4381,N_3848,N_3971);
nor U4382 (N_4382,N_3970,N_3686);
nand U4383 (N_4383,N_3168,N_3963);
nor U4384 (N_4384,N_3879,N_3604);
nand U4385 (N_4385,N_3824,N_3816);
or U4386 (N_4386,N_3267,N_3226);
nand U4387 (N_4387,N_3411,N_3227);
nand U4388 (N_4388,N_3829,N_3355);
nand U4389 (N_4389,N_3404,N_3671);
or U4390 (N_4390,N_3414,N_3235);
nor U4391 (N_4391,N_3360,N_3582);
nand U4392 (N_4392,N_3998,N_3463);
or U4393 (N_4393,N_3803,N_3996);
nand U4394 (N_4394,N_3023,N_3897);
nor U4395 (N_4395,N_3780,N_3783);
nor U4396 (N_4396,N_3171,N_3914);
xor U4397 (N_4397,N_3307,N_3353);
and U4398 (N_4398,N_3379,N_3808);
nor U4399 (N_4399,N_3822,N_3348);
nand U4400 (N_4400,N_3125,N_3903);
and U4401 (N_4401,N_3939,N_3244);
xnor U4402 (N_4402,N_3559,N_3748);
nor U4403 (N_4403,N_3569,N_3396);
and U4404 (N_4404,N_3645,N_3771);
nor U4405 (N_4405,N_3109,N_3074);
nor U4406 (N_4406,N_3734,N_3058);
nor U4407 (N_4407,N_3329,N_3471);
or U4408 (N_4408,N_3705,N_3926);
nand U4409 (N_4409,N_3057,N_3557);
xnor U4410 (N_4410,N_3878,N_3340);
xnor U4411 (N_4411,N_3723,N_3562);
nand U4412 (N_4412,N_3370,N_3357);
and U4413 (N_4413,N_3194,N_3456);
and U4414 (N_4414,N_3434,N_3526);
nand U4415 (N_4415,N_3967,N_3018);
or U4416 (N_4416,N_3788,N_3111);
nand U4417 (N_4417,N_3608,N_3432);
or U4418 (N_4418,N_3147,N_3283);
nor U4419 (N_4419,N_3007,N_3238);
nand U4420 (N_4420,N_3302,N_3835);
and U4421 (N_4421,N_3927,N_3862);
or U4422 (N_4422,N_3224,N_3773);
nor U4423 (N_4423,N_3095,N_3843);
nor U4424 (N_4424,N_3730,N_3937);
or U4425 (N_4425,N_3833,N_3444);
or U4426 (N_4426,N_3040,N_3146);
nand U4427 (N_4427,N_3610,N_3144);
nand U4428 (N_4428,N_3669,N_3181);
or U4429 (N_4429,N_3358,N_3480);
nor U4430 (N_4430,N_3028,N_3692);
nor U4431 (N_4431,N_3545,N_3496);
or U4432 (N_4432,N_3676,N_3846);
nand U4433 (N_4433,N_3214,N_3421);
nand U4434 (N_4434,N_3344,N_3813);
nor U4435 (N_4435,N_3027,N_3034);
and U4436 (N_4436,N_3995,N_3859);
nor U4437 (N_4437,N_3222,N_3795);
and U4438 (N_4438,N_3965,N_3202);
xnor U4439 (N_4439,N_3416,N_3273);
and U4440 (N_4440,N_3460,N_3852);
or U4441 (N_4441,N_3522,N_3667);
and U4442 (N_4442,N_3893,N_3543);
or U4443 (N_4443,N_3638,N_3781);
or U4444 (N_4444,N_3373,N_3984);
and U4445 (N_4445,N_3134,N_3112);
nor U4446 (N_4446,N_3285,N_3446);
and U4447 (N_4447,N_3555,N_3405);
nor U4448 (N_4448,N_3820,N_3420);
or U4449 (N_4449,N_3767,N_3113);
nor U4450 (N_4450,N_3586,N_3449);
and U4451 (N_4451,N_3666,N_3311);
or U4452 (N_4452,N_3272,N_3252);
and U4453 (N_4453,N_3025,N_3602);
nand U4454 (N_4454,N_3910,N_3193);
or U4455 (N_4455,N_3650,N_3149);
or U4456 (N_4456,N_3213,N_3450);
or U4457 (N_4457,N_3823,N_3477);
nand U4458 (N_4458,N_3241,N_3792);
or U4459 (N_4459,N_3106,N_3857);
nor U4460 (N_4460,N_3371,N_3429);
or U4461 (N_4461,N_3289,N_3197);
nand U4462 (N_4462,N_3758,N_3304);
or U4463 (N_4463,N_3749,N_3533);
nor U4464 (N_4464,N_3320,N_3296);
nand U4465 (N_4465,N_3142,N_3132);
and U4466 (N_4466,N_3455,N_3270);
or U4467 (N_4467,N_3389,N_3187);
and U4468 (N_4468,N_3512,N_3685);
or U4469 (N_4469,N_3486,N_3902);
nand U4470 (N_4470,N_3982,N_3673);
or U4471 (N_4471,N_3919,N_3760);
and U4472 (N_4472,N_3259,N_3135);
nand U4473 (N_4473,N_3055,N_3254);
nor U4474 (N_4474,N_3720,N_3407);
nand U4475 (N_4475,N_3679,N_3365);
nor U4476 (N_4476,N_3366,N_3081);
and U4477 (N_4477,N_3188,N_3419);
xnor U4478 (N_4478,N_3090,N_3306);
nor U4479 (N_4479,N_3615,N_3298);
and U4480 (N_4480,N_3909,N_3847);
nand U4481 (N_4481,N_3572,N_3487);
nand U4482 (N_4482,N_3189,N_3744);
nand U4483 (N_4483,N_3737,N_3506);
or U4484 (N_4484,N_3279,N_3341);
nand U4485 (N_4485,N_3535,N_3024);
and U4486 (N_4486,N_3158,N_3858);
xor U4487 (N_4487,N_3162,N_3075);
nor U4488 (N_4488,N_3942,N_3326);
nor U4489 (N_4489,N_3354,N_3039);
nor U4490 (N_4490,N_3649,N_3225);
xnor U4491 (N_4491,N_3485,N_3990);
nor U4492 (N_4492,N_3426,N_3670);
or U4493 (N_4493,N_3849,N_3678);
xnor U4494 (N_4494,N_3906,N_3960);
xnor U4495 (N_4495,N_3305,N_3581);
or U4496 (N_4496,N_3869,N_3084);
nand U4497 (N_4497,N_3174,N_3333);
or U4498 (N_4498,N_3475,N_3738);
and U4499 (N_4499,N_3755,N_3753);
or U4500 (N_4500,N_3001,N_3454);
or U4501 (N_4501,N_3249,N_3618);
nor U4502 (N_4502,N_3319,N_3168);
nand U4503 (N_4503,N_3649,N_3000);
nand U4504 (N_4504,N_3868,N_3254);
and U4505 (N_4505,N_3468,N_3950);
nor U4506 (N_4506,N_3195,N_3744);
and U4507 (N_4507,N_3038,N_3798);
nor U4508 (N_4508,N_3569,N_3867);
and U4509 (N_4509,N_3007,N_3500);
nand U4510 (N_4510,N_3859,N_3040);
xor U4511 (N_4511,N_3766,N_3930);
or U4512 (N_4512,N_3778,N_3458);
nand U4513 (N_4513,N_3087,N_3776);
and U4514 (N_4514,N_3356,N_3422);
xnor U4515 (N_4515,N_3110,N_3344);
nor U4516 (N_4516,N_3766,N_3294);
or U4517 (N_4517,N_3648,N_3978);
and U4518 (N_4518,N_3814,N_3584);
or U4519 (N_4519,N_3863,N_3455);
and U4520 (N_4520,N_3593,N_3685);
nor U4521 (N_4521,N_3970,N_3359);
nand U4522 (N_4522,N_3820,N_3273);
and U4523 (N_4523,N_3363,N_3967);
nor U4524 (N_4524,N_3292,N_3670);
and U4525 (N_4525,N_3270,N_3046);
or U4526 (N_4526,N_3730,N_3848);
nand U4527 (N_4527,N_3584,N_3993);
or U4528 (N_4528,N_3628,N_3332);
nor U4529 (N_4529,N_3006,N_3936);
nand U4530 (N_4530,N_3020,N_3238);
or U4531 (N_4531,N_3935,N_3133);
and U4532 (N_4532,N_3727,N_3494);
nor U4533 (N_4533,N_3887,N_3220);
nor U4534 (N_4534,N_3411,N_3325);
or U4535 (N_4535,N_3637,N_3256);
nand U4536 (N_4536,N_3159,N_3964);
nor U4537 (N_4537,N_3336,N_3493);
nand U4538 (N_4538,N_3624,N_3200);
xnor U4539 (N_4539,N_3314,N_3269);
nor U4540 (N_4540,N_3471,N_3714);
or U4541 (N_4541,N_3973,N_3183);
and U4542 (N_4542,N_3485,N_3447);
or U4543 (N_4543,N_3647,N_3694);
nor U4544 (N_4544,N_3779,N_3664);
or U4545 (N_4545,N_3673,N_3432);
nor U4546 (N_4546,N_3678,N_3716);
and U4547 (N_4547,N_3398,N_3634);
xor U4548 (N_4548,N_3926,N_3232);
nor U4549 (N_4549,N_3640,N_3916);
or U4550 (N_4550,N_3469,N_3963);
and U4551 (N_4551,N_3409,N_3363);
and U4552 (N_4552,N_3417,N_3794);
nand U4553 (N_4553,N_3801,N_3642);
nor U4554 (N_4554,N_3471,N_3861);
or U4555 (N_4555,N_3521,N_3083);
and U4556 (N_4556,N_3454,N_3631);
and U4557 (N_4557,N_3186,N_3444);
and U4558 (N_4558,N_3307,N_3407);
or U4559 (N_4559,N_3437,N_3293);
or U4560 (N_4560,N_3292,N_3917);
or U4561 (N_4561,N_3288,N_3013);
or U4562 (N_4562,N_3048,N_3329);
nand U4563 (N_4563,N_3648,N_3387);
nand U4564 (N_4564,N_3067,N_3880);
or U4565 (N_4565,N_3505,N_3897);
xnor U4566 (N_4566,N_3085,N_3961);
xor U4567 (N_4567,N_3974,N_3405);
and U4568 (N_4568,N_3460,N_3848);
or U4569 (N_4569,N_3294,N_3559);
and U4570 (N_4570,N_3898,N_3180);
nor U4571 (N_4571,N_3207,N_3978);
nand U4572 (N_4572,N_3406,N_3550);
nor U4573 (N_4573,N_3209,N_3915);
nor U4574 (N_4574,N_3866,N_3801);
and U4575 (N_4575,N_3404,N_3132);
or U4576 (N_4576,N_3216,N_3900);
and U4577 (N_4577,N_3923,N_3979);
nand U4578 (N_4578,N_3354,N_3152);
and U4579 (N_4579,N_3106,N_3305);
nor U4580 (N_4580,N_3097,N_3418);
nor U4581 (N_4581,N_3139,N_3807);
nor U4582 (N_4582,N_3560,N_3923);
nor U4583 (N_4583,N_3874,N_3096);
or U4584 (N_4584,N_3798,N_3569);
and U4585 (N_4585,N_3299,N_3079);
or U4586 (N_4586,N_3095,N_3744);
or U4587 (N_4587,N_3281,N_3027);
and U4588 (N_4588,N_3843,N_3003);
nand U4589 (N_4589,N_3258,N_3889);
or U4590 (N_4590,N_3199,N_3773);
nor U4591 (N_4591,N_3933,N_3892);
and U4592 (N_4592,N_3559,N_3488);
xnor U4593 (N_4593,N_3024,N_3107);
and U4594 (N_4594,N_3155,N_3768);
nor U4595 (N_4595,N_3162,N_3231);
xnor U4596 (N_4596,N_3063,N_3629);
nor U4597 (N_4597,N_3092,N_3868);
xnor U4598 (N_4598,N_3172,N_3595);
or U4599 (N_4599,N_3792,N_3250);
xor U4600 (N_4600,N_3429,N_3222);
or U4601 (N_4601,N_3092,N_3629);
nor U4602 (N_4602,N_3070,N_3491);
nand U4603 (N_4603,N_3526,N_3449);
nor U4604 (N_4604,N_3189,N_3307);
nand U4605 (N_4605,N_3257,N_3966);
or U4606 (N_4606,N_3634,N_3145);
and U4607 (N_4607,N_3863,N_3725);
nor U4608 (N_4608,N_3729,N_3706);
or U4609 (N_4609,N_3146,N_3817);
and U4610 (N_4610,N_3543,N_3058);
or U4611 (N_4611,N_3362,N_3115);
or U4612 (N_4612,N_3082,N_3734);
xor U4613 (N_4613,N_3440,N_3038);
nor U4614 (N_4614,N_3489,N_3397);
and U4615 (N_4615,N_3641,N_3587);
or U4616 (N_4616,N_3095,N_3508);
nor U4617 (N_4617,N_3868,N_3701);
or U4618 (N_4618,N_3535,N_3869);
nand U4619 (N_4619,N_3276,N_3060);
nor U4620 (N_4620,N_3042,N_3050);
nor U4621 (N_4621,N_3682,N_3976);
nor U4622 (N_4622,N_3132,N_3107);
nor U4623 (N_4623,N_3925,N_3798);
or U4624 (N_4624,N_3028,N_3001);
or U4625 (N_4625,N_3062,N_3556);
nand U4626 (N_4626,N_3590,N_3737);
or U4627 (N_4627,N_3248,N_3323);
or U4628 (N_4628,N_3848,N_3236);
nand U4629 (N_4629,N_3293,N_3427);
or U4630 (N_4630,N_3164,N_3094);
nor U4631 (N_4631,N_3948,N_3565);
nor U4632 (N_4632,N_3458,N_3255);
nor U4633 (N_4633,N_3981,N_3808);
xnor U4634 (N_4634,N_3058,N_3266);
or U4635 (N_4635,N_3558,N_3336);
nor U4636 (N_4636,N_3750,N_3590);
and U4637 (N_4637,N_3008,N_3086);
and U4638 (N_4638,N_3955,N_3644);
or U4639 (N_4639,N_3539,N_3904);
nand U4640 (N_4640,N_3868,N_3028);
nor U4641 (N_4641,N_3723,N_3077);
nor U4642 (N_4642,N_3200,N_3552);
or U4643 (N_4643,N_3403,N_3639);
nor U4644 (N_4644,N_3202,N_3734);
nand U4645 (N_4645,N_3342,N_3109);
nand U4646 (N_4646,N_3731,N_3861);
nor U4647 (N_4647,N_3284,N_3950);
nand U4648 (N_4648,N_3813,N_3129);
or U4649 (N_4649,N_3752,N_3279);
and U4650 (N_4650,N_3696,N_3335);
nand U4651 (N_4651,N_3741,N_3483);
nand U4652 (N_4652,N_3987,N_3109);
nor U4653 (N_4653,N_3888,N_3820);
nand U4654 (N_4654,N_3473,N_3074);
and U4655 (N_4655,N_3914,N_3611);
nor U4656 (N_4656,N_3616,N_3621);
or U4657 (N_4657,N_3298,N_3155);
or U4658 (N_4658,N_3638,N_3955);
and U4659 (N_4659,N_3172,N_3076);
nor U4660 (N_4660,N_3699,N_3020);
nand U4661 (N_4661,N_3028,N_3385);
nor U4662 (N_4662,N_3460,N_3032);
nor U4663 (N_4663,N_3486,N_3287);
or U4664 (N_4664,N_3273,N_3248);
nor U4665 (N_4665,N_3717,N_3501);
or U4666 (N_4666,N_3344,N_3912);
nand U4667 (N_4667,N_3514,N_3446);
and U4668 (N_4668,N_3986,N_3618);
nand U4669 (N_4669,N_3183,N_3273);
or U4670 (N_4670,N_3148,N_3781);
or U4671 (N_4671,N_3483,N_3994);
xnor U4672 (N_4672,N_3725,N_3642);
and U4673 (N_4673,N_3056,N_3223);
nor U4674 (N_4674,N_3517,N_3680);
nand U4675 (N_4675,N_3725,N_3929);
or U4676 (N_4676,N_3613,N_3678);
xnor U4677 (N_4677,N_3773,N_3189);
and U4678 (N_4678,N_3881,N_3764);
xnor U4679 (N_4679,N_3670,N_3789);
and U4680 (N_4680,N_3805,N_3507);
nor U4681 (N_4681,N_3993,N_3292);
nand U4682 (N_4682,N_3611,N_3413);
and U4683 (N_4683,N_3654,N_3742);
nor U4684 (N_4684,N_3244,N_3176);
xor U4685 (N_4685,N_3851,N_3197);
or U4686 (N_4686,N_3822,N_3860);
xor U4687 (N_4687,N_3626,N_3961);
xor U4688 (N_4688,N_3112,N_3377);
and U4689 (N_4689,N_3037,N_3536);
or U4690 (N_4690,N_3722,N_3476);
or U4691 (N_4691,N_3942,N_3415);
nand U4692 (N_4692,N_3561,N_3683);
nor U4693 (N_4693,N_3375,N_3094);
nand U4694 (N_4694,N_3923,N_3513);
nor U4695 (N_4695,N_3882,N_3005);
and U4696 (N_4696,N_3778,N_3052);
nand U4697 (N_4697,N_3031,N_3806);
xor U4698 (N_4698,N_3275,N_3868);
and U4699 (N_4699,N_3494,N_3703);
or U4700 (N_4700,N_3811,N_3238);
or U4701 (N_4701,N_3658,N_3130);
xor U4702 (N_4702,N_3860,N_3731);
nor U4703 (N_4703,N_3117,N_3975);
or U4704 (N_4704,N_3991,N_3539);
and U4705 (N_4705,N_3872,N_3363);
nor U4706 (N_4706,N_3480,N_3743);
nand U4707 (N_4707,N_3059,N_3016);
nand U4708 (N_4708,N_3868,N_3727);
or U4709 (N_4709,N_3724,N_3132);
nor U4710 (N_4710,N_3212,N_3513);
and U4711 (N_4711,N_3788,N_3548);
and U4712 (N_4712,N_3586,N_3572);
and U4713 (N_4713,N_3982,N_3312);
nand U4714 (N_4714,N_3350,N_3470);
and U4715 (N_4715,N_3332,N_3974);
nand U4716 (N_4716,N_3447,N_3251);
nand U4717 (N_4717,N_3499,N_3564);
nand U4718 (N_4718,N_3584,N_3332);
or U4719 (N_4719,N_3575,N_3270);
and U4720 (N_4720,N_3019,N_3695);
xnor U4721 (N_4721,N_3753,N_3688);
nand U4722 (N_4722,N_3936,N_3094);
or U4723 (N_4723,N_3692,N_3237);
nor U4724 (N_4724,N_3621,N_3257);
or U4725 (N_4725,N_3057,N_3946);
or U4726 (N_4726,N_3628,N_3789);
or U4727 (N_4727,N_3483,N_3240);
and U4728 (N_4728,N_3646,N_3044);
xnor U4729 (N_4729,N_3789,N_3386);
nor U4730 (N_4730,N_3820,N_3224);
nand U4731 (N_4731,N_3073,N_3480);
and U4732 (N_4732,N_3224,N_3857);
nand U4733 (N_4733,N_3494,N_3726);
nor U4734 (N_4734,N_3447,N_3506);
xnor U4735 (N_4735,N_3116,N_3961);
or U4736 (N_4736,N_3776,N_3467);
and U4737 (N_4737,N_3027,N_3410);
or U4738 (N_4738,N_3055,N_3230);
or U4739 (N_4739,N_3431,N_3619);
and U4740 (N_4740,N_3584,N_3853);
nor U4741 (N_4741,N_3667,N_3880);
and U4742 (N_4742,N_3589,N_3379);
xnor U4743 (N_4743,N_3574,N_3270);
nand U4744 (N_4744,N_3533,N_3625);
nor U4745 (N_4745,N_3282,N_3223);
nor U4746 (N_4746,N_3082,N_3492);
nor U4747 (N_4747,N_3791,N_3445);
or U4748 (N_4748,N_3327,N_3297);
nor U4749 (N_4749,N_3387,N_3298);
and U4750 (N_4750,N_3629,N_3515);
or U4751 (N_4751,N_3165,N_3662);
nor U4752 (N_4752,N_3448,N_3139);
nand U4753 (N_4753,N_3697,N_3653);
nor U4754 (N_4754,N_3909,N_3301);
nor U4755 (N_4755,N_3877,N_3149);
nor U4756 (N_4756,N_3971,N_3946);
nand U4757 (N_4757,N_3862,N_3811);
nand U4758 (N_4758,N_3628,N_3753);
nand U4759 (N_4759,N_3345,N_3871);
nand U4760 (N_4760,N_3104,N_3470);
or U4761 (N_4761,N_3082,N_3130);
and U4762 (N_4762,N_3453,N_3590);
nor U4763 (N_4763,N_3311,N_3166);
nand U4764 (N_4764,N_3189,N_3609);
or U4765 (N_4765,N_3356,N_3577);
or U4766 (N_4766,N_3833,N_3060);
nor U4767 (N_4767,N_3184,N_3870);
nand U4768 (N_4768,N_3780,N_3416);
nand U4769 (N_4769,N_3604,N_3266);
nand U4770 (N_4770,N_3609,N_3296);
and U4771 (N_4771,N_3706,N_3238);
and U4772 (N_4772,N_3369,N_3763);
and U4773 (N_4773,N_3495,N_3682);
nor U4774 (N_4774,N_3322,N_3877);
xnor U4775 (N_4775,N_3913,N_3524);
nand U4776 (N_4776,N_3975,N_3647);
or U4777 (N_4777,N_3400,N_3073);
nand U4778 (N_4778,N_3681,N_3114);
xnor U4779 (N_4779,N_3159,N_3075);
nor U4780 (N_4780,N_3241,N_3859);
and U4781 (N_4781,N_3658,N_3274);
and U4782 (N_4782,N_3350,N_3870);
nand U4783 (N_4783,N_3051,N_3378);
nor U4784 (N_4784,N_3495,N_3869);
or U4785 (N_4785,N_3754,N_3858);
xor U4786 (N_4786,N_3213,N_3053);
nand U4787 (N_4787,N_3313,N_3032);
or U4788 (N_4788,N_3659,N_3529);
and U4789 (N_4789,N_3001,N_3570);
and U4790 (N_4790,N_3283,N_3952);
nand U4791 (N_4791,N_3179,N_3485);
nor U4792 (N_4792,N_3267,N_3044);
nand U4793 (N_4793,N_3236,N_3494);
or U4794 (N_4794,N_3527,N_3634);
and U4795 (N_4795,N_3360,N_3260);
or U4796 (N_4796,N_3099,N_3775);
nand U4797 (N_4797,N_3416,N_3182);
or U4798 (N_4798,N_3774,N_3102);
nor U4799 (N_4799,N_3677,N_3121);
and U4800 (N_4800,N_3633,N_3838);
nand U4801 (N_4801,N_3410,N_3189);
or U4802 (N_4802,N_3502,N_3770);
or U4803 (N_4803,N_3284,N_3243);
or U4804 (N_4804,N_3266,N_3854);
nor U4805 (N_4805,N_3871,N_3326);
and U4806 (N_4806,N_3180,N_3437);
nand U4807 (N_4807,N_3228,N_3978);
or U4808 (N_4808,N_3151,N_3072);
nand U4809 (N_4809,N_3869,N_3309);
and U4810 (N_4810,N_3087,N_3747);
and U4811 (N_4811,N_3609,N_3567);
nand U4812 (N_4812,N_3715,N_3874);
and U4813 (N_4813,N_3284,N_3405);
or U4814 (N_4814,N_3881,N_3331);
and U4815 (N_4815,N_3949,N_3501);
or U4816 (N_4816,N_3749,N_3993);
nand U4817 (N_4817,N_3508,N_3465);
and U4818 (N_4818,N_3429,N_3208);
nand U4819 (N_4819,N_3912,N_3868);
and U4820 (N_4820,N_3276,N_3659);
nand U4821 (N_4821,N_3763,N_3414);
nand U4822 (N_4822,N_3491,N_3852);
xnor U4823 (N_4823,N_3505,N_3392);
and U4824 (N_4824,N_3823,N_3005);
and U4825 (N_4825,N_3412,N_3577);
xor U4826 (N_4826,N_3987,N_3421);
xor U4827 (N_4827,N_3071,N_3044);
nand U4828 (N_4828,N_3470,N_3447);
or U4829 (N_4829,N_3450,N_3734);
nor U4830 (N_4830,N_3284,N_3740);
and U4831 (N_4831,N_3664,N_3382);
nor U4832 (N_4832,N_3628,N_3827);
and U4833 (N_4833,N_3758,N_3515);
nor U4834 (N_4834,N_3444,N_3552);
or U4835 (N_4835,N_3429,N_3059);
or U4836 (N_4836,N_3531,N_3678);
nand U4837 (N_4837,N_3004,N_3512);
or U4838 (N_4838,N_3291,N_3346);
nand U4839 (N_4839,N_3495,N_3829);
and U4840 (N_4840,N_3000,N_3038);
nand U4841 (N_4841,N_3281,N_3185);
or U4842 (N_4842,N_3968,N_3300);
nor U4843 (N_4843,N_3156,N_3146);
or U4844 (N_4844,N_3697,N_3148);
or U4845 (N_4845,N_3066,N_3601);
nand U4846 (N_4846,N_3290,N_3199);
and U4847 (N_4847,N_3955,N_3570);
xnor U4848 (N_4848,N_3999,N_3143);
or U4849 (N_4849,N_3698,N_3894);
xnor U4850 (N_4850,N_3045,N_3108);
or U4851 (N_4851,N_3482,N_3211);
and U4852 (N_4852,N_3442,N_3853);
nor U4853 (N_4853,N_3377,N_3876);
xnor U4854 (N_4854,N_3150,N_3396);
nor U4855 (N_4855,N_3789,N_3179);
nand U4856 (N_4856,N_3157,N_3862);
nand U4857 (N_4857,N_3342,N_3325);
nor U4858 (N_4858,N_3051,N_3213);
and U4859 (N_4859,N_3726,N_3924);
nand U4860 (N_4860,N_3273,N_3964);
nor U4861 (N_4861,N_3571,N_3393);
nand U4862 (N_4862,N_3352,N_3597);
nor U4863 (N_4863,N_3945,N_3886);
nand U4864 (N_4864,N_3645,N_3065);
nand U4865 (N_4865,N_3889,N_3493);
and U4866 (N_4866,N_3910,N_3579);
nand U4867 (N_4867,N_3385,N_3615);
or U4868 (N_4868,N_3228,N_3557);
nand U4869 (N_4869,N_3407,N_3567);
nand U4870 (N_4870,N_3254,N_3625);
nand U4871 (N_4871,N_3011,N_3203);
and U4872 (N_4872,N_3729,N_3637);
and U4873 (N_4873,N_3459,N_3448);
xnor U4874 (N_4874,N_3602,N_3722);
and U4875 (N_4875,N_3104,N_3397);
or U4876 (N_4876,N_3213,N_3329);
nand U4877 (N_4877,N_3267,N_3843);
nor U4878 (N_4878,N_3396,N_3074);
and U4879 (N_4879,N_3219,N_3888);
or U4880 (N_4880,N_3788,N_3497);
nor U4881 (N_4881,N_3641,N_3491);
nor U4882 (N_4882,N_3630,N_3627);
nor U4883 (N_4883,N_3660,N_3088);
or U4884 (N_4884,N_3337,N_3556);
nor U4885 (N_4885,N_3841,N_3019);
xnor U4886 (N_4886,N_3001,N_3816);
nand U4887 (N_4887,N_3039,N_3592);
or U4888 (N_4888,N_3620,N_3551);
nor U4889 (N_4889,N_3187,N_3200);
and U4890 (N_4890,N_3835,N_3327);
nor U4891 (N_4891,N_3391,N_3943);
nand U4892 (N_4892,N_3558,N_3301);
or U4893 (N_4893,N_3533,N_3761);
and U4894 (N_4894,N_3570,N_3007);
xnor U4895 (N_4895,N_3771,N_3563);
or U4896 (N_4896,N_3896,N_3999);
and U4897 (N_4897,N_3616,N_3376);
nand U4898 (N_4898,N_3131,N_3645);
xor U4899 (N_4899,N_3815,N_3526);
nand U4900 (N_4900,N_3900,N_3656);
nor U4901 (N_4901,N_3752,N_3558);
nand U4902 (N_4902,N_3419,N_3117);
nand U4903 (N_4903,N_3915,N_3295);
nand U4904 (N_4904,N_3027,N_3048);
and U4905 (N_4905,N_3775,N_3109);
nor U4906 (N_4906,N_3456,N_3376);
and U4907 (N_4907,N_3702,N_3554);
or U4908 (N_4908,N_3010,N_3284);
or U4909 (N_4909,N_3676,N_3564);
and U4910 (N_4910,N_3556,N_3144);
nor U4911 (N_4911,N_3498,N_3182);
nor U4912 (N_4912,N_3503,N_3127);
nor U4913 (N_4913,N_3371,N_3682);
and U4914 (N_4914,N_3916,N_3784);
or U4915 (N_4915,N_3554,N_3662);
nand U4916 (N_4916,N_3093,N_3270);
or U4917 (N_4917,N_3752,N_3679);
or U4918 (N_4918,N_3968,N_3173);
or U4919 (N_4919,N_3622,N_3024);
and U4920 (N_4920,N_3729,N_3162);
nor U4921 (N_4921,N_3601,N_3240);
nor U4922 (N_4922,N_3310,N_3338);
and U4923 (N_4923,N_3248,N_3655);
nand U4924 (N_4924,N_3712,N_3193);
and U4925 (N_4925,N_3255,N_3158);
nand U4926 (N_4926,N_3884,N_3153);
or U4927 (N_4927,N_3956,N_3879);
and U4928 (N_4928,N_3769,N_3303);
or U4929 (N_4929,N_3441,N_3266);
and U4930 (N_4930,N_3273,N_3826);
or U4931 (N_4931,N_3424,N_3977);
or U4932 (N_4932,N_3358,N_3268);
xnor U4933 (N_4933,N_3691,N_3022);
nand U4934 (N_4934,N_3219,N_3796);
or U4935 (N_4935,N_3087,N_3624);
nand U4936 (N_4936,N_3284,N_3075);
or U4937 (N_4937,N_3545,N_3914);
nand U4938 (N_4938,N_3922,N_3481);
and U4939 (N_4939,N_3560,N_3872);
xnor U4940 (N_4940,N_3304,N_3358);
nand U4941 (N_4941,N_3660,N_3039);
and U4942 (N_4942,N_3566,N_3732);
nor U4943 (N_4943,N_3087,N_3281);
nand U4944 (N_4944,N_3145,N_3698);
or U4945 (N_4945,N_3233,N_3879);
or U4946 (N_4946,N_3146,N_3498);
or U4947 (N_4947,N_3530,N_3277);
and U4948 (N_4948,N_3602,N_3763);
and U4949 (N_4949,N_3561,N_3267);
xor U4950 (N_4950,N_3794,N_3412);
or U4951 (N_4951,N_3875,N_3536);
nand U4952 (N_4952,N_3530,N_3722);
and U4953 (N_4953,N_3084,N_3937);
nor U4954 (N_4954,N_3666,N_3609);
nand U4955 (N_4955,N_3201,N_3637);
or U4956 (N_4956,N_3599,N_3263);
or U4957 (N_4957,N_3553,N_3802);
or U4958 (N_4958,N_3374,N_3262);
nor U4959 (N_4959,N_3698,N_3676);
nand U4960 (N_4960,N_3742,N_3932);
or U4961 (N_4961,N_3677,N_3685);
nand U4962 (N_4962,N_3703,N_3109);
or U4963 (N_4963,N_3087,N_3343);
nand U4964 (N_4964,N_3510,N_3548);
nor U4965 (N_4965,N_3400,N_3268);
and U4966 (N_4966,N_3260,N_3822);
xnor U4967 (N_4967,N_3604,N_3774);
nor U4968 (N_4968,N_3094,N_3051);
or U4969 (N_4969,N_3200,N_3766);
xnor U4970 (N_4970,N_3192,N_3338);
nor U4971 (N_4971,N_3713,N_3255);
nor U4972 (N_4972,N_3607,N_3116);
nor U4973 (N_4973,N_3385,N_3382);
or U4974 (N_4974,N_3741,N_3951);
xnor U4975 (N_4975,N_3807,N_3946);
or U4976 (N_4976,N_3165,N_3171);
nand U4977 (N_4977,N_3767,N_3772);
nand U4978 (N_4978,N_3729,N_3518);
nand U4979 (N_4979,N_3911,N_3545);
or U4980 (N_4980,N_3944,N_3718);
nand U4981 (N_4981,N_3962,N_3139);
nor U4982 (N_4982,N_3519,N_3521);
or U4983 (N_4983,N_3225,N_3545);
nand U4984 (N_4984,N_3863,N_3873);
and U4985 (N_4985,N_3823,N_3071);
xnor U4986 (N_4986,N_3781,N_3850);
and U4987 (N_4987,N_3050,N_3774);
nand U4988 (N_4988,N_3012,N_3496);
nor U4989 (N_4989,N_3285,N_3684);
or U4990 (N_4990,N_3537,N_3503);
nand U4991 (N_4991,N_3868,N_3145);
or U4992 (N_4992,N_3932,N_3379);
nor U4993 (N_4993,N_3840,N_3468);
and U4994 (N_4994,N_3853,N_3711);
xor U4995 (N_4995,N_3531,N_3650);
or U4996 (N_4996,N_3975,N_3756);
nor U4997 (N_4997,N_3316,N_3666);
and U4998 (N_4998,N_3853,N_3517);
and U4999 (N_4999,N_3702,N_3003);
nand U5000 (N_5000,N_4387,N_4504);
nand U5001 (N_5001,N_4374,N_4862);
nand U5002 (N_5002,N_4984,N_4094);
nor U5003 (N_5003,N_4894,N_4695);
nor U5004 (N_5004,N_4304,N_4294);
or U5005 (N_5005,N_4740,N_4453);
and U5006 (N_5006,N_4745,N_4999);
nand U5007 (N_5007,N_4354,N_4156);
nor U5008 (N_5008,N_4035,N_4779);
or U5009 (N_5009,N_4781,N_4028);
nand U5010 (N_5010,N_4213,N_4340);
or U5011 (N_5011,N_4788,N_4001);
nor U5012 (N_5012,N_4382,N_4995);
or U5013 (N_5013,N_4088,N_4582);
or U5014 (N_5014,N_4112,N_4075);
or U5015 (N_5015,N_4404,N_4265);
nor U5016 (N_5016,N_4483,N_4957);
nand U5017 (N_5017,N_4746,N_4816);
and U5018 (N_5018,N_4978,N_4090);
and U5019 (N_5019,N_4983,N_4500);
or U5020 (N_5020,N_4197,N_4043);
and U5021 (N_5021,N_4542,N_4737);
or U5022 (N_5022,N_4425,N_4305);
or U5023 (N_5023,N_4365,N_4243);
nand U5024 (N_5024,N_4630,N_4282);
and U5025 (N_5025,N_4199,N_4108);
or U5026 (N_5026,N_4420,N_4981);
nand U5027 (N_5027,N_4553,N_4550);
nand U5028 (N_5028,N_4171,N_4661);
and U5029 (N_5029,N_4828,N_4878);
nor U5030 (N_5030,N_4893,N_4654);
nand U5031 (N_5031,N_4020,N_4705);
or U5032 (N_5032,N_4371,N_4008);
nand U5033 (N_5033,N_4384,N_4308);
or U5034 (N_5034,N_4170,N_4741);
and U5035 (N_5035,N_4306,N_4773);
and U5036 (N_5036,N_4857,N_4143);
and U5037 (N_5037,N_4877,N_4522);
and U5038 (N_5038,N_4520,N_4934);
and U5039 (N_5039,N_4208,N_4814);
nor U5040 (N_5040,N_4317,N_4244);
and U5041 (N_5041,N_4402,N_4458);
and U5042 (N_5042,N_4764,N_4687);
nand U5043 (N_5043,N_4846,N_4936);
and U5044 (N_5044,N_4168,N_4986);
nor U5045 (N_5045,N_4190,N_4449);
nor U5046 (N_5046,N_4896,N_4397);
and U5047 (N_5047,N_4296,N_4044);
and U5048 (N_5048,N_4355,N_4847);
or U5049 (N_5049,N_4884,N_4584);
and U5050 (N_5050,N_4937,N_4032);
and U5051 (N_5051,N_4069,N_4601);
nand U5052 (N_5052,N_4897,N_4845);
nand U5053 (N_5053,N_4395,N_4195);
nand U5054 (N_5054,N_4417,N_4637);
or U5055 (N_5055,N_4776,N_4376);
and U5056 (N_5056,N_4136,N_4126);
xnor U5057 (N_5057,N_4853,N_4875);
or U5058 (N_5058,N_4130,N_4172);
xor U5059 (N_5059,N_4639,N_4348);
xnor U5060 (N_5060,N_4519,N_4804);
nand U5061 (N_5061,N_4794,N_4971);
nand U5062 (N_5062,N_4769,N_4414);
nor U5063 (N_5063,N_4451,N_4876);
nand U5064 (N_5064,N_4347,N_4429);
and U5065 (N_5065,N_4501,N_4295);
nand U5066 (N_5066,N_4109,N_4714);
nor U5067 (N_5067,N_4569,N_4820);
nand U5068 (N_5068,N_4189,N_4408);
or U5069 (N_5069,N_4290,N_4611);
nand U5070 (N_5070,N_4167,N_4510);
and U5071 (N_5071,N_4092,N_4947);
or U5072 (N_5072,N_4754,N_4797);
and U5073 (N_5073,N_4855,N_4430);
or U5074 (N_5074,N_4410,N_4289);
or U5075 (N_5075,N_4874,N_4074);
xor U5076 (N_5076,N_4684,N_4386);
and U5077 (N_5077,N_4724,N_4676);
nor U5078 (N_5078,N_4956,N_4603);
and U5079 (N_5079,N_4716,N_4196);
nand U5080 (N_5080,N_4176,N_4352);
nand U5081 (N_5081,N_4800,N_4146);
xor U5082 (N_5082,N_4575,N_4907);
and U5083 (N_5083,N_4071,N_4629);
nor U5084 (N_5084,N_4481,N_4418);
nand U5085 (N_5085,N_4924,N_4585);
and U5086 (N_5086,N_4840,N_4186);
and U5087 (N_5087,N_4280,N_4600);
and U5088 (N_5088,N_4320,N_4202);
and U5089 (N_5089,N_4285,N_4318);
and U5090 (N_5090,N_4013,N_4729);
nor U5091 (N_5091,N_4632,N_4996);
nor U5092 (N_5092,N_4759,N_4762);
and U5093 (N_5093,N_4191,N_4682);
xnor U5094 (N_5094,N_4303,N_4822);
or U5095 (N_5095,N_4591,N_4938);
and U5096 (N_5096,N_4038,N_4330);
or U5097 (N_5097,N_4685,N_4061);
and U5098 (N_5098,N_4627,N_4065);
and U5099 (N_5099,N_4832,N_4882);
or U5100 (N_5100,N_4056,N_4660);
nor U5101 (N_5101,N_4771,N_4442);
nor U5102 (N_5102,N_4913,N_4619);
xnor U5103 (N_5103,N_4987,N_4713);
nand U5104 (N_5104,N_4149,N_4815);
nand U5105 (N_5105,N_4869,N_4512);
and U5106 (N_5106,N_4643,N_4666);
and U5107 (N_5107,N_4037,N_4113);
nor U5108 (N_5108,N_4014,N_4989);
or U5109 (N_5109,N_4139,N_4902);
and U5110 (N_5110,N_4283,N_4341);
nand U5111 (N_5111,N_4055,N_4612);
nor U5112 (N_5112,N_4726,N_4183);
or U5113 (N_5113,N_4889,N_4496);
nor U5114 (N_5114,N_4772,N_4091);
or U5115 (N_5115,N_4720,N_4653);
or U5116 (N_5116,N_4050,N_4419);
nor U5117 (N_5117,N_4710,N_4792);
nand U5118 (N_5118,N_4499,N_4524);
xor U5119 (N_5119,N_4187,N_4029);
and U5120 (N_5120,N_4669,N_4118);
nand U5121 (N_5121,N_4642,N_4002);
nor U5122 (N_5122,N_4239,N_4086);
and U5123 (N_5123,N_4329,N_4141);
and U5124 (N_5124,N_4751,N_4537);
nand U5125 (N_5125,N_4786,N_4473);
and U5126 (N_5126,N_4096,N_4678);
nand U5127 (N_5127,N_4604,N_4940);
nand U5128 (N_5128,N_4256,N_4595);
xnor U5129 (N_5129,N_4105,N_4085);
and U5130 (N_5130,N_4078,N_4502);
and U5131 (N_5131,N_4848,N_4058);
and U5132 (N_5132,N_4558,N_4858);
nand U5133 (N_5133,N_4272,N_4808);
or U5134 (N_5134,N_4045,N_4916);
and U5135 (N_5135,N_4931,N_4259);
or U5136 (N_5136,N_4439,N_4403);
and U5137 (N_5137,N_4332,N_4707);
and U5138 (N_5138,N_4556,N_4005);
or U5139 (N_5139,N_4333,N_4979);
or U5140 (N_5140,N_4470,N_4288);
and U5141 (N_5141,N_4150,N_4236);
and U5142 (N_5142,N_4153,N_4812);
nor U5143 (N_5143,N_4049,N_4689);
or U5144 (N_5144,N_4932,N_4227);
and U5145 (N_5145,N_4432,N_4825);
and U5146 (N_5146,N_4693,N_4129);
nand U5147 (N_5147,N_4904,N_4489);
and U5148 (N_5148,N_4818,N_4246);
or U5149 (N_5149,N_4593,N_4405);
or U5150 (N_5150,N_4250,N_4398);
nand U5151 (N_5151,N_4219,N_4515);
nor U5152 (N_5152,N_4588,N_4561);
nor U5153 (N_5153,N_4346,N_4162);
nand U5154 (N_5154,N_4928,N_4155);
nor U5155 (N_5155,N_4597,N_4727);
nand U5156 (N_5156,N_4943,N_4343);
or U5157 (N_5157,N_4444,N_4334);
and U5158 (N_5158,N_4018,N_4338);
nand U5159 (N_5159,N_4665,N_4734);
or U5160 (N_5160,N_4719,N_4253);
and U5161 (N_5161,N_4491,N_4448);
nor U5162 (N_5162,N_4973,N_4711);
or U5163 (N_5163,N_4966,N_4279);
or U5164 (N_5164,N_4933,N_4562);
nand U5165 (N_5165,N_4271,N_4803);
and U5166 (N_5166,N_4640,N_4712);
or U5167 (N_5167,N_4563,N_4704);
or U5168 (N_5168,N_4568,N_4454);
or U5169 (N_5169,N_4344,N_4264);
nor U5170 (N_5170,N_4663,N_4440);
or U5171 (N_5171,N_4472,N_4401);
nand U5172 (N_5172,N_4022,N_4099);
and U5173 (N_5173,N_4513,N_4586);
or U5174 (N_5174,N_4369,N_4854);
or U5175 (N_5175,N_4939,N_4675);
xnor U5176 (N_5176,N_4177,N_4089);
and U5177 (N_5177,N_4951,N_4117);
xor U5178 (N_5178,N_4217,N_4381);
nand U5179 (N_5179,N_4942,N_4421);
or U5180 (N_5180,N_4245,N_4813);
and U5181 (N_5181,N_4912,N_4948);
or U5182 (N_5182,N_4615,N_4976);
or U5183 (N_5183,N_4778,N_4363);
nand U5184 (N_5184,N_4610,N_4215);
nand U5185 (N_5185,N_4485,N_4131);
or U5186 (N_5186,N_4638,N_4645);
nor U5187 (N_5187,N_4165,N_4511);
nor U5188 (N_5188,N_4577,N_4380);
nand U5189 (N_5189,N_4681,N_4574);
nand U5190 (N_5190,N_4313,N_4205);
and U5191 (N_5191,N_4211,N_4406);
xor U5192 (N_5192,N_4154,N_4880);
or U5193 (N_5193,N_4564,N_4400);
nand U5194 (N_5194,N_4225,N_4521);
or U5195 (N_5195,N_4007,N_4337);
or U5196 (N_5196,N_4010,N_4016);
and U5197 (N_5197,N_4908,N_4415);
and U5198 (N_5198,N_4081,N_4378);
nor U5199 (N_5199,N_4635,N_4625);
and U5200 (N_5200,N_4962,N_4609);
and U5201 (N_5201,N_4409,N_4696);
and U5202 (N_5202,N_4624,N_4311);
and U5203 (N_5203,N_4534,N_4299);
and U5204 (N_5204,N_4242,N_4683);
nand U5205 (N_5205,N_4158,N_4443);
nor U5206 (N_5206,N_4752,N_4218);
or U5207 (N_5207,N_4662,N_4407);
or U5208 (N_5208,N_4652,N_4744);
nor U5209 (N_5209,N_4003,N_4412);
nand U5210 (N_5210,N_4068,N_4834);
nand U5211 (N_5211,N_4927,N_4426);
xor U5212 (N_5212,N_4514,N_4743);
or U5213 (N_5213,N_4810,N_4321);
nor U5214 (N_5214,N_4373,N_4900);
nor U5215 (N_5215,N_4025,N_4590);
nor U5216 (N_5216,N_4101,N_4503);
nor U5217 (N_5217,N_4839,N_4416);
and U5218 (N_5218,N_4677,N_4919);
and U5219 (N_5219,N_4230,N_4886);
xnor U5220 (N_5220,N_4709,N_4756);
or U5221 (N_5221,N_4431,N_4725);
nand U5222 (N_5222,N_4819,N_4768);
nand U5223 (N_5223,N_4184,N_4077);
nor U5224 (N_5224,N_4438,N_4326);
nand U5225 (N_5225,N_4671,N_4461);
nand U5226 (N_5226,N_4850,N_4888);
and U5227 (N_5227,N_4555,N_4396);
nand U5228 (N_5228,N_4673,N_4626);
nand U5229 (N_5229,N_4031,N_4132);
and U5230 (N_5230,N_4906,N_4536);
and U5231 (N_5231,N_4753,N_4668);
nand U5232 (N_5232,N_4210,N_4423);
nand U5233 (N_5233,N_4968,N_4982);
nor U5234 (N_5234,N_4004,N_4480);
nand U5235 (N_5235,N_4864,N_4749);
and U5236 (N_5236,N_4970,N_4292);
xor U5237 (N_5237,N_4268,N_4370);
or U5238 (N_5238,N_4809,N_4274);
and U5239 (N_5239,N_4990,N_4103);
or U5240 (N_5240,N_4067,N_4731);
and U5241 (N_5241,N_4861,N_4399);
or U5242 (N_5242,N_4617,N_4361);
nor U5243 (N_5243,N_4580,N_4469);
and U5244 (N_5244,N_4733,N_4770);
nand U5245 (N_5245,N_4391,N_4457);
and U5246 (N_5246,N_4674,N_4547);
or U5247 (N_5247,N_4173,N_4789);
nand U5248 (N_5248,N_4836,N_4234);
nor U5249 (N_5249,N_4841,N_4142);
nor U5250 (N_5250,N_4903,N_4873);
or U5251 (N_5251,N_4059,N_4124);
nor U5252 (N_5252,N_4507,N_4433);
xor U5253 (N_5253,N_4594,N_4284);
nand U5254 (N_5254,N_4508,N_4700);
or U5255 (N_5255,N_4307,N_4476);
and U5256 (N_5256,N_4083,N_4151);
or U5257 (N_5257,N_4080,N_4351);
or U5258 (N_5258,N_4048,N_4708);
or U5259 (N_5259,N_4212,N_4544);
or U5260 (N_5260,N_4528,N_4427);
nor U5261 (N_5261,N_4801,N_4918);
nand U5262 (N_5262,N_4910,N_4270);
nand U5263 (N_5263,N_4389,N_4699);
and U5264 (N_5264,N_4686,N_4765);
nor U5265 (N_5265,N_4623,N_4817);
or U5266 (N_5266,N_4350,N_4310);
xnor U5267 (N_5267,N_4961,N_4747);
nor U5268 (N_5268,N_4702,N_4929);
or U5269 (N_5269,N_4039,N_4249);
and U5270 (N_5270,N_4220,N_4941);
or U5271 (N_5271,N_4865,N_4297);
nand U5272 (N_5272,N_4505,N_4047);
nor U5273 (N_5273,N_4093,N_4204);
nand U5274 (N_5274,N_4763,N_4868);
or U5275 (N_5275,N_4179,N_4466);
xnor U5276 (N_5276,N_4267,N_4325);
nor U5277 (N_5277,N_4368,N_4286);
or U5278 (N_5278,N_4206,N_4484);
nor U5279 (N_5279,N_4698,N_4821);
nor U5280 (N_5280,N_4527,N_4336);
nor U5281 (N_5281,N_4015,N_4703);
nor U5282 (N_5282,N_4027,N_4863);
and U5283 (N_5283,N_4413,N_4488);
xor U5284 (N_5284,N_4164,N_4844);
or U5285 (N_5285,N_4881,N_4646);
xnor U5286 (N_5286,N_4070,N_4474);
or U5287 (N_5287,N_4766,N_4175);
or U5288 (N_5288,N_4023,N_4795);
nand U5289 (N_5289,N_4054,N_4435);
or U5290 (N_5290,N_4622,N_4620);
and U5291 (N_5291,N_4494,N_4920);
nor U5292 (N_5292,N_4636,N_4450);
and U5293 (N_5293,N_4833,N_4605);
nand U5294 (N_5294,N_4890,N_4921);
nand U5295 (N_5295,N_4144,N_4026);
nand U5296 (N_5296,N_4331,N_4867);
xor U5297 (N_5297,N_4988,N_4040);
nand U5298 (N_5298,N_4106,N_4214);
nor U5299 (N_5299,N_4159,N_4383);
nor U5300 (N_5300,N_4559,N_4885);
nor U5301 (N_5301,N_4166,N_4784);
and U5302 (N_5302,N_4656,N_4509);
nand U5303 (N_5303,N_4589,N_4255);
nand U5304 (N_5304,N_4967,N_4959);
or U5305 (N_5305,N_4538,N_4471);
and U5306 (N_5306,N_4830,N_4216);
or U5307 (N_5307,N_4180,N_4892);
or U5308 (N_5308,N_4372,N_4965);
and U5309 (N_5309,N_4935,N_4540);
or U5310 (N_5310,N_4963,N_4917);
nand U5311 (N_5311,N_4905,N_4257);
nand U5312 (N_5312,N_4339,N_4870);
nor U5313 (N_5313,N_4324,N_4994);
nor U5314 (N_5314,N_4360,N_4446);
nand U5315 (N_5315,N_4487,N_4262);
and U5316 (N_5316,N_4057,N_4525);
xor U5317 (N_5317,N_4260,N_4648);
and U5318 (N_5318,N_4923,N_4441);
nand U5319 (N_5319,N_4805,N_4121);
or U5320 (N_5320,N_4240,N_4802);
nand U5321 (N_5321,N_4241,N_4628);
nand U5322 (N_5322,N_4659,N_4084);
nand U5323 (N_5323,N_4377,N_4539);
or U5324 (N_5324,N_4621,N_4690);
nor U5325 (N_5325,N_4985,N_4053);
or U5326 (N_5326,N_4287,N_4277);
nor U5327 (N_5327,N_4335,N_4823);
xor U5328 (N_5328,N_4366,N_4060);
nand U5329 (N_5329,N_4276,N_4843);
nand U5330 (N_5330,N_4148,N_4024);
nand U5331 (N_5331,N_4342,N_4598);
or U5332 (N_5332,N_4479,N_4811);
and U5333 (N_5333,N_4757,N_4127);
xnor U5334 (N_5334,N_4530,N_4717);
nand U5335 (N_5335,N_4679,N_4879);
nor U5336 (N_5336,N_4644,N_4300);
and U5337 (N_5337,N_4315,N_4827);
or U5338 (N_5338,N_4796,N_4657);
nor U5339 (N_5339,N_4613,N_4718);
nor U5340 (N_5340,N_4356,N_4281);
or U5341 (N_5341,N_4883,N_4775);
xor U5342 (N_5342,N_4774,N_4152);
and U5343 (N_5343,N_4546,N_4898);
and U5344 (N_5344,N_4393,N_4571);
nor U5345 (N_5345,N_4455,N_4394);
and U5346 (N_5346,N_4664,N_4842);
xor U5347 (N_5347,N_4115,N_4533);
and U5348 (N_5348,N_4291,N_4076);
nor U5349 (N_5349,N_4838,N_4806);
nor U5350 (N_5350,N_4301,N_4871);
nand U5351 (N_5351,N_4506,N_4079);
nand U5352 (N_5352,N_4095,N_4163);
and U5353 (N_5353,N_4602,N_4447);
nand U5354 (N_5354,N_4730,N_4872);
xnor U5355 (N_5355,N_4535,N_4641);
nor U5356 (N_5356,N_4964,N_4736);
and U5357 (N_5357,N_4518,N_4799);
or U5358 (N_5358,N_4557,N_4181);
nand U5359 (N_5359,N_4114,N_4581);
nand U5360 (N_5360,N_4991,N_4478);
nor U5361 (N_5361,N_4082,N_4911);
nor U5362 (N_5362,N_4835,N_4949);
nor U5363 (N_5363,N_4437,N_4135);
or U5364 (N_5364,N_4523,N_4174);
or U5365 (N_5365,N_4345,N_4104);
and U5366 (N_5366,N_4647,N_4950);
xnor U5367 (N_5367,N_4616,N_4993);
nand U5368 (N_5368,N_4312,N_4790);
xnor U5369 (N_5369,N_4263,N_4651);
xnor U5370 (N_5370,N_4565,N_4266);
or U5371 (N_5371,N_4182,N_4761);
and U5372 (N_5372,N_4379,N_4314);
xor U5373 (N_5373,N_4701,N_4137);
nand U5374 (N_5374,N_4552,N_4614);
nand U5375 (N_5375,N_4517,N_4572);
nor U5376 (N_5376,N_4541,N_4021);
or U5377 (N_5377,N_4463,N_4691);
nand U5378 (N_5378,N_4969,N_4495);
or U5379 (N_5379,N_4100,N_4723);
xor U5380 (N_5380,N_4200,N_4477);
nand U5381 (N_5381,N_4178,N_4327);
and U5382 (N_5382,N_4992,N_4235);
xor U5383 (N_5383,N_4560,N_4033);
xor U5384 (N_5384,N_4493,N_4107);
or U5385 (N_5385,N_4098,N_4548);
nand U5386 (N_5386,N_4758,N_4247);
xor U5387 (N_5387,N_4551,N_4722);
nor U5388 (N_5388,N_4554,N_4516);
xnor U5389 (N_5389,N_4111,N_4697);
nor U5390 (N_5390,N_4302,N_4460);
and U5391 (N_5391,N_4490,N_4122);
and U5392 (N_5392,N_4207,N_4543);
xnor U5393 (N_5393,N_4465,N_4755);
xnor U5394 (N_5394,N_4424,N_4064);
nand U5395 (N_5395,N_4952,N_4618);
or U5396 (N_5396,N_4459,N_4787);
and U5397 (N_5397,N_4238,N_4566);
xnor U5398 (N_5398,N_4323,N_4309);
xnor U5399 (N_5399,N_4019,N_4051);
xor U5400 (N_5400,N_4468,N_4997);
nand U5401 (N_5401,N_4358,N_4852);
or U5402 (N_5402,N_4742,N_4599);
nand U5403 (N_5403,N_4120,N_4452);
nand U5404 (N_5404,N_4930,N_4667);
xnor U5405 (N_5405,N_4201,N_4357);
nor U5406 (N_5406,N_4634,N_4009);
and U5407 (N_5407,N_4782,N_4073);
nor U5408 (N_5408,N_4856,N_4607);
and U5409 (N_5409,N_4960,N_4860);
nor U5410 (N_5410,N_4072,N_4980);
nand U5411 (N_5411,N_4052,N_4316);
or U5412 (N_5412,N_4583,N_4233);
nand U5413 (N_5413,N_4128,N_4188);
or U5414 (N_5414,N_4102,N_4017);
and U5415 (N_5415,N_4133,N_4655);
and U5416 (N_5416,N_4251,N_4261);
nand U5417 (N_5417,N_4388,N_4851);
nand U5418 (N_5418,N_4977,N_4362);
nand U5419 (N_5419,N_4411,N_4694);
or U5420 (N_5420,N_4829,N_4209);
nand U5421 (N_5421,N_4946,N_4748);
nor U5422 (N_5422,N_4298,N_4062);
nand U5423 (N_5423,N_4649,N_4066);
nand U5424 (N_5424,N_4587,N_4909);
nor U5425 (N_5425,N_4608,N_4579);
and U5426 (N_5426,N_4231,N_4944);
and U5427 (N_5427,N_4807,N_4526);
nand U5428 (N_5428,N_4954,N_4570);
and U5429 (N_5429,N_4123,N_4467);
xnor U5430 (N_5430,N_4392,N_4780);
and U5431 (N_5431,N_4042,N_4576);
or U5432 (N_5432,N_4631,N_4269);
nand U5433 (N_5433,N_4953,N_4063);
and U5434 (N_5434,N_4293,N_4715);
and U5435 (N_5435,N_4041,N_4464);
or U5436 (N_5436,N_4750,N_4087);
nand U5437 (N_5437,N_4434,N_4958);
nand U5438 (N_5438,N_4732,N_4036);
and U5439 (N_5439,N_4498,N_4422);
nand U5440 (N_5440,N_4633,N_4322);
or U5441 (N_5441,N_4237,N_4739);
or U5442 (N_5442,N_4194,N_4573);
and U5443 (N_5443,N_4658,N_4606);
nor U5444 (N_5444,N_4532,N_4012);
and U5445 (N_5445,N_4436,N_4899);
or U5446 (N_5446,N_4364,N_4492);
and U5447 (N_5447,N_4011,N_4680);
nor U5448 (N_5448,N_4456,N_4169);
nor U5449 (N_5449,N_4945,N_4273);
or U5450 (N_5450,N_4914,N_4592);
or U5451 (N_5451,N_4134,N_4783);
nand U5452 (N_5452,N_4767,N_4831);
and U5453 (N_5453,N_4706,N_4116);
nor U5454 (N_5454,N_4193,N_4922);
xor U5455 (N_5455,N_4157,N_4475);
and U5456 (N_5456,N_4275,N_4895);
or U5457 (N_5457,N_4837,N_4887);
or U5458 (N_5458,N_4000,N_4578);
xnor U5459 (N_5459,N_4650,N_4258);
nor U5460 (N_5460,N_4596,N_4777);
xor U5461 (N_5461,N_4891,N_4486);
nand U5462 (N_5462,N_4760,N_4798);
nor U5463 (N_5463,N_4824,N_4901);
and U5464 (N_5464,N_4849,N_4226);
nand U5465 (N_5465,N_4791,N_4119);
nand U5466 (N_5466,N_4367,N_4926);
nor U5467 (N_5467,N_4254,N_4185);
nor U5468 (N_5468,N_4359,N_4955);
nor U5469 (N_5469,N_4145,N_4925);
nand U5470 (N_5470,N_4482,N_4147);
nor U5471 (N_5471,N_4125,N_4529);
or U5472 (N_5472,N_4531,N_4390);
nor U5473 (N_5473,N_4222,N_4998);
and U5474 (N_5474,N_4721,N_4006);
or U5475 (N_5475,N_4793,N_4975);
or U5476 (N_5476,N_4728,N_4497);
nor U5477 (N_5477,N_4140,N_4549);
nand U5478 (N_5478,N_4228,N_4328);
or U5479 (N_5479,N_4462,N_4428);
or U5480 (N_5480,N_4252,N_4223);
nand U5481 (N_5481,N_4034,N_4974);
and U5482 (N_5482,N_4738,N_4046);
nand U5483 (N_5483,N_4110,N_4445);
nor U5484 (N_5484,N_4688,N_4198);
nor U5485 (N_5485,N_4915,N_4353);
nand U5486 (N_5486,N_4672,N_4385);
or U5487 (N_5487,N_4785,N_4692);
nand U5488 (N_5488,N_4221,N_4278);
or U5489 (N_5489,N_4826,N_4229);
xnor U5490 (N_5490,N_4567,N_4161);
or U5491 (N_5491,N_4030,N_4097);
and U5492 (N_5492,N_4349,N_4232);
nand U5493 (N_5493,N_4319,N_4735);
or U5494 (N_5494,N_4248,N_4859);
nor U5495 (N_5495,N_4160,N_4866);
and U5496 (N_5496,N_4375,N_4138);
nand U5497 (N_5497,N_4972,N_4192);
and U5498 (N_5498,N_4670,N_4224);
nand U5499 (N_5499,N_4203,N_4545);
xnor U5500 (N_5500,N_4972,N_4969);
nor U5501 (N_5501,N_4426,N_4655);
and U5502 (N_5502,N_4070,N_4626);
nor U5503 (N_5503,N_4174,N_4734);
or U5504 (N_5504,N_4595,N_4797);
xor U5505 (N_5505,N_4485,N_4363);
and U5506 (N_5506,N_4441,N_4328);
nand U5507 (N_5507,N_4607,N_4314);
nand U5508 (N_5508,N_4490,N_4258);
and U5509 (N_5509,N_4345,N_4644);
and U5510 (N_5510,N_4354,N_4986);
or U5511 (N_5511,N_4132,N_4683);
and U5512 (N_5512,N_4097,N_4624);
nand U5513 (N_5513,N_4658,N_4925);
xor U5514 (N_5514,N_4337,N_4314);
nor U5515 (N_5515,N_4773,N_4832);
nand U5516 (N_5516,N_4592,N_4025);
and U5517 (N_5517,N_4385,N_4309);
nand U5518 (N_5518,N_4018,N_4698);
nor U5519 (N_5519,N_4318,N_4811);
nor U5520 (N_5520,N_4529,N_4918);
or U5521 (N_5521,N_4745,N_4438);
nand U5522 (N_5522,N_4398,N_4492);
and U5523 (N_5523,N_4878,N_4853);
and U5524 (N_5524,N_4354,N_4238);
nand U5525 (N_5525,N_4838,N_4581);
nor U5526 (N_5526,N_4322,N_4612);
nor U5527 (N_5527,N_4273,N_4483);
xnor U5528 (N_5528,N_4420,N_4641);
nand U5529 (N_5529,N_4459,N_4194);
nand U5530 (N_5530,N_4569,N_4898);
or U5531 (N_5531,N_4492,N_4607);
nor U5532 (N_5532,N_4460,N_4619);
nand U5533 (N_5533,N_4655,N_4367);
xnor U5534 (N_5534,N_4434,N_4932);
and U5535 (N_5535,N_4951,N_4141);
and U5536 (N_5536,N_4247,N_4376);
and U5537 (N_5537,N_4931,N_4817);
or U5538 (N_5538,N_4185,N_4204);
and U5539 (N_5539,N_4137,N_4187);
nand U5540 (N_5540,N_4486,N_4274);
and U5541 (N_5541,N_4366,N_4956);
nand U5542 (N_5542,N_4815,N_4869);
nand U5543 (N_5543,N_4965,N_4968);
or U5544 (N_5544,N_4671,N_4485);
or U5545 (N_5545,N_4709,N_4116);
and U5546 (N_5546,N_4661,N_4383);
nor U5547 (N_5547,N_4221,N_4273);
nand U5548 (N_5548,N_4521,N_4139);
nand U5549 (N_5549,N_4686,N_4327);
and U5550 (N_5550,N_4819,N_4370);
nor U5551 (N_5551,N_4145,N_4029);
xor U5552 (N_5552,N_4538,N_4411);
nand U5553 (N_5553,N_4789,N_4690);
nand U5554 (N_5554,N_4019,N_4185);
xnor U5555 (N_5555,N_4773,N_4637);
nand U5556 (N_5556,N_4023,N_4009);
or U5557 (N_5557,N_4867,N_4387);
nor U5558 (N_5558,N_4580,N_4398);
nor U5559 (N_5559,N_4651,N_4762);
and U5560 (N_5560,N_4261,N_4079);
nor U5561 (N_5561,N_4073,N_4876);
and U5562 (N_5562,N_4274,N_4721);
or U5563 (N_5563,N_4410,N_4824);
and U5564 (N_5564,N_4292,N_4907);
nand U5565 (N_5565,N_4634,N_4409);
nor U5566 (N_5566,N_4444,N_4616);
and U5567 (N_5567,N_4553,N_4433);
and U5568 (N_5568,N_4501,N_4926);
nand U5569 (N_5569,N_4668,N_4288);
and U5570 (N_5570,N_4041,N_4656);
and U5571 (N_5571,N_4224,N_4380);
nor U5572 (N_5572,N_4495,N_4185);
xor U5573 (N_5573,N_4117,N_4897);
nand U5574 (N_5574,N_4222,N_4750);
or U5575 (N_5575,N_4533,N_4248);
nand U5576 (N_5576,N_4813,N_4844);
or U5577 (N_5577,N_4532,N_4955);
or U5578 (N_5578,N_4625,N_4632);
nand U5579 (N_5579,N_4774,N_4494);
nor U5580 (N_5580,N_4472,N_4274);
and U5581 (N_5581,N_4270,N_4034);
and U5582 (N_5582,N_4582,N_4157);
and U5583 (N_5583,N_4117,N_4503);
nor U5584 (N_5584,N_4905,N_4321);
xor U5585 (N_5585,N_4726,N_4096);
and U5586 (N_5586,N_4412,N_4826);
nor U5587 (N_5587,N_4855,N_4747);
xor U5588 (N_5588,N_4438,N_4280);
or U5589 (N_5589,N_4909,N_4881);
nor U5590 (N_5590,N_4233,N_4095);
nor U5591 (N_5591,N_4495,N_4765);
nand U5592 (N_5592,N_4120,N_4783);
xnor U5593 (N_5593,N_4257,N_4627);
or U5594 (N_5594,N_4693,N_4787);
and U5595 (N_5595,N_4251,N_4937);
nor U5596 (N_5596,N_4595,N_4209);
nor U5597 (N_5597,N_4126,N_4324);
nand U5598 (N_5598,N_4562,N_4474);
xnor U5599 (N_5599,N_4226,N_4339);
xor U5600 (N_5600,N_4204,N_4535);
nand U5601 (N_5601,N_4441,N_4928);
and U5602 (N_5602,N_4492,N_4283);
xnor U5603 (N_5603,N_4406,N_4174);
xnor U5604 (N_5604,N_4220,N_4833);
and U5605 (N_5605,N_4662,N_4298);
nand U5606 (N_5606,N_4628,N_4697);
and U5607 (N_5607,N_4794,N_4582);
or U5608 (N_5608,N_4077,N_4102);
or U5609 (N_5609,N_4884,N_4504);
or U5610 (N_5610,N_4202,N_4536);
nor U5611 (N_5611,N_4567,N_4581);
nor U5612 (N_5612,N_4789,N_4648);
nor U5613 (N_5613,N_4080,N_4145);
nor U5614 (N_5614,N_4916,N_4631);
or U5615 (N_5615,N_4642,N_4896);
or U5616 (N_5616,N_4543,N_4579);
xor U5617 (N_5617,N_4678,N_4006);
and U5618 (N_5618,N_4230,N_4910);
nand U5619 (N_5619,N_4270,N_4391);
nand U5620 (N_5620,N_4800,N_4602);
or U5621 (N_5621,N_4535,N_4532);
nand U5622 (N_5622,N_4416,N_4847);
nor U5623 (N_5623,N_4785,N_4089);
nor U5624 (N_5624,N_4637,N_4149);
or U5625 (N_5625,N_4562,N_4332);
or U5626 (N_5626,N_4297,N_4856);
xor U5627 (N_5627,N_4210,N_4817);
or U5628 (N_5628,N_4090,N_4671);
nor U5629 (N_5629,N_4716,N_4372);
nor U5630 (N_5630,N_4111,N_4544);
nand U5631 (N_5631,N_4854,N_4069);
nor U5632 (N_5632,N_4487,N_4114);
nand U5633 (N_5633,N_4457,N_4003);
or U5634 (N_5634,N_4201,N_4528);
or U5635 (N_5635,N_4093,N_4580);
nand U5636 (N_5636,N_4706,N_4574);
nand U5637 (N_5637,N_4135,N_4865);
xnor U5638 (N_5638,N_4606,N_4729);
and U5639 (N_5639,N_4266,N_4734);
nor U5640 (N_5640,N_4573,N_4867);
or U5641 (N_5641,N_4203,N_4968);
nand U5642 (N_5642,N_4012,N_4937);
and U5643 (N_5643,N_4204,N_4887);
nand U5644 (N_5644,N_4461,N_4228);
or U5645 (N_5645,N_4416,N_4913);
or U5646 (N_5646,N_4857,N_4965);
nand U5647 (N_5647,N_4602,N_4270);
nand U5648 (N_5648,N_4103,N_4496);
and U5649 (N_5649,N_4555,N_4710);
xor U5650 (N_5650,N_4090,N_4160);
nor U5651 (N_5651,N_4284,N_4632);
nor U5652 (N_5652,N_4556,N_4246);
and U5653 (N_5653,N_4758,N_4252);
and U5654 (N_5654,N_4622,N_4979);
or U5655 (N_5655,N_4315,N_4481);
xor U5656 (N_5656,N_4712,N_4559);
nand U5657 (N_5657,N_4523,N_4443);
nor U5658 (N_5658,N_4362,N_4150);
or U5659 (N_5659,N_4258,N_4158);
xnor U5660 (N_5660,N_4680,N_4424);
and U5661 (N_5661,N_4287,N_4197);
nor U5662 (N_5662,N_4097,N_4806);
or U5663 (N_5663,N_4086,N_4688);
or U5664 (N_5664,N_4009,N_4336);
nand U5665 (N_5665,N_4434,N_4507);
xor U5666 (N_5666,N_4883,N_4489);
or U5667 (N_5667,N_4452,N_4617);
or U5668 (N_5668,N_4287,N_4525);
and U5669 (N_5669,N_4571,N_4179);
nand U5670 (N_5670,N_4731,N_4921);
xor U5671 (N_5671,N_4923,N_4798);
nor U5672 (N_5672,N_4923,N_4368);
nand U5673 (N_5673,N_4850,N_4670);
nor U5674 (N_5674,N_4340,N_4362);
and U5675 (N_5675,N_4058,N_4380);
and U5676 (N_5676,N_4005,N_4772);
and U5677 (N_5677,N_4053,N_4207);
nor U5678 (N_5678,N_4962,N_4118);
nor U5679 (N_5679,N_4384,N_4735);
and U5680 (N_5680,N_4522,N_4755);
nand U5681 (N_5681,N_4585,N_4632);
nor U5682 (N_5682,N_4347,N_4511);
xnor U5683 (N_5683,N_4626,N_4600);
nand U5684 (N_5684,N_4516,N_4607);
and U5685 (N_5685,N_4189,N_4233);
nand U5686 (N_5686,N_4799,N_4997);
or U5687 (N_5687,N_4239,N_4521);
or U5688 (N_5688,N_4234,N_4823);
and U5689 (N_5689,N_4752,N_4853);
or U5690 (N_5690,N_4506,N_4697);
nand U5691 (N_5691,N_4855,N_4573);
or U5692 (N_5692,N_4822,N_4509);
or U5693 (N_5693,N_4955,N_4856);
and U5694 (N_5694,N_4636,N_4979);
or U5695 (N_5695,N_4836,N_4497);
nor U5696 (N_5696,N_4050,N_4615);
nand U5697 (N_5697,N_4057,N_4329);
nor U5698 (N_5698,N_4371,N_4318);
and U5699 (N_5699,N_4504,N_4862);
xnor U5700 (N_5700,N_4015,N_4199);
nor U5701 (N_5701,N_4734,N_4323);
nor U5702 (N_5702,N_4753,N_4371);
or U5703 (N_5703,N_4342,N_4907);
nor U5704 (N_5704,N_4351,N_4232);
or U5705 (N_5705,N_4644,N_4332);
nand U5706 (N_5706,N_4286,N_4590);
and U5707 (N_5707,N_4282,N_4379);
nand U5708 (N_5708,N_4865,N_4985);
or U5709 (N_5709,N_4200,N_4849);
or U5710 (N_5710,N_4243,N_4710);
or U5711 (N_5711,N_4432,N_4555);
and U5712 (N_5712,N_4156,N_4572);
and U5713 (N_5713,N_4653,N_4262);
or U5714 (N_5714,N_4221,N_4077);
nor U5715 (N_5715,N_4291,N_4571);
and U5716 (N_5716,N_4920,N_4705);
and U5717 (N_5717,N_4233,N_4170);
and U5718 (N_5718,N_4195,N_4047);
or U5719 (N_5719,N_4950,N_4121);
and U5720 (N_5720,N_4005,N_4538);
nor U5721 (N_5721,N_4520,N_4621);
nor U5722 (N_5722,N_4812,N_4890);
xor U5723 (N_5723,N_4401,N_4486);
nor U5724 (N_5724,N_4554,N_4144);
or U5725 (N_5725,N_4067,N_4610);
and U5726 (N_5726,N_4715,N_4927);
nor U5727 (N_5727,N_4448,N_4489);
and U5728 (N_5728,N_4683,N_4043);
nand U5729 (N_5729,N_4901,N_4175);
or U5730 (N_5730,N_4076,N_4736);
xnor U5731 (N_5731,N_4703,N_4205);
or U5732 (N_5732,N_4882,N_4064);
and U5733 (N_5733,N_4070,N_4900);
nor U5734 (N_5734,N_4569,N_4883);
or U5735 (N_5735,N_4724,N_4110);
and U5736 (N_5736,N_4848,N_4403);
and U5737 (N_5737,N_4846,N_4370);
or U5738 (N_5738,N_4557,N_4133);
nor U5739 (N_5739,N_4811,N_4480);
nor U5740 (N_5740,N_4907,N_4429);
and U5741 (N_5741,N_4876,N_4335);
nand U5742 (N_5742,N_4108,N_4596);
nor U5743 (N_5743,N_4552,N_4191);
or U5744 (N_5744,N_4682,N_4628);
or U5745 (N_5745,N_4273,N_4774);
and U5746 (N_5746,N_4923,N_4533);
or U5747 (N_5747,N_4165,N_4116);
nor U5748 (N_5748,N_4887,N_4762);
nor U5749 (N_5749,N_4937,N_4759);
and U5750 (N_5750,N_4142,N_4553);
nand U5751 (N_5751,N_4734,N_4946);
and U5752 (N_5752,N_4769,N_4190);
and U5753 (N_5753,N_4258,N_4576);
nor U5754 (N_5754,N_4057,N_4736);
nand U5755 (N_5755,N_4245,N_4249);
or U5756 (N_5756,N_4371,N_4857);
or U5757 (N_5757,N_4536,N_4656);
or U5758 (N_5758,N_4055,N_4537);
and U5759 (N_5759,N_4017,N_4323);
nand U5760 (N_5760,N_4067,N_4867);
and U5761 (N_5761,N_4588,N_4445);
nand U5762 (N_5762,N_4281,N_4353);
and U5763 (N_5763,N_4201,N_4435);
nand U5764 (N_5764,N_4844,N_4045);
nand U5765 (N_5765,N_4371,N_4487);
xor U5766 (N_5766,N_4683,N_4362);
or U5767 (N_5767,N_4772,N_4394);
nand U5768 (N_5768,N_4822,N_4422);
nor U5769 (N_5769,N_4673,N_4234);
nand U5770 (N_5770,N_4773,N_4442);
nand U5771 (N_5771,N_4446,N_4795);
xnor U5772 (N_5772,N_4192,N_4199);
and U5773 (N_5773,N_4370,N_4790);
xor U5774 (N_5774,N_4836,N_4511);
nand U5775 (N_5775,N_4516,N_4712);
nand U5776 (N_5776,N_4892,N_4423);
and U5777 (N_5777,N_4138,N_4106);
or U5778 (N_5778,N_4338,N_4761);
or U5779 (N_5779,N_4255,N_4574);
and U5780 (N_5780,N_4856,N_4854);
or U5781 (N_5781,N_4920,N_4469);
or U5782 (N_5782,N_4376,N_4576);
and U5783 (N_5783,N_4494,N_4917);
nand U5784 (N_5784,N_4498,N_4014);
nor U5785 (N_5785,N_4428,N_4781);
or U5786 (N_5786,N_4646,N_4193);
nand U5787 (N_5787,N_4504,N_4879);
nand U5788 (N_5788,N_4859,N_4546);
nor U5789 (N_5789,N_4135,N_4460);
or U5790 (N_5790,N_4355,N_4498);
nor U5791 (N_5791,N_4138,N_4416);
nand U5792 (N_5792,N_4363,N_4781);
xor U5793 (N_5793,N_4182,N_4612);
or U5794 (N_5794,N_4654,N_4331);
and U5795 (N_5795,N_4575,N_4730);
nor U5796 (N_5796,N_4433,N_4534);
nor U5797 (N_5797,N_4905,N_4287);
or U5798 (N_5798,N_4245,N_4018);
nand U5799 (N_5799,N_4554,N_4125);
or U5800 (N_5800,N_4362,N_4133);
nand U5801 (N_5801,N_4282,N_4596);
nand U5802 (N_5802,N_4285,N_4241);
nand U5803 (N_5803,N_4260,N_4910);
nor U5804 (N_5804,N_4342,N_4030);
nor U5805 (N_5805,N_4608,N_4719);
nand U5806 (N_5806,N_4599,N_4286);
nand U5807 (N_5807,N_4692,N_4297);
nand U5808 (N_5808,N_4106,N_4600);
or U5809 (N_5809,N_4648,N_4502);
and U5810 (N_5810,N_4445,N_4726);
nor U5811 (N_5811,N_4410,N_4453);
or U5812 (N_5812,N_4802,N_4934);
or U5813 (N_5813,N_4502,N_4432);
nor U5814 (N_5814,N_4059,N_4735);
nand U5815 (N_5815,N_4653,N_4702);
and U5816 (N_5816,N_4644,N_4983);
xor U5817 (N_5817,N_4849,N_4671);
nand U5818 (N_5818,N_4246,N_4300);
xnor U5819 (N_5819,N_4009,N_4914);
or U5820 (N_5820,N_4398,N_4403);
nor U5821 (N_5821,N_4947,N_4400);
nor U5822 (N_5822,N_4178,N_4017);
nor U5823 (N_5823,N_4375,N_4603);
nor U5824 (N_5824,N_4631,N_4599);
nor U5825 (N_5825,N_4706,N_4989);
nor U5826 (N_5826,N_4706,N_4041);
and U5827 (N_5827,N_4572,N_4097);
nand U5828 (N_5828,N_4216,N_4904);
nand U5829 (N_5829,N_4892,N_4639);
and U5830 (N_5830,N_4816,N_4421);
nor U5831 (N_5831,N_4980,N_4221);
or U5832 (N_5832,N_4350,N_4807);
nand U5833 (N_5833,N_4831,N_4374);
nor U5834 (N_5834,N_4922,N_4077);
xnor U5835 (N_5835,N_4238,N_4458);
nor U5836 (N_5836,N_4581,N_4278);
nor U5837 (N_5837,N_4377,N_4069);
and U5838 (N_5838,N_4747,N_4452);
and U5839 (N_5839,N_4711,N_4709);
nand U5840 (N_5840,N_4621,N_4425);
nand U5841 (N_5841,N_4100,N_4383);
and U5842 (N_5842,N_4929,N_4971);
or U5843 (N_5843,N_4509,N_4680);
nor U5844 (N_5844,N_4528,N_4646);
nor U5845 (N_5845,N_4503,N_4313);
and U5846 (N_5846,N_4790,N_4230);
nor U5847 (N_5847,N_4310,N_4475);
nand U5848 (N_5848,N_4624,N_4633);
nor U5849 (N_5849,N_4287,N_4151);
xnor U5850 (N_5850,N_4249,N_4092);
nor U5851 (N_5851,N_4507,N_4537);
xnor U5852 (N_5852,N_4716,N_4594);
nand U5853 (N_5853,N_4226,N_4360);
nor U5854 (N_5854,N_4410,N_4484);
or U5855 (N_5855,N_4959,N_4277);
nand U5856 (N_5856,N_4097,N_4066);
or U5857 (N_5857,N_4570,N_4260);
or U5858 (N_5858,N_4964,N_4371);
or U5859 (N_5859,N_4107,N_4411);
or U5860 (N_5860,N_4871,N_4748);
or U5861 (N_5861,N_4730,N_4114);
nand U5862 (N_5862,N_4508,N_4155);
nor U5863 (N_5863,N_4646,N_4802);
nand U5864 (N_5864,N_4309,N_4391);
or U5865 (N_5865,N_4477,N_4314);
nand U5866 (N_5866,N_4349,N_4043);
nor U5867 (N_5867,N_4817,N_4102);
nand U5868 (N_5868,N_4190,N_4342);
and U5869 (N_5869,N_4761,N_4022);
or U5870 (N_5870,N_4672,N_4734);
xnor U5871 (N_5871,N_4931,N_4049);
or U5872 (N_5872,N_4278,N_4319);
nor U5873 (N_5873,N_4340,N_4826);
nand U5874 (N_5874,N_4304,N_4768);
nor U5875 (N_5875,N_4535,N_4433);
and U5876 (N_5876,N_4646,N_4056);
nand U5877 (N_5877,N_4099,N_4195);
and U5878 (N_5878,N_4655,N_4927);
and U5879 (N_5879,N_4668,N_4875);
and U5880 (N_5880,N_4090,N_4822);
and U5881 (N_5881,N_4510,N_4013);
or U5882 (N_5882,N_4396,N_4310);
or U5883 (N_5883,N_4202,N_4904);
or U5884 (N_5884,N_4204,N_4301);
and U5885 (N_5885,N_4456,N_4998);
nor U5886 (N_5886,N_4915,N_4820);
nor U5887 (N_5887,N_4373,N_4860);
nor U5888 (N_5888,N_4079,N_4309);
xnor U5889 (N_5889,N_4032,N_4705);
and U5890 (N_5890,N_4977,N_4983);
or U5891 (N_5891,N_4318,N_4914);
or U5892 (N_5892,N_4922,N_4664);
nor U5893 (N_5893,N_4577,N_4843);
xnor U5894 (N_5894,N_4274,N_4085);
or U5895 (N_5895,N_4830,N_4552);
nor U5896 (N_5896,N_4450,N_4433);
and U5897 (N_5897,N_4501,N_4251);
or U5898 (N_5898,N_4434,N_4005);
or U5899 (N_5899,N_4071,N_4686);
nand U5900 (N_5900,N_4013,N_4938);
and U5901 (N_5901,N_4751,N_4876);
and U5902 (N_5902,N_4920,N_4603);
and U5903 (N_5903,N_4686,N_4774);
and U5904 (N_5904,N_4456,N_4691);
nor U5905 (N_5905,N_4404,N_4655);
and U5906 (N_5906,N_4910,N_4949);
nor U5907 (N_5907,N_4917,N_4519);
and U5908 (N_5908,N_4561,N_4192);
nand U5909 (N_5909,N_4313,N_4093);
nor U5910 (N_5910,N_4598,N_4023);
and U5911 (N_5911,N_4068,N_4737);
and U5912 (N_5912,N_4691,N_4484);
nor U5913 (N_5913,N_4433,N_4333);
and U5914 (N_5914,N_4843,N_4354);
or U5915 (N_5915,N_4220,N_4099);
nor U5916 (N_5916,N_4050,N_4336);
or U5917 (N_5917,N_4910,N_4866);
and U5918 (N_5918,N_4923,N_4231);
or U5919 (N_5919,N_4624,N_4963);
and U5920 (N_5920,N_4391,N_4315);
xnor U5921 (N_5921,N_4449,N_4308);
nor U5922 (N_5922,N_4982,N_4981);
nor U5923 (N_5923,N_4071,N_4868);
nand U5924 (N_5924,N_4176,N_4288);
or U5925 (N_5925,N_4439,N_4317);
nand U5926 (N_5926,N_4215,N_4170);
nor U5927 (N_5927,N_4558,N_4282);
nand U5928 (N_5928,N_4632,N_4438);
and U5929 (N_5929,N_4236,N_4148);
and U5930 (N_5930,N_4776,N_4447);
or U5931 (N_5931,N_4768,N_4886);
nor U5932 (N_5932,N_4630,N_4068);
and U5933 (N_5933,N_4837,N_4067);
and U5934 (N_5934,N_4586,N_4486);
or U5935 (N_5935,N_4789,N_4546);
and U5936 (N_5936,N_4643,N_4569);
nor U5937 (N_5937,N_4242,N_4024);
or U5938 (N_5938,N_4894,N_4793);
nand U5939 (N_5939,N_4933,N_4930);
and U5940 (N_5940,N_4446,N_4980);
nor U5941 (N_5941,N_4038,N_4846);
and U5942 (N_5942,N_4694,N_4756);
nand U5943 (N_5943,N_4043,N_4575);
nor U5944 (N_5944,N_4953,N_4826);
and U5945 (N_5945,N_4319,N_4422);
or U5946 (N_5946,N_4187,N_4875);
or U5947 (N_5947,N_4130,N_4279);
nand U5948 (N_5948,N_4215,N_4192);
and U5949 (N_5949,N_4556,N_4776);
nand U5950 (N_5950,N_4478,N_4538);
or U5951 (N_5951,N_4699,N_4652);
and U5952 (N_5952,N_4478,N_4838);
or U5953 (N_5953,N_4163,N_4667);
nor U5954 (N_5954,N_4994,N_4347);
nand U5955 (N_5955,N_4300,N_4764);
or U5956 (N_5956,N_4250,N_4115);
or U5957 (N_5957,N_4315,N_4352);
nor U5958 (N_5958,N_4631,N_4193);
nor U5959 (N_5959,N_4956,N_4204);
nor U5960 (N_5960,N_4607,N_4041);
and U5961 (N_5961,N_4673,N_4897);
nand U5962 (N_5962,N_4815,N_4089);
or U5963 (N_5963,N_4407,N_4647);
or U5964 (N_5964,N_4356,N_4308);
nand U5965 (N_5965,N_4376,N_4996);
nand U5966 (N_5966,N_4723,N_4486);
nand U5967 (N_5967,N_4209,N_4497);
nor U5968 (N_5968,N_4001,N_4205);
and U5969 (N_5969,N_4369,N_4359);
or U5970 (N_5970,N_4824,N_4636);
nand U5971 (N_5971,N_4913,N_4541);
nand U5972 (N_5972,N_4659,N_4579);
and U5973 (N_5973,N_4686,N_4201);
xnor U5974 (N_5974,N_4343,N_4946);
nor U5975 (N_5975,N_4431,N_4346);
nor U5976 (N_5976,N_4929,N_4810);
nand U5977 (N_5977,N_4316,N_4152);
nor U5978 (N_5978,N_4440,N_4498);
nor U5979 (N_5979,N_4258,N_4595);
nand U5980 (N_5980,N_4345,N_4940);
nand U5981 (N_5981,N_4391,N_4568);
xnor U5982 (N_5982,N_4079,N_4662);
and U5983 (N_5983,N_4444,N_4607);
or U5984 (N_5984,N_4022,N_4741);
nor U5985 (N_5985,N_4401,N_4806);
and U5986 (N_5986,N_4498,N_4562);
nor U5987 (N_5987,N_4420,N_4980);
or U5988 (N_5988,N_4138,N_4449);
xor U5989 (N_5989,N_4228,N_4941);
or U5990 (N_5990,N_4592,N_4651);
and U5991 (N_5991,N_4066,N_4756);
nand U5992 (N_5992,N_4712,N_4594);
xnor U5993 (N_5993,N_4868,N_4773);
and U5994 (N_5994,N_4871,N_4521);
and U5995 (N_5995,N_4970,N_4968);
or U5996 (N_5996,N_4779,N_4560);
nand U5997 (N_5997,N_4797,N_4297);
nand U5998 (N_5998,N_4735,N_4518);
nand U5999 (N_5999,N_4497,N_4927);
and U6000 (N_6000,N_5085,N_5956);
or U6001 (N_6001,N_5747,N_5122);
and U6002 (N_6002,N_5182,N_5276);
nand U6003 (N_6003,N_5681,N_5277);
or U6004 (N_6004,N_5469,N_5318);
or U6005 (N_6005,N_5661,N_5119);
and U6006 (N_6006,N_5636,N_5320);
nand U6007 (N_6007,N_5211,N_5598);
nor U6008 (N_6008,N_5768,N_5654);
or U6009 (N_6009,N_5214,N_5310);
nand U6010 (N_6010,N_5080,N_5256);
nand U6011 (N_6011,N_5857,N_5787);
nand U6012 (N_6012,N_5088,N_5039);
nand U6013 (N_6013,N_5795,N_5835);
nand U6014 (N_6014,N_5359,N_5018);
nor U6015 (N_6015,N_5626,N_5035);
xnor U6016 (N_6016,N_5806,N_5130);
xnor U6017 (N_6017,N_5943,N_5838);
nand U6018 (N_6018,N_5351,N_5413);
nand U6019 (N_6019,N_5764,N_5184);
xor U6020 (N_6020,N_5819,N_5341);
nand U6021 (N_6021,N_5307,N_5760);
or U6022 (N_6022,N_5763,N_5027);
nand U6023 (N_6023,N_5492,N_5890);
or U6024 (N_6024,N_5178,N_5345);
nand U6025 (N_6025,N_5172,N_5059);
and U6026 (N_6026,N_5308,N_5421);
and U6027 (N_6027,N_5632,N_5954);
nand U6028 (N_6028,N_5199,N_5190);
nor U6029 (N_6029,N_5232,N_5311);
or U6030 (N_6030,N_5804,N_5081);
nand U6031 (N_6031,N_5571,N_5121);
nand U6032 (N_6032,N_5669,N_5432);
or U6033 (N_6033,N_5519,N_5065);
nor U6034 (N_6034,N_5301,N_5040);
and U6035 (N_6035,N_5921,N_5614);
nand U6036 (N_6036,N_5961,N_5185);
and U6037 (N_6037,N_5937,N_5775);
and U6038 (N_6038,N_5319,N_5837);
nor U6039 (N_6039,N_5309,N_5832);
nand U6040 (N_6040,N_5297,N_5370);
and U6041 (N_6041,N_5471,N_5445);
and U6042 (N_6042,N_5493,N_5842);
or U6043 (N_6043,N_5322,N_5673);
or U6044 (N_6044,N_5602,N_5828);
or U6045 (N_6045,N_5132,N_5484);
and U6046 (N_6046,N_5267,N_5970);
xnor U6047 (N_6047,N_5019,N_5639);
or U6048 (N_6048,N_5540,N_5316);
and U6049 (N_6049,N_5758,N_5118);
nor U6050 (N_6050,N_5642,N_5062);
and U6051 (N_6051,N_5658,N_5176);
or U6052 (N_6052,N_5048,N_5706);
or U6053 (N_6053,N_5175,N_5079);
and U6054 (N_6054,N_5762,N_5227);
nand U6055 (N_6055,N_5955,N_5414);
and U6056 (N_6056,N_5449,N_5818);
or U6057 (N_6057,N_5913,N_5399);
nand U6058 (N_6058,N_5047,N_5982);
nand U6059 (N_6059,N_5503,N_5774);
nor U6060 (N_6060,N_5847,N_5367);
and U6061 (N_6061,N_5146,N_5126);
or U6062 (N_6062,N_5011,N_5587);
nor U6063 (N_6063,N_5247,N_5558);
and U6064 (N_6064,N_5567,N_5284);
and U6065 (N_6065,N_5701,N_5957);
nor U6066 (N_6066,N_5253,N_5254);
and U6067 (N_6067,N_5848,N_5083);
nand U6068 (N_6068,N_5691,N_5325);
nor U6069 (N_6069,N_5148,N_5724);
and U6070 (N_6070,N_5507,N_5700);
and U6071 (N_6071,N_5874,N_5565);
or U6072 (N_6072,N_5996,N_5672);
nand U6073 (N_6073,N_5482,N_5850);
xnor U6074 (N_6074,N_5332,N_5574);
and U6075 (N_6075,N_5456,N_5866);
nand U6076 (N_6076,N_5511,N_5902);
and U6077 (N_6077,N_5486,N_5530);
nand U6078 (N_6078,N_5221,N_5106);
nor U6079 (N_6079,N_5811,N_5055);
nor U6080 (N_6080,N_5293,N_5885);
xor U6081 (N_6081,N_5139,N_5689);
and U6082 (N_6082,N_5860,N_5645);
nor U6083 (N_6083,N_5749,N_5077);
nor U6084 (N_6084,N_5594,N_5167);
nor U6085 (N_6085,N_5057,N_5999);
and U6086 (N_6086,N_5873,N_5128);
xnor U6087 (N_6087,N_5069,N_5676);
and U6088 (N_6088,N_5726,N_5495);
xnor U6089 (N_6089,N_5329,N_5708);
or U6090 (N_6090,N_5222,N_5534);
or U6091 (N_6091,N_5515,N_5712);
nor U6092 (N_6092,N_5878,N_5422);
or U6093 (N_6093,N_5058,N_5340);
nor U6094 (N_6094,N_5289,N_5647);
or U6095 (N_6095,N_5285,N_5907);
nor U6096 (N_6096,N_5366,N_5997);
or U6097 (N_6097,N_5191,N_5305);
nand U6098 (N_6098,N_5922,N_5521);
nor U6099 (N_6099,N_5829,N_5382);
and U6100 (N_6100,N_5485,N_5513);
or U6101 (N_6101,N_5536,N_5737);
nand U6102 (N_6102,N_5667,N_5776);
xor U6103 (N_6103,N_5434,N_5797);
xor U6104 (N_6104,N_5010,N_5420);
nor U6105 (N_6105,N_5117,N_5459);
nand U6106 (N_6106,N_5028,N_5024);
nand U6107 (N_6107,N_5923,N_5753);
nor U6108 (N_6108,N_5555,N_5635);
and U6109 (N_6109,N_5827,N_5962);
xnor U6110 (N_6110,N_5692,N_5568);
nor U6111 (N_6111,N_5723,N_5824);
or U6112 (N_6112,N_5280,N_5431);
and U6113 (N_6113,N_5554,N_5110);
nand U6114 (N_6114,N_5801,N_5634);
nor U6115 (N_6115,N_5882,N_5008);
nand U6116 (N_6116,N_5089,N_5531);
and U6117 (N_6117,N_5444,N_5049);
or U6118 (N_6118,N_5389,N_5759);
nor U6119 (N_6119,N_5241,N_5385);
nand U6120 (N_6120,N_5064,N_5391);
and U6121 (N_6121,N_5446,N_5695);
xnor U6122 (N_6122,N_5727,N_5900);
or U6123 (N_6123,N_5985,N_5966);
and U6124 (N_6124,N_5685,N_5757);
and U6125 (N_6125,N_5538,N_5196);
xnor U6126 (N_6126,N_5076,N_5053);
and U6127 (N_6127,N_5153,N_5936);
nand U6128 (N_6128,N_5520,N_5663);
xor U6129 (N_6129,N_5638,N_5711);
xor U6130 (N_6130,N_5968,N_5816);
and U6131 (N_6131,N_5694,N_5911);
or U6132 (N_6132,N_5353,N_5440);
nand U6133 (N_6133,N_5977,N_5326);
nand U6134 (N_6134,N_5271,N_5561);
nor U6135 (N_6135,N_5780,N_5508);
and U6136 (N_6136,N_5983,N_5948);
nor U6137 (N_6137,N_5286,N_5138);
or U6138 (N_6138,N_5361,N_5651);
or U6139 (N_6139,N_5164,N_5916);
or U6140 (N_6140,N_5836,N_5075);
and U6141 (N_6141,N_5032,N_5670);
or U6142 (N_6142,N_5617,N_5107);
nor U6143 (N_6143,N_5496,N_5260);
or U6144 (N_6144,N_5250,N_5718);
nand U6145 (N_6145,N_5817,N_5887);
or U6146 (N_6146,N_5633,N_5452);
xor U6147 (N_6147,N_5406,N_5805);
nor U6148 (N_6148,N_5240,N_5037);
nor U6149 (N_6149,N_5335,N_5073);
xor U6150 (N_6150,N_5147,N_5810);
nor U6151 (N_6151,N_5901,N_5500);
nor U6152 (N_6152,N_5543,N_5579);
nor U6153 (N_6153,N_5171,N_5597);
nand U6154 (N_6154,N_5282,N_5671);
or U6155 (N_6155,N_5441,N_5821);
or U6156 (N_6156,N_5397,N_5514);
nand U6157 (N_6157,N_5109,N_5363);
nor U6158 (N_6158,N_5161,N_5417);
or U6159 (N_6159,N_5595,N_5721);
nor U6160 (N_6160,N_5551,N_5262);
nand U6161 (N_6161,N_5570,N_5732);
nor U6162 (N_6162,N_5845,N_5195);
xnor U6163 (N_6163,N_5330,N_5583);
or U6164 (N_6164,N_5858,N_5296);
xor U6165 (N_6165,N_5879,N_5814);
and U6166 (N_6166,N_5497,N_5272);
nor U6167 (N_6167,N_5269,N_5914);
nand U6168 (N_6168,N_5905,N_5853);
nor U6169 (N_6169,N_5662,N_5581);
xnor U6170 (N_6170,N_5499,N_5575);
or U6171 (N_6171,N_5294,N_5577);
nand U6172 (N_6172,N_5934,N_5168);
nor U6173 (N_6173,N_5462,N_5944);
nand U6174 (N_6174,N_5388,N_5210);
or U6175 (N_6175,N_5736,N_5355);
or U6176 (N_6176,N_5609,N_5984);
and U6177 (N_6177,N_5084,N_5742);
nand U6178 (N_6178,N_5186,N_5022);
or U6179 (N_6179,N_5830,N_5523);
or U6180 (N_6180,N_5105,N_5339);
nand U6181 (N_6181,N_5864,N_5349);
nand U6182 (N_6182,N_5321,N_5187);
nand U6183 (N_6183,N_5502,N_5722);
nor U6184 (N_6184,N_5012,N_5738);
nor U6185 (N_6185,N_5283,N_5061);
nor U6186 (N_6186,N_5549,N_5090);
nand U6187 (N_6187,N_5584,N_5665);
or U6188 (N_6188,N_5849,N_5745);
xnor U6189 (N_6189,N_5468,N_5933);
or U6190 (N_6190,N_5615,N_5133);
nand U6191 (N_6191,N_5798,N_5157);
or U6192 (N_6192,N_5398,N_5884);
and U6193 (N_6193,N_5401,N_5789);
nand U6194 (N_6194,N_5599,N_5149);
or U6195 (N_6195,N_5546,N_5931);
nand U6196 (N_6196,N_5051,N_5238);
or U6197 (N_6197,N_5627,N_5165);
nand U6198 (N_6198,N_5248,N_5003);
nand U6199 (N_6199,N_5160,N_5664);
nor U6200 (N_6200,N_5404,N_5266);
nor U6201 (N_6201,N_5347,N_5435);
xor U6202 (N_6202,N_5964,N_5116);
and U6203 (N_6203,N_5125,N_5637);
nor U6204 (N_6204,N_5539,N_5033);
xnor U6205 (N_6205,N_5877,N_5994);
nand U6206 (N_6206,N_5682,N_5337);
and U6207 (N_6207,N_5640,N_5342);
nand U6208 (N_6208,N_5043,N_5244);
and U6209 (N_6209,N_5331,N_5920);
and U6210 (N_6210,N_5453,N_5155);
and U6211 (N_6211,N_5292,N_5739);
and U6212 (N_6212,N_5300,N_5201);
and U6213 (N_6213,N_5628,N_5387);
and U6214 (N_6214,N_5924,N_5429);
or U6215 (N_6215,N_5717,N_5899);
nand U6216 (N_6216,N_5257,N_5564);
nand U6217 (N_6217,N_5365,N_5591);
nor U6218 (N_6218,N_5437,N_5976);
or U6219 (N_6219,N_5772,N_5972);
or U6220 (N_6220,N_5120,N_5610);
nor U6221 (N_6221,N_5725,N_5078);
nand U6222 (N_6222,N_5181,N_5973);
xor U6223 (N_6223,N_5518,N_5291);
or U6224 (N_6224,N_5872,N_5713);
nand U6225 (N_6225,N_5173,N_5754);
and U6226 (N_6226,N_5483,N_5782);
nand U6227 (N_6227,N_5451,N_5590);
nand U6228 (N_6228,N_5263,N_5140);
and U6229 (N_6229,N_5707,N_5228);
nand U6230 (N_6230,N_5481,N_5034);
or U6231 (N_6231,N_5041,N_5402);
nor U6232 (N_6232,N_5655,N_5526);
and U6233 (N_6233,N_5755,N_5200);
nor U6234 (N_6234,N_5074,N_5137);
nor U6235 (N_6235,N_5215,N_5831);
or U6236 (N_6236,N_5846,N_5478);
and U6237 (N_6237,N_5490,N_5897);
xnor U6238 (N_6238,N_5969,N_5807);
nor U6239 (N_6239,N_5094,N_5392);
and U6240 (N_6240,N_5940,N_5218);
or U6241 (N_6241,N_5231,N_5312);
nor U6242 (N_6242,N_5825,N_5588);
nand U6243 (N_6243,N_5573,N_5224);
nor U6244 (N_6244,N_5056,N_5455);
nand U6245 (N_6245,N_5792,N_5005);
or U6246 (N_6246,N_5833,N_5416);
nor U6247 (N_6247,N_5491,N_5674);
nand U6248 (N_6248,N_5710,N_5927);
or U6249 (N_6249,N_5188,N_5871);
nor U6250 (N_6250,N_5423,N_5270);
nor U6251 (N_6251,N_5910,N_5629);
or U6252 (N_6252,N_5593,N_5103);
and U6253 (N_6253,N_5863,N_5623);
nand U6254 (N_6254,N_5093,N_5225);
nand U6255 (N_6255,N_5142,N_5448);
xor U6256 (N_6256,N_5442,N_5031);
or U6257 (N_6257,N_5101,N_5427);
nor U6258 (N_6258,N_5652,N_5025);
nor U6259 (N_6259,N_5170,N_5261);
or U6260 (N_6260,N_5773,N_5714);
xor U6261 (N_6261,N_5941,N_5589);
nand U6262 (N_6262,N_5314,N_5875);
nor U6263 (N_6263,N_5192,N_5208);
nor U6264 (N_6264,N_5802,N_5386);
or U6265 (N_6265,N_5791,N_5613);
nor U6266 (N_6266,N_5766,N_5562);
xnor U6267 (N_6267,N_5553,N_5631);
or U6268 (N_6268,N_5544,N_5368);
nor U6269 (N_6269,N_5946,N_5799);
or U6270 (N_6270,N_5021,N_5380);
or U6271 (N_6271,N_5891,N_5381);
and U6272 (N_6272,N_5249,N_5418);
or U6273 (N_6273,N_5236,N_5438);
nor U6274 (N_6274,N_5046,N_5067);
nand U6275 (N_6275,N_5566,N_5229);
xor U6276 (N_6276,N_5656,N_5362);
nand U6277 (N_6277,N_5660,N_5136);
nand U6278 (N_6278,N_5971,N_5781);
nand U6279 (N_6279,N_5528,N_5313);
nor U6280 (N_6280,N_5790,N_5302);
or U6281 (N_6281,N_5487,N_5425);
or U6282 (N_6282,N_5883,N_5358);
and U6283 (N_6283,N_5400,N_5881);
and U6284 (N_6284,N_5052,N_5141);
and U6285 (N_6285,N_5744,N_5895);
xor U6286 (N_6286,N_5778,N_5653);
nand U6287 (N_6287,N_5524,N_5771);
nor U6288 (N_6288,N_5258,N_5108);
nor U6289 (N_6289,N_5219,N_5334);
and U6290 (N_6290,N_5488,N_5686);
nand U6291 (N_6291,N_5621,N_5364);
nand U6292 (N_6292,N_5794,N_5317);
nor U6293 (N_6293,N_5823,N_5981);
or U6294 (N_6294,N_5752,N_5505);
or U6295 (N_6295,N_5162,N_5060);
nor U6296 (N_6296,N_5324,N_5552);
and U6297 (N_6297,N_5454,N_5619);
and U6298 (N_6298,N_5865,N_5949);
xor U6299 (N_6299,N_5068,N_5123);
nand U6300 (N_6300,N_5988,N_5489);
and U6301 (N_6301,N_5680,N_5226);
nor U6302 (N_6302,N_5207,N_5467);
and U6303 (N_6303,N_5586,N_5926);
and U6304 (N_6304,N_5177,N_5379);
nand U6305 (N_6305,N_5273,N_5151);
nand U6306 (N_6306,N_5158,N_5113);
and U6307 (N_6307,N_5777,N_5851);
nand U6308 (N_6308,N_5287,N_5473);
nand U6309 (N_6309,N_5992,N_5690);
and U6310 (N_6310,N_5705,N_5697);
xor U6311 (N_6311,N_5014,N_5004);
xnor U6312 (N_6312,N_5072,N_5447);
nand U6313 (N_6313,N_5939,N_5541);
nand U6314 (N_6314,N_5995,N_5243);
nor U6315 (N_6315,N_5159,N_5115);
nand U6316 (N_6316,N_5393,N_5384);
and U6317 (N_6317,N_5720,N_5369);
nand U6318 (N_6318,N_5868,N_5470);
or U6319 (N_6319,N_5278,N_5841);
nand U6320 (N_6320,N_5044,N_5246);
or U6321 (N_6321,N_5684,N_5111);
nor U6322 (N_6322,N_5740,N_5563);
nand U6323 (N_6323,N_5843,N_5114);
nand U6324 (N_6324,N_5327,N_5741);
and U6325 (N_6325,N_5086,N_5788);
nand U6326 (N_6326,N_5183,N_5784);
nand U6327 (N_6327,N_5054,N_5683);
nor U6328 (N_6328,N_5731,N_5336);
xor U6329 (N_6329,N_5346,N_5396);
nor U6330 (N_6330,N_5769,N_5516);
xor U6331 (N_6331,N_5578,N_5016);
nor U6332 (N_6332,N_5649,N_5426);
or U6333 (N_6333,N_5194,N_5750);
and U6334 (N_6334,N_5815,N_5730);
and U6335 (N_6335,N_5405,N_5793);
and U6336 (N_6336,N_5252,N_5099);
or U6337 (N_6337,N_5071,N_5585);
nand U6338 (N_6338,N_5092,N_5709);
nand U6339 (N_6339,N_5965,N_5251);
nor U6340 (N_6340,N_5703,N_5436);
or U6341 (N_6341,N_5102,N_5978);
and U6342 (N_6342,N_5506,N_5622);
nand U6343 (N_6343,N_5306,N_5087);
nand U6344 (N_6344,N_5888,N_5394);
and U6345 (N_6345,N_5840,N_5702);
and U6346 (N_6346,N_5929,N_5026);
nor U6347 (N_6347,N_5770,N_5197);
or U6348 (N_6348,N_5198,N_5217);
or U6349 (N_6349,N_5315,N_5129);
nand U6350 (N_6350,N_5374,N_5980);
nor U6351 (N_6351,N_5403,N_5604);
nor U6352 (N_6352,N_5693,N_5098);
nor U6353 (N_6353,N_5372,N_5535);
or U6354 (N_6354,N_5274,N_5457);
or U6355 (N_6355,N_5063,N_5698);
and U6356 (N_6356,N_5268,N_5522);
nand U6357 (N_6357,N_5687,N_5958);
or U6358 (N_6358,N_5904,N_5839);
nand U6359 (N_6359,N_5020,N_5233);
xnor U6360 (N_6360,N_5428,N_5156);
xnor U6361 (N_6361,N_5889,N_5951);
or U6362 (N_6362,N_5696,N_5082);
or U6363 (N_6363,N_5668,N_5480);
nand U6364 (N_6364,N_5463,N_5230);
nor U6365 (N_6365,N_5279,N_5288);
or U6366 (N_6366,N_5859,N_5748);
nor U6367 (N_6367,N_5704,N_5127);
nand U6368 (N_6368,N_5960,N_5134);
or U6369 (N_6369,N_5245,N_5017);
and U6370 (N_6370,N_5699,N_5935);
nor U6371 (N_6371,N_5007,N_5216);
nor U6372 (N_6372,N_5650,N_5834);
nor U6373 (N_6373,N_5677,N_5281);
xnor U6374 (N_6374,N_5193,N_5932);
nor U6375 (N_6375,N_5206,N_5813);
nor U6376 (N_6376,N_5298,N_5861);
or U6377 (N_6377,N_5477,N_5135);
xnor U6378 (N_6378,N_5343,N_5611);
and U6379 (N_6379,N_5765,N_5356);
nor U6380 (N_6380,N_5360,N_5154);
and U6381 (N_6381,N_5800,N_5509);
nand U6382 (N_6382,N_5424,N_5433);
nand U6383 (N_6383,N_5180,N_5204);
nor U6384 (N_6384,N_5152,N_5378);
nor U6385 (N_6385,N_5786,N_5894);
nor U6386 (N_6386,N_5569,N_5265);
nor U6387 (N_6387,N_5930,N_5550);
or U6388 (N_6388,N_5678,N_5517);
nor U6389 (N_6389,N_5812,N_5991);
and U6390 (N_6390,N_5179,N_5559);
or U6391 (N_6391,N_5338,N_5472);
nand U6392 (N_6392,N_5419,N_5646);
and U6393 (N_6393,N_5856,N_5323);
and U6394 (N_6394,N_5494,N_5557);
xnor U6395 (N_6395,N_5352,N_5909);
nor U6396 (N_6396,N_5659,N_5371);
nand U6397 (N_6397,N_5855,N_5715);
nand U6398 (N_6398,N_5666,N_5430);
nor U6399 (N_6399,N_5091,N_5783);
nor U6400 (N_6400,N_5002,N_5242);
nor U6401 (N_6401,N_5820,N_5202);
nor U6402 (N_6402,N_5045,N_5290);
nor U6403 (N_6403,N_5601,N_5915);
and U6404 (N_6404,N_5808,N_5189);
and U6405 (N_6405,N_5560,N_5620);
xor U6406 (N_6406,N_5328,N_5532);
and U6407 (N_6407,N_5919,N_5163);
nor U6408 (N_6408,N_5213,N_5906);
or U6409 (N_6409,N_5303,N_5036);
and U6410 (N_6410,N_5854,N_5908);
and U6411 (N_6411,N_5112,N_5892);
nand U6412 (N_6412,N_5785,N_5675);
xor U6413 (N_6413,N_5605,N_5603);
nor U6414 (N_6414,N_5479,N_5600);
and U6415 (N_6415,N_5030,N_5761);
nor U6416 (N_6416,N_5144,N_5461);
xor U6417 (N_6417,N_5938,N_5796);
xnor U6418 (N_6418,N_5734,N_5409);
nor U6419 (N_6419,N_5383,N_5410);
and U6420 (N_6420,N_5537,N_5203);
nand U6421 (N_6421,N_5716,N_5844);
and U6422 (N_6422,N_5474,N_5050);
and U6423 (N_6423,N_5735,N_5869);
or U6424 (N_6424,N_5023,N_5928);
or U6425 (N_6425,N_5466,N_5411);
or U6426 (N_6426,N_5862,N_5679);
or U6427 (N_6427,N_5476,N_5606);
nor U6428 (N_6428,N_5886,N_5643);
or U6429 (N_6429,N_5918,N_5344);
xnor U6430 (N_6430,N_5357,N_5333);
nor U6431 (N_6431,N_5350,N_5822);
xor U6432 (N_6432,N_5624,N_5898);
and U6433 (N_6433,N_5408,N_5987);
and U6434 (N_6434,N_5377,N_5967);
and U6435 (N_6435,N_5458,N_5104);
nor U6436 (N_6436,N_5746,N_5751);
nand U6437 (N_6437,N_5264,N_5150);
or U6438 (N_6438,N_5042,N_5596);
or U6439 (N_6439,N_5950,N_5464);
or U6440 (N_6440,N_5545,N_5959);
nand U6441 (N_6441,N_5612,N_5625);
or U6442 (N_6442,N_5648,N_5450);
nor U6443 (N_6443,N_5618,N_5354);
xor U6444 (N_6444,N_5616,N_5006);
nand U6445 (N_6445,N_5501,N_5407);
and U6446 (N_6446,N_5504,N_5223);
xnor U6447 (N_6447,N_5893,N_5896);
and U6448 (N_6448,N_5096,N_5644);
or U6449 (N_6449,N_5512,N_5529);
nand U6450 (N_6450,N_5826,N_5013);
nand U6451 (N_6451,N_5767,N_5974);
nor U6452 (N_6452,N_5475,N_5641);
or U6453 (N_6453,N_5000,N_5169);
or U6454 (N_6454,N_5867,N_5912);
nor U6455 (N_6455,N_5963,N_5220);
xnor U6456 (N_6456,N_5299,N_5209);
nor U6457 (N_6457,N_5498,N_5556);
or U6458 (N_6458,N_5743,N_5131);
nor U6459 (N_6459,N_5395,N_5876);
and U6460 (N_6460,N_5803,N_5234);
nand U6461 (N_6461,N_5998,N_5237);
and U6462 (N_6462,N_5582,N_5576);
xor U6463 (N_6463,N_5009,N_5510);
or U6464 (N_6464,N_5095,N_5756);
nor U6465 (N_6465,N_5975,N_5439);
nor U6466 (N_6466,N_5412,N_5145);
nand U6467 (N_6467,N_5990,N_5572);
xnor U6468 (N_6468,N_5001,N_5143);
or U6469 (N_6469,N_5070,N_5729);
or U6470 (N_6470,N_5235,N_5870);
nor U6471 (N_6471,N_5275,N_5592);
xor U6472 (N_6472,N_5945,N_5852);
nand U6473 (N_6473,N_5986,N_5880);
or U6474 (N_6474,N_5952,N_5688);
and U6475 (N_6475,N_5630,N_5903);
or U6476 (N_6476,N_5205,N_5212);
and U6477 (N_6477,N_5979,N_5993);
nor U6478 (N_6478,N_5608,N_5525);
xor U6479 (N_6479,N_5917,N_5542);
nand U6480 (N_6480,N_5376,N_5390);
nand U6481 (N_6481,N_5029,N_5809);
nor U6482 (N_6482,N_5304,N_5239);
nor U6483 (N_6483,N_5259,N_5373);
and U6484 (N_6484,N_5657,N_5989);
or U6485 (N_6485,N_5533,N_5443);
nand U6486 (N_6486,N_5295,N_5255);
and U6487 (N_6487,N_5015,N_5465);
or U6488 (N_6488,N_5100,N_5166);
and U6489 (N_6489,N_5607,N_5947);
or U6490 (N_6490,N_5548,N_5953);
nor U6491 (N_6491,N_5174,N_5066);
nand U6492 (N_6492,N_5460,N_5097);
and U6493 (N_6493,N_5038,N_5375);
nand U6494 (N_6494,N_5580,N_5348);
and U6495 (N_6495,N_5547,N_5124);
nand U6496 (N_6496,N_5942,N_5728);
and U6497 (N_6497,N_5733,N_5415);
nor U6498 (N_6498,N_5527,N_5779);
and U6499 (N_6499,N_5719,N_5925);
and U6500 (N_6500,N_5307,N_5336);
nand U6501 (N_6501,N_5863,N_5100);
or U6502 (N_6502,N_5800,N_5733);
xor U6503 (N_6503,N_5896,N_5507);
nor U6504 (N_6504,N_5525,N_5677);
and U6505 (N_6505,N_5343,N_5780);
nor U6506 (N_6506,N_5579,N_5174);
or U6507 (N_6507,N_5351,N_5193);
and U6508 (N_6508,N_5333,N_5420);
nand U6509 (N_6509,N_5141,N_5461);
xnor U6510 (N_6510,N_5194,N_5088);
nand U6511 (N_6511,N_5663,N_5596);
xor U6512 (N_6512,N_5270,N_5929);
and U6513 (N_6513,N_5370,N_5847);
xor U6514 (N_6514,N_5764,N_5335);
or U6515 (N_6515,N_5347,N_5345);
nor U6516 (N_6516,N_5022,N_5112);
xor U6517 (N_6517,N_5719,N_5325);
nor U6518 (N_6518,N_5864,N_5666);
nor U6519 (N_6519,N_5664,N_5599);
nand U6520 (N_6520,N_5528,N_5016);
xnor U6521 (N_6521,N_5992,N_5421);
and U6522 (N_6522,N_5524,N_5033);
and U6523 (N_6523,N_5021,N_5983);
or U6524 (N_6524,N_5541,N_5209);
nor U6525 (N_6525,N_5408,N_5915);
nand U6526 (N_6526,N_5961,N_5522);
nor U6527 (N_6527,N_5235,N_5582);
or U6528 (N_6528,N_5464,N_5396);
and U6529 (N_6529,N_5522,N_5492);
xnor U6530 (N_6530,N_5993,N_5311);
or U6531 (N_6531,N_5220,N_5612);
and U6532 (N_6532,N_5472,N_5962);
xor U6533 (N_6533,N_5203,N_5222);
or U6534 (N_6534,N_5012,N_5485);
nor U6535 (N_6535,N_5297,N_5755);
and U6536 (N_6536,N_5120,N_5677);
nand U6537 (N_6537,N_5725,N_5015);
or U6538 (N_6538,N_5127,N_5751);
and U6539 (N_6539,N_5367,N_5677);
nand U6540 (N_6540,N_5458,N_5318);
nor U6541 (N_6541,N_5577,N_5169);
and U6542 (N_6542,N_5338,N_5543);
or U6543 (N_6543,N_5518,N_5979);
nand U6544 (N_6544,N_5431,N_5091);
nand U6545 (N_6545,N_5484,N_5238);
and U6546 (N_6546,N_5348,N_5986);
or U6547 (N_6547,N_5054,N_5227);
or U6548 (N_6548,N_5012,N_5064);
or U6549 (N_6549,N_5906,N_5766);
nor U6550 (N_6550,N_5928,N_5954);
nand U6551 (N_6551,N_5614,N_5358);
and U6552 (N_6552,N_5635,N_5059);
or U6553 (N_6553,N_5115,N_5371);
xor U6554 (N_6554,N_5586,N_5566);
nand U6555 (N_6555,N_5788,N_5428);
and U6556 (N_6556,N_5602,N_5134);
xnor U6557 (N_6557,N_5928,N_5999);
and U6558 (N_6558,N_5725,N_5905);
and U6559 (N_6559,N_5449,N_5491);
and U6560 (N_6560,N_5662,N_5290);
or U6561 (N_6561,N_5971,N_5214);
or U6562 (N_6562,N_5853,N_5431);
or U6563 (N_6563,N_5932,N_5120);
nor U6564 (N_6564,N_5913,N_5900);
and U6565 (N_6565,N_5515,N_5898);
or U6566 (N_6566,N_5181,N_5515);
or U6567 (N_6567,N_5118,N_5323);
and U6568 (N_6568,N_5429,N_5534);
nor U6569 (N_6569,N_5018,N_5692);
nand U6570 (N_6570,N_5898,N_5411);
and U6571 (N_6571,N_5928,N_5415);
nand U6572 (N_6572,N_5233,N_5449);
nand U6573 (N_6573,N_5938,N_5161);
nand U6574 (N_6574,N_5820,N_5446);
and U6575 (N_6575,N_5137,N_5662);
nand U6576 (N_6576,N_5789,N_5520);
and U6577 (N_6577,N_5697,N_5832);
nor U6578 (N_6578,N_5410,N_5456);
or U6579 (N_6579,N_5213,N_5290);
and U6580 (N_6580,N_5704,N_5825);
nor U6581 (N_6581,N_5753,N_5688);
xor U6582 (N_6582,N_5277,N_5670);
and U6583 (N_6583,N_5165,N_5559);
nand U6584 (N_6584,N_5662,N_5596);
or U6585 (N_6585,N_5295,N_5002);
or U6586 (N_6586,N_5216,N_5854);
nand U6587 (N_6587,N_5842,N_5132);
xor U6588 (N_6588,N_5706,N_5832);
nand U6589 (N_6589,N_5813,N_5414);
nor U6590 (N_6590,N_5385,N_5135);
nand U6591 (N_6591,N_5617,N_5834);
nor U6592 (N_6592,N_5284,N_5565);
xor U6593 (N_6593,N_5703,N_5421);
nand U6594 (N_6594,N_5570,N_5751);
or U6595 (N_6595,N_5531,N_5471);
or U6596 (N_6596,N_5334,N_5665);
and U6597 (N_6597,N_5425,N_5498);
nor U6598 (N_6598,N_5556,N_5127);
nand U6599 (N_6599,N_5722,N_5588);
nand U6600 (N_6600,N_5420,N_5119);
xnor U6601 (N_6601,N_5558,N_5686);
nor U6602 (N_6602,N_5450,N_5485);
and U6603 (N_6603,N_5983,N_5895);
and U6604 (N_6604,N_5223,N_5757);
nor U6605 (N_6605,N_5246,N_5913);
and U6606 (N_6606,N_5426,N_5503);
nand U6607 (N_6607,N_5275,N_5642);
or U6608 (N_6608,N_5509,N_5066);
or U6609 (N_6609,N_5623,N_5757);
nand U6610 (N_6610,N_5168,N_5724);
and U6611 (N_6611,N_5363,N_5149);
and U6612 (N_6612,N_5441,N_5834);
nor U6613 (N_6613,N_5291,N_5902);
and U6614 (N_6614,N_5296,N_5916);
nor U6615 (N_6615,N_5605,N_5734);
or U6616 (N_6616,N_5093,N_5258);
nand U6617 (N_6617,N_5177,N_5123);
or U6618 (N_6618,N_5521,N_5040);
nor U6619 (N_6619,N_5337,N_5206);
nor U6620 (N_6620,N_5115,N_5818);
or U6621 (N_6621,N_5976,N_5816);
nand U6622 (N_6622,N_5521,N_5773);
and U6623 (N_6623,N_5747,N_5526);
and U6624 (N_6624,N_5411,N_5167);
and U6625 (N_6625,N_5148,N_5938);
or U6626 (N_6626,N_5892,N_5358);
xor U6627 (N_6627,N_5775,N_5960);
nor U6628 (N_6628,N_5115,N_5521);
or U6629 (N_6629,N_5780,N_5776);
and U6630 (N_6630,N_5575,N_5331);
nand U6631 (N_6631,N_5922,N_5711);
and U6632 (N_6632,N_5367,N_5109);
and U6633 (N_6633,N_5676,N_5402);
and U6634 (N_6634,N_5466,N_5386);
nand U6635 (N_6635,N_5886,N_5180);
nor U6636 (N_6636,N_5935,N_5518);
nand U6637 (N_6637,N_5591,N_5135);
nand U6638 (N_6638,N_5534,N_5227);
nor U6639 (N_6639,N_5356,N_5750);
or U6640 (N_6640,N_5750,N_5247);
nor U6641 (N_6641,N_5500,N_5424);
or U6642 (N_6642,N_5732,N_5610);
nor U6643 (N_6643,N_5100,N_5337);
nand U6644 (N_6644,N_5597,N_5930);
xnor U6645 (N_6645,N_5785,N_5504);
nand U6646 (N_6646,N_5095,N_5843);
or U6647 (N_6647,N_5667,N_5492);
nor U6648 (N_6648,N_5010,N_5363);
or U6649 (N_6649,N_5298,N_5502);
and U6650 (N_6650,N_5561,N_5696);
or U6651 (N_6651,N_5048,N_5279);
xnor U6652 (N_6652,N_5596,N_5364);
and U6653 (N_6653,N_5044,N_5776);
nor U6654 (N_6654,N_5798,N_5565);
nand U6655 (N_6655,N_5648,N_5687);
or U6656 (N_6656,N_5528,N_5275);
and U6657 (N_6657,N_5246,N_5461);
nor U6658 (N_6658,N_5860,N_5725);
or U6659 (N_6659,N_5915,N_5459);
and U6660 (N_6660,N_5921,N_5187);
nand U6661 (N_6661,N_5450,N_5941);
xnor U6662 (N_6662,N_5597,N_5234);
nor U6663 (N_6663,N_5756,N_5706);
or U6664 (N_6664,N_5310,N_5989);
nor U6665 (N_6665,N_5218,N_5760);
nor U6666 (N_6666,N_5149,N_5425);
nor U6667 (N_6667,N_5439,N_5768);
xnor U6668 (N_6668,N_5293,N_5150);
and U6669 (N_6669,N_5453,N_5258);
nand U6670 (N_6670,N_5524,N_5938);
nor U6671 (N_6671,N_5185,N_5642);
or U6672 (N_6672,N_5083,N_5280);
xor U6673 (N_6673,N_5333,N_5120);
or U6674 (N_6674,N_5021,N_5927);
nor U6675 (N_6675,N_5135,N_5357);
nand U6676 (N_6676,N_5032,N_5138);
and U6677 (N_6677,N_5491,N_5770);
nor U6678 (N_6678,N_5225,N_5253);
nor U6679 (N_6679,N_5376,N_5098);
or U6680 (N_6680,N_5427,N_5262);
and U6681 (N_6681,N_5346,N_5501);
or U6682 (N_6682,N_5171,N_5068);
and U6683 (N_6683,N_5980,N_5078);
nor U6684 (N_6684,N_5860,N_5480);
and U6685 (N_6685,N_5506,N_5761);
and U6686 (N_6686,N_5867,N_5035);
and U6687 (N_6687,N_5471,N_5488);
nand U6688 (N_6688,N_5008,N_5938);
xor U6689 (N_6689,N_5373,N_5170);
and U6690 (N_6690,N_5220,N_5677);
nand U6691 (N_6691,N_5645,N_5771);
or U6692 (N_6692,N_5812,N_5804);
and U6693 (N_6693,N_5456,N_5275);
nor U6694 (N_6694,N_5266,N_5805);
and U6695 (N_6695,N_5816,N_5913);
and U6696 (N_6696,N_5361,N_5664);
nor U6697 (N_6697,N_5301,N_5323);
or U6698 (N_6698,N_5206,N_5647);
and U6699 (N_6699,N_5032,N_5567);
xor U6700 (N_6700,N_5815,N_5501);
or U6701 (N_6701,N_5786,N_5366);
and U6702 (N_6702,N_5486,N_5305);
and U6703 (N_6703,N_5547,N_5973);
nor U6704 (N_6704,N_5538,N_5180);
xnor U6705 (N_6705,N_5737,N_5543);
nor U6706 (N_6706,N_5544,N_5818);
nor U6707 (N_6707,N_5076,N_5332);
and U6708 (N_6708,N_5545,N_5479);
and U6709 (N_6709,N_5307,N_5397);
and U6710 (N_6710,N_5380,N_5866);
or U6711 (N_6711,N_5872,N_5420);
and U6712 (N_6712,N_5842,N_5641);
nor U6713 (N_6713,N_5179,N_5780);
nor U6714 (N_6714,N_5784,N_5809);
or U6715 (N_6715,N_5780,N_5389);
or U6716 (N_6716,N_5580,N_5158);
and U6717 (N_6717,N_5840,N_5645);
or U6718 (N_6718,N_5167,N_5812);
nand U6719 (N_6719,N_5789,N_5208);
nand U6720 (N_6720,N_5430,N_5979);
nand U6721 (N_6721,N_5897,N_5709);
and U6722 (N_6722,N_5858,N_5378);
and U6723 (N_6723,N_5055,N_5507);
nand U6724 (N_6724,N_5488,N_5888);
nand U6725 (N_6725,N_5611,N_5745);
and U6726 (N_6726,N_5896,N_5869);
or U6727 (N_6727,N_5775,N_5665);
nor U6728 (N_6728,N_5598,N_5028);
nor U6729 (N_6729,N_5274,N_5683);
xor U6730 (N_6730,N_5304,N_5766);
and U6731 (N_6731,N_5104,N_5471);
xnor U6732 (N_6732,N_5218,N_5125);
nand U6733 (N_6733,N_5332,N_5160);
and U6734 (N_6734,N_5713,N_5015);
nand U6735 (N_6735,N_5191,N_5934);
nor U6736 (N_6736,N_5357,N_5370);
xnor U6737 (N_6737,N_5036,N_5355);
or U6738 (N_6738,N_5241,N_5428);
or U6739 (N_6739,N_5141,N_5921);
nand U6740 (N_6740,N_5573,N_5244);
nand U6741 (N_6741,N_5733,N_5288);
nor U6742 (N_6742,N_5132,N_5771);
and U6743 (N_6743,N_5859,N_5587);
or U6744 (N_6744,N_5049,N_5599);
or U6745 (N_6745,N_5284,N_5276);
nor U6746 (N_6746,N_5901,N_5916);
nor U6747 (N_6747,N_5665,N_5061);
nand U6748 (N_6748,N_5677,N_5949);
nand U6749 (N_6749,N_5133,N_5245);
and U6750 (N_6750,N_5153,N_5413);
and U6751 (N_6751,N_5656,N_5077);
xor U6752 (N_6752,N_5327,N_5040);
and U6753 (N_6753,N_5379,N_5645);
nor U6754 (N_6754,N_5741,N_5714);
and U6755 (N_6755,N_5470,N_5452);
nand U6756 (N_6756,N_5799,N_5199);
nand U6757 (N_6757,N_5393,N_5826);
nor U6758 (N_6758,N_5892,N_5238);
nor U6759 (N_6759,N_5972,N_5136);
nand U6760 (N_6760,N_5690,N_5044);
nor U6761 (N_6761,N_5397,N_5555);
nand U6762 (N_6762,N_5749,N_5956);
and U6763 (N_6763,N_5976,N_5011);
and U6764 (N_6764,N_5958,N_5680);
nor U6765 (N_6765,N_5674,N_5147);
xnor U6766 (N_6766,N_5592,N_5453);
and U6767 (N_6767,N_5186,N_5030);
nand U6768 (N_6768,N_5011,N_5802);
xor U6769 (N_6769,N_5083,N_5303);
and U6770 (N_6770,N_5108,N_5304);
nor U6771 (N_6771,N_5578,N_5745);
nor U6772 (N_6772,N_5885,N_5053);
xnor U6773 (N_6773,N_5511,N_5084);
and U6774 (N_6774,N_5077,N_5601);
nand U6775 (N_6775,N_5298,N_5178);
and U6776 (N_6776,N_5232,N_5068);
xor U6777 (N_6777,N_5061,N_5071);
and U6778 (N_6778,N_5059,N_5447);
or U6779 (N_6779,N_5209,N_5486);
or U6780 (N_6780,N_5726,N_5860);
and U6781 (N_6781,N_5259,N_5539);
nor U6782 (N_6782,N_5446,N_5588);
xnor U6783 (N_6783,N_5312,N_5846);
or U6784 (N_6784,N_5263,N_5410);
nand U6785 (N_6785,N_5183,N_5050);
nor U6786 (N_6786,N_5556,N_5460);
or U6787 (N_6787,N_5797,N_5567);
nor U6788 (N_6788,N_5146,N_5130);
nand U6789 (N_6789,N_5493,N_5988);
and U6790 (N_6790,N_5150,N_5375);
xnor U6791 (N_6791,N_5553,N_5435);
or U6792 (N_6792,N_5181,N_5664);
nand U6793 (N_6793,N_5382,N_5053);
or U6794 (N_6794,N_5877,N_5600);
and U6795 (N_6795,N_5647,N_5857);
and U6796 (N_6796,N_5344,N_5106);
nand U6797 (N_6797,N_5336,N_5137);
nor U6798 (N_6798,N_5440,N_5573);
nand U6799 (N_6799,N_5073,N_5856);
nand U6800 (N_6800,N_5151,N_5847);
nor U6801 (N_6801,N_5644,N_5796);
and U6802 (N_6802,N_5502,N_5692);
and U6803 (N_6803,N_5987,N_5486);
or U6804 (N_6804,N_5040,N_5168);
nor U6805 (N_6805,N_5387,N_5908);
and U6806 (N_6806,N_5581,N_5807);
nor U6807 (N_6807,N_5011,N_5037);
nand U6808 (N_6808,N_5318,N_5902);
nor U6809 (N_6809,N_5311,N_5760);
or U6810 (N_6810,N_5813,N_5673);
nor U6811 (N_6811,N_5205,N_5043);
xor U6812 (N_6812,N_5728,N_5561);
and U6813 (N_6813,N_5776,N_5332);
and U6814 (N_6814,N_5064,N_5450);
and U6815 (N_6815,N_5223,N_5629);
nor U6816 (N_6816,N_5327,N_5264);
nor U6817 (N_6817,N_5650,N_5938);
and U6818 (N_6818,N_5783,N_5449);
and U6819 (N_6819,N_5826,N_5188);
nand U6820 (N_6820,N_5631,N_5421);
and U6821 (N_6821,N_5836,N_5593);
nor U6822 (N_6822,N_5751,N_5052);
nor U6823 (N_6823,N_5673,N_5554);
nand U6824 (N_6824,N_5483,N_5309);
or U6825 (N_6825,N_5243,N_5367);
and U6826 (N_6826,N_5402,N_5298);
nand U6827 (N_6827,N_5041,N_5241);
or U6828 (N_6828,N_5818,N_5795);
or U6829 (N_6829,N_5627,N_5118);
and U6830 (N_6830,N_5525,N_5897);
or U6831 (N_6831,N_5011,N_5971);
and U6832 (N_6832,N_5870,N_5625);
or U6833 (N_6833,N_5883,N_5509);
nor U6834 (N_6834,N_5600,N_5496);
and U6835 (N_6835,N_5813,N_5082);
and U6836 (N_6836,N_5398,N_5689);
xor U6837 (N_6837,N_5817,N_5184);
or U6838 (N_6838,N_5143,N_5054);
or U6839 (N_6839,N_5565,N_5482);
nand U6840 (N_6840,N_5663,N_5267);
nand U6841 (N_6841,N_5599,N_5858);
nor U6842 (N_6842,N_5128,N_5716);
and U6843 (N_6843,N_5731,N_5521);
nand U6844 (N_6844,N_5706,N_5866);
nand U6845 (N_6845,N_5315,N_5458);
and U6846 (N_6846,N_5329,N_5537);
or U6847 (N_6847,N_5327,N_5766);
nand U6848 (N_6848,N_5594,N_5712);
nand U6849 (N_6849,N_5006,N_5132);
nand U6850 (N_6850,N_5318,N_5504);
nor U6851 (N_6851,N_5786,N_5646);
nand U6852 (N_6852,N_5019,N_5961);
nand U6853 (N_6853,N_5109,N_5127);
or U6854 (N_6854,N_5754,N_5389);
nor U6855 (N_6855,N_5235,N_5368);
and U6856 (N_6856,N_5485,N_5858);
nand U6857 (N_6857,N_5464,N_5871);
and U6858 (N_6858,N_5684,N_5763);
nand U6859 (N_6859,N_5846,N_5436);
and U6860 (N_6860,N_5447,N_5694);
or U6861 (N_6861,N_5948,N_5786);
nor U6862 (N_6862,N_5224,N_5285);
xnor U6863 (N_6863,N_5201,N_5908);
and U6864 (N_6864,N_5422,N_5616);
or U6865 (N_6865,N_5544,N_5764);
or U6866 (N_6866,N_5517,N_5016);
nand U6867 (N_6867,N_5154,N_5150);
nor U6868 (N_6868,N_5379,N_5689);
or U6869 (N_6869,N_5529,N_5930);
and U6870 (N_6870,N_5112,N_5276);
nand U6871 (N_6871,N_5341,N_5822);
nand U6872 (N_6872,N_5668,N_5469);
or U6873 (N_6873,N_5508,N_5632);
or U6874 (N_6874,N_5914,N_5128);
nor U6875 (N_6875,N_5971,N_5659);
nand U6876 (N_6876,N_5288,N_5881);
and U6877 (N_6877,N_5486,N_5130);
nand U6878 (N_6878,N_5139,N_5068);
or U6879 (N_6879,N_5250,N_5733);
nor U6880 (N_6880,N_5884,N_5546);
and U6881 (N_6881,N_5855,N_5173);
or U6882 (N_6882,N_5986,N_5442);
and U6883 (N_6883,N_5884,N_5907);
nor U6884 (N_6884,N_5908,N_5016);
xor U6885 (N_6885,N_5494,N_5594);
nor U6886 (N_6886,N_5649,N_5159);
xor U6887 (N_6887,N_5368,N_5462);
nor U6888 (N_6888,N_5470,N_5953);
or U6889 (N_6889,N_5181,N_5462);
nand U6890 (N_6890,N_5411,N_5864);
nand U6891 (N_6891,N_5728,N_5919);
and U6892 (N_6892,N_5293,N_5854);
or U6893 (N_6893,N_5421,N_5448);
or U6894 (N_6894,N_5453,N_5313);
nor U6895 (N_6895,N_5114,N_5773);
and U6896 (N_6896,N_5509,N_5197);
and U6897 (N_6897,N_5929,N_5273);
or U6898 (N_6898,N_5265,N_5450);
nand U6899 (N_6899,N_5609,N_5842);
nand U6900 (N_6900,N_5288,N_5250);
or U6901 (N_6901,N_5144,N_5369);
or U6902 (N_6902,N_5903,N_5823);
and U6903 (N_6903,N_5746,N_5686);
nand U6904 (N_6904,N_5178,N_5108);
nor U6905 (N_6905,N_5998,N_5381);
or U6906 (N_6906,N_5759,N_5739);
and U6907 (N_6907,N_5328,N_5227);
nor U6908 (N_6908,N_5731,N_5176);
nor U6909 (N_6909,N_5730,N_5296);
nand U6910 (N_6910,N_5125,N_5467);
xor U6911 (N_6911,N_5918,N_5626);
and U6912 (N_6912,N_5554,N_5742);
nor U6913 (N_6913,N_5906,N_5298);
or U6914 (N_6914,N_5184,N_5108);
and U6915 (N_6915,N_5368,N_5730);
and U6916 (N_6916,N_5999,N_5537);
nor U6917 (N_6917,N_5725,N_5870);
nor U6918 (N_6918,N_5563,N_5832);
nor U6919 (N_6919,N_5407,N_5457);
xnor U6920 (N_6920,N_5191,N_5266);
nand U6921 (N_6921,N_5273,N_5898);
and U6922 (N_6922,N_5837,N_5429);
nor U6923 (N_6923,N_5533,N_5213);
nand U6924 (N_6924,N_5357,N_5652);
nor U6925 (N_6925,N_5378,N_5834);
or U6926 (N_6926,N_5962,N_5245);
xor U6927 (N_6927,N_5360,N_5376);
or U6928 (N_6928,N_5797,N_5943);
and U6929 (N_6929,N_5941,N_5151);
nand U6930 (N_6930,N_5925,N_5814);
xor U6931 (N_6931,N_5049,N_5269);
and U6932 (N_6932,N_5642,N_5135);
xor U6933 (N_6933,N_5842,N_5787);
nand U6934 (N_6934,N_5548,N_5435);
nor U6935 (N_6935,N_5972,N_5395);
or U6936 (N_6936,N_5805,N_5749);
or U6937 (N_6937,N_5853,N_5197);
and U6938 (N_6938,N_5782,N_5143);
or U6939 (N_6939,N_5701,N_5817);
nor U6940 (N_6940,N_5990,N_5005);
nand U6941 (N_6941,N_5156,N_5581);
nand U6942 (N_6942,N_5355,N_5224);
nor U6943 (N_6943,N_5620,N_5837);
nor U6944 (N_6944,N_5961,N_5084);
and U6945 (N_6945,N_5890,N_5828);
nor U6946 (N_6946,N_5033,N_5440);
or U6947 (N_6947,N_5090,N_5331);
or U6948 (N_6948,N_5038,N_5909);
and U6949 (N_6949,N_5677,N_5965);
nand U6950 (N_6950,N_5359,N_5993);
xor U6951 (N_6951,N_5803,N_5293);
or U6952 (N_6952,N_5265,N_5109);
or U6953 (N_6953,N_5697,N_5387);
or U6954 (N_6954,N_5552,N_5941);
nor U6955 (N_6955,N_5087,N_5585);
xor U6956 (N_6956,N_5263,N_5186);
xor U6957 (N_6957,N_5705,N_5007);
nor U6958 (N_6958,N_5950,N_5996);
and U6959 (N_6959,N_5600,N_5292);
nor U6960 (N_6960,N_5848,N_5893);
xor U6961 (N_6961,N_5776,N_5998);
xor U6962 (N_6962,N_5546,N_5175);
nor U6963 (N_6963,N_5232,N_5763);
nand U6964 (N_6964,N_5429,N_5882);
or U6965 (N_6965,N_5741,N_5275);
nor U6966 (N_6966,N_5787,N_5976);
and U6967 (N_6967,N_5396,N_5003);
xor U6968 (N_6968,N_5472,N_5507);
and U6969 (N_6969,N_5722,N_5517);
nor U6970 (N_6970,N_5162,N_5380);
or U6971 (N_6971,N_5510,N_5000);
and U6972 (N_6972,N_5727,N_5206);
nand U6973 (N_6973,N_5025,N_5289);
or U6974 (N_6974,N_5443,N_5418);
xor U6975 (N_6975,N_5445,N_5996);
nand U6976 (N_6976,N_5475,N_5275);
nor U6977 (N_6977,N_5732,N_5377);
nand U6978 (N_6978,N_5128,N_5839);
nor U6979 (N_6979,N_5836,N_5196);
xor U6980 (N_6980,N_5874,N_5573);
or U6981 (N_6981,N_5320,N_5297);
nor U6982 (N_6982,N_5505,N_5778);
or U6983 (N_6983,N_5777,N_5774);
and U6984 (N_6984,N_5806,N_5934);
xnor U6985 (N_6985,N_5071,N_5316);
nor U6986 (N_6986,N_5781,N_5752);
and U6987 (N_6987,N_5615,N_5955);
or U6988 (N_6988,N_5225,N_5464);
or U6989 (N_6989,N_5958,N_5757);
xor U6990 (N_6990,N_5543,N_5074);
nor U6991 (N_6991,N_5521,N_5052);
and U6992 (N_6992,N_5224,N_5815);
or U6993 (N_6993,N_5563,N_5537);
or U6994 (N_6994,N_5353,N_5064);
nor U6995 (N_6995,N_5890,N_5863);
xor U6996 (N_6996,N_5806,N_5830);
and U6997 (N_6997,N_5088,N_5177);
nor U6998 (N_6998,N_5344,N_5204);
nor U6999 (N_6999,N_5306,N_5777);
nor U7000 (N_7000,N_6187,N_6443);
xor U7001 (N_7001,N_6118,N_6981);
nand U7002 (N_7002,N_6344,N_6907);
or U7003 (N_7003,N_6918,N_6915);
and U7004 (N_7004,N_6507,N_6682);
or U7005 (N_7005,N_6246,N_6942);
and U7006 (N_7006,N_6498,N_6331);
and U7007 (N_7007,N_6342,N_6808);
xnor U7008 (N_7008,N_6862,N_6822);
nor U7009 (N_7009,N_6031,N_6400);
and U7010 (N_7010,N_6112,N_6480);
and U7011 (N_7011,N_6529,N_6912);
nor U7012 (N_7012,N_6626,N_6855);
nor U7013 (N_7013,N_6766,N_6100);
nand U7014 (N_7014,N_6490,N_6913);
and U7015 (N_7015,N_6817,N_6253);
xnor U7016 (N_7016,N_6420,N_6314);
or U7017 (N_7017,N_6273,N_6572);
or U7018 (N_7018,N_6271,N_6881);
nor U7019 (N_7019,N_6738,N_6160);
nand U7020 (N_7020,N_6235,N_6526);
nor U7021 (N_7021,N_6302,N_6208);
or U7022 (N_7022,N_6047,N_6362);
nand U7023 (N_7023,N_6773,N_6295);
nand U7024 (N_7024,N_6565,N_6110);
or U7025 (N_7025,N_6413,N_6081);
nor U7026 (N_7026,N_6838,N_6592);
nand U7027 (N_7027,N_6461,N_6122);
and U7028 (N_7028,N_6183,N_6045);
and U7029 (N_7029,N_6414,N_6537);
or U7030 (N_7030,N_6111,N_6501);
nand U7031 (N_7031,N_6230,N_6806);
or U7032 (N_7032,N_6554,N_6860);
and U7033 (N_7033,N_6466,N_6904);
and U7034 (N_7034,N_6582,N_6388);
nor U7035 (N_7035,N_6865,N_6527);
and U7036 (N_7036,N_6758,N_6555);
nor U7037 (N_7037,N_6624,N_6812);
or U7038 (N_7038,N_6611,N_6159);
and U7039 (N_7039,N_6444,N_6158);
or U7040 (N_7040,N_6004,N_6930);
xnor U7041 (N_7041,N_6963,N_6757);
or U7042 (N_7042,N_6712,N_6177);
nand U7043 (N_7043,N_6902,N_6458);
or U7044 (N_7044,N_6182,N_6946);
or U7045 (N_7045,N_6002,N_6686);
and U7046 (N_7046,N_6240,N_6746);
and U7047 (N_7047,N_6108,N_6109);
or U7048 (N_7048,N_6630,N_6654);
and U7049 (N_7049,N_6416,N_6660);
or U7050 (N_7050,N_6628,N_6327);
xor U7051 (N_7051,N_6759,N_6368);
xor U7052 (N_7052,N_6538,N_6714);
nor U7053 (N_7053,N_6186,N_6745);
nor U7054 (N_7054,N_6222,N_6509);
or U7055 (N_7055,N_6672,N_6882);
nand U7056 (N_7056,N_6429,N_6154);
and U7057 (N_7057,N_6434,N_6959);
xor U7058 (N_7058,N_6581,N_6439);
xnor U7059 (N_7059,N_6023,N_6851);
nor U7060 (N_7060,N_6695,N_6528);
and U7061 (N_7061,N_6237,N_6995);
nor U7062 (N_7062,N_6141,N_6561);
nand U7063 (N_7063,N_6503,N_6929);
or U7064 (N_7064,N_6784,N_6477);
and U7065 (N_7065,N_6536,N_6329);
nor U7066 (N_7066,N_6417,N_6608);
and U7067 (N_7067,N_6793,N_6026);
nor U7068 (N_7068,N_6427,N_6489);
or U7069 (N_7069,N_6857,N_6917);
or U7070 (N_7070,N_6203,N_6966);
or U7071 (N_7071,N_6653,N_6078);
nand U7072 (N_7072,N_6722,N_6632);
nand U7073 (N_7073,N_6681,N_6209);
or U7074 (N_7074,N_6927,N_6409);
or U7075 (N_7075,N_6623,N_6188);
nor U7076 (N_7076,N_6175,N_6127);
or U7077 (N_7077,N_6522,N_6949);
or U7078 (N_7078,N_6598,N_6114);
nor U7079 (N_7079,N_6625,N_6768);
nand U7080 (N_7080,N_6832,N_6986);
nand U7081 (N_7081,N_6433,N_6000);
nor U7082 (N_7082,N_6303,N_6576);
xor U7083 (N_7083,N_6866,N_6506);
or U7084 (N_7084,N_6980,N_6039);
and U7085 (N_7085,N_6496,N_6853);
nand U7086 (N_7086,N_6559,N_6059);
or U7087 (N_7087,N_6150,N_6394);
or U7088 (N_7088,N_6063,N_6261);
or U7089 (N_7089,N_6666,N_6070);
xnor U7090 (N_7090,N_6631,N_6962);
and U7091 (N_7091,N_6890,N_6322);
xor U7092 (N_7092,N_6234,N_6622);
and U7093 (N_7093,N_6014,N_6820);
and U7094 (N_7094,N_6337,N_6316);
and U7095 (N_7095,N_6874,N_6541);
nand U7096 (N_7096,N_6618,N_6492);
and U7097 (N_7097,N_6025,N_6854);
nor U7098 (N_7098,N_6763,N_6104);
or U7099 (N_7099,N_6084,N_6192);
nor U7100 (N_7100,N_6066,N_6367);
nor U7101 (N_7101,N_6015,N_6574);
nor U7102 (N_7102,N_6391,N_6201);
or U7103 (N_7103,N_6934,N_6162);
nand U7104 (N_7104,N_6356,N_6479);
nor U7105 (N_7105,N_6494,N_6871);
or U7106 (N_7106,N_6258,N_6062);
or U7107 (N_7107,N_6021,N_6837);
or U7108 (N_7108,N_6969,N_6087);
xor U7109 (N_7109,N_6842,N_6055);
or U7110 (N_7110,N_6558,N_6397);
and U7111 (N_7111,N_6782,N_6487);
xnor U7112 (N_7112,N_6846,N_6795);
or U7113 (N_7113,N_6992,N_6291);
nand U7114 (N_7114,N_6245,N_6741);
and U7115 (N_7115,N_6221,N_6277);
xor U7116 (N_7116,N_6334,N_6484);
nand U7117 (N_7117,N_6613,N_6449);
and U7118 (N_7118,N_6824,N_6032);
nor U7119 (N_7119,N_6550,N_6580);
and U7120 (N_7120,N_6977,N_6844);
and U7121 (N_7121,N_6596,N_6923);
and U7122 (N_7122,N_6715,N_6885);
or U7123 (N_7123,N_6470,N_6423);
nor U7124 (N_7124,N_6553,N_6473);
nand U7125 (N_7125,N_6620,N_6199);
or U7126 (N_7126,N_6131,N_6048);
nor U7127 (N_7127,N_6785,N_6251);
nand U7128 (N_7128,N_6105,N_6691);
xnor U7129 (N_7129,N_6034,N_6914);
or U7130 (N_7130,N_6556,N_6442);
and U7131 (N_7131,N_6260,N_6732);
or U7132 (N_7132,N_6872,N_6140);
and U7133 (N_7133,N_6644,N_6614);
and U7134 (N_7134,N_6970,N_6119);
nor U7135 (N_7135,N_6074,N_6174);
and U7136 (N_7136,N_6249,N_6733);
or U7137 (N_7137,N_6826,N_6481);
and U7138 (N_7138,N_6121,N_6769);
and U7139 (N_7139,N_6223,N_6530);
nor U7140 (N_7140,N_6134,N_6410);
and U7141 (N_7141,N_6508,N_6560);
and U7142 (N_7142,N_6751,N_6462);
or U7143 (N_7143,N_6756,N_6577);
nor U7144 (N_7144,N_6279,N_6272);
nand U7145 (N_7145,N_6964,N_6373);
xnor U7146 (N_7146,N_6752,N_6340);
nand U7147 (N_7147,N_6798,N_6378);
or U7148 (N_7148,N_6856,N_6057);
and U7149 (N_7149,N_6950,N_6350);
or U7150 (N_7150,N_6876,N_6116);
or U7151 (N_7151,N_6094,N_6786);
or U7152 (N_7152,N_6886,N_6850);
xor U7153 (N_7153,N_6285,N_6266);
nor U7154 (N_7154,N_6597,N_6667);
or U7155 (N_7155,N_6248,N_6892);
nor U7156 (N_7156,N_6376,N_6369);
and U7157 (N_7157,N_6190,N_6478);
and U7158 (N_7158,N_6288,N_6586);
or U7159 (N_7159,N_6326,N_6859);
nand U7160 (N_7160,N_6009,N_6287);
and U7161 (N_7161,N_6901,N_6197);
or U7162 (N_7162,N_6713,N_6041);
nand U7163 (N_7163,N_6848,N_6728);
nand U7164 (N_7164,N_6130,N_6772);
nand U7165 (N_7165,N_6241,N_6475);
nor U7166 (N_7166,N_6309,N_6293);
nand U7167 (N_7167,N_6520,N_6379);
and U7168 (N_7168,N_6973,N_6879);
nand U7169 (N_7169,N_6424,N_6765);
nor U7170 (N_7170,N_6744,N_6339);
and U7171 (N_7171,N_6778,N_6435);
and U7172 (N_7172,N_6007,N_6431);
nand U7173 (N_7173,N_6767,N_6263);
nand U7174 (N_7174,N_6899,N_6357);
and U7175 (N_7175,N_6145,N_6402);
and U7176 (N_7176,N_6944,N_6583);
or U7177 (N_7177,N_6384,N_6552);
nor U7178 (N_7178,N_6286,N_6707);
nor U7179 (N_7179,N_6587,N_6079);
xnor U7180 (N_7180,N_6038,N_6775);
or U7181 (N_7181,N_6858,N_6148);
or U7182 (N_7182,N_6422,N_6562);
nor U7183 (N_7183,N_6155,N_6016);
or U7184 (N_7184,N_6210,N_6521);
or U7185 (N_7185,N_6485,N_6042);
nand U7186 (N_7186,N_6705,N_6090);
and U7187 (N_7187,N_6894,N_6983);
nand U7188 (N_7188,N_6067,N_6893);
xor U7189 (N_7189,N_6953,N_6954);
nand U7190 (N_7190,N_6493,N_6284);
nor U7191 (N_7191,N_6568,N_6227);
or U7192 (N_7192,N_6779,N_6801);
nand U7193 (N_7193,N_6701,N_6610);
and U7194 (N_7194,N_6697,N_6441);
and U7195 (N_7195,N_6430,N_6651);
nor U7196 (N_7196,N_6138,N_6979);
nor U7197 (N_7197,N_6703,N_6336);
nand U7198 (N_7198,N_6505,N_6688);
xor U7199 (N_7199,N_6957,N_6179);
or U7200 (N_7200,N_6276,N_6975);
or U7201 (N_7201,N_6510,N_6925);
nand U7202 (N_7202,N_6236,N_6107);
nor U7203 (N_7203,N_6264,N_6711);
or U7204 (N_7204,N_6564,N_6147);
and U7205 (N_7205,N_6684,N_6120);
and U7206 (N_7206,N_6377,N_6920);
nand U7207 (N_7207,N_6557,N_6952);
or U7208 (N_7208,N_6244,N_6810);
nand U7209 (N_7209,N_6198,N_6634);
nand U7210 (N_7210,N_6500,N_6319);
and U7211 (N_7211,N_6787,N_6513);
and U7212 (N_7212,N_6972,N_6019);
nor U7213 (N_7213,N_6152,N_6013);
nor U7214 (N_7214,N_6143,N_6621);
and U7215 (N_7215,N_6432,N_6867);
nand U7216 (N_7216,N_6821,N_6464);
xnor U7217 (N_7217,N_6076,N_6324);
nand U7218 (N_7218,N_6616,N_6807);
and U7219 (N_7219,N_6392,N_6495);
nand U7220 (N_7220,N_6095,N_6370);
nor U7221 (N_7221,N_6290,N_6948);
xnor U7222 (N_7222,N_6615,N_6551);
and U7223 (N_7223,N_6092,N_6774);
nand U7224 (N_7224,N_6217,N_6818);
nor U7225 (N_7225,N_6664,N_6990);
and U7226 (N_7226,N_6171,N_6135);
nand U7227 (N_7227,N_6005,N_6156);
or U7228 (N_7228,N_6659,N_6730);
and U7229 (N_7229,N_6643,N_6547);
xor U7230 (N_7230,N_6411,N_6106);
or U7231 (N_7231,N_6670,N_6839);
and U7232 (N_7232,N_6191,N_6678);
nor U7233 (N_7233,N_6897,N_6657);
xnor U7234 (N_7234,N_6870,N_6884);
nor U7235 (N_7235,N_6231,N_6233);
xnor U7236 (N_7236,N_6305,N_6069);
and U7237 (N_7237,N_6612,N_6663);
nand U7238 (N_7238,N_6447,N_6593);
nor U7239 (N_7239,N_6649,N_6180);
and U7240 (N_7240,N_6096,N_6993);
xnor U7241 (N_7241,N_6803,N_6709);
xnor U7242 (N_7242,N_6534,N_6457);
nor U7243 (N_7243,N_6566,N_6265);
or U7244 (N_7244,N_6542,N_6421);
and U7245 (N_7245,N_6931,N_6298);
nand U7246 (N_7246,N_6259,N_6989);
nand U7247 (N_7247,N_6671,N_6184);
and U7248 (N_7248,N_6700,N_6648);
nand U7249 (N_7249,N_6242,N_6679);
and U7250 (N_7250,N_6533,N_6900);
nor U7251 (N_7251,N_6082,N_6652);
nor U7252 (N_7252,N_6365,N_6910);
nand U7253 (N_7253,N_6304,N_6816);
nand U7254 (N_7254,N_6933,N_6283);
or U7255 (N_7255,N_6656,N_6735);
nor U7256 (N_7256,N_6073,N_6219);
and U7257 (N_7257,N_6737,N_6532);
nand U7258 (N_7258,N_6381,N_6861);
or U7259 (N_7259,N_6163,N_6908);
nor U7260 (N_7260,N_6777,N_6905);
or U7261 (N_7261,N_6804,N_6012);
nand U7262 (N_7262,N_6463,N_6633);
or U7263 (N_7263,N_6517,N_6525);
nand U7264 (N_7264,N_6301,N_6835);
nand U7265 (N_7265,N_6717,N_6888);
or U7266 (N_7266,N_6997,N_6022);
nor U7267 (N_7267,N_6407,N_6157);
nand U7268 (N_7268,N_6776,N_6205);
nor U7269 (N_7269,N_6575,N_6406);
nor U7270 (N_7270,N_6911,N_6988);
nor U7271 (N_7271,N_6352,N_6440);
xnor U7272 (N_7272,N_6307,N_6764);
nor U7273 (N_7273,N_6998,N_6640);
xor U7274 (N_7274,N_6142,N_6448);
nor U7275 (N_7275,N_6571,N_6702);
or U7276 (N_7276,N_6056,N_6708);
and U7277 (N_7277,N_6405,N_6602);
or U7278 (N_7278,N_6573,N_6828);
and U7279 (N_7279,N_6146,N_6468);
nand U7280 (N_7280,N_6178,N_6325);
nor U7281 (N_7281,N_6515,N_6987);
or U7282 (N_7282,N_6451,N_6491);
nand U7283 (N_7283,N_6252,N_6836);
nand U7284 (N_7284,N_6635,N_6315);
nand U7285 (N_7285,N_6945,N_6060);
or U7286 (N_7286,N_6172,N_6321);
and U7287 (N_7287,N_6723,N_6348);
xor U7288 (N_7288,N_6961,N_6743);
nand U7289 (N_7289,N_6788,N_6408);
or U7290 (N_7290,N_6212,N_6386);
nand U7291 (N_7291,N_6166,N_6229);
nand U7292 (N_7292,N_6124,N_6133);
and U7293 (N_7293,N_6418,N_6225);
nor U7294 (N_7294,N_6880,N_6830);
and U7295 (N_7295,N_6721,N_6010);
xor U7296 (N_7296,N_6097,N_6514);
or U7297 (N_7297,N_6875,N_6898);
and U7298 (N_7298,N_6465,N_6218);
and U7299 (N_7299,N_6289,N_6349);
nand U7300 (N_7300,N_6740,N_6941);
nand U7301 (N_7301,N_6694,N_6058);
nand U7302 (N_7302,N_6488,N_6051);
or U7303 (N_7303,N_6512,N_6976);
nand U7304 (N_7304,N_6086,N_6650);
nand U7305 (N_7305,N_6922,N_6794);
nand U7306 (N_7306,N_6877,N_6932);
or U7307 (N_7307,N_6578,N_6518);
or U7308 (N_7308,N_6690,N_6761);
and U7309 (N_7309,N_6359,N_6300);
or U7310 (N_7310,N_6061,N_6570);
nor U7311 (N_7311,N_6139,N_6661);
nand U7312 (N_7312,N_6499,N_6629);
nand U7313 (N_7313,N_6318,N_6841);
and U7314 (N_7314,N_6594,N_6030);
and U7315 (N_7315,N_6967,N_6200);
nand U7316 (N_7316,N_6294,N_6044);
or U7317 (N_7317,N_6165,N_6792);
or U7318 (N_7318,N_6254,N_6125);
and U7319 (N_7319,N_6668,N_6275);
and U7320 (N_7320,N_6590,N_6206);
nor U7321 (N_7321,N_6239,N_6207);
and U7322 (N_7322,N_6719,N_6641);
and U7323 (N_7323,N_6168,N_6805);
nor U7324 (N_7324,N_6358,N_6675);
nand U7325 (N_7325,N_6412,N_6589);
and U7326 (N_7326,N_6008,N_6226);
or U7327 (N_7327,N_6718,N_6049);
xor U7328 (N_7328,N_6372,N_6739);
or U7329 (N_7329,N_6683,N_6167);
or U7330 (N_7330,N_6313,N_6296);
nand U7331 (N_7331,N_6068,N_6585);
nand U7332 (N_7332,N_6991,N_6003);
nor U7333 (N_7333,N_6129,N_6863);
and U7334 (N_7334,N_6374,N_6437);
nor U7335 (N_7335,N_6364,N_6036);
or U7336 (N_7336,N_6789,N_6809);
or U7337 (N_7337,N_6891,N_6878);
or U7338 (N_7338,N_6760,N_6696);
xor U7339 (N_7339,N_6591,N_6999);
or U7340 (N_7340,N_6332,N_6445);
or U7341 (N_7341,N_6968,N_6033);
or U7342 (N_7342,N_6323,N_6627);
nor U7343 (N_7343,N_6943,N_6928);
and U7344 (N_7344,N_6452,N_6698);
and U7345 (N_7345,N_6539,N_6831);
nor U7346 (N_7346,N_6726,N_6843);
nand U7347 (N_7347,N_6028,N_6011);
nand U7348 (N_7348,N_6543,N_6873);
and U7349 (N_7349,N_6742,N_6791);
or U7350 (N_7350,N_6482,N_6799);
xor U7351 (N_7351,N_6687,N_6396);
and U7352 (N_7352,N_6662,N_6921);
nand U7353 (N_7353,N_6647,N_6375);
xor U7354 (N_7354,N_6256,N_6238);
nand U7355 (N_7355,N_6604,N_6639);
and U7356 (N_7356,N_6729,N_6269);
and U7357 (N_7357,N_6755,N_6747);
xor U7358 (N_7358,N_6619,N_6366);
xor U7359 (N_7359,N_6813,N_6748);
nor U7360 (N_7360,N_6869,N_6415);
nor U7361 (N_7361,N_6796,N_6382);
and U7362 (N_7362,N_6247,N_6354);
nand U7363 (N_7363,N_6919,N_6136);
nand U7364 (N_7364,N_6338,N_6312);
nand U7365 (N_7365,N_6161,N_6404);
xnor U7366 (N_7366,N_6371,N_6658);
or U7367 (N_7367,N_6540,N_6689);
and U7368 (N_7368,N_6642,N_6669);
xor U7369 (N_7369,N_6393,N_6545);
nand U7370 (N_7370,N_6895,N_6706);
nor U7371 (N_7371,N_6502,N_6438);
nor U7372 (N_7372,N_6335,N_6486);
nand U7373 (N_7373,N_6909,N_6924);
nand U7374 (N_7374,N_6645,N_6072);
and U7375 (N_7375,N_6262,N_6117);
and U7376 (N_7376,N_6308,N_6144);
or U7377 (N_7377,N_6232,N_6310);
nand U7378 (N_7378,N_6753,N_6523);
and U7379 (N_7379,N_6017,N_6535);
nand U7380 (N_7380,N_6250,N_6781);
and U7381 (N_7381,N_6194,N_6020);
nand U7382 (N_7382,N_6345,N_6398);
nor U7383 (N_7383,N_6214,N_6454);
and U7384 (N_7384,N_6280,N_6720);
nand U7385 (N_7385,N_6137,N_6815);
nor U7386 (N_7386,N_6965,N_6896);
and U7387 (N_7387,N_6029,N_6926);
or U7388 (N_7388,N_6189,N_6460);
or U7389 (N_7389,N_6385,N_6985);
and U7390 (N_7390,N_6754,N_6617);
and U7391 (N_7391,N_6951,N_6149);
or U7392 (N_7392,N_6224,N_6903);
or U7393 (N_7393,N_6603,N_6204);
nand U7394 (N_7394,N_6071,N_6202);
nand U7395 (N_7395,N_6693,N_6845);
and U7396 (N_7396,N_6299,N_6834);
nor U7397 (N_7397,N_6089,N_6827);
nor U7398 (N_7398,N_6347,N_6646);
xor U7399 (N_7399,N_6099,N_6947);
or U7400 (N_7400,N_6292,N_6749);
nor U7401 (N_7401,N_6243,N_6680);
and U7402 (N_7402,N_6800,N_6220);
nor U7403 (N_7403,N_6390,N_6027);
or U7404 (N_7404,N_6955,N_6636);
and U7405 (N_7405,N_6588,N_6906);
nor U7406 (N_7406,N_6053,N_6333);
nand U7407 (N_7407,N_6710,N_6363);
xor U7408 (N_7408,N_6734,N_6883);
nor U7409 (N_7409,N_6637,N_6052);
or U7410 (N_7410,N_6077,N_6823);
xor U7411 (N_7411,N_6497,N_6193);
or U7412 (N_7412,N_6088,N_6126);
and U7413 (N_7413,N_6436,N_6297);
or U7414 (N_7414,N_6054,N_6783);
nor U7415 (N_7415,N_6790,N_6387);
xnor U7416 (N_7416,N_6426,N_6196);
nand U7417 (N_7417,N_6982,N_6380);
nor U7418 (N_7418,N_6403,N_6504);
and U7419 (N_7419,N_6270,N_6001);
and U7420 (N_7420,N_6864,N_6083);
nand U7421 (N_7421,N_6994,N_6609);
nand U7422 (N_7422,N_6123,N_6164);
and U7423 (N_7423,N_6101,N_6228);
nand U7424 (N_7424,N_6724,N_6544);
nor U7425 (N_7425,N_6257,N_6361);
and U7426 (N_7426,N_6050,N_6456);
xor U7427 (N_7427,N_6814,N_6213);
or U7428 (N_7428,N_6132,N_6974);
and U7429 (N_7429,N_6211,N_6673);
xnor U7430 (N_7430,N_6852,N_6731);
nand U7431 (N_7431,N_6692,N_6546);
and U7432 (N_7432,N_6455,N_6531);
nand U7433 (N_7433,N_6064,N_6511);
xor U7434 (N_7434,N_6353,N_6018);
nor U7435 (N_7435,N_6677,N_6330);
or U7436 (N_7436,N_6770,N_6476);
xor U7437 (N_7437,N_6939,N_6889);
and U7438 (N_7438,N_6006,N_6868);
nor U7439 (N_7439,N_6936,N_6549);
nor U7440 (N_7440,N_6195,N_6916);
nor U7441 (N_7441,N_6040,N_6780);
nor U7442 (N_7442,N_6762,N_6599);
and U7443 (N_7443,N_6401,N_6419);
nand U7444 (N_7444,N_6153,N_6483);
nand U7445 (N_7445,N_6043,N_6080);
nand U7446 (N_7446,N_6113,N_6736);
nand U7447 (N_7447,N_6459,N_6847);
nor U7448 (N_7448,N_6024,N_6956);
and U7449 (N_7449,N_6797,N_6065);
nand U7450 (N_7450,N_6085,N_6173);
and U7451 (N_7451,N_6524,N_6268);
nand U7452 (N_7452,N_6725,N_6978);
nand U7453 (N_7453,N_6355,N_6607);
or U7454 (N_7454,N_6840,N_6601);
xor U7455 (N_7455,N_6467,N_6819);
and U7456 (N_7456,N_6395,N_6399);
nand U7457 (N_7457,N_6035,N_6169);
or U7458 (N_7458,N_6311,N_6935);
nand U7459 (N_7459,N_6185,N_6605);
and U7460 (N_7460,N_6519,N_6802);
nor U7461 (N_7461,N_6958,N_6699);
or U7462 (N_7462,N_6428,N_6115);
and U7463 (N_7463,N_6674,N_6771);
nand U7464 (N_7464,N_6472,N_6037);
xor U7465 (N_7465,N_6446,N_6267);
and U7466 (N_7466,N_6093,N_6274);
and U7467 (N_7467,N_6128,N_6940);
xnor U7468 (N_7468,N_6849,N_6606);
or U7469 (N_7469,N_6548,N_6389);
xor U7470 (N_7470,N_6453,N_6727);
or U7471 (N_7471,N_6563,N_6750);
nor U7472 (N_7472,N_6984,N_6937);
nand U7473 (N_7473,N_6685,N_6960);
and U7474 (N_7474,N_6716,N_6425);
or U7475 (N_7475,N_6278,N_6046);
nand U7476 (N_7476,N_6655,N_6595);
or U7477 (N_7477,N_6665,N_6170);
or U7478 (N_7478,N_6360,N_6569);
xnor U7479 (N_7479,N_6474,N_6102);
nor U7480 (N_7480,N_6829,N_6971);
nor U7481 (N_7481,N_6450,N_6579);
nor U7482 (N_7482,N_6343,N_6281);
nand U7483 (N_7483,N_6282,N_6075);
nor U7484 (N_7484,N_6471,N_6215);
or U7485 (N_7485,N_6833,N_6600);
nand U7486 (N_7486,N_6181,N_6704);
and U7487 (N_7487,N_6317,N_6346);
nand U7488 (N_7488,N_6996,N_6383);
or U7489 (N_7489,N_6091,N_6469);
or U7490 (N_7490,N_6320,N_6351);
and U7491 (N_7491,N_6328,N_6103);
xnor U7492 (N_7492,N_6098,N_6938);
or U7493 (N_7493,N_6638,N_6306);
nand U7494 (N_7494,N_6176,N_6825);
or U7495 (N_7495,N_6216,N_6151);
and U7496 (N_7496,N_6516,N_6567);
and U7497 (N_7497,N_6255,N_6584);
nand U7498 (N_7498,N_6341,N_6676);
or U7499 (N_7499,N_6887,N_6811);
or U7500 (N_7500,N_6380,N_6838);
and U7501 (N_7501,N_6330,N_6780);
or U7502 (N_7502,N_6112,N_6006);
and U7503 (N_7503,N_6388,N_6959);
and U7504 (N_7504,N_6384,N_6041);
nand U7505 (N_7505,N_6503,N_6711);
or U7506 (N_7506,N_6650,N_6670);
nor U7507 (N_7507,N_6146,N_6688);
nor U7508 (N_7508,N_6423,N_6820);
and U7509 (N_7509,N_6817,N_6150);
nor U7510 (N_7510,N_6188,N_6789);
and U7511 (N_7511,N_6764,N_6719);
nor U7512 (N_7512,N_6081,N_6950);
and U7513 (N_7513,N_6806,N_6901);
xnor U7514 (N_7514,N_6171,N_6082);
xnor U7515 (N_7515,N_6148,N_6984);
and U7516 (N_7516,N_6527,N_6511);
nor U7517 (N_7517,N_6987,N_6908);
nor U7518 (N_7518,N_6868,N_6017);
xor U7519 (N_7519,N_6500,N_6823);
xor U7520 (N_7520,N_6723,N_6750);
nor U7521 (N_7521,N_6999,N_6421);
nand U7522 (N_7522,N_6051,N_6058);
nor U7523 (N_7523,N_6675,N_6327);
xnor U7524 (N_7524,N_6914,N_6758);
xnor U7525 (N_7525,N_6283,N_6964);
or U7526 (N_7526,N_6954,N_6883);
and U7527 (N_7527,N_6049,N_6928);
nand U7528 (N_7528,N_6504,N_6077);
nand U7529 (N_7529,N_6043,N_6692);
nand U7530 (N_7530,N_6885,N_6033);
nor U7531 (N_7531,N_6859,N_6644);
and U7532 (N_7532,N_6675,N_6621);
nand U7533 (N_7533,N_6105,N_6131);
xnor U7534 (N_7534,N_6440,N_6377);
nor U7535 (N_7535,N_6207,N_6126);
xnor U7536 (N_7536,N_6619,N_6327);
or U7537 (N_7537,N_6382,N_6592);
nand U7538 (N_7538,N_6564,N_6755);
nand U7539 (N_7539,N_6628,N_6274);
and U7540 (N_7540,N_6358,N_6786);
nand U7541 (N_7541,N_6979,N_6261);
nand U7542 (N_7542,N_6941,N_6254);
nand U7543 (N_7543,N_6249,N_6358);
nand U7544 (N_7544,N_6964,N_6456);
nand U7545 (N_7545,N_6429,N_6042);
nand U7546 (N_7546,N_6445,N_6032);
or U7547 (N_7547,N_6455,N_6242);
or U7548 (N_7548,N_6259,N_6398);
nand U7549 (N_7549,N_6780,N_6092);
nor U7550 (N_7550,N_6577,N_6525);
nand U7551 (N_7551,N_6394,N_6928);
nor U7552 (N_7552,N_6897,N_6492);
nor U7553 (N_7553,N_6141,N_6612);
nand U7554 (N_7554,N_6578,N_6234);
and U7555 (N_7555,N_6751,N_6028);
nor U7556 (N_7556,N_6657,N_6292);
or U7557 (N_7557,N_6537,N_6699);
or U7558 (N_7558,N_6367,N_6721);
and U7559 (N_7559,N_6959,N_6775);
and U7560 (N_7560,N_6094,N_6531);
and U7561 (N_7561,N_6649,N_6851);
nor U7562 (N_7562,N_6004,N_6664);
nand U7563 (N_7563,N_6441,N_6370);
xnor U7564 (N_7564,N_6876,N_6544);
nor U7565 (N_7565,N_6015,N_6488);
nor U7566 (N_7566,N_6153,N_6760);
nand U7567 (N_7567,N_6315,N_6476);
or U7568 (N_7568,N_6131,N_6726);
nand U7569 (N_7569,N_6239,N_6636);
or U7570 (N_7570,N_6322,N_6380);
nor U7571 (N_7571,N_6145,N_6001);
or U7572 (N_7572,N_6941,N_6142);
or U7573 (N_7573,N_6907,N_6756);
nand U7574 (N_7574,N_6612,N_6914);
nand U7575 (N_7575,N_6268,N_6551);
and U7576 (N_7576,N_6776,N_6600);
or U7577 (N_7577,N_6276,N_6554);
and U7578 (N_7578,N_6396,N_6143);
nand U7579 (N_7579,N_6625,N_6475);
nand U7580 (N_7580,N_6157,N_6868);
nand U7581 (N_7581,N_6548,N_6675);
nand U7582 (N_7582,N_6095,N_6941);
nand U7583 (N_7583,N_6739,N_6839);
xnor U7584 (N_7584,N_6581,N_6246);
and U7585 (N_7585,N_6519,N_6745);
xnor U7586 (N_7586,N_6201,N_6636);
nand U7587 (N_7587,N_6362,N_6279);
or U7588 (N_7588,N_6112,N_6945);
or U7589 (N_7589,N_6583,N_6435);
or U7590 (N_7590,N_6250,N_6611);
and U7591 (N_7591,N_6169,N_6633);
and U7592 (N_7592,N_6380,N_6456);
nor U7593 (N_7593,N_6656,N_6579);
xnor U7594 (N_7594,N_6852,N_6346);
nor U7595 (N_7595,N_6779,N_6087);
and U7596 (N_7596,N_6449,N_6593);
xor U7597 (N_7597,N_6297,N_6998);
nor U7598 (N_7598,N_6670,N_6775);
xor U7599 (N_7599,N_6685,N_6146);
nand U7600 (N_7600,N_6283,N_6887);
and U7601 (N_7601,N_6691,N_6081);
or U7602 (N_7602,N_6579,N_6814);
nand U7603 (N_7603,N_6784,N_6546);
nor U7604 (N_7604,N_6259,N_6460);
nor U7605 (N_7605,N_6622,N_6282);
nor U7606 (N_7606,N_6284,N_6015);
nand U7607 (N_7607,N_6571,N_6814);
xnor U7608 (N_7608,N_6802,N_6586);
and U7609 (N_7609,N_6208,N_6516);
or U7610 (N_7610,N_6086,N_6006);
xor U7611 (N_7611,N_6124,N_6275);
and U7612 (N_7612,N_6503,N_6261);
and U7613 (N_7613,N_6576,N_6209);
nand U7614 (N_7614,N_6938,N_6126);
and U7615 (N_7615,N_6590,N_6075);
xnor U7616 (N_7616,N_6634,N_6421);
xnor U7617 (N_7617,N_6804,N_6896);
and U7618 (N_7618,N_6434,N_6362);
or U7619 (N_7619,N_6357,N_6851);
or U7620 (N_7620,N_6776,N_6079);
and U7621 (N_7621,N_6469,N_6680);
nor U7622 (N_7622,N_6238,N_6205);
and U7623 (N_7623,N_6800,N_6564);
and U7624 (N_7624,N_6024,N_6242);
and U7625 (N_7625,N_6443,N_6459);
and U7626 (N_7626,N_6440,N_6295);
and U7627 (N_7627,N_6911,N_6608);
nor U7628 (N_7628,N_6390,N_6466);
nand U7629 (N_7629,N_6438,N_6367);
nand U7630 (N_7630,N_6975,N_6312);
nand U7631 (N_7631,N_6834,N_6489);
or U7632 (N_7632,N_6422,N_6237);
xnor U7633 (N_7633,N_6121,N_6302);
nand U7634 (N_7634,N_6161,N_6000);
xnor U7635 (N_7635,N_6563,N_6014);
nor U7636 (N_7636,N_6782,N_6519);
nand U7637 (N_7637,N_6654,N_6887);
or U7638 (N_7638,N_6625,N_6718);
nor U7639 (N_7639,N_6848,N_6807);
and U7640 (N_7640,N_6813,N_6948);
and U7641 (N_7641,N_6071,N_6404);
xnor U7642 (N_7642,N_6422,N_6401);
or U7643 (N_7643,N_6307,N_6869);
nor U7644 (N_7644,N_6906,N_6824);
nand U7645 (N_7645,N_6335,N_6688);
xor U7646 (N_7646,N_6184,N_6960);
or U7647 (N_7647,N_6423,N_6716);
and U7648 (N_7648,N_6344,N_6366);
or U7649 (N_7649,N_6903,N_6400);
xor U7650 (N_7650,N_6466,N_6163);
nand U7651 (N_7651,N_6776,N_6707);
nor U7652 (N_7652,N_6751,N_6752);
nand U7653 (N_7653,N_6388,N_6548);
nand U7654 (N_7654,N_6810,N_6677);
and U7655 (N_7655,N_6170,N_6509);
nand U7656 (N_7656,N_6720,N_6920);
nand U7657 (N_7657,N_6587,N_6985);
or U7658 (N_7658,N_6005,N_6678);
or U7659 (N_7659,N_6857,N_6753);
nand U7660 (N_7660,N_6067,N_6630);
and U7661 (N_7661,N_6113,N_6887);
nor U7662 (N_7662,N_6719,N_6184);
xnor U7663 (N_7663,N_6858,N_6618);
nor U7664 (N_7664,N_6125,N_6571);
nor U7665 (N_7665,N_6060,N_6385);
or U7666 (N_7666,N_6717,N_6867);
or U7667 (N_7667,N_6960,N_6610);
and U7668 (N_7668,N_6372,N_6706);
or U7669 (N_7669,N_6845,N_6700);
nor U7670 (N_7670,N_6991,N_6916);
nand U7671 (N_7671,N_6242,N_6548);
nand U7672 (N_7672,N_6477,N_6792);
and U7673 (N_7673,N_6865,N_6795);
nand U7674 (N_7674,N_6043,N_6195);
nor U7675 (N_7675,N_6575,N_6146);
and U7676 (N_7676,N_6689,N_6060);
nor U7677 (N_7677,N_6886,N_6940);
and U7678 (N_7678,N_6149,N_6061);
xor U7679 (N_7679,N_6679,N_6091);
xor U7680 (N_7680,N_6942,N_6533);
or U7681 (N_7681,N_6193,N_6061);
xor U7682 (N_7682,N_6421,N_6133);
and U7683 (N_7683,N_6847,N_6169);
or U7684 (N_7684,N_6544,N_6299);
nand U7685 (N_7685,N_6846,N_6967);
or U7686 (N_7686,N_6749,N_6829);
nor U7687 (N_7687,N_6857,N_6289);
or U7688 (N_7688,N_6575,N_6817);
or U7689 (N_7689,N_6357,N_6464);
xor U7690 (N_7690,N_6124,N_6465);
xor U7691 (N_7691,N_6179,N_6827);
nor U7692 (N_7692,N_6094,N_6047);
nand U7693 (N_7693,N_6991,N_6168);
or U7694 (N_7694,N_6259,N_6900);
and U7695 (N_7695,N_6609,N_6133);
or U7696 (N_7696,N_6594,N_6097);
nand U7697 (N_7697,N_6635,N_6645);
or U7698 (N_7698,N_6825,N_6838);
or U7699 (N_7699,N_6363,N_6995);
nor U7700 (N_7700,N_6594,N_6406);
or U7701 (N_7701,N_6521,N_6913);
nor U7702 (N_7702,N_6176,N_6550);
or U7703 (N_7703,N_6397,N_6606);
or U7704 (N_7704,N_6192,N_6391);
or U7705 (N_7705,N_6525,N_6785);
xor U7706 (N_7706,N_6635,N_6613);
nand U7707 (N_7707,N_6112,N_6927);
and U7708 (N_7708,N_6711,N_6037);
xor U7709 (N_7709,N_6187,N_6628);
nor U7710 (N_7710,N_6547,N_6483);
nand U7711 (N_7711,N_6982,N_6482);
and U7712 (N_7712,N_6714,N_6094);
or U7713 (N_7713,N_6647,N_6585);
nand U7714 (N_7714,N_6287,N_6363);
and U7715 (N_7715,N_6566,N_6558);
and U7716 (N_7716,N_6848,N_6077);
nor U7717 (N_7717,N_6655,N_6037);
nor U7718 (N_7718,N_6677,N_6968);
nand U7719 (N_7719,N_6687,N_6036);
and U7720 (N_7720,N_6588,N_6758);
nand U7721 (N_7721,N_6253,N_6218);
or U7722 (N_7722,N_6262,N_6478);
nand U7723 (N_7723,N_6126,N_6637);
or U7724 (N_7724,N_6405,N_6558);
and U7725 (N_7725,N_6486,N_6305);
or U7726 (N_7726,N_6200,N_6563);
and U7727 (N_7727,N_6750,N_6618);
xor U7728 (N_7728,N_6324,N_6120);
and U7729 (N_7729,N_6430,N_6597);
nor U7730 (N_7730,N_6181,N_6451);
or U7731 (N_7731,N_6562,N_6744);
or U7732 (N_7732,N_6047,N_6569);
nand U7733 (N_7733,N_6359,N_6056);
and U7734 (N_7734,N_6740,N_6328);
or U7735 (N_7735,N_6571,N_6022);
or U7736 (N_7736,N_6724,N_6489);
and U7737 (N_7737,N_6873,N_6733);
or U7738 (N_7738,N_6441,N_6231);
nand U7739 (N_7739,N_6500,N_6714);
nand U7740 (N_7740,N_6581,N_6629);
and U7741 (N_7741,N_6969,N_6262);
or U7742 (N_7742,N_6950,N_6034);
or U7743 (N_7743,N_6924,N_6448);
and U7744 (N_7744,N_6320,N_6802);
and U7745 (N_7745,N_6751,N_6840);
nand U7746 (N_7746,N_6603,N_6067);
nand U7747 (N_7747,N_6298,N_6935);
or U7748 (N_7748,N_6010,N_6295);
and U7749 (N_7749,N_6793,N_6511);
xnor U7750 (N_7750,N_6539,N_6719);
nand U7751 (N_7751,N_6194,N_6180);
or U7752 (N_7752,N_6651,N_6747);
or U7753 (N_7753,N_6118,N_6207);
or U7754 (N_7754,N_6124,N_6347);
nand U7755 (N_7755,N_6061,N_6815);
xnor U7756 (N_7756,N_6334,N_6858);
nand U7757 (N_7757,N_6172,N_6741);
nor U7758 (N_7758,N_6103,N_6547);
or U7759 (N_7759,N_6246,N_6031);
nor U7760 (N_7760,N_6453,N_6704);
nor U7761 (N_7761,N_6238,N_6654);
nand U7762 (N_7762,N_6568,N_6592);
nor U7763 (N_7763,N_6172,N_6807);
nand U7764 (N_7764,N_6511,N_6924);
nand U7765 (N_7765,N_6893,N_6600);
nand U7766 (N_7766,N_6746,N_6380);
nand U7767 (N_7767,N_6911,N_6133);
and U7768 (N_7768,N_6826,N_6104);
nor U7769 (N_7769,N_6454,N_6699);
nor U7770 (N_7770,N_6831,N_6540);
nor U7771 (N_7771,N_6940,N_6397);
nor U7772 (N_7772,N_6134,N_6592);
and U7773 (N_7773,N_6073,N_6685);
or U7774 (N_7774,N_6818,N_6776);
nor U7775 (N_7775,N_6887,N_6525);
and U7776 (N_7776,N_6672,N_6148);
or U7777 (N_7777,N_6980,N_6055);
nand U7778 (N_7778,N_6842,N_6985);
nor U7779 (N_7779,N_6849,N_6120);
xor U7780 (N_7780,N_6733,N_6905);
or U7781 (N_7781,N_6634,N_6650);
or U7782 (N_7782,N_6037,N_6102);
or U7783 (N_7783,N_6448,N_6720);
and U7784 (N_7784,N_6013,N_6714);
xor U7785 (N_7785,N_6484,N_6102);
nor U7786 (N_7786,N_6319,N_6022);
xnor U7787 (N_7787,N_6213,N_6872);
nand U7788 (N_7788,N_6491,N_6626);
xnor U7789 (N_7789,N_6347,N_6267);
nor U7790 (N_7790,N_6863,N_6182);
nand U7791 (N_7791,N_6796,N_6095);
xor U7792 (N_7792,N_6216,N_6518);
xnor U7793 (N_7793,N_6475,N_6031);
nand U7794 (N_7794,N_6985,N_6271);
and U7795 (N_7795,N_6626,N_6148);
nand U7796 (N_7796,N_6634,N_6332);
nand U7797 (N_7797,N_6467,N_6025);
and U7798 (N_7798,N_6023,N_6073);
xnor U7799 (N_7799,N_6772,N_6919);
or U7800 (N_7800,N_6701,N_6474);
or U7801 (N_7801,N_6496,N_6577);
and U7802 (N_7802,N_6290,N_6468);
or U7803 (N_7803,N_6016,N_6028);
nand U7804 (N_7804,N_6606,N_6148);
nor U7805 (N_7805,N_6456,N_6066);
nand U7806 (N_7806,N_6299,N_6310);
and U7807 (N_7807,N_6745,N_6828);
nor U7808 (N_7808,N_6894,N_6818);
xor U7809 (N_7809,N_6565,N_6220);
or U7810 (N_7810,N_6038,N_6813);
nand U7811 (N_7811,N_6089,N_6672);
and U7812 (N_7812,N_6749,N_6093);
nor U7813 (N_7813,N_6144,N_6787);
or U7814 (N_7814,N_6343,N_6026);
or U7815 (N_7815,N_6294,N_6914);
xor U7816 (N_7816,N_6677,N_6287);
nand U7817 (N_7817,N_6644,N_6103);
or U7818 (N_7818,N_6432,N_6378);
nand U7819 (N_7819,N_6649,N_6086);
xnor U7820 (N_7820,N_6316,N_6395);
and U7821 (N_7821,N_6657,N_6100);
nor U7822 (N_7822,N_6941,N_6479);
xor U7823 (N_7823,N_6444,N_6321);
nor U7824 (N_7824,N_6287,N_6452);
nand U7825 (N_7825,N_6266,N_6486);
xor U7826 (N_7826,N_6817,N_6785);
or U7827 (N_7827,N_6589,N_6790);
nand U7828 (N_7828,N_6179,N_6089);
and U7829 (N_7829,N_6306,N_6129);
or U7830 (N_7830,N_6263,N_6200);
nand U7831 (N_7831,N_6799,N_6854);
and U7832 (N_7832,N_6013,N_6964);
nand U7833 (N_7833,N_6739,N_6746);
nand U7834 (N_7834,N_6674,N_6511);
xnor U7835 (N_7835,N_6970,N_6441);
nand U7836 (N_7836,N_6475,N_6310);
xor U7837 (N_7837,N_6948,N_6996);
or U7838 (N_7838,N_6826,N_6723);
or U7839 (N_7839,N_6995,N_6520);
nand U7840 (N_7840,N_6037,N_6010);
nand U7841 (N_7841,N_6306,N_6805);
nand U7842 (N_7842,N_6686,N_6064);
and U7843 (N_7843,N_6678,N_6831);
nor U7844 (N_7844,N_6848,N_6925);
and U7845 (N_7845,N_6643,N_6819);
or U7846 (N_7846,N_6290,N_6821);
nor U7847 (N_7847,N_6993,N_6726);
nand U7848 (N_7848,N_6910,N_6991);
xnor U7849 (N_7849,N_6829,N_6574);
and U7850 (N_7850,N_6097,N_6592);
nand U7851 (N_7851,N_6071,N_6507);
nand U7852 (N_7852,N_6609,N_6166);
or U7853 (N_7853,N_6812,N_6691);
and U7854 (N_7854,N_6569,N_6936);
xnor U7855 (N_7855,N_6911,N_6828);
and U7856 (N_7856,N_6513,N_6239);
or U7857 (N_7857,N_6626,N_6445);
nand U7858 (N_7858,N_6466,N_6542);
xnor U7859 (N_7859,N_6461,N_6745);
nor U7860 (N_7860,N_6327,N_6284);
nor U7861 (N_7861,N_6189,N_6464);
nor U7862 (N_7862,N_6281,N_6017);
and U7863 (N_7863,N_6676,N_6876);
nand U7864 (N_7864,N_6128,N_6212);
nor U7865 (N_7865,N_6086,N_6019);
nor U7866 (N_7866,N_6032,N_6120);
and U7867 (N_7867,N_6696,N_6263);
or U7868 (N_7868,N_6767,N_6251);
nor U7869 (N_7869,N_6012,N_6780);
or U7870 (N_7870,N_6048,N_6694);
and U7871 (N_7871,N_6105,N_6464);
or U7872 (N_7872,N_6764,N_6644);
xor U7873 (N_7873,N_6499,N_6259);
xor U7874 (N_7874,N_6453,N_6345);
nor U7875 (N_7875,N_6551,N_6456);
nand U7876 (N_7876,N_6975,N_6177);
nand U7877 (N_7877,N_6161,N_6321);
and U7878 (N_7878,N_6636,N_6718);
nor U7879 (N_7879,N_6600,N_6377);
nor U7880 (N_7880,N_6394,N_6583);
nor U7881 (N_7881,N_6830,N_6407);
nand U7882 (N_7882,N_6749,N_6972);
and U7883 (N_7883,N_6259,N_6022);
and U7884 (N_7884,N_6693,N_6409);
and U7885 (N_7885,N_6912,N_6805);
or U7886 (N_7886,N_6256,N_6336);
and U7887 (N_7887,N_6580,N_6094);
xnor U7888 (N_7888,N_6177,N_6447);
and U7889 (N_7889,N_6397,N_6774);
nand U7890 (N_7890,N_6361,N_6528);
and U7891 (N_7891,N_6546,N_6246);
and U7892 (N_7892,N_6578,N_6637);
and U7893 (N_7893,N_6456,N_6526);
or U7894 (N_7894,N_6283,N_6214);
xnor U7895 (N_7895,N_6569,N_6349);
nor U7896 (N_7896,N_6706,N_6743);
or U7897 (N_7897,N_6588,N_6004);
and U7898 (N_7898,N_6463,N_6957);
nor U7899 (N_7899,N_6514,N_6363);
or U7900 (N_7900,N_6459,N_6931);
nor U7901 (N_7901,N_6830,N_6353);
and U7902 (N_7902,N_6444,N_6234);
or U7903 (N_7903,N_6620,N_6059);
or U7904 (N_7904,N_6169,N_6929);
xor U7905 (N_7905,N_6564,N_6071);
nor U7906 (N_7906,N_6886,N_6333);
nor U7907 (N_7907,N_6332,N_6108);
nand U7908 (N_7908,N_6178,N_6442);
nand U7909 (N_7909,N_6941,N_6743);
nor U7910 (N_7910,N_6074,N_6786);
or U7911 (N_7911,N_6967,N_6008);
and U7912 (N_7912,N_6712,N_6277);
nor U7913 (N_7913,N_6150,N_6504);
or U7914 (N_7914,N_6523,N_6740);
nand U7915 (N_7915,N_6678,N_6021);
xnor U7916 (N_7916,N_6602,N_6766);
and U7917 (N_7917,N_6940,N_6546);
and U7918 (N_7918,N_6967,N_6607);
or U7919 (N_7919,N_6572,N_6841);
xor U7920 (N_7920,N_6789,N_6579);
and U7921 (N_7921,N_6464,N_6979);
or U7922 (N_7922,N_6015,N_6853);
nand U7923 (N_7923,N_6654,N_6218);
and U7924 (N_7924,N_6077,N_6630);
nand U7925 (N_7925,N_6876,N_6805);
and U7926 (N_7926,N_6701,N_6295);
or U7927 (N_7927,N_6981,N_6444);
nor U7928 (N_7928,N_6143,N_6095);
and U7929 (N_7929,N_6088,N_6635);
or U7930 (N_7930,N_6391,N_6433);
or U7931 (N_7931,N_6380,N_6855);
nand U7932 (N_7932,N_6966,N_6383);
or U7933 (N_7933,N_6196,N_6643);
xnor U7934 (N_7934,N_6572,N_6281);
and U7935 (N_7935,N_6079,N_6456);
nor U7936 (N_7936,N_6740,N_6228);
nor U7937 (N_7937,N_6890,N_6310);
nor U7938 (N_7938,N_6621,N_6230);
xor U7939 (N_7939,N_6378,N_6921);
nor U7940 (N_7940,N_6056,N_6136);
nand U7941 (N_7941,N_6442,N_6160);
nand U7942 (N_7942,N_6036,N_6705);
xor U7943 (N_7943,N_6739,N_6950);
and U7944 (N_7944,N_6559,N_6712);
nand U7945 (N_7945,N_6391,N_6954);
xnor U7946 (N_7946,N_6779,N_6800);
or U7947 (N_7947,N_6312,N_6672);
or U7948 (N_7948,N_6807,N_6163);
or U7949 (N_7949,N_6436,N_6755);
nand U7950 (N_7950,N_6444,N_6419);
nand U7951 (N_7951,N_6260,N_6355);
or U7952 (N_7952,N_6059,N_6853);
or U7953 (N_7953,N_6064,N_6515);
nor U7954 (N_7954,N_6109,N_6503);
nor U7955 (N_7955,N_6560,N_6862);
or U7956 (N_7956,N_6697,N_6790);
or U7957 (N_7957,N_6722,N_6068);
and U7958 (N_7958,N_6450,N_6580);
and U7959 (N_7959,N_6087,N_6473);
or U7960 (N_7960,N_6287,N_6170);
and U7961 (N_7961,N_6401,N_6812);
nor U7962 (N_7962,N_6600,N_6421);
nand U7963 (N_7963,N_6021,N_6034);
xnor U7964 (N_7964,N_6509,N_6379);
nor U7965 (N_7965,N_6321,N_6903);
nand U7966 (N_7966,N_6991,N_6297);
nor U7967 (N_7967,N_6018,N_6617);
and U7968 (N_7968,N_6064,N_6902);
nand U7969 (N_7969,N_6317,N_6598);
xor U7970 (N_7970,N_6085,N_6693);
nor U7971 (N_7971,N_6256,N_6420);
nor U7972 (N_7972,N_6053,N_6836);
or U7973 (N_7973,N_6057,N_6396);
nand U7974 (N_7974,N_6132,N_6290);
nor U7975 (N_7975,N_6075,N_6555);
or U7976 (N_7976,N_6794,N_6515);
and U7977 (N_7977,N_6122,N_6164);
and U7978 (N_7978,N_6184,N_6170);
xnor U7979 (N_7979,N_6105,N_6785);
and U7980 (N_7980,N_6649,N_6521);
nor U7981 (N_7981,N_6396,N_6974);
or U7982 (N_7982,N_6869,N_6288);
and U7983 (N_7983,N_6107,N_6010);
and U7984 (N_7984,N_6445,N_6813);
and U7985 (N_7985,N_6150,N_6280);
nor U7986 (N_7986,N_6911,N_6565);
and U7987 (N_7987,N_6801,N_6968);
and U7988 (N_7988,N_6377,N_6551);
nand U7989 (N_7989,N_6549,N_6516);
or U7990 (N_7990,N_6813,N_6069);
nor U7991 (N_7991,N_6906,N_6914);
nor U7992 (N_7992,N_6249,N_6993);
nor U7993 (N_7993,N_6464,N_6543);
or U7994 (N_7994,N_6291,N_6081);
and U7995 (N_7995,N_6214,N_6983);
or U7996 (N_7996,N_6844,N_6101);
and U7997 (N_7997,N_6709,N_6778);
nor U7998 (N_7998,N_6958,N_6478);
and U7999 (N_7999,N_6741,N_6081);
and U8000 (N_8000,N_7326,N_7190);
nor U8001 (N_8001,N_7896,N_7490);
or U8002 (N_8002,N_7953,N_7753);
nand U8003 (N_8003,N_7881,N_7290);
nand U8004 (N_8004,N_7076,N_7540);
nand U8005 (N_8005,N_7462,N_7372);
and U8006 (N_8006,N_7447,N_7364);
nor U8007 (N_8007,N_7343,N_7066);
or U8008 (N_8008,N_7198,N_7743);
or U8009 (N_8009,N_7432,N_7093);
nor U8010 (N_8010,N_7107,N_7439);
xor U8011 (N_8011,N_7413,N_7787);
or U8012 (N_8012,N_7717,N_7480);
nand U8013 (N_8013,N_7919,N_7534);
and U8014 (N_8014,N_7758,N_7228);
and U8015 (N_8015,N_7176,N_7120);
or U8016 (N_8016,N_7634,N_7530);
or U8017 (N_8017,N_7659,N_7960);
and U8018 (N_8018,N_7279,N_7169);
nand U8019 (N_8019,N_7848,N_7003);
nand U8020 (N_8020,N_7360,N_7218);
and U8021 (N_8021,N_7523,N_7351);
nand U8022 (N_8022,N_7217,N_7824);
nand U8023 (N_8023,N_7974,N_7177);
xnor U8024 (N_8024,N_7297,N_7903);
xor U8025 (N_8025,N_7786,N_7150);
xor U8026 (N_8026,N_7792,N_7132);
and U8027 (N_8027,N_7681,N_7819);
and U8028 (N_8028,N_7053,N_7330);
or U8029 (N_8029,N_7238,N_7453);
or U8030 (N_8030,N_7261,N_7844);
or U8031 (N_8031,N_7492,N_7160);
or U8032 (N_8032,N_7564,N_7780);
nor U8033 (N_8033,N_7603,N_7438);
nor U8034 (N_8034,N_7155,N_7508);
and U8035 (N_8035,N_7986,N_7361);
nand U8036 (N_8036,N_7934,N_7752);
and U8037 (N_8037,N_7312,N_7663);
nor U8038 (N_8038,N_7018,N_7902);
and U8039 (N_8039,N_7460,N_7166);
nand U8040 (N_8040,N_7158,N_7631);
nand U8041 (N_8041,N_7365,N_7377);
nor U8042 (N_8042,N_7324,N_7253);
and U8043 (N_8043,N_7382,N_7957);
and U8044 (N_8044,N_7207,N_7011);
and U8045 (N_8045,N_7989,N_7212);
or U8046 (N_8046,N_7715,N_7452);
and U8047 (N_8047,N_7455,N_7032);
or U8048 (N_8048,N_7461,N_7767);
or U8049 (N_8049,N_7676,N_7916);
and U8050 (N_8050,N_7882,N_7674);
nand U8051 (N_8051,N_7867,N_7707);
nand U8052 (N_8052,N_7313,N_7146);
nand U8053 (N_8053,N_7282,N_7337);
nor U8054 (N_8054,N_7251,N_7259);
xnor U8055 (N_8055,N_7315,N_7426);
or U8056 (N_8056,N_7839,N_7179);
or U8057 (N_8057,N_7005,N_7936);
and U8058 (N_8058,N_7021,N_7976);
nand U8059 (N_8059,N_7933,N_7850);
nand U8060 (N_8060,N_7857,N_7802);
nor U8061 (N_8061,N_7174,N_7098);
nor U8062 (N_8062,N_7449,N_7651);
and U8063 (N_8063,N_7777,N_7255);
and U8064 (N_8064,N_7551,N_7996);
xnor U8065 (N_8065,N_7489,N_7940);
or U8066 (N_8066,N_7376,N_7849);
nor U8067 (N_8067,N_7263,N_7770);
nand U8068 (N_8068,N_7615,N_7646);
and U8069 (N_8069,N_7944,N_7947);
or U8070 (N_8070,N_7287,N_7878);
nor U8071 (N_8071,N_7955,N_7069);
nor U8072 (N_8072,N_7214,N_7143);
or U8073 (N_8073,N_7749,N_7359);
or U8074 (N_8074,N_7227,N_7733);
nand U8075 (N_8075,N_7039,N_7062);
nor U8076 (N_8076,N_7528,N_7347);
nor U8077 (N_8077,N_7532,N_7549);
xor U8078 (N_8078,N_7864,N_7982);
xor U8079 (N_8079,N_7684,N_7584);
xnor U8080 (N_8080,N_7704,N_7072);
xnor U8081 (N_8081,N_7224,N_7473);
and U8082 (N_8082,N_7090,N_7593);
xor U8083 (N_8083,N_7642,N_7070);
nor U8084 (N_8084,N_7156,N_7956);
xnor U8085 (N_8085,N_7379,N_7741);
and U8086 (N_8086,N_7772,N_7429);
xnor U8087 (N_8087,N_7428,N_7022);
nor U8088 (N_8088,N_7325,N_7952);
nand U8089 (N_8089,N_7249,N_7052);
or U8090 (N_8090,N_7973,N_7856);
nor U8091 (N_8091,N_7084,N_7766);
xnor U8092 (N_8092,N_7464,N_7804);
or U8093 (N_8093,N_7424,N_7135);
nor U8094 (N_8094,N_7133,N_7478);
or U8095 (N_8095,N_7998,N_7242);
nor U8096 (N_8096,N_7191,N_7025);
nand U8097 (N_8097,N_7840,N_7927);
or U8098 (N_8098,N_7581,N_7421);
nor U8099 (N_8099,N_7513,N_7123);
nand U8100 (N_8100,N_7204,N_7703);
or U8101 (N_8101,N_7122,N_7307);
nand U8102 (N_8102,N_7127,N_7496);
nand U8103 (N_8103,N_7291,N_7789);
and U8104 (N_8104,N_7740,N_7983);
or U8105 (N_8105,N_7170,N_7946);
or U8106 (N_8106,N_7285,N_7451);
or U8107 (N_8107,N_7892,N_7813);
and U8108 (N_8108,N_7153,N_7689);
nor U8109 (N_8109,N_7491,N_7109);
or U8110 (N_8110,N_7951,N_7163);
and U8111 (N_8111,N_7275,N_7550);
and U8112 (N_8112,N_7334,N_7724);
nor U8113 (N_8113,N_7001,N_7614);
nor U8114 (N_8114,N_7806,N_7474);
nor U8115 (N_8115,N_7654,N_7873);
nand U8116 (N_8116,N_7706,N_7535);
nand U8117 (N_8117,N_7638,N_7537);
nor U8118 (N_8118,N_7725,N_7798);
nand U8119 (N_8119,N_7510,N_7055);
and U8120 (N_8120,N_7157,N_7722);
nand U8121 (N_8121,N_7697,N_7696);
nor U8122 (N_8122,N_7346,N_7463);
nor U8123 (N_8123,N_7609,N_7517);
and U8124 (N_8124,N_7292,N_7682);
and U8125 (N_8125,N_7695,N_7583);
and U8126 (N_8126,N_7754,N_7041);
and U8127 (N_8127,N_7845,N_7412);
nor U8128 (N_8128,N_7992,N_7814);
nand U8129 (N_8129,N_7110,N_7876);
nand U8130 (N_8130,N_7827,N_7056);
nor U8131 (N_8131,N_7173,N_7736);
xor U8132 (N_8132,N_7941,N_7723);
nand U8133 (N_8133,N_7495,N_7137);
nor U8134 (N_8134,N_7437,N_7991);
xor U8135 (N_8135,N_7771,N_7942);
nand U8136 (N_8136,N_7289,N_7580);
nand U8137 (N_8137,N_7807,N_7795);
nor U8138 (N_8138,N_7327,N_7811);
or U8139 (N_8139,N_7081,N_7910);
or U8140 (N_8140,N_7546,N_7196);
xnor U8141 (N_8141,N_7082,N_7899);
and U8142 (N_8142,N_7618,N_7044);
nand U8143 (N_8143,N_7295,N_7430);
nor U8144 (N_8144,N_7433,N_7860);
nand U8145 (N_8145,N_7504,N_7250);
and U8146 (N_8146,N_7643,N_7685);
nand U8147 (N_8147,N_7559,N_7907);
or U8148 (N_8148,N_7590,N_7310);
and U8149 (N_8149,N_7086,N_7677);
or U8150 (N_8150,N_7928,N_7125);
or U8151 (N_8151,N_7821,N_7594);
nor U8152 (N_8152,N_7019,N_7416);
and U8153 (N_8153,N_7775,N_7639);
and U8154 (N_8154,N_7620,N_7768);
nand U8155 (N_8155,N_7932,N_7230);
xnor U8156 (N_8156,N_7653,N_7512);
xnor U8157 (N_8157,N_7678,N_7183);
or U8158 (N_8158,N_7317,N_7605);
nand U8159 (N_8159,N_7818,N_7656);
and U8160 (N_8160,N_7894,N_7900);
nor U8161 (N_8161,N_7094,N_7755);
or U8162 (N_8162,N_7990,N_7624);
nor U8163 (N_8163,N_7661,N_7893);
or U8164 (N_8164,N_7505,N_7929);
xnor U8165 (N_8165,N_7306,N_7471);
or U8166 (N_8166,N_7141,N_7344);
or U8167 (N_8167,N_7843,N_7050);
and U8168 (N_8168,N_7048,N_7200);
nor U8169 (N_8169,N_7995,N_7621);
nor U8170 (N_8170,N_7381,N_7063);
nor U8171 (N_8171,N_7318,N_7494);
nor U8172 (N_8172,N_7920,N_7035);
xnor U8173 (N_8173,N_7260,N_7533);
or U8174 (N_8174,N_7144,N_7554);
or U8175 (N_8175,N_7977,N_7467);
xnor U8176 (N_8176,N_7553,N_7014);
and U8177 (N_8177,N_7288,N_7193);
nand U8178 (N_8178,N_7465,N_7031);
and U8179 (N_8179,N_7375,N_7872);
xnor U8180 (N_8180,N_7906,N_7617);
nor U8181 (N_8181,N_7908,N_7162);
nor U8182 (N_8182,N_7104,N_7272);
nor U8183 (N_8183,N_7924,N_7411);
or U8184 (N_8184,N_7672,N_7585);
nor U8185 (N_8185,N_7869,N_7889);
or U8186 (N_8186,N_7138,N_7130);
nor U8187 (N_8187,N_7520,N_7536);
or U8188 (N_8188,N_7409,N_7475);
nor U8189 (N_8189,N_7809,N_7484);
nand U8190 (N_8190,N_7599,N_7264);
and U8191 (N_8191,N_7274,N_7506);
xor U8192 (N_8192,N_7950,N_7633);
nand U8193 (N_8193,N_7610,N_7579);
and U8194 (N_8194,N_7403,N_7277);
nand U8195 (N_8195,N_7219,N_7443);
nand U8196 (N_8196,N_7229,N_7825);
nand U8197 (N_8197,N_7516,N_7943);
or U8198 (N_8198,N_7338,N_7577);
and U8199 (N_8199,N_7362,N_7834);
nor U8200 (N_8200,N_7525,N_7801);
nor U8201 (N_8201,N_7636,N_7606);
and U8202 (N_8202,N_7008,N_7803);
or U8203 (N_8203,N_7859,N_7124);
and U8204 (N_8204,N_7572,N_7458);
nor U8205 (N_8205,N_7978,N_7342);
and U8206 (N_8206,N_7963,N_7009);
nand U8207 (N_8207,N_7912,N_7959);
nor U8208 (N_8208,N_7435,N_7734);
or U8209 (N_8209,N_7100,N_7855);
xnor U8210 (N_8210,N_7367,N_7891);
nor U8211 (N_8211,N_7040,N_7222);
and U8212 (N_8212,N_7024,N_7791);
or U8213 (N_8213,N_7886,N_7033);
xor U8214 (N_8214,N_7023,N_7149);
and U8215 (N_8215,N_7237,N_7061);
and U8216 (N_8216,N_7628,N_7842);
nor U8217 (N_8217,N_7108,N_7895);
and U8218 (N_8218,N_7975,N_7175);
nand U8219 (N_8219,N_7988,N_7105);
and U8220 (N_8220,N_7640,N_7917);
and U8221 (N_8221,N_7765,N_7391);
nor U8222 (N_8222,N_7923,N_7254);
xor U8223 (N_8223,N_7357,N_7838);
and U8224 (N_8224,N_7673,N_7984);
nor U8225 (N_8225,N_7748,N_7232);
nand U8226 (N_8226,N_7485,N_7797);
or U8227 (N_8227,N_7454,N_7737);
and U8228 (N_8228,N_7388,N_7374);
nand U8229 (N_8229,N_7392,N_7119);
and U8230 (N_8230,N_7262,N_7664);
nand U8231 (N_8231,N_7225,N_7178);
xor U8232 (N_8232,N_7914,N_7587);
or U8233 (N_8233,N_7657,N_7356);
or U8234 (N_8234,N_7300,N_7000);
or U8235 (N_8235,N_7199,N_7373);
and U8236 (N_8236,N_7397,N_7529);
and U8237 (N_8237,N_7964,N_7853);
and U8238 (N_8238,N_7761,N_7233);
nand U8239 (N_8239,N_7999,N_7721);
nor U8240 (N_8240,N_7680,N_7210);
nand U8241 (N_8241,N_7383,N_7500);
or U8242 (N_8242,N_7836,N_7258);
nand U8243 (N_8243,N_7880,N_7414);
nand U8244 (N_8244,N_7060,N_7472);
nand U8245 (N_8245,N_7563,N_7139);
nor U8246 (N_8246,N_7519,N_7997);
or U8247 (N_8247,N_7547,N_7700);
and U8248 (N_8248,N_7187,N_7235);
nand U8249 (N_8249,N_7099,N_7817);
or U8250 (N_8250,N_7284,N_7476);
and U8251 (N_8251,N_7305,N_7220);
nand U8252 (N_8252,N_7442,N_7687);
nand U8253 (N_8253,N_7469,N_7625);
or U8254 (N_8254,N_7562,N_7102);
nor U8255 (N_8255,N_7875,N_7425);
nand U8256 (N_8256,N_7029,N_7405);
nand U8257 (N_8257,N_7152,N_7582);
xnor U8258 (N_8258,N_7402,N_7764);
nand U8259 (N_8259,N_7714,N_7650);
nor U8260 (N_8260,N_7962,N_7189);
and U8261 (N_8261,N_7064,N_7742);
and U8262 (N_8262,N_7065,N_7726);
xnor U8263 (N_8263,N_7637,N_7556);
or U8264 (N_8264,N_7241,N_7822);
or U8265 (N_8265,N_7349,N_7870);
nor U8266 (N_8266,N_7016,N_7799);
and U8267 (N_8267,N_7406,N_7783);
and U8268 (N_8268,N_7215,N_7710);
nand U8269 (N_8269,N_7479,N_7731);
nand U8270 (N_8270,N_7745,N_7800);
or U8271 (N_8271,N_7598,N_7322);
nor U8272 (N_8272,N_7969,N_7006);
nor U8273 (N_8273,N_7883,N_7404);
and U8274 (N_8274,N_7611,N_7201);
xor U8275 (N_8275,N_7779,N_7091);
and U8276 (N_8276,N_7954,N_7206);
or U8277 (N_8277,N_7552,N_7134);
nor U8278 (N_8278,N_7925,N_7885);
nor U8279 (N_8279,N_7622,N_7441);
or U8280 (N_8280,N_7395,N_7419);
nand U8281 (N_8281,N_7970,N_7645);
nor U8282 (N_8282,N_7862,N_7269);
nor U8283 (N_8283,N_7569,N_7560);
and U8284 (N_8284,N_7159,N_7320);
or U8285 (N_8285,N_7221,N_7036);
nand U8286 (N_8286,N_7340,N_7281);
and U8287 (N_8287,N_7352,N_7145);
or U8288 (N_8288,N_7888,N_7702);
nand U8289 (N_8289,N_7470,N_7126);
and U8290 (N_8290,N_7252,N_7167);
nor U8291 (N_8291,N_7666,N_7884);
nor U8292 (N_8292,N_7165,N_7705);
or U8293 (N_8293,N_7851,N_7161);
and U8294 (N_8294,N_7732,N_7223);
or U8295 (N_8295,N_7117,N_7348);
xor U8296 (N_8296,N_7660,N_7142);
xnor U8297 (N_8297,N_7945,N_7431);
nand U8298 (N_8298,N_7012,N_7450);
xor U8299 (N_8299,N_7810,N_7905);
or U8300 (N_8300,N_7283,N_7151);
and U8301 (N_8301,N_7314,N_7597);
nand U8302 (N_8302,N_7180,N_7887);
nand U8303 (N_8303,N_7616,N_7667);
nand U8304 (N_8304,N_7332,N_7698);
nand U8305 (N_8305,N_7762,N_7482);
or U8306 (N_8306,N_7539,N_7101);
nor U8307 (N_8307,N_7020,N_7243);
and U8308 (N_8308,N_7852,N_7820);
nand U8309 (N_8309,N_7046,N_7445);
and U8310 (N_8310,N_7607,N_7353);
nand U8311 (N_8311,N_7497,N_7400);
nand U8312 (N_8312,N_7586,N_7909);
xnor U8313 (N_8313,N_7747,N_7493);
nor U8314 (N_8314,N_7877,N_7648);
or U8315 (N_8315,N_7502,N_7985);
or U8316 (N_8316,N_7034,N_7466);
xnor U8317 (N_8317,N_7655,N_7566);
nor U8318 (N_8318,N_7387,N_7042);
xor U8319 (N_8319,N_7711,N_7693);
xnor U8320 (N_8320,N_7623,N_7075);
or U8321 (N_8321,N_7576,N_7632);
and U8322 (N_8322,N_7627,N_7694);
nand U8323 (N_8323,N_7074,N_7708);
nor U8324 (N_8324,N_7949,N_7776);
nor U8325 (N_8325,N_7863,N_7613);
nand U8326 (N_8326,N_7004,N_7182);
and U8327 (N_8327,N_7319,N_7841);
nand U8328 (N_8328,N_7097,N_7369);
or U8329 (N_8329,N_7796,N_7358);
and U8330 (N_8330,N_7668,N_7498);
nand U8331 (N_8331,N_7027,N_7541);
nand U8332 (N_8332,N_7037,N_7647);
nand U8333 (N_8333,N_7136,N_7394);
nand U8334 (N_8334,N_7823,N_7380);
or U8335 (N_8335,N_7833,N_7140);
or U8336 (N_8336,N_7446,N_7879);
or U8337 (N_8337,N_7602,N_7756);
nand U8338 (N_8338,N_7298,N_7937);
nand U8339 (N_8339,N_7837,N_7926);
xnor U8340 (N_8340,N_7782,N_7026);
nor U8341 (N_8341,N_7423,N_7600);
nand U8342 (N_8342,N_7267,N_7874);
xor U8343 (N_8343,N_7257,N_7930);
xnor U8344 (N_8344,N_7720,N_7612);
or U8345 (N_8345,N_7378,N_7270);
nor U8346 (N_8346,N_7578,N_7662);
nor U8347 (N_8347,N_7831,N_7538);
nor U8348 (N_8348,N_7709,N_7299);
and U8349 (N_8349,N_7911,N_7209);
or U8350 (N_8350,N_7354,N_7398);
xor U8351 (N_8351,N_7194,N_7979);
and U8352 (N_8352,N_7366,N_7861);
nand U8353 (N_8353,N_7993,N_7244);
or U8354 (N_8354,N_7172,N_7106);
or U8355 (N_8355,N_7015,N_7865);
or U8356 (N_8356,N_7331,N_7192);
nand U8357 (N_8357,N_7521,N_7812);
nor U8358 (N_8358,N_7418,N_7245);
and U8359 (N_8359,N_7363,N_7746);
or U8360 (N_8360,N_7316,N_7088);
nor U8361 (N_8361,N_7670,N_7321);
nand U8362 (N_8362,N_7280,N_7049);
or U8363 (N_8363,N_7045,N_7308);
xor U8364 (N_8364,N_7067,N_7047);
nor U8365 (N_8365,N_7077,N_7236);
xnor U8366 (N_8366,N_7701,N_7486);
nor U8367 (N_8367,N_7248,N_7339);
and U8368 (N_8368,N_7630,N_7759);
and U8369 (N_8369,N_7328,N_7246);
xnor U8370 (N_8370,N_7526,N_7728);
nor U8371 (N_8371,N_7488,N_7644);
or U8372 (N_8372,N_7760,N_7483);
or U8373 (N_8373,N_7071,N_7401);
nand U8374 (N_8374,N_7738,N_7781);
nand U8375 (N_8375,N_7866,N_7545);
nand U8376 (N_8376,N_7095,N_7750);
nor U8377 (N_8377,N_7213,N_7769);
or U8378 (N_8378,N_7571,N_7835);
xor U8379 (N_8379,N_7968,N_7719);
or U8380 (N_8380,N_7128,N_7116);
or U8381 (N_8381,N_7785,N_7931);
and U8382 (N_8382,N_7436,N_7739);
nor U8383 (N_8383,N_7211,N_7635);
and U8384 (N_8384,N_7846,N_7448);
nor U8385 (N_8385,N_7309,N_7002);
or U8386 (N_8386,N_7068,N_7350);
xor U8387 (N_8387,N_7871,N_7591);
nand U8388 (N_8388,N_7188,N_7980);
nand U8389 (N_8389,N_7113,N_7816);
and U8390 (N_8390,N_7202,N_7092);
or U8391 (N_8391,N_7972,N_7345);
nand U8392 (N_8392,N_7273,N_7010);
or U8393 (N_8393,N_7778,N_7981);
nor U8394 (N_8394,N_7057,N_7303);
and U8395 (N_8395,N_7399,N_7509);
nand U8396 (N_8396,N_7858,N_7440);
or U8397 (N_8397,N_7341,N_7078);
and U8398 (N_8398,N_7692,N_7573);
nor U8399 (N_8399,N_7481,N_7575);
and U8400 (N_8400,N_7649,N_7103);
and U8401 (N_8401,N_7958,N_7051);
or U8402 (N_8402,N_7794,N_7393);
and U8403 (N_8403,N_7131,N_7115);
nand U8404 (N_8404,N_7548,N_7080);
or U8405 (N_8405,N_7205,N_7168);
or U8406 (N_8406,N_7890,N_7589);
and U8407 (N_8407,N_7386,N_7712);
nand U8408 (N_8408,N_7389,N_7181);
xor U8409 (N_8409,N_7355,N_7408);
nor U8410 (N_8410,N_7574,N_7456);
and U8411 (N_8411,N_7531,N_7118);
nand U8412 (N_8412,N_7604,N_7522);
or U8413 (N_8413,N_7544,N_7396);
nand U8414 (N_8414,N_7336,N_7240);
or U8415 (N_8415,N_7757,N_7938);
or U8416 (N_8416,N_7477,N_7868);
or U8417 (N_8417,N_7567,N_7058);
and U8418 (N_8418,N_7265,N_7971);
nor U8419 (N_8419,N_7671,N_7921);
or U8420 (N_8420,N_7017,N_7247);
nor U8421 (N_8421,N_7730,N_7744);
nand U8422 (N_8422,N_7987,N_7415);
nor U8423 (N_8423,N_7301,N_7608);
and U8424 (N_8424,N_7059,N_7901);
or U8425 (N_8425,N_7333,N_7729);
nor U8426 (N_8426,N_7713,N_7718);
nand U8427 (N_8427,N_7568,N_7089);
and U8428 (N_8428,N_7966,N_7407);
nor U8429 (N_8429,N_7043,N_7028);
nand U8430 (N_8430,N_7007,N_7335);
and U8431 (N_8431,N_7679,N_7847);
nor U8432 (N_8432,N_7268,N_7129);
nor U8433 (N_8433,N_7555,N_7371);
nor U8434 (N_8434,N_7427,N_7185);
and U8435 (N_8435,N_7276,N_7967);
or U8436 (N_8436,N_7417,N_7524);
nor U8437 (N_8437,N_7370,N_7826);
xor U8438 (N_8438,N_7790,N_7208);
nor U8439 (N_8439,N_7296,N_7897);
or U8440 (N_8440,N_7773,N_7186);
or U8441 (N_8441,N_7385,N_7154);
nor U8442 (N_8442,N_7683,N_7501);
nor U8443 (N_8443,N_7716,N_7234);
or U8444 (N_8444,N_7751,N_7898);
nor U8445 (N_8445,N_7691,N_7558);
nand U8446 (N_8446,N_7266,N_7961);
nand U8447 (N_8447,N_7256,N_7763);
nand U8448 (N_8448,N_7457,N_7808);
xnor U8449 (N_8449,N_7079,N_7148);
nor U8450 (N_8450,N_7514,N_7829);
or U8451 (N_8451,N_7570,N_7216);
nand U8452 (N_8452,N_7686,N_7652);
nor U8453 (N_8453,N_7965,N_7619);
nand U8454 (N_8454,N_7278,N_7085);
or U8455 (N_8455,N_7669,N_7294);
xor U8456 (N_8456,N_7390,N_7727);
nand U8457 (N_8457,N_7422,N_7420);
nand U8458 (N_8458,N_7323,N_7304);
nand U8459 (N_8459,N_7195,N_7164);
or U8460 (N_8460,N_7592,N_7410);
and U8461 (N_8461,N_7557,N_7784);
nor U8462 (N_8462,N_7830,N_7239);
nor U8463 (N_8463,N_7913,N_7527);
nor U8464 (N_8464,N_7832,N_7658);
nand U8465 (N_8465,N_7459,N_7226);
and U8466 (N_8466,N_7629,N_7147);
nand U8467 (N_8467,N_7293,N_7073);
or U8468 (N_8468,N_7507,N_7588);
and U8469 (N_8469,N_7915,N_7302);
nand U8470 (N_8470,N_7688,N_7096);
nand U8471 (N_8471,N_7774,N_7595);
xor U8472 (N_8472,N_7854,N_7935);
xnor U8473 (N_8473,N_7596,N_7565);
or U8474 (N_8474,N_7499,N_7111);
or U8475 (N_8475,N_7184,N_7038);
xnor U8476 (N_8476,N_7329,N_7815);
nor U8477 (N_8477,N_7286,N_7114);
nand U8478 (N_8478,N_7054,N_7626);
and U8479 (N_8479,N_7203,N_7434);
nor U8480 (N_8480,N_7083,N_7690);
and U8481 (N_8481,N_7675,N_7793);
or U8482 (N_8482,N_7121,N_7543);
xor U8483 (N_8483,N_7561,N_7665);
nor U8484 (N_8484,N_7271,N_7904);
and U8485 (N_8485,N_7468,N_7542);
nand U8486 (N_8486,N_7013,N_7699);
nand U8487 (N_8487,N_7641,N_7384);
nand U8488 (N_8488,N_7030,N_7112);
nor U8489 (N_8489,N_7311,N_7511);
or U8490 (N_8490,N_7948,N_7939);
and U8491 (N_8491,N_7503,N_7922);
xnor U8492 (N_8492,N_7444,N_7487);
or U8493 (N_8493,N_7515,N_7197);
or U8494 (N_8494,N_7994,N_7805);
nand U8495 (N_8495,N_7171,N_7601);
nor U8496 (N_8496,N_7828,N_7788);
or U8497 (N_8497,N_7518,N_7735);
nand U8498 (N_8498,N_7231,N_7087);
and U8499 (N_8499,N_7918,N_7368);
xor U8500 (N_8500,N_7363,N_7762);
nand U8501 (N_8501,N_7489,N_7011);
and U8502 (N_8502,N_7871,N_7464);
or U8503 (N_8503,N_7973,N_7116);
or U8504 (N_8504,N_7115,N_7721);
nor U8505 (N_8505,N_7549,N_7450);
or U8506 (N_8506,N_7142,N_7077);
or U8507 (N_8507,N_7375,N_7533);
or U8508 (N_8508,N_7849,N_7514);
nor U8509 (N_8509,N_7889,N_7428);
or U8510 (N_8510,N_7664,N_7305);
xor U8511 (N_8511,N_7174,N_7211);
nor U8512 (N_8512,N_7319,N_7903);
or U8513 (N_8513,N_7389,N_7376);
nand U8514 (N_8514,N_7827,N_7903);
xor U8515 (N_8515,N_7090,N_7610);
nand U8516 (N_8516,N_7428,N_7409);
nand U8517 (N_8517,N_7963,N_7710);
nand U8518 (N_8518,N_7837,N_7779);
and U8519 (N_8519,N_7579,N_7158);
nor U8520 (N_8520,N_7761,N_7854);
nand U8521 (N_8521,N_7186,N_7948);
nor U8522 (N_8522,N_7017,N_7970);
and U8523 (N_8523,N_7030,N_7358);
xor U8524 (N_8524,N_7568,N_7060);
or U8525 (N_8525,N_7654,N_7333);
or U8526 (N_8526,N_7062,N_7734);
and U8527 (N_8527,N_7133,N_7376);
nand U8528 (N_8528,N_7644,N_7832);
or U8529 (N_8529,N_7612,N_7231);
or U8530 (N_8530,N_7736,N_7490);
nand U8531 (N_8531,N_7710,N_7927);
xnor U8532 (N_8532,N_7386,N_7257);
xnor U8533 (N_8533,N_7159,N_7909);
nor U8534 (N_8534,N_7781,N_7303);
nor U8535 (N_8535,N_7588,N_7373);
and U8536 (N_8536,N_7486,N_7372);
or U8537 (N_8537,N_7279,N_7812);
and U8538 (N_8538,N_7604,N_7026);
or U8539 (N_8539,N_7282,N_7744);
nand U8540 (N_8540,N_7316,N_7664);
nand U8541 (N_8541,N_7201,N_7164);
or U8542 (N_8542,N_7548,N_7491);
nand U8543 (N_8543,N_7956,N_7487);
or U8544 (N_8544,N_7694,N_7747);
and U8545 (N_8545,N_7476,N_7381);
or U8546 (N_8546,N_7413,N_7433);
or U8547 (N_8547,N_7316,N_7502);
nand U8548 (N_8548,N_7772,N_7338);
nor U8549 (N_8549,N_7732,N_7294);
nor U8550 (N_8550,N_7321,N_7348);
nor U8551 (N_8551,N_7438,N_7104);
and U8552 (N_8552,N_7132,N_7594);
and U8553 (N_8553,N_7631,N_7222);
nor U8554 (N_8554,N_7227,N_7157);
nor U8555 (N_8555,N_7967,N_7735);
or U8556 (N_8556,N_7185,N_7744);
and U8557 (N_8557,N_7130,N_7228);
or U8558 (N_8558,N_7750,N_7973);
nor U8559 (N_8559,N_7432,N_7694);
and U8560 (N_8560,N_7352,N_7514);
and U8561 (N_8561,N_7832,N_7236);
or U8562 (N_8562,N_7380,N_7873);
or U8563 (N_8563,N_7524,N_7440);
nor U8564 (N_8564,N_7671,N_7862);
nand U8565 (N_8565,N_7709,N_7082);
or U8566 (N_8566,N_7586,N_7016);
nor U8567 (N_8567,N_7715,N_7283);
nor U8568 (N_8568,N_7733,N_7505);
nor U8569 (N_8569,N_7163,N_7001);
nor U8570 (N_8570,N_7307,N_7947);
and U8571 (N_8571,N_7826,N_7583);
nor U8572 (N_8572,N_7553,N_7387);
nand U8573 (N_8573,N_7605,N_7935);
or U8574 (N_8574,N_7098,N_7991);
and U8575 (N_8575,N_7143,N_7027);
nand U8576 (N_8576,N_7324,N_7667);
nand U8577 (N_8577,N_7076,N_7225);
or U8578 (N_8578,N_7544,N_7167);
nor U8579 (N_8579,N_7903,N_7793);
xor U8580 (N_8580,N_7845,N_7734);
nand U8581 (N_8581,N_7950,N_7877);
or U8582 (N_8582,N_7648,N_7268);
or U8583 (N_8583,N_7019,N_7497);
xor U8584 (N_8584,N_7464,N_7985);
nor U8585 (N_8585,N_7365,N_7507);
nor U8586 (N_8586,N_7553,N_7417);
and U8587 (N_8587,N_7651,N_7135);
nor U8588 (N_8588,N_7087,N_7630);
nand U8589 (N_8589,N_7966,N_7815);
xnor U8590 (N_8590,N_7185,N_7632);
nor U8591 (N_8591,N_7236,N_7797);
and U8592 (N_8592,N_7460,N_7526);
and U8593 (N_8593,N_7239,N_7606);
nand U8594 (N_8594,N_7631,N_7220);
or U8595 (N_8595,N_7319,N_7952);
or U8596 (N_8596,N_7890,N_7282);
nand U8597 (N_8597,N_7210,N_7877);
nand U8598 (N_8598,N_7806,N_7188);
or U8599 (N_8599,N_7018,N_7401);
nor U8600 (N_8600,N_7403,N_7723);
nand U8601 (N_8601,N_7274,N_7481);
or U8602 (N_8602,N_7148,N_7939);
xor U8603 (N_8603,N_7261,N_7428);
or U8604 (N_8604,N_7728,N_7558);
nor U8605 (N_8605,N_7380,N_7187);
nand U8606 (N_8606,N_7919,N_7662);
nor U8607 (N_8607,N_7523,N_7376);
nor U8608 (N_8608,N_7834,N_7312);
nor U8609 (N_8609,N_7324,N_7258);
xor U8610 (N_8610,N_7880,N_7789);
or U8611 (N_8611,N_7173,N_7662);
nand U8612 (N_8612,N_7762,N_7999);
nor U8613 (N_8613,N_7341,N_7393);
nor U8614 (N_8614,N_7478,N_7983);
and U8615 (N_8615,N_7991,N_7610);
or U8616 (N_8616,N_7743,N_7693);
and U8617 (N_8617,N_7674,N_7859);
or U8618 (N_8618,N_7081,N_7921);
nor U8619 (N_8619,N_7337,N_7652);
nor U8620 (N_8620,N_7421,N_7049);
nor U8621 (N_8621,N_7959,N_7931);
nand U8622 (N_8622,N_7295,N_7573);
nor U8623 (N_8623,N_7275,N_7661);
or U8624 (N_8624,N_7149,N_7364);
and U8625 (N_8625,N_7767,N_7572);
or U8626 (N_8626,N_7828,N_7724);
and U8627 (N_8627,N_7131,N_7737);
and U8628 (N_8628,N_7371,N_7872);
nor U8629 (N_8629,N_7140,N_7232);
nand U8630 (N_8630,N_7314,N_7289);
nand U8631 (N_8631,N_7567,N_7098);
nor U8632 (N_8632,N_7681,N_7377);
or U8633 (N_8633,N_7569,N_7203);
nand U8634 (N_8634,N_7882,N_7307);
or U8635 (N_8635,N_7999,N_7368);
nand U8636 (N_8636,N_7171,N_7781);
nor U8637 (N_8637,N_7170,N_7091);
or U8638 (N_8638,N_7365,N_7601);
nand U8639 (N_8639,N_7285,N_7630);
or U8640 (N_8640,N_7876,N_7339);
or U8641 (N_8641,N_7494,N_7323);
nor U8642 (N_8642,N_7911,N_7795);
or U8643 (N_8643,N_7552,N_7469);
nand U8644 (N_8644,N_7052,N_7524);
nor U8645 (N_8645,N_7048,N_7023);
and U8646 (N_8646,N_7087,N_7802);
nor U8647 (N_8647,N_7692,N_7707);
or U8648 (N_8648,N_7932,N_7079);
nor U8649 (N_8649,N_7211,N_7333);
nand U8650 (N_8650,N_7054,N_7151);
and U8651 (N_8651,N_7673,N_7164);
and U8652 (N_8652,N_7813,N_7509);
or U8653 (N_8653,N_7976,N_7970);
nor U8654 (N_8654,N_7574,N_7748);
nand U8655 (N_8655,N_7979,N_7412);
and U8656 (N_8656,N_7546,N_7797);
nor U8657 (N_8657,N_7036,N_7708);
nand U8658 (N_8658,N_7882,N_7973);
or U8659 (N_8659,N_7462,N_7501);
nand U8660 (N_8660,N_7255,N_7564);
nor U8661 (N_8661,N_7102,N_7633);
nand U8662 (N_8662,N_7576,N_7655);
and U8663 (N_8663,N_7620,N_7921);
xnor U8664 (N_8664,N_7803,N_7484);
nor U8665 (N_8665,N_7101,N_7851);
and U8666 (N_8666,N_7670,N_7398);
nor U8667 (N_8667,N_7533,N_7699);
nor U8668 (N_8668,N_7851,N_7145);
nand U8669 (N_8669,N_7045,N_7469);
nand U8670 (N_8670,N_7872,N_7991);
or U8671 (N_8671,N_7864,N_7388);
and U8672 (N_8672,N_7436,N_7049);
xnor U8673 (N_8673,N_7859,N_7502);
nand U8674 (N_8674,N_7385,N_7613);
nand U8675 (N_8675,N_7392,N_7391);
xnor U8676 (N_8676,N_7155,N_7801);
nand U8677 (N_8677,N_7266,N_7559);
or U8678 (N_8678,N_7271,N_7755);
or U8679 (N_8679,N_7176,N_7782);
or U8680 (N_8680,N_7497,N_7786);
and U8681 (N_8681,N_7877,N_7239);
nor U8682 (N_8682,N_7707,N_7098);
nand U8683 (N_8683,N_7458,N_7013);
nor U8684 (N_8684,N_7059,N_7135);
xor U8685 (N_8685,N_7954,N_7548);
or U8686 (N_8686,N_7037,N_7571);
nand U8687 (N_8687,N_7611,N_7488);
nor U8688 (N_8688,N_7486,N_7888);
nor U8689 (N_8689,N_7149,N_7868);
nor U8690 (N_8690,N_7447,N_7862);
and U8691 (N_8691,N_7051,N_7566);
nand U8692 (N_8692,N_7007,N_7673);
nor U8693 (N_8693,N_7671,N_7251);
xor U8694 (N_8694,N_7089,N_7639);
and U8695 (N_8695,N_7104,N_7489);
or U8696 (N_8696,N_7626,N_7386);
nand U8697 (N_8697,N_7590,N_7253);
or U8698 (N_8698,N_7116,N_7549);
or U8699 (N_8699,N_7062,N_7156);
and U8700 (N_8700,N_7942,N_7131);
and U8701 (N_8701,N_7009,N_7842);
and U8702 (N_8702,N_7372,N_7005);
and U8703 (N_8703,N_7968,N_7113);
nor U8704 (N_8704,N_7932,N_7757);
xnor U8705 (N_8705,N_7195,N_7904);
nand U8706 (N_8706,N_7725,N_7625);
nor U8707 (N_8707,N_7947,N_7926);
nand U8708 (N_8708,N_7411,N_7683);
nor U8709 (N_8709,N_7715,N_7069);
nor U8710 (N_8710,N_7442,N_7592);
nand U8711 (N_8711,N_7989,N_7550);
nor U8712 (N_8712,N_7289,N_7012);
nand U8713 (N_8713,N_7083,N_7503);
nand U8714 (N_8714,N_7404,N_7243);
and U8715 (N_8715,N_7058,N_7513);
nor U8716 (N_8716,N_7304,N_7167);
nor U8717 (N_8717,N_7275,N_7434);
nand U8718 (N_8718,N_7571,N_7128);
and U8719 (N_8719,N_7864,N_7528);
or U8720 (N_8720,N_7520,N_7886);
nand U8721 (N_8721,N_7941,N_7849);
nor U8722 (N_8722,N_7678,N_7598);
or U8723 (N_8723,N_7384,N_7127);
and U8724 (N_8724,N_7489,N_7639);
and U8725 (N_8725,N_7937,N_7841);
xnor U8726 (N_8726,N_7429,N_7980);
and U8727 (N_8727,N_7834,N_7498);
nand U8728 (N_8728,N_7625,N_7774);
nor U8729 (N_8729,N_7435,N_7047);
nor U8730 (N_8730,N_7072,N_7423);
or U8731 (N_8731,N_7772,N_7986);
and U8732 (N_8732,N_7039,N_7359);
and U8733 (N_8733,N_7609,N_7922);
or U8734 (N_8734,N_7393,N_7293);
or U8735 (N_8735,N_7621,N_7276);
nor U8736 (N_8736,N_7639,N_7218);
nor U8737 (N_8737,N_7892,N_7346);
nand U8738 (N_8738,N_7389,N_7284);
nor U8739 (N_8739,N_7463,N_7526);
nand U8740 (N_8740,N_7440,N_7525);
or U8741 (N_8741,N_7442,N_7697);
or U8742 (N_8742,N_7130,N_7923);
or U8743 (N_8743,N_7050,N_7115);
nor U8744 (N_8744,N_7992,N_7863);
nor U8745 (N_8745,N_7913,N_7158);
and U8746 (N_8746,N_7092,N_7181);
and U8747 (N_8747,N_7504,N_7759);
or U8748 (N_8748,N_7883,N_7505);
or U8749 (N_8749,N_7672,N_7968);
nor U8750 (N_8750,N_7736,N_7928);
or U8751 (N_8751,N_7041,N_7113);
nand U8752 (N_8752,N_7519,N_7473);
nor U8753 (N_8753,N_7377,N_7413);
nand U8754 (N_8754,N_7956,N_7262);
nor U8755 (N_8755,N_7446,N_7582);
and U8756 (N_8756,N_7541,N_7457);
nor U8757 (N_8757,N_7699,N_7385);
nand U8758 (N_8758,N_7816,N_7380);
nand U8759 (N_8759,N_7267,N_7440);
nand U8760 (N_8760,N_7307,N_7019);
nor U8761 (N_8761,N_7664,N_7688);
nand U8762 (N_8762,N_7363,N_7108);
nor U8763 (N_8763,N_7602,N_7263);
nor U8764 (N_8764,N_7406,N_7878);
xnor U8765 (N_8765,N_7706,N_7598);
or U8766 (N_8766,N_7035,N_7727);
or U8767 (N_8767,N_7247,N_7022);
or U8768 (N_8768,N_7860,N_7324);
nor U8769 (N_8769,N_7594,N_7457);
nand U8770 (N_8770,N_7225,N_7588);
nand U8771 (N_8771,N_7912,N_7087);
nand U8772 (N_8772,N_7992,N_7716);
or U8773 (N_8773,N_7889,N_7987);
or U8774 (N_8774,N_7250,N_7147);
and U8775 (N_8775,N_7537,N_7798);
and U8776 (N_8776,N_7657,N_7809);
xor U8777 (N_8777,N_7185,N_7271);
and U8778 (N_8778,N_7691,N_7508);
and U8779 (N_8779,N_7448,N_7028);
and U8780 (N_8780,N_7147,N_7472);
and U8781 (N_8781,N_7120,N_7602);
nor U8782 (N_8782,N_7325,N_7611);
nor U8783 (N_8783,N_7063,N_7847);
or U8784 (N_8784,N_7991,N_7893);
and U8785 (N_8785,N_7736,N_7953);
and U8786 (N_8786,N_7848,N_7635);
nand U8787 (N_8787,N_7682,N_7828);
and U8788 (N_8788,N_7983,N_7476);
nor U8789 (N_8789,N_7488,N_7388);
nand U8790 (N_8790,N_7341,N_7436);
and U8791 (N_8791,N_7599,N_7463);
nand U8792 (N_8792,N_7766,N_7000);
or U8793 (N_8793,N_7144,N_7896);
nor U8794 (N_8794,N_7098,N_7283);
nor U8795 (N_8795,N_7399,N_7999);
or U8796 (N_8796,N_7649,N_7485);
or U8797 (N_8797,N_7917,N_7773);
or U8798 (N_8798,N_7867,N_7138);
nand U8799 (N_8799,N_7833,N_7610);
xor U8800 (N_8800,N_7600,N_7053);
nor U8801 (N_8801,N_7325,N_7391);
and U8802 (N_8802,N_7453,N_7666);
and U8803 (N_8803,N_7778,N_7044);
xnor U8804 (N_8804,N_7374,N_7113);
and U8805 (N_8805,N_7968,N_7536);
or U8806 (N_8806,N_7232,N_7492);
or U8807 (N_8807,N_7172,N_7575);
or U8808 (N_8808,N_7160,N_7154);
nor U8809 (N_8809,N_7613,N_7302);
nand U8810 (N_8810,N_7236,N_7228);
nand U8811 (N_8811,N_7874,N_7569);
nand U8812 (N_8812,N_7255,N_7136);
xor U8813 (N_8813,N_7421,N_7155);
or U8814 (N_8814,N_7243,N_7689);
nand U8815 (N_8815,N_7035,N_7010);
nor U8816 (N_8816,N_7867,N_7409);
or U8817 (N_8817,N_7863,N_7745);
and U8818 (N_8818,N_7852,N_7677);
or U8819 (N_8819,N_7074,N_7544);
and U8820 (N_8820,N_7307,N_7987);
or U8821 (N_8821,N_7881,N_7274);
and U8822 (N_8822,N_7949,N_7743);
or U8823 (N_8823,N_7344,N_7244);
and U8824 (N_8824,N_7703,N_7630);
or U8825 (N_8825,N_7673,N_7620);
nand U8826 (N_8826,N_7620,N_7500);
nand U8827 (N_8827,N_7737,N_7015);
or U8828 (N_8828,N_7288,N_7953);
nand U8829 (N_8829,N_7696,N_7423);
or U8830 (N_8830,N_7619,N_7612);
nand U8831 (N_8831,N_7466,N_7195);
xnor U8832 (N_8832,N_7149,N_7729);
nor U8833 (N_8833,N_7853,N_7606);
and U8834 (N_8834,N_7297,N_7551);
or U8835 (N_8835,N_7745,N_7261);
nand U8836 (N_8836,N_7391,N_7377);
xor U8837 (N_8837,N_7997,N_7176);
and U8838 (N_8838,N_7960,N_7629);
or U8839 (N_8839,N_7266,N_7788);
and U8840 (N_8840,N_7421,N_7223);
or U8841 (N_8841,N_7978,N_7633);
nand U8842 (N_8842,N_7751,N_7745);
or U8843 (N_8843,N_7953,N_7291);
nor U8844 (N_8844,N_7380,N_7858);
and U8845 (N_8845,N_7038,N_7178);
nand U8846 (N_8846,N_7178,N_7545);
or U8847 (N_8847,N_7161,N_7790);
and U8848 (N_8848,N_7636,N_7055);
xor U8849 (N_8849,N_7801,N_7799);
or U8850 (N_8850,N_7530,N_7150);
nand U8851 (N_8851,N_7823,N_7936);
or U8852 (N_8852,N_7415,N_7882);
or U8853 (N_8853,N_7284,N_7713);
nor U8854 (N_8854,N_7074,N_7462);
nor U8855 (N_8855,N_7847,N_7953);
or U8856 (N_8856,N_7164,N_7324);
and U8857 (N_8857,N_7028,N_7418);
and U8858 (N_8858,N_7013,N_7804);
nand U8859 (N_8859,N_7899,N_7231);
and U8860 (N_8860,N_7640,N_7610);
nand U8861 (N_8861,N_7093,N_7919);
nand U8862 (N_8862,N_7709,N_7467);
nand U8863 (N_8863,N_7030,N_7891);
nor U8864 (N_8864,N_7502,N_7217);
xnor U8865 (N_8865,N_7144,N_7663);
nor U8866 (N_8866,N_7551,N_7376);
nand U8867 (N_8867,N_7196,N_7104);
nor U8868 (N_8868,N_7022,N_7780);
or U8869 (N_8869,N_7990,N_7913);
and U8870 (N_8870,N_7105,N_7107);
nor U8871 (N_8871,N_7345,N_7845);
nor U8872 (N_8872,N_7961,N_7285);
nor U8873 (N_8873,N_7207,N_7634);
and U8874 (N_8874,N_7898,N_7365);
or U8875 (N_8875,N_7339,N_7079);
or U8876 (N_8876,N_7404,N_7341);
and U8877 (N_8877,N_7079,N_7821);
or U8878 (N_8878,N_7791,N_7089);
nor U8879 (N_8879,N_7448,N_7905);
nor U8880 (N_8880,N_7533,N_7426);
or U8881 (N_8881,N_7216,N_7773);
nor U8882 (N_8882,N_7123,N_7363);
and U8883 (N_8883,N_7231,N_7072);
or U8884 (N_8884,N_7280,N_7090);
nand U8885 (N_8885,N_7899,N_7189);
nor U8886 (N_8886,N_7652,N_7561);
xor U8887 (N_8887,N_7544,N_7668);
nor U8888 (N_8888,N_7170,N_7161);
or U8889 (N_8889,N_7159,N_7736);
nor U8890 (N_8890,N_7555,N_7084);
and U8891 (N_8891,N_7794,N_7374);
and U8892 (N_8892,N_7009,N_7918);
and U8893 (N_8893,N_7963,N_7576);
nand U8894 (N_8894,N_7379,N_7954);
nor U8895 (N_8895,N_7293,N_7413);
xor U8896 (N_8896,N_7458,N_7684);
and U8897 (N_8897,N_7260,N_7654);
xor U8898 (N_8898,N_7902,N_7779);
nor U8899 (N_8899,N_7360,N_7537);
nand U8900 (N_8900,N_7227,N_7913);
or U8901 (N_8901,N_7267,N_7161);
and U8902 (N_8902,N_7543,N_7120);
and U8903 (N_8903,N_7625,N_7947);
xor U8904 (N_8904,N_7732,N_7515);
nor U8905 (N_8905,N_7667,N_7691);
and U8906 (N_8906,N_7911,N_7818);
nor U8907 (N_8907,N_7914,N_7597);
nand U8908 (N_8908,N_7522,N_7051);
or U8909 (N_8909,N_7529,N_7176);
and U8910 (N_8910,N_7556,N_7352);
nor U8911 (N_8911,N_7209,N_7355);
nor U8912 (N_8912,N_7330,N_7527);
nor U8913 (N_8913,N_7051,N_7671);
and U8914 (N_8914,N_7213,N_7451);
nor U8915 (N_8915,N_7438,N_7795);
and U8916 (N_8916,N_7701,N_7218);
nor U8917 (N_8917,N_7616,N_7471);
and U8918 (N_8918,N_7028,N_7711);
or U8919 (N_8919,N_7113,N_7741);
or U8920 (N_8920,N_7354,N_7787);
xor U8921 (N_8921,N_7632,N_7389);
and U8922 (N_8922,N_7433,N_7530);
xnor U8923 (N_8923,N_7016,N_7414);
nand U8924 (N_8924,N_7767,N_7165);
xor U8925 (N_8925,N_7782,N_7086);
and U8926 (N_8926,N_7068,N_7235);
or U8927 (N_8927,N_7940,N_7714);
nand U8928 (N_8928,N_7830,N_7868);
nor U8929 (N_8929,N_7217,N_7478);
nor U8930 (N_8930,N_7630,N_7601);
or U8931 (N_8931,N_7704,N_7926);
and U8932 (N_8932,N_7305,N_7179);
nand U8933 (N_8933,N_7721,N_7495);
nor U8934 (N_8934,N_7394,N_7102);
xor U8935 (N_8935,N_7933,N_7480);
xor U8936 (N_8936,N_7169,N_7317);
nand U8937 (N_8937,N_7024,N_7916);
or U8938 (N_8938,N_7617,N_7932);
nor U8939 (N_8939,N_7408,N_7947);
nor U8940 (N_8940,N_7227,N_7510);
nand U8941 (N_8941,N_7833,N_7179);
nor U8942 (N_8942,N_7320,N_7699);
nor U8943 (N_8943,N_7762,N_7473);
or U8944 (N_8944,N_7016,N_7155);
nand U8945 (N_8945,N_7999,N_7385);
nand U8946 (N_8946,N_7868,N_7535);
nand U8947 (N_8947,N_7278,N_7271);
nor U8948 (N_8948,N_7926,N_7487);
and U8949 (N_8949,N_7099,N_7664);
or U8950 (N_8950,N_7019,N_7538);
and U8951 (N_8951,N_7173,N_7684);
nor U8952 (N_8952,N_7149,N_7528);
nand U8953 (N_8953,N_7183,N_7474);
and U8954 (N_8954,N_7086,N_7290);
or U8955 (N_8955,N_7726,N_7469);
nor U8956 (N_8956,N_7836,N_7963);
nand U8957 (N_8957,N_7907,N_7839);
nor U8958 (N_8958,N_7512,N_7114);
xnor U8959 (N_8959,N_7684,N_7482);
nand U8960 (N_8960,N_7073,N_7646);
nor U8961 (N_8961,N_7495,N_7783);
or U8962 (N_8962,N_7993,N_7251);
or U8963 (N_8963,N_7044,N_7674);
and U8964 (N_8964,N_7900,N_7567);
and U8965 (N_8965,N_7141,N_7162);
nand U8966 (N_8966,N_7697,N_7831);
and U8967 (N_8967,N_7148,N_7495);
nand U8968 (N_8968,N_7443,N_7218);
nor U8969 (N_8969,N_7698,N_7230);
xor U8970 (N_8970,N_7453,N_7501);
nand U8971 (N_8971,N_7052,N_7477);
nor U8972 (N_8972,N_7016,N_7474);
nand U8973 (N_8973,N_7969,N_7275);
or U8974 (N_8974,N_7445,N_7711);
xnor U8975 (N_8975,N_7783,N_7553);
nand U8976 (N_8976,N_7001,N_7580);
and U8977 (N_8977,N_7895,N_7171);
nor U8978 (N_8978,N_7020,N_7096);
nor U8979 (N_8979,N_7670,N_7195);
nand U8980 (N_8980,N_7849,N_7980);
nand U8981 (N_8981,N_7145,N_7454);
nor U8982 (N_8982,N_7765,N_7716);
xor U8983 (N_8983,N_7491,N_7514);
and U8984 (N_8984,N_7857,N_7540);
or U8985 (N_8985,N_7719,N_7750);
and U8986 (N_8986,N_7707,N_7288);
and U8987 (N_8987,N_7138,N_7001);
nand U8988 (N_8988,N_7432,N_7928);
nand U8989 (N_8989,N_7013,N_7026);
nor U8990 (N_8990,N_7242,N_7439);
and U8991 (N_8991,N_7544,N_7214);
or U8992 (N_8992,N_7403,N_7912);
nor U8993 (N_8993,N_7081,N_7747);
and U8994 (N_8994,N_7603,N_7036);
or U8995 (N_8995,N_7044,N_7977);
nor U8996 (N_8996,N_7254,N_7338);
nor U8997 (N_8997,N_7723,N_7557);
nor U8998 (N_8998,N_7262,N_7483);
xnor U8999 (N_8999,N_7352,N_7020);
or U9000 (N_9000,N_8577,N_8545);
nor U9001 (N_9001,N_8310,N_8556);
nand U9002 (N_9002,N_8026,N_8932);
xor U9003 (N_9003,N_8790,N_8377);
or U9004 (N_9004,N_8595,N_8172);
nand U9005 (N_9005,N_8159,N_8430);
nor U9006 (N_9006,N_8114,N_8324);
nor U9007 (N_9007,N_8848,N_8519);
nor U9008 (N_9008,N_8135,N_8754);
nor U9009 (N_9009,N_8220,N_8130);
or U9010 (N_9010,N_8642,N_8063);
nand U9011 (N_9011,N_8668,N_8024);
nor U9012 (N_9012,N_8355,N_8516);
and U9013 (N_9013,N_8412,N_8550);
nor U9014 (N_9014,N_8100,N_8632);
or U9015 (N_9015,N_8131,N_8404);
and U9016 (N_9016,N_8524,N_8558);
nand U9017 (N_9017,N_8985,N_8546);
and U9018 (N_9018,N_8693,N_8168);
or U9019 (N_9019,N_8941,N_8098);
nor U9020 (N_9020,N_8515,N_8297);
nor U9021 (N_9021,N_8224,N_8249);
xnor U9022 (N_9022,N_8443,N_8768);
nand U9023 (N_9023,N_8036,N_8256);
nor U9024 (N_9024,N_8433,N_8648);
and U9025 (N_9025,N_8822,N_8806);
and U9026 (N_9026,N_8216,N_8846);
nor U9027 (N_9027,N_8299,N_8563);
nand U9028 (N_9028,N_8839,N_8285);
nand U9029 (N_9029,N_8939,N_8905);
nor U9030 (N_9030,N_8475,N_8230);
nand U9031 (N_9031,N_8749,N_8725);
nand U9032 (N_9032,N_8920,N_8597);
nor U9033 (N_9033,N_8145,N_8742);
nor U9034 (N_9034,N_8535,N_8434);
nand U9035 (N_9035,N_8554,N_8091);
or U9036 (N_9036,N_8007,N_8841);
or U9037 (N_9037,N_8010,N_8469);
nor U9038 (N_9038,N_8017,N_8808);
and U9039 (N_9039,N_8077,N_8620);
and U9040 (N_9040,N_8153,N_8513);
or U9041 (N_9041,N_8237,N_8779);
or U9042 (N_9042,N_8660,N_8275);
xnor U9043 (N_9043,N_8991,N_8925);
nor U9044 (N_9044,N_8122,N_8889);
nand U9045 (N_9045,N_8626,N_8734);
and U9046 (N_9046,N_8700,N_8963);
nor U9047 (N_9047,N_8094,N_8476);
nand U9048 (N_9048,N_8041,N_8803);
xor U9049 (N_9049,N_8990,N_8858);
nor U9050 (N_9050,N_8929,N_8025);
nand U9051 (N_9051,N_8784,N_8820);
or U9052 (N_9052,N_8013,N_8246);
nand U9053 (N_9053,N_8138,N_8681);
and U9054 (N_9054,N_8588,N_8346);
nand U9055 (N_9055,N_8093,N_8211);
or U9056 (N_9056,N_8188,N_8079);
nand U9057 (N_9057,N_8793,N_8829);
or U9058 (N_9058,N_8951,N_8067);
and U9059 (N_9059,N_8826,N_8508);
or U9060 (N_9060,N_8694,N_8395);
and U9061 (N_9061,N_8902,N_8279);
nand U9062 (N_9062,N_8251,N_8520);
nor U9063 (N_9063,N_8360,N_8802);
or U9064 (N_9064,N_8402,N_8092);
nor U9065 (N_9065,N_8399,N_8727);
and U9066 (N_9066,N_8765,N_8776);
nand U9067 (N_9067,N_8591,N_8761);
nand U9068 (N_9068,N_8290,N_8322);
or U9069 (N_9069,N_8560,N_8181);
xor U9070 (N_9070,N_8624,N_8947);
nor U9071 (N_9071,N_8072,N_8193);
nand U9072 (N_9072,N_8612,N_8305);
and U9073 (N_9073,N_8328,N_8259);
and U9074 (N_9074,N_8167,N_8045);
nand U9075 (N_9075,N_8596,N_8174);
nand U9076 (N_9076,N_8446,N_8273);
nor U9077 (N_9077,N_8073,N_8052);
nor U9078 (N_9078,N_8622,N_8084);
or U9079 (N_9079,N_8277,N_8064);
or U9080 (N_9080,N_8125,N_8490);
nand U9081 (N_9081,N_8065,N_8762);
or U9082 (N_9082,N_8101,N_8325);
nor U9083 (N_9083,N_8018,N_8148);
and U9084 (N_9084,N_8714,N_8049);
nor U9085 (N_9085,N_8766,N_8787);
nor U9086 (N_9086,N_8182,N_8532);
nand U9087 (N_9087,N_8447,N_8382);
nand U9088 (N_9088,N_8928,N_8097);
or U9089 (N_9089,N_8995,N_8816);
and U9090 (N_9090,N_8547,N_8183);
and U9091 (N_9091,N_8175,N_8191);
and U9092 (N_9092,N_8002,N_8659);
and U9093 (N_9093,N_8397,N_8435);
and U9094 (N_9094,N_8926,N_8268);
and U9095 (N_9095,N_8239,N_8486);
and U9096 (N_9096,N_8702,N_8302);
nand U9097 (N_9097,N_8893,N_8599);
or U9098 (N_9098,N_8289,N_8194);
or U9099 (N_9099,N_8294,N_8717);
and U9100 (N_9100,N_8112,N_8387);
or U9101 (N_9101,N_8374,N_8407);
nor U9102 (N_9102,N_8497,N_8616);
or U9103 (N_9103,N_8821,N_8317);
xor U9104 (N_9104,N_8190,N_8150);
or U9105 (N_9105,N_8592,N_8353);
nand U9106 (N_9106,N_8804,N_8977);
and U9107 (N_9107,N_8605,N_8165);
nand U9108 (N_9108,N_8284,N_8772);
and U9109 (N_9109,N_8916,N_8785);
or U9110 (N_9110,N_8957,N_8586);
and U9111 (N_9111,N_8260,N_8186);
and U9112 (N_9112,N_8813,N_8640);
nor U9113 (N_9113,N_8738,N_8336);
nor U9114 (N_9114,N_8955,N_8223);
nand U9115 (N_9115,N_8231,N_8836);
or U9116 (N_9116,N_8937,N_8661);
nor U9117 (N_9117,N_8401,N_8933);
and U9118 (N_9118,N_8729,N_8409);
and U9119 (N_9119,N_8057,N_8488);
nand U9120 (N_9120,N_8370,N_8979);
nor U9121 (N_9121,N_8891,N_8931);
and U9122 (N_9122,N_8307,N_8743);
nor U9123 (N_9123,N_8048,N_8966);
nor U9124 (N_9124,N_8087,N_8202);
nor U9125 (N_9125,N_8033,N_8894);
nand U9126 (N_9126,N_8203,N_8365);
xnor U9127 (N_9127,N_8144,N_8917);
and U9128 (N_9128,N_8332,N_8060);
or U9129 (N_9129,N_8562,N_8993);
xnor U9130 (N_9130,N_8958,N_8467);
and U9131 (N_9131,N_8451,N_8671);
and U9132 (N_9132,N_8331,N_8236);
nor U9133 (N_9133,N_8831,N_8865);
or U9134 (N_9134,N_8528,N_8206);
nor U9135 (N_9135,N_8016,N_8716);
nand U9136 (N_9136,N_8031,N_8732);
and U9137 (N_9137,N_8089,N_8708);
xor U9138 (N_9138,N_8484,N_8980);
nand U9139 (N_9139,N_8021,N_8276);
or U9140 (N_9140,N_8567,N_8267);
nand U9141 (N_9141,N_8767,N_8509);
nor U9142 (N_9142,N_8908,N_8350);
and U9143 (N_9143,N_8898,N_8888);
nor U9144 (N_9144,N_8326,N_8684);
and U9145 (N_9145,N_8054,N_8911);
xnor U9146 (N_9146,N_8915,N_8868);
and U9147 (N_9147,N_8924,N_8886);
xor U9148 (N_9148,N_8649,N_8870);
or U9149 (N_9149,N_8356,N_8169);
nand U9150 (N_9150,N_8644,N_8495);
xnor U9151 (N_9151,N_8300,N_8359);
or U9152 (N_9152,N_8835,N_8587);
nor U9153 (N_9153,N_8003,N_8367);
and U9154 (N_9154,N_8158,N_8847);
nand U9155 (N_9155,N_8358,N_8436);
nor U9156 (N_9156,N_8155,N_8132);
nand U9157 (N_9157,N_8631,N_8071);
nand U9158 (N_9158,N_8949,N_8780);
or U9159 (N_9159,N_8306,N_8243);
nand U9160 (N_9160,N_8537,N_8456);
nand U9161 (N_9161,N_8964,N_8445);
nand U9162 (N_9162,N_8895,N_8424);
nand U9163 (N_9163,N_8873,N_8383);
nor U9164 (N_9164,N_8050,N_8037);
or U9165 (N_9165,N_8076,N_8976);
nand U9166 (N_9166,N_8565,N_8392);
nor U9167 (N_9167,N_8861,N_8697);
or U9168 (N_9168,N_8857,N_8498);
or U9169 (N_9169,N_8607,N_8335);
and U9170 (N_9170,N_8971,N_8248);
nand U9171 (N_9171,N_8162,N_8914);
nor U9172 (N_9172,N_8582,N_8102);
and U9173 (N_9173,N_8442,N_8126);
nand U9174 (N_9174,N_8166,N_8099);
xnor U9175 (N_9175,N_8735,N_8280);
nand U9176 (N_9176,N_8313,N_8968);
nand U9177 (N_9177,N_8584,N_8421);
xnor U9178 (N_9178,N_8856,N_8386);
or U9179 (N_9179,N_8349,N_8000);
nand U9180 (N_9180,N_8849,N_8919);
and U9181 (N_9181,N_8011,N_8176);
nand U9182 (N_9182,N_8111,N_8090);
nand U9183 (N_9183,N_8527,N_8628);
nor U9184 (N_9184,N_8363,N_8461);
nand U9185 (N_9185,N_8217,N_8163);
and U9186 (N_9186,N_8376,N_8266);
nor U9187 (N_9187,N_8879,N_8777);
and U9188 (N_9188,N_8636,N_8759);
and U9189 (N_9189,N_8811,N_8773);
nor U9190 (N_9190,N_8637,N_8380);
nor U9191 (N_9191,N_8238,N_8338);
or U9192 (N_9192,N_8627,N_8311);
nor U9193 (N_9193,N_8405,N_8487);
or U9194 (N_9194,N_8687,N_8062);
or U9195 (N_9195,N_8798,N_8227);
nand U9196 (N_9196,N_8910,N_8196);
nand U9197 (N_9197,N_8385,N_8746);
nand U9198 (N_9198,N_8723,N_8701);
nand U9199 (N_9199,N_8411,N_8420);
and U9200 (N_9200,N_8470,N_8719);
nand U9201 (N_9201,N_8264,N_8344);
and U9202 (N_9202,N_8579,N_8250);
and U9203 (N_9203,N_8680,N_8974);
and U9204 (N_9204,N_8157,N_8593);
and U9205 (N_9205,N_8568,N_8432);
and U9206 (N_9206,N_8789,N_8786);
and U9207 (N_9207,N_8333,N_8117);
or U9208 (N_9208,N_8666,N_8427);
or U9209 (N_9209,N_8140,N_8345);
or U9210 (N_9210,N_8123,N_8676);
nor U9211 (N_9211,N_8961,N_8733);
nand U9212 (N_9212,N_8118,N_8909);
or U9213 (N_9213,N_8161,N_8526);
or U9214 (N_9214,N_8113,N_8160);
or U9215 (N_9215,N_8828,N_8884);
and U9216 (N_9216,N_8241,N_8748);
or U9217 (N_9217,N_8457,N_8270);
and U9218 (N_9218,N_8598,N_8507);
and U9219 (N_9219,N_8896,N_8996);
nand U9220 (N_9220,N_8988,N_8199);
nand U9221 (N_9221,N_8824,N_8388);
xnor U9222 (N_9222,N_8418,N_8055);
nand U9223 (N_9223,N_8146,N_8935);
or U9224 (N_9224,N_8170,N_8540);
nor U9225 (N_9225,N_8617,N_8791);
and U9226 (N_9226,N_8450,N_8219);
or U9227 (N_9227,N_8136,N_8070);
or U9228 (N_9228,N_8110,N_8818);
or U9229 (N_9229,N_8066,N_8959);
and U9230 (N_9230,N_8542,N_8492);
nor U9231 (N_9231,N_8291,N_8690);
xnor U9232 (N_9232,N_8726,N_8274);
nand U9233 (N_9233,N_8827,N_8329);
nand U9234 (N_9234,N_8878,N_8288);
xor U9235 (N_9235,N_8585,N_8533);
nor U9236 (N_9236,N_8269,N_8623);
xnor U9237 (N_9237,N_8272,N_8778);
nor U9238 (N_9238,N_8023,N_8473);
xor U9239 (N_9239,N_8678,N_8496);
nor U9240 (N_9240,N_8244,N_8059);
or U9241 (N_9241,N_8752,N_8453);
nor U9242 (N_9242,N_8390,N_8679);
nand U9243 (N_9243,N_8147,N_8788);
or U9244 (N_9244,N_8740,N_8711);
nor U9245 (N_9245,N_8866,N_8107);
or U9246 (N_9246,N_8214,N_8830);
nand U9247 (N_9247,N_8369,N_8208);
nand U9248 (N_9248,N_8463,N_8225);
nand U9249 (N_9249,N_8531,N_8423);
or U9250 (N_9250,N_8757,N_8795);
xnor U9251 (N_9251,N_8658,N_8228);
and U9252 (N_9252,N_8232,N_8669);
xor U9253 (N_9253,N_8173,N_8521);
xnor U9254 (N_9254,N_8095,N_8954);
and U9255 (N_9255,N_8152,N_8184);
nand U9256 (N_9256,N_8698,N_8695);
nand U9257 (N_9257,N_8403,N_8863);
nor U9258 (N_9258,N_8664,N_8321);
nor U9259 (N_9259,N_8200,N_8364);
and U9260 (N_9260,N_8728,N_8984);
nand U9261 (N_9261,N_8298,N_8722);
xnor U9262 (N_9262,N_8887,N_8471);
or U9263 (N_9263,N_8851,N_8852);
nor U9264 (N_9264,N_8938,N_8794);
or U9265 (N_9265,N_8536,N_8969);
and U9266 (N_9266,N_8154,N_8769);
or U9267 (N_9267,N_8549,N_8685);
nand U9268 (N_9268,N_8215,N_8973);
nor U9269 (N_9269,N_8553,N_8005);
nand U9270 (N_9270,N_8361,N_8141);
and U9271 (N_9271,N_8569,N_8682);
nor U9272 (N_9272,N_8602,N_8396);
xnor U9273 (N_9273,N_8192,N_8337);
and U9274 (N_9274,N_8647,N_8750);
nor U9275 (N_9275,N_8718,N_8240);
and U9276 (N_9276,N_8234,N_8096);
nor U9277 (N_9277,N_8201,N_8559);
or U9278 (N_9278,N_8491,N_8982);
nand U9279 (N_9279,N_8665,N_8815);
and U9280 (N_9280,N_8384,N_8633);
xnor U9281 (N_9281,N_8730,N_8775);
nand U9282 (N_9282,N_8229,N_8737);
xor U9283 (N_9283,N_8872,N_8838);
xnor U9284 (N_9284,N_8254,N_8198);
nand U9285 (N_9285,N_8667,N_8663);
or U9286 (N_9286,N_8416,N_8843);
nor U9287 (N_9287,N_8946,N_8504);
or U9288 (N_9288,N_8810,N_8572);
and U9289 (N_9289,N_8673,N_8287);
xnor U9290 (N_9290,N_8061,N_8656);
nor U9291 (N_9291,N_8575,N_8342);
nand U9292 (N_9292,N_8340,N_8389);
and U9293 (N_9293,N_8652,N_8137);
or U9294 (N_9294,N_8373,N_8871);
or U9295 (N_9295,N_8869,N_8736);
xor U9296 (N_9296,N_8247,N_8797);
and U9297 (N_9297,N_8042,N_8253);
nor U9298 (N_9298,N_8109,N_8987);
or U9299 (N_9299,N_8371,N_8850);
nor U9300 (N_9300,N_8124,N_8712);
nand U9301 (N_9301,N_8429,N_8792);
nand U9302 (N_9302,N_8195,N_8295);
nand U9303 (N_9303,N_8756,N_8960);
and U9304 (N_9304,N_8004,N_8043);
nor U9305 (N_9305,N_8417,N_8413);
or U9306 (N_9306,N_8760,N_8351);
and U9307 (N_9307,N_8372,N_8603);
nand U9308 (N_9308,N_8710,N_8594);
and U9309 (N_9309,N_8845,N_8468);
xor U9310 (N_9310,N_8012,N_8511);
and U9311 (N_9311,N_8460,N_8454);
and U9312 (N_9312,N_8561,N_8103);
nand U9313 (N_9313,N_8581,N_8543);
nor U9314 (N_9314,N_8842,N_8529);
nor U9315 (N_9315,N_8482,N_8720);
xnor U9316 (N_9316,N_8352,N_8844);
and U9317 (N_9317,N_8641,N_8539);
and U9318 (N_9318,N_8178,N_8621);
or U9319 (N_9319,N_8989,N_8151);
or U9320 (N_9320,N_8518,N_8945);
or U9321 (N_9321,N_8781,N_8994);
nand U9322 (N_9322,N_8783,N_8271);
or U9323 (N_9323,N_8962,N_8292);
nor U9324 (N_9324,N_8646,N_8483);
or U9325 (N_9325,N_8278,N_8880);
nand U9326 (N_9326,N_8944,N_8771);
and U9327 (N_9327,N_8213,N_8907);
nor U9328 (N_9328,N_8601,N_8020);
xor U9329 (N_9329,N_8009,N_8505);
nor U9330 (N_9330,N_8134,N_8265);
and U9331 (N_9331,N_8751,N_8035);
nand U9332 (N_9332,N_8398,N_8943);
or U9333 (N_9333,N_8502,N_8323);
or U9334 (N_9334,N_8721,N_8108);
and U9335 (N_9335,N_8840,N_8799);
nand U9336 (N_9336,N_8674,N_8221);
nor U9337 (N_9337,N_8431,N_8205);
or U9338 (N_9338,N_8347,N_8074);
nor U9339 (N_9339,N_8747,N_8449);
nor U9340 (N_9340,N_8304,N_8653);
and U9341 (N_9341,N_8997,N_8800);
and U9342 (N_9342,N_8044,N_8530);
nor U9343 (N_9343,N_8867,N_8245);
or U9344 (N_9344,N_8466,N_8686);
nor U9345 (N_9345,N_8948,N_8334);
xor U9346 (N_9346,N_8032,N_8881);
nor U9347 (N_9347,N_8222,N_8480);
or U9348 (N_9348,N_8606,N_8139);
and U9349 (N_9349,N_8426,N_8316);
xnor U9350 (N_9350,N_8801,N_8459);
nor U9351 (N_9351,N_8741,N_8876);
nand U9352 (N_9352,N_8282,N_8814);
nand U9353 (N_9353,N_8512,N_8499);
or U9354 (N_9354,N_8164,N_8904);
or U9355 (N_9355,N_8327,N_8986);
nand U9356 (N_9356,N_8051,N_8934);
and U9357 (N_9357,N_8923,N_8312);
and U9358 (N_9358,N_8992,N_8551);
or U9359 (N_9359,N_8864,N_8489);
nor U9360 (N_9360,N_8083,N_8209);
or U9361 (N_9361,N_8133,N_8825);
and U9362 (N_9362,N_8918,N_8913);
xnor U9363 (N_9363,N_8308,N_8422);
xnor U9364 (N_9364,N_8315,N_8912);
nand U9365 (N_9365,N_8252,N_8437);
or U9366 (N_9366,N_8425,N_8029);
or U9367 (N_9367,N_8303,N_8465);
or U9368 (N_9368,N_8823,N_8877);
nor U9369 (N_9369,N_8862,N_8544);
and U9370 (N_9370,N_8965,N_8391);
and U9371 (N_9371,N_8998,N_8441);
xor U9372 (N_9372,N_8807,N_8408);
nand U9373 (N_9373,N_8739,N_8809);
nand U9374 (N_9374,N_8854,N_8406);
nand U9375 (N_9375,N_8650,N_8745);
xor U9376 (N_9376,N_8981,N_8900);
or U9377 (N_9377,N_8080,N_8474);
and U9378 (N_9378,N_8655,N_8040);
nor U9379 (N_9379,N_8242,N_8218);
or U9380 (N_9380,N_8506,N_8187);
and U9381 (N_9381,N_8683,N_8419);
nand U9382 (N_9382,N_8930,N_8853);
and U9383 (N_9383,N_8263,N_8571);
nand U9384 (N_9384,N_8613,N_8635);
nand U9385 (N_9385,N_8614,N_8258);
nor U9386 (N_9386,N_8534,N_8782);
nand U9387 (N_9387,N_8953,N_8705);
and U9388 (N_9388,N_8608,N_8481);
or U9389 (N_9389,N_8501,N_8378);
and U9390 (N_9390,N_8262,N_8833);
or U9391 (N_9391,N_8672,N_8039);
nand U9392 (N_9392,N_8204,N_8197);
nor U9393 (N_9393,N_8610,N_8257);
nand U9394 (N_9394,N_8611,N_8691);
nor U9395 (N_9395,N_8022,N_8715);
xor U9396 (N_9396,N_8662,N_8086);
and U9397 (N_9397,N_8458,N_8975);
or U9398 (N_9398,N_8006,N_8983);
xor U9399 (N_9399,N_8171,N_8320);
nand U9400 (N_9400,N_8566,N_8514);
or U9401 (N_9401,N_8106,N_8675);
nor U9402 (N_9402,N_8921,N_8015);
or U9403 (N_9403,N_8085,N_8970);
nor U9404 (N_9404,N_8127,N_8394);
and U9405 (N_9405,N_8882,N_8819);
or U9406 (N_9406,N_8341,N_8770);
nor U9407 (N_9407,N_8455,N_8570);
nor U9408 (N_9408,N_8576,N_8834);
nor U9409 (N_9409,N_8281,N_8428);
nor U9410 (N_9410,N_8942,N_8552);
nand U9411 (N_9411,N_8899,N_8261);
and U9412 (N_9412,N_8523,N_8817);
or U9413 (N_9413,N_8859,N_8143);
nor U9414 (N_9414,N_8081,N_8255);
nor U9415 (N_9415,N_8439,N_8479);
and U9416 (N_9416,N_8472,N_8517);
nand U9417 (N_9417,N_8967,N_8699);
and U9418 (N_9418,N_8615,N_8522);
and U9419 (N_9419,N_8314,N_8832);
or U9420 (N_9420,N_8589,N_8047);
nand U9421 (N_9421,N_8645,N_8703);
nand U9422 (N_9422,N_8058,N_8286);
or U9423 (N_9423,N_8758,N_8713);
xor U9424 (N_9424,N_8226,N_8573);
nor U9425 (N_9425,N_8115,N_8046);
nand U9426 (N_9426,N_8555,N_8812);
nand U9427 (N_9427,N_8643,N_8557);
nor U9428 (N_9428,N_8903,N_8019);
or U9429 (N_9429,N_8874,N_8452);
and U9430 (N_9430,N_8574,N_8142);
nor U9431 (N_9431,N_8189,N_8906);
and U9432 (N_9432,N_8008,N_8319);
nand U9433 (N_9433,N_8330,N_8493);
nand U9434 (N_9434,N_8283,N_8583);
xnor U9435 (N_9435,N_8548,N_8120);
nor U9436 (N_9436,N_8414,N_8477);
or U9437 (N_9437,N_8901,N_8056);
xnor U9438 (N_9438,N_8538,N_8972);
xnor U9439 (N_9439,N_8639,N_8707);
nor U9440 (N_9440,N_8897,N_8410);
nand U9441 (N_9441,N_8485,N_8510);
nor U9442 (N_9442,N_8379,N_8580);
and U9443 (N_9443,N_8805,N_8128);
nor U9444 (N_9444,N_8600,N_8689);
nor U9445 (N_9445,N_8922,N_8235);
nand U9446 (N_9446,N_8629,N_8354);
and U9447 (N_9447,N_8651,N_8415);
and U9448 (N_9448,N_8233,N_8362);
nor U9449 (N_9449,N_8860,N_8619);
nor U9450 (N_9450,N_8952,N_8440);
nand U9451 (N_9451,N_8375,N_8069);
or U9452 (N_9452,N_8696,N_8001);
nand U9453 (N_9453,N_8763,N_8940);
nor U9454 (N_9454,N_8503,N_8654);
nor U9455 (N_9455,N_8119,N_8692);
and U9456 (N_9456,N_8706,N_8764);
nor U9457 (N_9457,N_8885,N_8149);
nor U9458 (N_9458,N_8630,N_8053);
and U9459 (N_9459,N_8883,N_8014);
xnor U9460 (N_9460,N_8293,N_8634);
nand U9461 (N_9461,N_8709,N_8731);
nor U9462 (N_9462,N_8936,N_8744);
or U9463 (N_9463,N_8500,N_8366);
nand U9464 (N_9464,N_8381,N_8075);
nand U9465 (N_9465,N_8185,N_8927);
nand U9466 (N_9466,N_8724,N_8339);
xnor U9467 (N_9467,N_8638,N_8564);
or U9468 (N_9468,N_8301,N_8950);
nand U9469 (N_9469,N_8670,N_8525);
or U9470 (N_9470,N_8027,N_8400);
nand U9471 (N_9471,N_8179,N_8755);
or U9472 (N_9472,N_8657,N_8541);
nand U9473 (N_9473,N_8688,N_8774);
xor U9474 (N_9474,N_8393,N_8448);
nand U9475 (N_9475,N_8038,N_8590);
xnor U9476 (N_9476,N_8104,N_8494);
or U9477 (N_9477,N_8978,N_8875);
nor U9478 (N_9478,N_8892,N_8604);
and U9479 (N_9479,N_8890,N_8343);
and U9480 (N_9480,N_8082,N_8704);
or U9481 (N_9481,N_8034,N_8156);
or U9482 (N_9482,N_8677,N_8368);
xnor U9483 (N_9483,N_8309,N_8444);
and U9484 (N_9484,N_8121,N_8129);
nor U9485 (N_9485,N_8068,N_8207);
xnor U9486 (N_9486,N_8028,N_8478);
xnor U9487 (N_9487,N_8855,N_8625);
nor U9488 (N_9488,N_8999,N_8212);
nor U9489 (N_9489,N_8464,N_8357);
xnor U9490 (N_9490,N_8796,N_8618);
and U9491 (N_9491,N_8105,N_8116);
or U9492 (N_9492,N_8030,N_8753);
and U9493 (N_9493,N_8078,N_8609);
and U9494 (N_9494,N_8177,N_8348);
nor U9495 (N_9495,N_8210,N_8578);
or U9496 (N_9496,N_8438,N_8088);
or U9497 (N_9497,N_8296,N_8318);
nor U9498 (N_9498,N_8180,N_8462);
nor U9499 (N_9499,N_8837,N_8956);
or U9500 (N_9500,N_8433,N_8478);
nor U9501 (N_9501,N_8388,N_8427);
xor U9502 (N_9502,N_8646,N_8757);
nor U9503 (N_9503,N_8510,N_8556);
nand U9504 (N_9504,N_8612,N_8596);
and U9505 (N_9505,N_8121,N_8891);
nand U9506 (N_9506,N_8998,N_8054);
and U9507 (N_9507,N_8172,N_8221);
or U9508 (N_9508,N_8249,N_8939);
nand U9509 (N_9509,N_8875,N_8691);
nand U9510 (N_9510,N_8058,N_8682);
nand U9511 (N_9511,N_8564,N_8800);
xnor U9512 (N_9512,N_8003,N_8815);
and U9513 (N_9513,N_8331,N_8514);
nand U9514 (N_9514,N_8103,N_8741);
nor U9515 (N_9515,N_8611,N_8820);
or U9516 (N_9516,N_8655,N_8008);
and U9517 (N_9517,N_8013,N_8617);
nor U9518 (N_9518,N_8224,N_8566);
or U9519 (N_9519,N_8809,N_8828);
xor U9520 (N_9520,N_8722,N_8674);
and U9521 (N_9521,N_8830,N_8720);
nand U9522 (N_9522,N_8322,N_8054);
and U9523 (N_9523,N_8329,N_8155);
nor U9524 (N_9524,N_8743,N_8774);
or U9525 (N_9525,N_8846,N_8551);
or U9526 (N_9526,N_8538,N_8278);
xnor U9527 (N_9527,N_8369,N_8213);
or U9528 (N_9528,N_8644,N_8477);
nor U9529 (N_9529,N_8764,N_8716);
and U9530 (N_9530,N_8969,N_8232);
xor U9531 (N_9531,N_8820,N_8208);
and U9532 (N_9532,N_8006,N_8531);
nor U9533 (N_9533,N_8710,N_8301);
nand U9534 (N_9534,N_8576,N_8700);
nand U9535 (N_9535,N_8089,N_8959);
nand U9536 (N_9536,N_8769,N_8919);
nor U9537 (N_9537,N_8407,N_8375);
nor U9538 (N_9538,N_8579,N_8108);
or U9539 (N_9539,N_8378,N_8478);
nor U9540 (N_9540,N_8181,N_8352);
xor U9541 (N_9541,N_8792,N_8575);
and U9542 (N_9542,N_8670,N_8227);
nand U9543 (N_9543,N_8800,N_8809);
xor U9544 (N_9544,N_8079,N_8148);
nor U9545 (N_9545,N_8635,N_8077);
nor U9546 (N_9546,N_8982,N_8929);
nand U9547 (N_9547,N_8871,N_8281);
and U9548 (N_9548,N_8470,N_8288);
and U9549 (N_9549,N_8794,N_8066);
nand U9550 (N_9550,N_8722,N_8120);
and U9551 (N_9551,N_8880,N_8403);
nand U9552 (N_9552,N_8995,N_8751);
nand U9553 (N_9553,N_8417,N_8999);
and U9554 (N_9554,N_8551,N_8966);
xnor U9555 (N_9555,N_8590,N_8985);
nand U9556 (N_9556,N_8784,N_8258);
nor U9557 (N_9557,N_8570,N_8249);
or U9558 (N_9558,N_8581,N_8196);
or U9559 (N_9559,N_8860,N_8190);
nand U9560 (N_9560,N_8762,N_8466);
nand U9561 (N_9561,N_8099,N_8522);
and U9562 (N_9562,N_8266,N_8801);
or U9563 (N_9563,N_8768,N_8618);
nand U9564 (N_9564,N_8170,N_8793);
or U9565 (N_9565,N_8090,N_8634);
nor U9566 (N_9566,N_8974,N_8909);
xnor U9567 (N_9567,N_8142,N_8278);
or U9568 (N_9568,N_8331,N_8191);
xor U9569 (N_9569,N_8089,N_8752);
nor U9570 (N_9570,N_8314,N_8548);
or U9571 (N_9571,N_8266,N_8013);
xnor U9572 (N_9572,N_8314,N_8907);
and U9573 (N_9573,N_8139,N_8757);
or U9574 (N_9574,N_8778,N_8025);
or U9575 (N_9575,N_8141,N_8197);
xnor U9576 (N_9576,N_8895,N_8434);
nand U9577 (N_9577,N_8321,N_8753);
and U9578 (N_9578,N_8437,N_8722);
and U9579 (N_9579,N_8295,N_8182);
or U9580 (N_9580,N_8361,N_8456);
or U9581 (N_9581,N_8524,N_8251);
and U9582 (N_9582,N_8612,N_8310);
nor U9583 (N_9583,N_8895,N_8346);
and U9584 (N_9584,N_8358,N_8557);
nor U9585 (N_9585,N_8372,N_8706);
or U9586 (N_9586,N_8316,N_8073);
nor U9587 (N_9587,N_8986,N_8323);
nand U9588 (N_9588,N_8020,N_8737);
nor U9589 (N_9589,N_8345,N_8041);
nor U9590 (N_9590,N_8657,N_8506);
nand U9591 (N_9591,N_8161,N_8485);
or U9592 (N_9592,N_8134,N_8778);
nor U9593 (N_9593,N_8988,N_8909);
or U9594 (N_9594,N_8742,N_8164);
nand U9595 (N_9595,N_8452,N_8270);
and U9596 (N_9596,N_8361,N_8261);
nor U9597 (N_9597,N_8709,N_8116);
or U9598 (N_9598,N_8317,N_8331);
xor U9599 (N_9599,N_8358,N_8710);
and U9600 (N_9600,N_8321,N_8045);
and U9601 (N_9601,N_8343,N_8201);
and U9602 (N_9602,N_8029,N_8228);
or U9603 (N_9603,N_8187,N_8988);
nor U9604 (N_9604,N_8226,N_8788);
and U9605 (N_9605,N_8992,N_8257);
or U9606 (N_9606,N_8666,N_8764);
or U9607 (N_9607,N_8249,N_8900);
and U9608 (N_9608,N_8116,N_8435);
and U9609 (N_9609,N_8791,N_8349);
or U9610 (N_9610,N_8655,N_8518);
or U9611 (N_9611,N_8011,N_8418);
or U9612 (N_9612,N_8703,N_8052);
nor U9613 (N_9613,N_8401,N_8450);
nand U9614 (N_9614,N_8203,N_8102);
xor U9615 (N_9615,N_8088,N_8010);
and U9616 (N_9616,N_8980,N_8110);
nor U9617 (N_9617,N_8146,N_8772);
and U9618 (N_9618,N_8442,N_8720);
and U9619 (N_9619,N_8180,N_8110);
or U9620 (N_9620,N_8946,N_8774);
nor U9621 (N_9621,N_8750,N_8766);
and U9622 (N_9622,N_8317,N_8241);
and U9623 (N_9623,N_8221,N_8604);
or U9624 (N_9624,N_8830,N_8843);
or U9625 (N_9625,N_8979,N_8771);
nor U9626 (N_9626,N_8068,N_8642);
nor U9627 (N_9627,N_8169,N_8517);
nand U9628 (N_9628,N_8536,N_8661);
nand U9629 (N_9629,N_8620,N_8081);
nand U9630 (N_9630,N_8096,N_8416);
nor U9631 (N_9631,N_8871,N_8745);
nor U9632 (N_9632,N_8777,N_8818);
nand U9633 (N_9633,N_8179,N_8688);
and U9634 (N_9634,N_8666,N_8069);
xnor U9635 (N_9635,N_8579,N_8772);
nand U9636 (N_9636,N_8850,N_8608);
or U9637 (N_9637,N_8185,N_8300);
and U9638 (N_9638,N_8020,N_8544);
nand U9639 (N_9639,N_8004,N_8358);
nand U9640 (N_9640,N_8159,N_8326);
nor U9641 (N_9641,N_8507,N_8817);
and U9642 (N_9642,N_8037,N_8151);
nor U9643 (N_9643,N_8421,N_8945);
or U9644 (N_9644,N_8630,N_8551);
nand U9645 (N_9645,N_8394,N_8807);
nand U9646 (N_9646,N_8686,N_8645);
nand U9647 (N_9647,N_8304,N_8218);
nor U9648 (N_9648,N_8096,N_8106);
nor U9649 (N_9649,N_8424,N_8218);
nor U9650 (N_9650,N_8320,N_8110);
and U9651 (N_9651,N_8854,N_8484);
nand U9652 (N_9652,N_8657,N_8233);
nor U9653 (N_9653,N_8564,N_8213);
nor U9654 (N_9654,N_8437,N_8788);
nand U9655 (N_9655,N_8067,N_8318);
or U9656 (N_9656,N_8329,N_8126);
nand U9657 (N_9657,N_8388,N_8744);
and U9658 (N_9658,N_8742,N_8571);
and U9659 (N_9659,N_8379,N_8324);
xor U9660 (N_9660,N_8583,N_8302);
nor U9661 (N_9661,N_8403,N_8727);
and U9662 (N_9662,N_8634,N_8789);
nand U9663 (N_9663,N_8144,N_8824);
nor U9664 (N_9664,N_8392,N_8995);
and U9665 (N_9665,N_8737,N_8489);
or U9666 (N_9666,N_8833,N_8322);
or U9667 (N_9667,N_8080,N_8112);
and U9668 (N_9668,N_8983,N_8895);
and U9669 (N_9669,N_8624,N_8509);
nand U9670 (N_9670,N_8866,N_8974);
and U9671 (N_9671,N_8006,N_8612);
nor U9672 (N_9672,N_8459,N_8221);
and U9673 (N_9673,N_8957,N_8699);
or U9674 (N_9674,N_8640,N_8594);
or U9675 (N_9675,N_8433,N_8578);
nand U9676 (N_9676,N_8229,N_8709);
nor U9677 (N_9677,N_8328,N_8340);
and U9678 (N_9678,N_8076,N_8378);
and U9679 (N_9679,N_8382,N_8728);
nand U9680 (N_9680,N_8452,N_8124);
nor U9681 (N_9681,N_8083,N_8861);
and U9682 (N_9682,N_8602,N_8423);
nand U9683 (N_9683,N_8650,N_8532);
xnor U9684 (N_9684,N_8832,N_8105);
and U9685 (N_9685,N_8525,N_8936);
nand U9686 (N_9686,N_8170,N_8226);
nor U9687 (N_9687,N_8525,N_8449);
or U9688 (N_9688,N_8404,N_8840);
nor U9689 (N_9689,N_8066,N_8145);
or U9690 (N_9690,N_8130,N_8899);
nor U9691 (N_9691,N_8355,N_8013);
nand U9692 (N_9692,N_8952,N_8939);
or U9693 (N_9693,N_8469,N_8062);
nor U9694 (N_9694,N_8002,N_8354);
or U9695 (N_9695,N_8405,N_8534);
nand U9696 (N_9696,N_8702,N_8319);
and U9697 (N_9697,N_8014,N_8433);
nor U9698 (N_9698,N_8674,N_8469);
xor U9699 (N_9699,N_8780,N_8140);
nor U9700 (N_9700,N_8103,N_8510);
xor U9701 (N_9701,N_8786,N_8453);
nor U9702 (N_9702,N_8968,N_8374);
and U9703 (N_9703,N_8321,N_8938);
nand U9704 (N_9704,N_8704,N_8517);
nor U9705 (N_9705,N_8392,N_8174);
or U9706 (N_9706,N_8479,N_8518);
and U9707 (N_9707,N_8036,N_8613);
nor U9708 (N_9708,N_8035,N_8689);
or U9709 (N_9709,N_8322,N_8162);
or U9710 (N_9710,N_8426,N_8711);
nor U9711 (N_9711,N_8141,N_8348);
and U9712 (N_9712,N_8325,N_8516);
and U9713 (N_9713,N_8367,N_8140);
nand U9714 (N_9714,N_8364,N_8190);
nor U9715 (N_9715,N_8059,N_8980);
and U9716 (N_9716,N_8567,N_8717);
or U9717 (N_9717,N_8560,N_8498);
nand U9718 (N_9718,N_8625,N_8500);
nand U9719 (N_9719,N_8467,N_8914);
and U9720 (N_9720,N_8776,N_8873);
and U9721 (N_9721,N_8168,N_8853);
or U9722 (N_9722,N_8457,N_8894);
nor U9723 (N_9723,N_8147,N_8196);
and U9724 (N_9724,N_8772,N_8602);
or U9725 (N_9725,N_8940,N_8050);
and U9726 (N_9726,N_8982,N_8337);
nor U9727 (N_9727,N_8551,N_8009);
or U9728 (N_9728,N_8543,N_8326);
nand U9729 (N_9729,N_8364,N_8529);
or U9730 (N_9730,N_8277,N_8402);
nand U9731 (N_9731,N_8701,N_8666);
or U9732 (N_9732,N_8301,N_8952);
and U9733 (N_9733,N_8868,N_8394);
and U9734 (N_9734,N_8798,N_8283);
nand U9735 (N_9735,N_8238,N_8430);
nor U9736 (N_9736,N_8481,N_8234);
nand U9737 (N_9737,N_8027,N_8046);
and U9738 (N_9738,N_8266,N_8574);
nand U9739 (N_9739,N_8489,N_8705);
or U9740 (N_9740,N_8154,N_8148);
nor U9741 (N_9741,N_8409,N_8656);
or U9742 (N_9742,N_8409,N_8714);
and U9743 (N_9743,N_8082,N_8667);
or U9744 (N_9744,N_8272,N_8922);
nand U9745 (N_9745,N_8952,N_8513);
nor U9746 (N_9746,N_8751,N_8274);
nand U9747 (N_9747,N_8016,N_8912);
or U9748 (N_9748,N_8782,N_8751);
and U9749 (N_9749,N_8730,N_8379);
or U9750 (N_9750,N_8794,N_8669);
nand U9751 (N_9751,N_8020,N_8099);
nand U9752 (N_9752,N_8888,N_8737);
xnor U9753 (N_9753,N_8442,N_8875);
nand U9754 (N_9754,N_8862,N_8389);
or U9755 (N_9755,N_8518,N_8252);
nor U9756 (N_9756,N_8628,N_8022);
and U9757 (N_9757,N_8324,N_8218);
xor U9758 (N_9758,N_8454,N_8464);
and U9759 (N_9759,N_8123,N_8946);
nand U9760 (N_9760,N_8406,N_8600);
or U9761 (N_9761,N_8780,N_8036);
and U9762 (N_9762,N_8418,N_8812);
nor U9763 (N_9763,N_8975,N_8796);
xnor U9764 (N_9764,N_8338,N_8011);
nor U9765 (N_9765,N_8247,N_8149);
nor U9766 (N_9766,N_8786,N_8812);
and U9767 (N_9767,N_8004,N_8366);
xnor U9768 (N_9768,N_8988,N_8951);
nand U9769 (N_9769,N_8628,N_8765);
nand U9770 (N_9770,N_8982,N_8368);
nand U9771 (N_9771,N_8659,N_8692);
or U9772 (N_9772,N_8108,N_8548);
nand U9773 (N_9773,N_8492,N_8546);
nor U9774 (N_9774,N_8295,N_8051);
nand U9775 (N_9775,N_8207,N_8319);
nand U9776 (N_9776,N_8171,N_8381);
nand U9777 (N_9777,N_8976,N_8029);
or U9778 (N_9778,N_8435,N_8106);
nor U9779 (N_9779,N_8953,N_8927);
xor U9780 (N_9780,N_8245,N_8025);
or U9781 (N_9781,N_8049,N_8351);
nor U9782 (N_9782,N_8689,N_8576);
or U9783 (N_9783,N_8896,N_8047);
or U9784 (N_9784,N_8455,N_8502);
nor U9785 (N_9785,N_8436,N_8142);
nor U9786 (N_9786,N_8385,N_8806);
nor U9787 (N_9787,N_8810,N_8373);
nand U9788 (N_9788,N_8716,N_8615);
nand U9789 (N_9789,N_8333,N_8192);
nor U9790 (N_9790,N_8238,N_8765);
and U9791 (N_9791,N_8085,N_8582);
nand U9792 (N_9792,N_8533,N_8323);
or U9793 (N_9793,N_8478,N_8349);
nand U9794 (N_9794,N_8745,N_8683);
or U9795 (N_9795,N_8481,N_8692);
or U9796 (N_9796,N_8556,N_8992);
nor U9797 (N_9797,N_8032,N_8217);
nor U9798 (N_9798,N_8734,N_8467);
nor U9799 (N_9799,N_8950,N_8288);
nand U9800 (N_9800,N_8609,N_8702);
and U9801 (N_9801,N_8866,N_8864);
and U9802 (N_9802,N_8285,N_8739);
or U9803 (N_9803,N_8776,N_8200);
and U9804 (N_9804,N_8919,N_8694);
nand U9805 (N_9805,N_8047,N_8412);
or U9806 (N_9806,N_8097,N_8154);
nand U9807 (N_9807,N_8826,N_8065);
xnor U9808 (N_9808,N_8915,N_8267);
or U9809 (N_9809,N_8753,N_8627);
nor U9810 (N_9810,N_8316,N_8797);
nor U9811 (N_9811,N_8636,N_8623);
or U9812 (N_9812,N_8220,N_8258);
or U9813 (N_9813,N_8009,N_8358);
xor U9814 (N_9814,N_8804,N_8475);
and U9815 (N_9815,N_8347,N_8539);
and U9816 (N_9816,N_8490,N_8396);
and U9817 (N_9817,N_8774,N_8540);
nand U9818 (N_9818,N_8180,N_8901);
and U9819 (N_9819,N_8934,N_8302);
xnor U9820 (N_9820,N_8992,N_8285);
and U9821 (N_9821,N_8256,N_8051);
or U9822 (N_9822,N_8033,N_8647);
xor U9823 (N_9823,N_8679,N_8275);
nand U9824 (N_9824,N_8846,N_8717);
nor U9825 (N_9825,N_8378,N_8442);
nand U9826 (N_9826,N_8954,N_8149);
nand U9827 (N_9827,N_8261,N_8137);
nand U9828 (N_9828,N_8036,N_8881);
and U9829 (N_9829,N_8876,N_8039);
or U9830 (N_9830,N_8801,N_8538);
or U9831 (N_9831,N_8625,N_8435);
nor U9832 (N_9832,N_8161,N_8308);
and U9833 (N_9833,N_8177,N_8223);
or U9834 (N_9834,N_8553,N_8523);
and U9835 (N_9835,N_8373,N_8231);
nor U9836 (N_9836,N_8001,N_8399);
nor U9837 (N_9837,N_8016,N_8058);
and U9838 (N_9838,N_8851,N_8039);
nor U9839 (N_9839,N_8026,N_8704);
or U9840 (N_9840,N_8143,N_8058);
nand U9841 (N_9841,N_8403,N_8283);
or U9842 (N_9842,N_8382,N_8279);
xnor U9843 (N_9843,N_8919,N_8698);
nor U9844 (N_9844,N_8966,N_8182);
and U9845 (N_9845,N_8427,N_8601);
nor U9846 (N_9846,N_8875,N_8453);
or U9847 (N_9847,N_8864,N_8088);
xnor U9848 (N_9848,N_8152,N_8564);
nor U9849 (N_9849,N_8318,N_8417);
nor U9850 (N_9850,N_8132,N_8303);
nand U9851 (N_9851,N_8431,N_8908);
nand U9852 (N_9852,N_8746,N_8808);
xor U9853 (N_9853,N_8448,N_8063);
nor U9854 (N_9854,N_8689,N_8210);
or U9855 (N_9855,N_8093,N_8718);
and U9856 (N_9856,N_8081,N_8151);
or U9857 (N_9857,N_8212,N_8356);
and U9858 (N_9858,N_8715,N_8501);
xor U9859 (N_9859,N_8335,N_8163);
nor U9860 (N_9860,N_8042,N_8776);
and U9861 (N_9861,N_8613,N_8281);
nor U9862 (N_9862,N_8924,N_8120);
xor U9863 (N_9863,N_8888,N_8300);
nand U9864 (N_9864,N_8421,N_8092);
nand U9865 (N_9865,N_8748,N_8969);
and U9866 (N_9866,N_8684,N_8481);
or U9867 (N_9867,N_8984,N_8074);
nand U9868 (N_9868,N_8941,N_8927);
and U9869 (N_9869,N_8841,N_8162);
nand U9870 (N_9870,N_8479,N_8273);
or U9871 (N_9871,N_8667,N_8906);
or U9872 (N_9872,N_8318,N_8688);
xor U9873 (N_9873,N_8931,N_8379);
nor U9874 (N_9874,N_8702,N_8010);
nor U9875 (N_9875,N_8954,N_8714);
nand U9876 (N_9876,N_8461,N_8081);
nand U9877 (N_9877,N_8184,N_8536);
nand U9878 (N_9878,N_8270,N_8265);
nand U9879 (N_9879,N_8095,N_8626);
or U9880 (N_9880,N_8786,N_8474);
and U9881 (N_9881,N_8601,N_8218);
and U9882 (N_9882,N_8932,N_8017);
and U9883 (N_9883,N_8424,N_8897);
or U9884 (N_9884,N_8183,N_8618);
and U9885 (N_9885,N_8493,N_8486);
or U9886 (N_9886,N_8097,N_8881);
or U9887 (N_9887,N_8757,N_8870);
or U9888 (N_9888,N_8838,N_8796);
nor U9889 (N_9889,N_8144,N_8287);
and U9890 (N_9890,N_8407,N_8996);
nor U9891 (N_9891,N_8582,N_8330);
or U9892 (N_9892,N_8114,N_8944);
nor U9893 (N_9893,N_8948,N_8048);
nor U9894 (N_9894,N_8620,N_8006);
xor U9895 (N_9895,N_8566,N_8721);
nand U9896 (N_9896,N_8091,N_8331);
nand U9897 (N_9897,N_8998,N_8743);
nand U9898 (N_9898,N_8598,N_8778);
nor U9899 (N_9899,N_8343,N_8623);
nor U9900 (N_9900,N_8551,N_8213);
and U9901 (N_9901,N_8741,N_8236);
or U9902 (N_9902,N_8170,N_8872);
xor U9903 (N_9903,N_8584,N_8499);
and U9904 (N_9904,N_8665,N_8993);
or U9905 (N_9905,N_8538,N_8750);
nor U9906 (N_9906,N_8369,N_8070);
and U9907 (N_9907,N_8526,N_8369);
xnor U9908 (N_9908,N_8459,N_8442);
xor U9909 (N_9909,N_8918,N_8125);
and U9910 (N_9910,N_8698,N_8396);
and U9911 (N_9911,N_8574,N_8662);
and U9912 (N_9912,N_8450,N_8954);
nand U9913 (N_9913,N_8592,N_8421);
xor U9914 (N_9914,N_8672,N_8311);
nor U9915 (N_9915,N_8380,N_8868);
nand U9916 (N_9916,N_8938,N_8154);
nor U9917 (N_9917,N_8199,N_8534);
and U9918 (N_9918,N_8771,N_8846);
xnor U9919 (N_9919,N_8335,N_8093);
xor U9920 (N_9920,N_8894,N_8147);
nand U9921 (N_9921,N_8628,N_8877);
or U9922 (N_9922,N_8478,N_8179);
nor U9923 (N_9923,N_8112,N_8738);
xnor U9924 (N_9924,N_8913,N_8633);
and U9925 (N_9925,N_8008,N_8563);
and U9926 (N_9926,N_8964,N_8906);
and U9927 (N_9927,N_8471,N_8446);
nor U9928 (N_9928,N_8159,N_8989);
and U9929 (N_9929,N_8354,N_8601);
or U9930 (N_9930,N_8954,N_8197);
or U9931 (N_9931,N_8999,N_8458);
nand U9932 (N_9932,N_8712,N_8357);
or U9933 (N_9933,N_8900,N_8768);
nand U9934 (N_9934,N_8287,N_8942);
nand U9935 (N_9935,N_8881,N_8028);
or U9936 (N_9936,N_8383,N_8358);
and U9937 (N_9937,N_8963,N_8485);
xnor U9938 (N_9938,N_8551,N_8969);
nand U9939 (N_9939,N_8360,N_8813);
or U9940 (N_9940,N_8450,N_8471);
nor U9941 (N_9941,N_8524,N_8739);
nand U9942 (N_9942,N_8676,N_8727);
and U9943 (N_9943,N_8286,N_8306);
and U9944 (N_9944,N_8474,N_8970);
and U9945 (N_9945,N_8932,N_8577);
nand U9946 (N_9946,N_8536,N_8199);
nor U9947 (N_9947,N_8078,N_8566);
nand U9948 (N_9948,N_8704,N_8088);
nor U9949 (N_9949,N_8966,N_8518);
xnor U9950 (N_9950,N_8778,N_8901);
nor U9951 (N_9951,N_8331,N_8378);
or U9952 (N_9952,N_8117,N_8432);
nand U9953 (N_9953,N_8647,N_8831);
and U9954 (N_9954,N_8882,N_8873);
nor U9955 (N_9955,N_8305,N_8655);
xor U9956 (N_9956,N_8153,N_8141);
xnor U9957 (N_9957,N_8689,N_8947);
and U9958 (N_9958,N_8014,N_8539);
nand U9959 (N_9959,N_8462,N_8988);
and U9960 (N_9960,N_8019,N_8848);
nor U9961 (N_9961,N_8009,N_8497);
or U9962 (N_9962,N_8314,N_8032);
and U9963 (N_9963,N_8841,N_8040);
xnor U9964 (N_9964,N_8475,N_8881);
and U9965 (N_9965,N_8663,N_8273);
or U9966 (N_9966,N_8473,N_8071);
or U9967 (N_9967,N_8723,N_8193);
nand U9968 (N_9968,N_8258,N_8872);
or U9969 (N_9969,N_8746,N_8640);
nand U9970 (N_9970,N_8485,N_8977);
nor U9971 (N_9971,N_8248,N_8514);
and U9972 (N_9972,N_8191,N_8416);
and U9973 (N_9973,N_8659,N_8965);
nor U9974 (N_9974,N_8966,N_8499);
nor U9975 (N_9975,N_8025,N_8422);
and U9976 (N_9976,N_8463,N_8935);
xor U9977 (N_9977,N_8773,N_8222);
or U9978 (N_9978,N_8345,N_8672);
and U9979 (N_9979,N_8979,N_8382);
or U9980 (N_9980,N_8253,N_8407);
nor U9981 (N_9981,N_8816,N_8243);
or U9982 (N_9982,N_8717,N_8768);
xnor U9983 (N_9983,N_8287,N_8313);
and U9984 (N_9984,N_8905,N_8544);
xnor U9985 (N_9985,N_8836,N_8433);
and U9986 (N_9986,N_8202,N_8792);
nand U9987 (N_9987,N_8341,N_8744);
xnor U9988 (N_9988,N_8313,N_8193);
and U9989 (N_9989,N_8258,N_8189);
and U9990 (N_9990,N_8129,N_8934);
nand U9991 (N_9991,N_8907,N_8649);
xnor U9992 (N_9992,N_8072,N_8154);
nand U9993 (N_9993,N_8357,N_8124);
nand U9994 (N_9994,N_8371,N_8676);
nand U9995 (N_9995,N_8212,N_8265);
xnor U9996 (N_9996,N_8777,N_8143);
or U9997 (N_9997,N_8714,N_8508);
or U9998 (N_9998,N_8887,N_8624);
nand U9999 (N_9999,N_8757,N_8357);
nor U10000 (N_10000,N_9119,N_9011);
nor U10001 (N_10001,N_9106,N_9688);
and U10002 (N_10002,N_9653,N_9853);
or U10003 (N_10003,N_9708,N_9901);
or U10004 (N_10004,N_9750,N_9188);
nand U10005 (N_10005,N_9087,N_9310);
or U10006 (N_10006,N_9848,N_9291);
nor U10007 (N_10007,N_9949,N_9892);
or U10008 (N_10008,N_9387,N_9487);
nand U10009 (N_10009,N_9572,N_9711);
or U10010 (N_10010,N_9797,N_9546);
or U10011 (N_10011,N_9985,N_9615);
nor U10012 (N_10012,N_9918,N_9331);
xor U10013 (N_10013,N_9995,N_9164);
nor U10014 (N_10014,N_9667,N_9607);
nand U10015 (N_10015,N_9184,N_9143);
xnor U10016 (N_10016,N_9495,N_9760);
nor U10017 (N_10017,N_9506,N_9254);
and U10018 (N_10018,N_9896,N_9205);
nor U10019 (N_10019,N_9062,N_9174);
nor U10020 (N_10020,N_9260,N_9704);
nand U10021 (N_10021,N_9695,N_9656);
and U10022 (N_10022,N_9341,N_9083);
nor U10023 (N_10023,N_9592,N_9599);
or U10024 (N_10024,N_9794,N_9420);
and U10025 (N_10025,N_9966,N_9044);
and U10026 (N_10026,N_9872,N_9582);
nor U10027 (N_10027,N_9718,N_9632);
nand U10028 (N_10028,N_9402,N_9281);
nor U10029 (N_10029,N_9411,N_9317);
nand U10030 (N_10030,N_9661,N_9746);
and U10031 (N_10031,N_9127,N_9871);
or U10032 (N_10032,N_9927,N_9752);
nor U10033 (N_10033,N_9758,N_9154);
nor U10034 (N_10034,N_9978,N_9518);
nor U10035 (N_10035,N_9601,N_9443);
and U10036 (N_10036,N_9404,N_9105);
nor U10037 (N_10037,N_9280,N_9671);
or U10038 (N_10038,N_9467,N_9771);
or U10039 (N_10039,N_9251,N_9041);
nor U10040 (N_10040,N_9840,N_9971);
or U10041 (N_10041,N_9496,N_9237);
or U10042 (N_10042,N_9815,N_9814);
and U10043 (N_10043,N_9446,N_9198);
nand U10044 (N_10044,N_9064,N_9159);
nand U10045 (N_10045,N_9297,N_9576);
nor U10046 (N_10046,N_9183,N_9456);
and U10047 (N_10047,N_9561,N_9086);
or U10048 (N_10048,N_9075,N_9644);
xnor U10049 (N_10049,N_9868,N_9444);
or U10050 (N_10050,N_9861,N_9664);
xnor U10051 (N_10051,N_9436,N_9415);
nor U10052 (N_10052,N_9318,N_9680);
nand U10053 (N_10053,N_9034,N_9977);
xor U10054 (N_10054,N_9604,N_9994);
nor U10055 (N_10055,N_9358,N_9796);
xnor U10056 (N_10056,N_9755,N_9545);
nand U10057 (N_10057,N_9395,N_9491);
nand U10058 (N_10058,N_9320,N_9278);
or U10059 (N_10059,N_9469,N_9339);
nand U10060 (N_10060,N_9306,N_9928);
nand U10061 (N_10061,N_9158,N_9334);
nor U10062 (N_10062,N_9267,N_9906);
xor U10063 (N_10063,N_9293,N_9890);
nand U10064 (N_10064,N_9922,N_9807);
nand U10065 (N_10065,N_9740,N_9130);
or U10066 (N_10066,N_9118,N_9882);
and U10067 (N_10067,N_9563,N_9282);
nand U10068 (N_10068,N_9145,N_9766);
and U10069 (N_10069,N_9846,N_9363);
xor U10070 (N_10070,N_9634,N_9388);
nor U10071 (N_10071,N_9976,N_9385);
nand U10072 (N_10072,N_9490,N_9253);
and U10073 (N_10073,N_9274,N_9960);
xnor U10074 (N_10074,N_9108,N_9213);
nor U10075 (N_10075,N_9268,N_9975);
nand U10076 (N_10076,N_9517,N_9246);
and U10077 (N_10077,N_9231,N_9125);
nor U10078 (N_10078,N_9991,N_9519);
or U10079 (N_10079,N_9099,N_9353);
nor U10080 (N_10080,N_9998,N_9825);
or U10081 (N_10081,N_9193,N_9612);
nand U10082 (N_10082,N_9935,N_9275);
and U10083 (N_10083,N_9453,N_9177);
or U10084 (N_10084,N_9379,N_9012);
or U10085 (N_10085,N_9539,N_9004);
nand U10086 (N_10086,N_9197,N_9629);
and U10087 (N_10087,N_9494,N_9273);
nand U10088 (N_10088,N_9532,N_9878);
nor U10089 (N_10089,N_9515,N_9685);
nor U10090 (N_10090,N_9191,N_9527);
nand U10091 (N_10091,N_9630,N_9945);
and U10092 (N_10092,N_9400,N_9781);
nand U10093 (N_10093,N_9575,N_9228);
xnor U10094 (N_10094,N_9031,N_9970);
nor U10095 (N_10095,N_9859,N_9431);
xor U10096 (N_10096,N_9899,N_9390);
or U10097 (N_10097,N_9126,N_9889);
or U10098 (N_10098,N_9298,N_9723);
and U10099 (N_10099,N_9556,N_9731);
xor U10100 (N_10100,N_9806,N_9510);
nor U10101 (N_10101,N_9397,N_9170);
nand U10102 (N_10102,N_9803,N_9425);
or U10103 (N_10103,N_9466,N_9157);
nor U10104 (N_10104,N_9732,N_9696);
and U10105 (N_10105,N_9788,N_9300);
and U10106 (N_10106,N_9547,N_9903);
and U10107 (N_10107,N_9951,N_9623);
nand U10108 (N_10108,N_9422,N_9015);
or U10109 (N_10109,N_9504,N_9429);
and U10110 (N_10110,N_9131,N_9920);
nor U10111 (N_10111,N_9374,N_9478);
and U10112 (N_10112,N_9335,N_9533);
nor U10113 (N_10113,N_9810,N_9540);
nand U10114 (N_10114,N_9338,N_9881);
nor U10115 (N_10115,N_9484,N_9912);
nand U10116 (N_10116,N_9659,N_9176);
or U10117 (N_10117,N_9663,N_9016);
nand U10118 (N_10118,N_9121,N_9964);
nand U10119 (N_10119,N_9097,N_9790);
or U10120 (N_10120,N_9409,N_9028);
and U10121 (N_10121,N_9835,N_9250);
xnor U10122 (N_10122,N_9285,N_9943);
xnor U10123 (N_10123,N_9590,N_9591);
nor U10124 (N_10124,N_9181,N_9324);
or U10125 (N_10125,N_9078,N_9336);
or U10126 (N_10126,N_9311,N_9203);
or U10127 (N_10127,N_9513,N_9141);
or U10128 (N_10128,N_9597,N_9873);
xor U10129 (N_10129,N_9096,N_9669);
or U10130 (N_10130,N_9554,N_9241);
or U10131 (N_10131,N_9081,N_9475);
nor U10132 (N_10132,N_9691,N_9401);
and U10133 (N_10133,N_9295,N_9089);
nand U10134 (N_10134,N_9212,N_9678);
nor U10135 (N_10135,N_9742,N_9812);
or U10136 (N_10136,N_9869,N_9646);
nor U10137 (N_10137,N_9792,N_9344);
xnor U10138 (N_10138,N_9931,N_9693);
nor U10139 (N_10139,N_9407,N_9703);
or U10140 (N_10140,N_9862,N_9548);
nor U10141 (N_10141,N_9571,N_9270);
nand U10142 (N_10142,N_9789,N_9464);
nor U10143 (N_10143,N_9944,N_9608);
and U10144 (N_10144,N_9000,N_9272);
and U10145 (N_10145,N_9541,N_9365);
or U10146 (N_10146,N_9216,N_9819);
or U10147 (N_10147,N_9486,N_9114);
or U10148 (N_10148,N_9018,N_9208);
nor U10149 (N_10149,N_9229,N_9783);
or U10150 (N_10150,N_9833,N_9605);
nand U10151 (N_10151,N_9117,N_9930);
or U10152 (N_10152,N_9969,N_9946);
nor U10153 (N_10153,N_9182,N_9025);
or U10154 (N_10154,N_9598,N_9611);
xor U10155 (N_10155,N_9152,N_9643);
and U10156 (N_10156,N_9354,N_9033);
xor U10157 (N_10157,N_9879,N_9776);
xor U10158 (N_10158,N_9080,N_9277);
nor U10159 (N_10159,N_9002,N_9568);
nor U10160 (N_10160,N_9479,N_9230);
xor U10161 (N_10161,N_9907,N_9256);
nand U10162 (N_10162,N_9367,N_9290);
xnor U10163 (N_10163,N_9116,N_9974);
or U10164 (N_10164,N_9902,N_9657);
nor U10165 (N_10165,N_9919,N_9037);
nand U10166 (N_10166,N_9304,N_9832);
xor U10167 (N_10167,N_9701,N_9574);
or U10168 (N_10168,N_9070,N_9512);
or U10169 (N_10169,N_9753,N_9421);
nand U10170 (N_10170,N_9606,N_9001);
nor U10171 (N_10171,N_9979,N_9150);
or U10172 (N_10172,N_9501,N_9850);
xor U10173 (N_10173,N_9102,N_9063);
or U10174 (N_10174,N_9795,N_9350);
nor U10175 (N_10175,N_9264,N_9791);
or U10176 (N_10176,N_9923,N_9124);
nand U10177 (N_10177,N_9136,N_9817);
nor U10178 (N_10178,N_9910,N_9968);
and U10179 (N_10179,N_9595,N_9639);
xnor U10180 (N_10180,N_9189,N_9507);
and U10181 (N_10181,N_9095,N_9645);
nor U10182 (N_10182,N_9067,N_9206);
nor U10183 (N_10183,N_9955,N_9594);
xnor U10184 (N_10184,N_9252,N_9628);
nand U10185 (N_10185,N_9244,N_9061);
xnor U10186 (N_10186,N_9477,N_9348);
nand U10187 (N_10187,N_9455,N_9148);
nand U10188 (N_10188,N_9900,N_9535);
nand U10189 (N_10189,N_9288,N_9043);
nor U10190 (N_10190,N_9194,N_9079);
and U10191 (N_10191,N_9305,N_9077);
xor U10192 (N_10192,N_9316,N_9356);
nor U10193 (N_10193,N_9508,N_9585);
nand U10194 (N_10194,N_9614,N_9672);
and U10195 (N_10195,N_9171,N_9658);
nand U10196 (N_10196,N_9555,N_9722);
and U10197 (N_10197,N_9523,N_9146);
or U10198 (N_10198,N_9626,N_9525);
nand U10199 (N_10199,N_9557,N_9567);
and U10200 (N_10200,N_9472,N_9550);
nor U10201 (N_10201,N_9767,N_9403);
and U10202 (N_10202,N_9471,N_9312);
nand U10203 (N_10203,N_9827,N_9751);
nand U10204 (N_10204,N_9168,N_9509);
and U10205 (N_10205,N_9874,N_9459);
or U10206 (N_10206,N_9588,N_9068);
nand U10207 (N_10207,N_9500,N_9824);
or U10208 (N_10208,N_9593,N_9738);
or U10209 (N_10209,N_9586,N_9142);
nor U10210 (N_10210,N_9589,N_9728);
and U10211 (N_10211,N_9552,N_9065);
nor U10212 (N_10212,N_9651,N_9497);
nand U10213 (N_10213,N_9138,N_9761);
nor U10214 (N_10214,N_9802,N_9689);
or U10215 (N_10215,N_9389,N_9670);
nor U10216 (N_10216,N_9715,N_9262);
nand U10217 (N_10217,N_9329,N_9377);
xnor U10218 (N_10218,N_9021,N_9369);
and U10219 (N_10219,N_9682,N_9036);
xor U10220 (N_10220,N_9725,N_9744);
nor U10221 (N_10221,N_9940,N_9035);
or U10222 (N_10222,N_9223,N_9772);
or U10223 (N_10223,N_9381,N_9294);
and U10224 (N_10224,N_9609,N_9449);
or U10225 (N_10225,N_9019,N_9332);
nand U10226 (N_10226,N_9424,N_9764);
and U10227 (N_10227,N_9573,N_9782);
and U10228 (N_10228,N_9352,N_9362);
and U10229 (N_10229,N_9405,N_9343);
nor U10230 (N_10230,N_9351,N_9112);
nand U10231 (N_10231,N_9877,N_9690);
nand U10232 (N_10232,N_9412,N_9768);
nand U10233 (N_10233,N_9104,N_9522);
and U10234 (N_10234,N_9747,N_9323);
nand U10235 (N_10235,N_9993,N_9855);
nand U10236 (N_10236,N_9992,N_9937);
xor U10237 (N_10237,N_9393,N_9844);
or U10238 (N_10238,N_9109,N_9876);
or U10239 (N_10239,N_9060,N_9898);
or U10240 (N_10240,N_9330,N_9382);
and U10241 (N_10241,N_9925,N_9866);
nand U10242 (N_10242,N_9683,N_9559);
nor U10243 (N_10243,N_9613,N_9132);
and U10244 (N_10244,N_9534,N_9973);
or U10245 (N_10245,N_9983,N_9739);
or U10246 (N_10246,N_9837,N_9238);
nor U10247 (N_10247,N_9885,N_9638);
xor U10248 (N_10248,N_9838,N_9406);
or U10249 (N_10249,N_9886,N_9745);
xnor U10250 (N_10250,N_9129,N_9423);
and U10251 (N_10251,N_9697,N_9313);
or U10252 (N_10252,N_9161,N_9435);
nor U10253 (N_10253,N_9648,N_9531);
or U10254 (N_10254,N_9702,N_9327);
or U10255 (N_10255,N_9470,N_9709);
xnor U10256 (N_10256,N_9637,N_9987);
nand U10257 (N_10257,N_9953,N_9749);
nor U10258 (N_10258,N_9636,N_9845);
or U10259 (N_10259,N_9823,N_9014);
nand U10260 (N_10260,N_9056,N_9911);
or U10261 (N_10261,N_9924,N_9337);
nand U10262 (N_10262,N_9774,N_9071);
and U10263 (N_10263,N_9936,N_9982);
and U10264 (N_10264,N_9058,N_9514);
nor U10265 (N_10265,N_9726,N_9769);
and U10266 (N_10266,N_9166,N_9360);
xor U10267 (N_10267,N_9618,N_9675);
and U10268 (N_10268,N_9679,N_9088);
nand U10269 (N_10269,N_9596,N_9100);
or U10270 (N_10270,N_9565,N_9858);
or U10271 (N_10271,N_9242,N_9520);
nor U10272 (N_10272,N_9811,N_9511);
nor U10273 (N_10273,N_9483,N_9660);
and U10274 (N_10274,N_9202,N_9932);
or U10275 (N_10275,N_9816,N_9624);
and U10276 (N_10276,N_9649,N_9743);
and U10277 (N_10277,N_9737,N_9529);
nor U10278 (N_10278,N_9110,N_9765);
xnor U10279 (N_10279,N_9448,N_9492);
nor U10280 (N_10280,N_9642,N_9357);
nor U10281 (N_10281,N_9888,N_9144);
nand U10282 (N_10282,N_9706,N_9383);
or U10283 (N_10283,N_9149,N_9717);
or U10284 (N_10284,N_9502,N_9439);
or U10285 (N_10285,N_9450,N_9913);
nor U10286 (N_10286,N_9829,N_9939);
or U10287 (N_10287,N_9773,N_9536);
or U10288 (N_10288,N_9286,N_9214);
nand U10289 (N_10289,N_9059,N_9053);
nor U10290 (N_10290,N_9528,N_9505);
nand U10291 (N_10291,N_9347,N_9372);
and U10292 (N_10292,N_9631,N_9447);
or U10293 (N_10293,N_9309,N_9849);
nor U10294 (N_10294,N_9570,N_9349);
nor U10295 (N_10295,N_9160,N_9107);
or U10296 (N_10296,N_9042,N_9140);
nand U10297 (N_10297,N_9210,N_9584);
xor U10298 (N_10298,N_9219,N_9926);
nor U10299 (N_10299,N_9894,N_9451);
or U10300 (N_10300,N_9895,N_9375);
and U10301 (N_10301,N_9271,N_9261);
nand U10302 (N_10302,N_9024,N_9516);
nor U10303 (N_10303,N_9699,N_9799);
and U10304 (N_10304,N_9284,N_9719);
xor U10305 (N_10305,N_9754,N_9185);
nand U10306 (N_10306,N_9676,N_9049);
nor U10307 (N_10307,N_9569,N_9707);
nand U10308 (N_10308,N_9359,N_9867);
nand U10309 (N_10309,N_9437,N_9763);
nor U10310 (N_10310,N_9538,N_9396);
nor U10311 (N_10311,N_9625,N_9074);
nor U10312 (N_10312,N_9694,N_9003);
nor U10313 (N_10313,N_9958,N_9333);
and U10314 (N_10314,N_9038,N_9371);
and U10315 (N_10315,N_9801,N_9884);
xor U10316 (N_10316,N_9713,N_9153);
or U10317 (N_10317,N_9526,N_9779);
xor U10318 (N_10318,N_9440,N_9370);
and U10319 (N_10319,N_9820,N_9462);
nand U10320 (N_10320,N_9342,N_9759);
or U10321 (N_10321,N_9716,N_9319);
nor U10322 (N_10322,N_9468,N_9736);
or U10323 (N_10323,N_9865,N_9169);
nor U10324 (N_10324,N_9010,N_9050);
nor U10325 (N_10325,N_9733,N_9340);
nor U10326 (N_10326,N_9581,N_9551);
nand U10327 (N_10327,N_9163,N_9013);
nor U10328 (N_10328,N_9735,N_9410);
or U10329 (N_10329,N_9066,N_9997);
and U10330 (N_10330,N_9988,N_9748);
and U10331 (N_10331,N_9222,N_9419);
nor U10332 (N_10332,N_9091,N_9072);
and U10333 (N_10333,N_9980,N_9916);
or U10334 (N_10334,N_9635,N_9209);
or U10335 (N_10335,N_9965,N_9564);
nand U10336 (N_10336,N_9215,N_9938);
nand U10337 (N_10337,N_9784,N_9101);
nor U10338 (N_10338,N_9133,N_9345);
xnor U10339 (N_10339,N_9654,N_9627);
nor U10340 (N_10340,N_9134,N_9195);
nand U10341 (N_10341,N_9055,N_9828);
nand U10342 (N_10342,N_9887,N_9677);
nand U10343 (N_10343,N_9263,N_9499);
nor U10344 (N_10344,N_9947,N_9778);
nand U10345 (N_10345,N_9257,N_9287);
nand U10346 (N_10346,N_9941,N_9674);
and U10347 (N_10347,N_9135,N_9962);
and U10348 (N_10348,N_9245,N_9493);
nand U10349 (N_10349,N_9583,N_9180);
and U10350 (N_10350,N_9255,N_9793);
xor U10351 (N_10351,N_9839,N_9549);
or U10352 (N_10352,N_9005,N_9269);
nor U10353 (N_10353,N_9179,N_9204);
and U10354 (N_10354,N_9673,N_9247);
nor U10355 (N_10355,N_9990,N_9452);
xor U10356 (N_10356,N_9211,N_9380);
xor U10357 (N_10357,N_9921,N_9813);
xnor U10358 (N_10358,N_9457,N_9756);
or U10359 (N_10359,N_9577,N_9640);
and U10360 (N_10360,N_9265,N_9875);
nor U10361 (N_10361,N_9843,N_9384);
and U10362 (N_10362,N_9432,N_9243);
nor U10363 (N_10363,N_9199,N_9200);
or U10364 (N_10364,N_9301,N_9240);
nand U10365 (N_10365,N_9805,N_9299);
nor U10366 (N_10366,N_9326,N_9933);
nor U10367 (N_10367,N_9558,N_9428);
nor U10368 (N_10368,N_9460,N_9984);
and U10369 (N_10369,N_9818,N_9705);
and U10370 (N_10370,N_9650,N_9580);
nand U10371 (N_10371,N_9948,N_9227);
or U10372 (N_10372,N_9022,N_9863);
nand U10373 (N_10373,N_9378,N_9220);
or U10374 (N_10374,N_9307,N_9259);
nand U10375 (N_10375,N_9308,N_9542);
or U10376 (N_10376,N_9655,N_9999);
nor U10377 (N_10377,N_9929,N_9616);
nor U10378 (N_10378,N_9831,N_9620);
and U10379 (N_10379,N_9610,N_9489);
nand U10380 (N_10380,N_9905,N_9173);
xnor U10381 (N_10381,N_9780,N_9821);
nand U10382 (N_10382,N_9020,N_9248);
or U10383 (N_10383,N_9026,N_9600);
and U10384 (N_10384,N_9376,N_9503);
nand U10385 (N_10385,N_9891,N_9762);
nor U10386 (N_10386,N_9120,N_9714);
or U10387 (N_10387,N_9239,N_9076);
and U10388 (N_10388,N_9399,N_9785);
nor U10389 (N_10389,N_9617,N_9809);
and U10390 (N_10390,N_9007,N_9434);
or U10391 (N_10391,N_9647,N_9668);
nand U10392 (N_10392,N_9417,N_9413);
and U10393 (N_10393,N_9430,N_9235);
and U10394 (N_10394,N_9017,N_9621);
or U10395 (N_10395,N_9137,N_9289);
nor U10396 (N_10396,N_9880,N_9934);
and U10397 (N_10397,N_9221,N_9155);
nand U10398 (N_10398,N_9553,N_9314);
nor U10399 (N_10399,N_9686,N_9734);
or U10400 (N_10400,N_9842,N_9952);
xnor U10401 (N_10401,N_9115,N_9315);
and U10402 (N_10402,N_9092,N_9266);
nand U10403 (N_10403,N_9027,N_9461);
nand U10404 (N_10404,N_9622,N_9729);
nor U10405 (N_10405,N_9302,N_9303);
and U10406 (N_10406,N_9602,N_9908);
nand U10407 (N_10407,N_9394,N_9454);
nand U10408 (N_10408,N_9963,N_9172);
xor U10409 (N_10409,N_9972,N_9391);
nor U10410 (N_10410,N_9954,N_9040);
or U10411 (N_10411,N_9128,N_9445);
nand U10412 (N_10412,N_9684,N_9950);
or U10413 (N_10413,N_9093,N_9398);
nor U10414 (N_10414,N_9488,N_9048);
or U10415 (N_10415,N_9392,N_9864);
or U10416 (N_10416,N_9724,N_9959);
and U10417 (N_10417,N_9652,N_9852);
nor U10418 (N_10418,N_9915,N_9860);
nand U10419 (N_10419,N_9741,N_9560);
or U10420 (N_10420,N_9757,N_9989);
nor U10421 (N_10421,N_9619,N_9296);
nand U10422 (N_10422,N_9700,N_9854);
nand U10423 (N_10423,N_9914,N_9433);
xnor U10424 (N_10424,N_9069,N_9720);
nor U10425 (N_10425,N_9057,N_9178);
nor U10426 (N_10426,N_9480,N_9851);
and U10427 (N_10427,N_9687,N_9603);
or U10428 (N_10428,N_9201,N_9721);
and U10429 (N_10429,N_9322,N_9662);
xor U10430 (N_10430,N_9162,N_9346);
and U10431 (N_10431,N_9029,N_9463);
and U10432 (N_10432,N_9770,N_9481);
xnor U10433 (N_10433,N_9054,N_9710);
nand U10434 (N_10434,N_9368,N_9692);
nand U10435 (N_10435,N_9052,N_9051);
nor U10436 (N_10436,N_9957,N_9834);
or U10437 (N_10437,N_9482,N_9904);
or U10438 (N_10438,N_9122,N_9225);
xnor U10439 (N_10439,N_9175,N_9416);
nand U10440 (N_10440,N_9418,N_9847);
nand U10441 (N_10441,N_9537,N_9804);
nand U10442 (N_10442,N_9325,N_9283);
or U10443 (N_10443,N_9666,N_9961);
nor U10444 (N_10444,N_9442,N_9094);
nand U10445 (N_10445,N_9543,N_9113);
and U10446 (N_10446,N_9800,N_9373);
or U10447 (N_10447,N_9826,N_9217);
and U10448 (N_10448,N_9579,N_9476);
nand U10449 (N_10449,N_9226,N_9986);
nor U10450 (N_10450,N_9258,N_9787);
nor U10451 (N_10451,N_9521,N_9386);
and U10452 (N_10452,N_9897,N_9473);
nand U10453 (N_10453,N_9956,N_9187);
and U10454 (N_10454,N_9578,N_9366);
or U10455 (N_10455,N_9321,N_9836);
nor U10456 (N_10456,N_9167,N_9712);
nand U10457 (N_10457,N_9045,N_9233);
and U10458 (N_10458,N_9798,N_9165);
xor U10459 (N_10459,N_9073,N_9566);
nand U10460 (N_10460,N_9364,N_9355);
or U10461 (N_10461,N_9474,N_9996);
nand U10462 (N_10462,N_9084,N_9156);
and U10463 (N_10463,N_9893,N_9917);
xor U10464 (N_10464,N_9730,N_9328);
xnor U10465 (N_10465,N_9046,N_9414);
nand U10466 (N_10466,N_9006,N_9023);
and U10467 (N_10467,N_9981,N_9441);
xnor U10468 (N_10468,N_9111,N_9857);
xor U10469 (N_10469,N_9151,N_9681);
nor U10470 (N_10470,N_9276,N_9438);
or U10471 (N_10471,N_9047,N_9408);
nand U10472 (N_10472,N_9103,N_9292);
nor U10473 (N_10473,N_9218,N_9186);
nor U10474 (N_10474,N_9498,N_9942);
and U10475 (N_10475,N_9665,N_9587);
xor U10476 (N_10476,N_9727,N_9147);
and U10477 (N_10477,N_9830,N_9224);
nor U10478 (N_10478,N_9485,N_9279);
nand U10479 (N_10479,N_9236,N_9883);
or U10480 (N_10480,N_9524,N_9426);
nor U10481 (N_10481,N_9190,N_9234);
nor U10482 (N_10482,N_9032,N_9530);
xnor U10483 (N_10483,N_9967,N_9641);
and U10484 (N_10484,N_9207,N_9192);
nand U10485 (N_10485,N_9039,N_9775);
and U10486 (N_10486,N_9822,N_9777);
nand U10487 (N_10487,N_9082,N_9562);
nor U10488 (N_10488,N_9458,N_9196);
or U10489 (N_10489,N_9009,N_9698);
nor U10490 (N_10490,N_9856,N_9841);
or U10491 (N_10491,N_9090,N_9030);
and U10492 (N_10492,N_9098,N_9427);
nor U10493 (N_10493,N_9085,N_9808);
or U10494 (N_10494,N_9633,N_9870);
and U10495 (N_10495,N_9544,N_9909);
or U10496 (N_10496,N_9008,N_9786);
nor U10497 (N_10497,N_9465,N_9139);
nor U10498 (N_10498,N_9361,N_9249);
nor U10499 (N_10499,N_9123,N_9232);
nand U10500 (N_10500,N_9692,N_9223);
nand U10501 (N_10501,N_9083,N_9361);
nand U10502 (N_10502,N_9512,N_9646);
or U10503 (N_10503,N_9833,N_9746);
nand U10504 (N_10504,N_9614,N_9572);
and U10505 (N_10505,N_9680,N_9405);
nor U10506 (N_10506,N_9819,N_9094);
nand U10507 (N_10507,N_9027,N_9515);
and U10508 (N_10508,N_9722,N_9942);
xor U10509 (N_10509,N_9964,N_9915);
and U10510 (N_10510,N_9063,N_9965);
nor U10511 (N_10511,N_9509,N_9656);
nand U10512 (N_10512,N_9265,N_9225);
and U10513 (N_10513,N_9688,N_9217);
nand U10514 (N_10514,N_9581,N_9465);
or U10515 (N_10515,N_9719,N_9959);
and U10516 (N_10516,N_9802,N_9031);
nand U10517 (N_10517,N_9425,N_9685);
and U10518 (N_10518,N_9291,N_9303);
nand U10519 (N_10519,N_9559,N_9224);
nor U10520 (N_10520,N_9956,N_9546);
and U10521 (N_10521,N_9277,N_9104);
nand U10522 (N_10522,N_9801,N_9479);
nor U10523 (N_10523,N_9222,N_9035);
xnor U10524 (N_10524,N_9921,N_9676);
and U10525 (N_10525,N_9632,N_9242);
nor U10526 (N_10526,N_9055,N_9606);
xnor U10527 (N_10527,N_9564,N_9811);
nor U10528 (N_10528,N_9635,N_9168);
nor U10529 (N_10529,N_9910,N_9209);
nor U10530 (N_10530,N_9141,N_9059);
or U10531 (N_10531,N_9309,N_9506);
or U10532 (N_10532,N_9905,N_9308);
nor U10533 (N_10533,N_9637,N_9954);
xor U10534 (N_10534,N_9102,N_9118);
and U10535 (N_10535,N_9647,N_9137);
xnor U10536 (N_10536,N_9389,N_9147);
and U10537 (N_10537,N_9319,N_9937);
nand U10538 (N_10538,N_9457,N_9497);
nor U10539 (N_10539,N_9793,N_9493);
xor U10540 (N_10540,N_9348,N_9878);
nor U10541 (N_10541,N_9036,N_9506);
nor U10542 (N_10542,N_9007,N_9987);
nor U10543 (N_10543,N_9883,N_9031);
and U10544 (N_10544,N_9683,N_9298);
or U10545 (N_10545,N_9952,N_9963);
or U10546 (N_10546,N_9076,N_9538);
or U10547 (N_10547,N_9926,N_9960);
or U10548 (N_10548,N_9560,N_9727);
nor U10549 (N_10549,N_9060,N_9289);
nand U10550 (N_10550,N_9523,N_9680);
nor U10551 (N_10551,N_9186,N_9277);
and U10552 (N_10552,N_9340,N_9754);
xnor U10553 (N_10553,N_9827,N_9707);
xnor U10554 (N_10554,N_9667,N_9108);
and U10555 (N_10555,N_9860,N_9727);
and U10556 (N_10556,N_9199,N_9446);
and U10557 (N_10557,N_9577,N_9825);
nand U10558 (N_10558,N_9283,N_9866);
and U10559 (N_10559,N_9319,N_9469);
or U10560 (N_10560,N_9820,N_9716);
nor U10561 (N_10561,N_9369,N_9143);
and U10562 (N_10562,N_9938,N_9458);
nand U10563 (N_10563,N_9723,N_9877);
nor U10564 (N_10564,N_9652,N_9833);
nor U10565 (N_10565,N_9385,N_9991);
nor U10566 (N_10566,N_9871,N_9096);
and U10567 (N_10567,N_9346,N_9029);
and U10568 (N_10568,N_9518,N_9446);
nand U10569 (N_10569,N_9444,N_9189);
nand U10570 (N_10570,N_9813,N_9844);
nor U10571 (N_10571,N_9723,N_9563);
nor U10572 (N_10572,N_9387,N_9728);
nand U10573 (N_10573,N_9062,N_9003);
or U10574 (N_10574,N_9834,N_9540);
or U10575 (N_10575,N_9844,N_9640);
and U10576 (N_10576,N_9459,N_9173);
and U10577 (N_10577,N_9175,N_9030);
and U10578 (N_10578,N_9124,N_9040);
or U10579 (N_10579,N_9982,N_9123);
and U10580 (N_10580,N_9755,N_9800);
and U10581 (N_10581,N_9884,N_9792);
nand U10582 (N_10582,N_9649,N_9576);
and U10583 (N_10583,N_9925,N_9438);
or U10584 (N_10584,N_9271,N_9953);
or U10585 (N_10585,N_9127,N_9314);
and U10586 (N_10586,N_9937,N_9340);
nand U10587 (N_10587,N_9027,N_9726);
and U10588 (N_10588,N_9280,N_9002);
xnor U10589 (N_10589,N_9081,N_9425);
or U10590 (N_10590,N_9849,N_9250);
nand U10591 (N_10591,N_9438,N_9565);
nor U10592 (N_10592,N_9005,N_9197);
and U10593 (N_10593,N_9645,N_9193);
or U10594 (N_10594,N_9294,N_9207);
nand U10595 (N_10595,N_9731,N_9857);
and U10596 (N_10596,N_9799,N_9421);
nand U10597 (N_10597,N_9196,N_9794);
and U10598 (N_10598,N_9697,N_9628);
nand U10599 (N_10599,N_9901,N_9427);
nand U10600 (N_10600,N_9211,N_9097);
and U10601 (N_10601,N_9636,N_9337);
nor U10602 (N_10602,N_9283,N_9569);
or U10603 (N_10603,N_9309,N_9601);
or U10604 (N_10604,N_9770,N_9446);
or U10605 (N_10605,N_9842,N_9460);
or U10606 (N_10606,N_9568,N_9603);
xor U10607 (N_10607,N_9249,N_9237);
nor U10608 (N_10608,N_9421,N_9066);
nand U10609 (N_10609,N_9319,N_9678);
nor U10610 (N_10610,N_9672,N_9621);
and U10611 (N_10611,N_9332,N_9185);
nand U10612 (N_10612,N_9954,N_9906);
nor U10613 (N_10613,N_9437,N_9333);
nor U10614 (N_10614,N_9413,N_9862);
xnor U10615 (N_10615,N_9812,N_9246);
nand U10616 (N_10616,N_9765,N_9506);
nand U10617 (N_10617,N_9895,N_9989);
nor U10618 (N_10618,N_9339,N_9054);
nand U10619 (N_10619,N_9677,N_9942);
nor U10620 (N_10620,N_9435,N_9825);
nand U10621 (N_10621,N_9800,N_9059);
nor U10622 (N_10622,N_9611,N_9675);
nand U10623 (N_10623,N_9897,N_9849);
nor U10624 (N_10624,N_9466,N_9112);
nor U10625 (N_10625,N_9067,N_9504);
nand U10626 (N_10626,N_9070,N_9857);
nand U10627 (N_10627,N_9671,N_9446);
nand U10628 (N_10628,N_9205,N_9607);
or U10629 (N_10629,N_9597,N_9781);
and U10630 (N_10630,N_9575,N_9693);
or U10631 (N_10631,N_9778,N_9170);
nor U10632 (N_10632,N_9761,N_9938);
or U10633 (N_10633,N_9137,N_9713);
xor U10634 (N_10634,N_9816,N_9238);
or U10635 (N_10635,N_9880,N_9752);
nor U10636 (N_10636,N_9872,N_9939);
nand U10637 (N_10637,N_9876,N_9028);
and U10638 (N_10638,N_9557,N_9959);
or U10639 (N_10639,N_9940,N_9790);
nor U10640 (N_10640,N_9289,N_9770);
and U10641 (N_10641,N_9527,N_9839);
and U10642 (N_10642,N_9769,N_9492);
or U10643 (N_10643,N_9815,N_9807);
or U10644 (N_10644,N_9127,N_9181);
nor U10645 (N_10645,N_9792,N_9982);
nand U10646 (N_10646,N_9283,N_9737);
nor U10647 (N_10647,N_9245,N_9016);
nand U10648 (N_10648,N_9002,N_9686);
nor U10649 (N_10649,N_9650,N_9345);
and U10650 (N_10650,N_9446,N_9530);
nand U10651 (N_10651,N_9066,N_9802);
or U10652 (N_10652,N_9149,N_9960);
nor U10653 (N_10653,N_9005,N_9736);
nand U10654 (N_10654,N_9722,N_9565);
and U10655 (N_10655,N_9692,N_9783);
or U10656 (N_10656,N_9914,N_9057);
or U10657 (N_10657,N_9314,N_9352);
nor U10658 (N_10658,N_9226,N_9060);
nand U10659 (N_10659,N_9263,N_9315);
nor U10660 (N_10660,N_9956,N_9575);
and U10661 (N_10661,N_9834,N_9287);
or U10662 (N_10662,N_9474,N_9002);
nand U10663 (N_10663,N_9319,N_9104);
nor U10664 (N_10664,N_9493,N_9834);
and U10665 (N_10665,N_9295,N_9831);
nand U10666 (N_10666,N_9066,N_9722);
nand U10667 (N_10667,N_9109,N_9658);
nor U10668 (N_10668,N_9026,N_9223);
or U10669 (N_10669,N_9085,N_9922);
or U10670 (N_10670,N_9343,N_9860);
nor U10671 (N_10671,N_9019,N_9850);
nor U10672 (N_10672,N_9215,N_9593);
xor U10673 (N_10673,N_9487,N_9832);
nor U10674 (N_10674,N_9443,N_9348);
or U10675 (N_10675,N_9495,N_9840);
nand U10676 (N_10676,N_9614,N_9807);
and U10677 (N_10677,N_9828,N_9457);
and U10678 (N_10678,N_9781,N_9963);
and U10679 (N_10679,N_9296,N_9024);
nor U10680 (N_10680,N_9419,N_9475);
nor U10681 (N_10681,N_9504,N_9720);
or U10682 (N_10682,N_9031,N_9149);
and U10683 (N_10683,N_9127,N_9885);
nor U10684 (N_10684,N_9581,N_9995);
or U10685 (N_10685,N_9128,N_9091);
nor U10686 (N_10686,N_9832,N_9155);
and U10687 (N_10687,N_9838,N_9174);
nand U10688 (N_10688,N_9206,N_9419);
nand U10689 (N_10689,N_9474,N_9540);
or U10690 (N_10690,N_9160,N_9718);
nand U10691 (N_10691,N_9118,N_9638);
nand U10692 (N_10692,N_9380,N_9168);
and U10693 (N_10693,N_9594,N_9990);
nand U10694 (N_10694,N_9750,N_9246);
xor U10695 (N_10695,N_9343,N_9288);
and U10696 (N_10696,N_9991,N_9174);
xor U10697 (N_10697,N_9857,N_9212);
nor U10698 (N_10698,N_9083,N_9983);
and U10699 (N_10699,N_9047,N_9515);
nor U10700 (N_10700,N_9178,N_9070);
and U10701 (N_10701,N_9208,N_9364);
nand U10702 (N_10702,N_9808,N_9901);
and U10703 (N_10703,N_9852,N_9268);
xor U10704 (N_10704,N_9423,N_9870);
or U10705 (N_10705,N_9197,N_9764);
nor U10706 (N_10706,N_9944,N_9401);
or U10707 (N_10707,N_9825,N_9003);
nor U10708 (N_10708,N_9308,N_9490);
nor U10709 (N_10709,N_9570,N_9741);
or U10710 (N_10710,N_9995,N_9529);
xnor U10711 (N_10711,N_9389,N_9962);
and U10712 (N_10712,N_9960,N_9909);
nor U10713 (N_10713,N_9880,N_9195);
or U10714 (N_10714,N_9151,N_9588);
or U10715 (N_10715,N_9324,N_9970);
and U10716 (N_10716,N_9045,N_9212);
nand U10717 (N_10717,N_9459,N_9375);
nand U10718 (N_10718,N_9019,N_9104);
nand U10719 (N_10719,N_9549,N_9509);
and U10720 (N_10720,N_9745,N_9449);
and U10721 (N_10721,N_9200,N_9861);
nor U10722 (N_10722,N_9806,N_9476);
or U10723 (N_10723,N_9882,N_9448);
xnor U10724 (N_10724,N_9123,N_9432);
or U10725 (N_10725,N_9879,N_9921);
nand U10726 (N_10726,N_9127,N_9331);
nand U10727 (N_10727,N_9876,N_9617);
nor U10728 (N_10728,N_9482,N_9834);
and U10729 (N_10729,N_9892,N_9602);
nand U10730 (N_10730,N_9401,N_9065);
xor U10731 (N_10731,N_9440,N_9571);
and U10732 (N_10732,N_9278,N_9075);
or U10733 (N_10733,N_9120,N_9706);
or U10734 (N_10734,N_9631,N_9723);
nor U10735 (N_10735,N_9658,N_9996);
xnor U10736 (N_10736,N_9512,N_9520);
nor U10737 (N_10737,N_9810,N_9662);
or U10738 (N_10738,N_9368,N_9613);
xnor U10739 (N_10739,N_9758,N_9823);
nor U10740 (N_10740,N_9195,N_9925);
xor U10741 (N_10741,N_9056,N_9483);
xnor U10742 (N_10742,N_9437,N_9615);
or U10743 (N_10743,N_9307,N_9827);
and U10744 (N_10744,N_9297,N_9081);
xnor U10745 (N_10745,N_9167,N_9919);
nor U10746 (N_10746,N_9510,N_9555);
nand U10747 (N_10747,N_9522,N_9086);
nor U10748 (N_10748,N_9721,N_9468);
and U10749 (N_10749,N_9381,N_9270);
nor U10750 (N_10750,N_9988,N_9010);
and U10751 (N_10751,N_9977,N_9096);
xor U10752 (N_10752,N_9923,N_9043);
nand U10753 (N_10753,N_9511,N_9401);
nand U10754 (N_10754,N_9350,N_9097);
xor U10755 (N_10755,N_9487,N_9670);
nor U10756 (N_10756,N_9298,N_9557);
and U10757 (N_10757,N_9380,N_9888);
or U10758 (N_10758,N_9031,N_9796);
and U10759 (N_10759,N_9393,N_9922);
and U10760 (N_10760,N_9155,N_9031);
nor U10761 (N_10761,N_9395,N_9377);
xor U10762 (N_10762,N_9181,N_9342);
nor U10763 (N_10763,N_9739,N_9142);
nand U10764 (N_10764,N_9458,N_9703);
nand U10765 (N_10765,N_9023,N_9508);
and U10766 (N_10766,N_9630,N_9413);
or U10767 (N_10767,N_9574,N_9327);
or U10768 (N_10768,N_9588,N_9019);
or U10769 (N_10769,N_9343,N_9845);
or U10770 (N_10770,N_9204,N_9328);
or U10771 (N_10771,N_9220,N_9830);
and U10772 (N_10772,N_9618,N_9681);
and U10773 (N_10773,N_9748,N_9942);
xnor U10774 (N_10774,N_9312,N_9605);
or U10775 (N_10775,N_9007,N_9628);
xnor U10776 (N_10776,N_9459,N_9668);
nor U10777 (N_10777,N_9374,N_9028);
or U10778 (N_10778,N_9069,N_9793);
nand U10779 (N_10779,N_9413,N_9728);
nor U10780 (N_10780,N_9236,N_9961);
nand U10781 (N_10781,N_9351,N_9590);
nand U10782 (N_10782,N_9578,N_9754);
nor U10783 (N_10783,N_9905,N_9121);
or U10784 (N_10784,N_9144,N_9254);
nand U10785 (N_10785,N_9597,N_9588);
or U10786 (N_10786,N_9372,N_9808);
nor U10787 (N_10787,N_9901,N_9875);
or U10788 (N_10788,N_9307,N_9633);
nor U10789 (N_10789,N_9371,N_9492);
nor U10790 (N_10790,N_9876,N_9526);
or U10791 (N_10791,N_9304,N_9521);
nand U10792 (N_10792,N_9152,N_9189);
nand U10793 (N_10793,N_9868,N_9559);
or U10794 (N_10794,N_9006,N_9959);
and U10795 (N_10795,N_9334,N_9165);
or U10796 (N_10796,N_9229,N_9225);
or U10797 (N_10797,N_9423,N_9948);
or U10798 (N_10798,N_9061,N_9192);
nor U10799 (N_10799,N_9933,N_9872);
and U10800 (N_10800,N_9087,N_9326);
or U10801 (N_10801,N_9060,N_9215);
and U10802 (N_10802,N_9449,N_9731);
xnor U10803 (N_10803,N_9184,N_9547);
and U10804 (N_10804,N_9583,N_9565);
or U10805 (N_10805,N_9888,N_9868);
nor U10806 (N_10806,N_9345,N_9611);
xnor U10807 (N_10807,N_9708,N_9570);
and U10808 (N_10808,N_9968,N_9935);
or U10809 (N_10809,N_9064,N_9922);
nor U10810 (N_10810,N_9090,N_9672);
nor U10811 (N_10811,N_9608,N_9341);
xnor U10812 (N_10812,N_9629,N_9949);
nand U10813 (N_10813,N_9281,N_9462);
nor U10814 (N_10814,N_9958,N_9876);
or U10815 (N_10815,N_9178,N_9873);
nor U10816 (N_10816,N_9648,N_9150);
or U10817 (N_10817,N_9338,N_9580);
and U10818 (N_10818,N_9236,N_9021);
or U10819 (N_10819,N_9944,N_9725);
nor U10820 (N_10820,N_9199,N_9623);
and U10821 (N_10821,N_9351,N_9852);
and U10822 (N_10822,N_9027,N_9765);
or U10823 (N_10823,N_9407,N_9221);
nor U10824 (N_10824,N_9303,N_9769);
and U10825 (N_10825,N_9756,N_9411);
nor U10826 (N_10826,N_9721,N_9739);
nand U10827 (N_10827,N_9170,N_9752);
nand U10828 (N_10828,N_9368,N_9987);
nand U10829 (N_10829,N_9036,N_9727);
nor U10830 (N_10830,N_9057,N_9584);
xor U10831 (N_10831,N_9608,N_9580);
or U10832 (N_10832,N_9407,N_9168);
and U10833 (N_10833,N_9913,N_9953);
or U10834 (N_10834,N_9743,N_9579);
and U10835 (N_10835,N_9243,N_9690);
nor U10836 (N_10836,N_9623,N_9655);
and U10837 (N_10837,N_9682,N_9204);
nand U10838 (N_10838,N_9606,N_9847);
and U10839 (N_10839,N_9155,N_9335);
or U10840 (N_10840,N_9683,N_9997);
nand U10841 (N_10841,N_9697,N_9280);
nand U10842 (N_10842,N_9146,N_9220);
and U10843 (N_10843,N_9580,N_9502);
nor U10844 (N_10844,N_9804,N_9970);
and U10845 (N_10845,N_9039,N_9637);
nor U10846 (N_10846,N_9085,N_9757);
xor U10847 (N_10847,N_9957,N_9576);
nand U10848 (N_10848,N_9329,N_9883);
nand U10849 (N_10849,N_9911,N_9522);
or U10850 (N_10850,N_9542,N_9800);
nor U10851 (N_10851,N_9270,N_9219);
and U10852 (N_10852,N_9280,N_9971);
and U10853 (N_10853,N_9191,N_9418);
or U10854 (N_10854,N_9372,N_9398);
xor U10855 (N_10855,N_9429,N_9917);
xnor U10856 (N_10856,N_9439,N_9586);
and U10857 (N_10857,N_9714,N_9851);
nor U10858 (N_10858,N_9776,N_9353);
or U10859 (N_10859,N_9863,N_9798);
nor U10860 (N_10860,N_9155,N_9873);
nand U10861 (N_10861,N_9789,N_9387);
xnor U10862 (N_10862,N_9961,N_9237);
nor U10863 (N_10863,N_9778,N_9624);
nand U10864 (N_10864,N_9431,N_9692);
xnor U10865 (N_10865,N_9246,N_9479);
nor U10866 (N_10866,N_9924,N_9945);
nor U10867 (N_10867,N_9880,N_9733);
and U10868 (N_10868,N_9568,N_9170);
nand U10869 (N_10869,N_9886,N_9418);
nor U10870 (N_10870,N_9644,N_9795);
xnor U10871 (N_10871,N_9754,N_9597);
nor U10872 (N_10872,N_9051,N_9938);
nand U10873 (N_10873,N_9104,N_9672);
or U10874 (N_10874,N_9561,N_9516);
or U10875 (N_10875,N_9993,N_9323);
or U10876 (N_10876,N_9689,N_9974);
or U10877 (N_10877,N_9282,N_9168);
and U10878 (N_10878,N_9530,N_9623);
or U10879 (N_10879,N_9775,N_9323);
and U10880 (N_10880,N_9117,N_9867);
nand U10881 (N_10881,N_9031,N_9334);
and U10882 (N_10882,N_9917,N_9013);
nor U10883 (N_10883,N_9336,N_9353);
or U10884 (N_10884,N_9869,N_9488);
and U10885 (N_10885,N_9879,N_9054);
nand U10886 (N_10886,N_9380,N_9560);
or U10887 (N_10887,N_9333,N_9225);
or U10888 (N_10888,N_9339,N_9926);
nand U10889 (N_10889,N_9836,N_9330);
nand U10890 (N_10890,N_9526,N_9306);
and U10891 (N_10891,N_9292,N_9752);
or U10892 (N_10892,N_9248,N_9902);
nor U10893 (N_10893,N_9139,N_9371);
xnor U10894 (N_10894,N_9592,N_9412);
nand U10895 (N_10895,N_9394,N_9739);
nand U10896 (N_10896,N_9553,N_9068);
xor U10897 (N_10897,N_9734,N_9504);
nand U10898 (N_10898,N_9206,N_9813);
nand U10899 (N_10899,N_9107,N_9922);
and U10900 (N_10900,N_9817,N_9157);
nor U10901 (N_10901,N_9816,N_9431);
or U10902 (N_10902,N_9335,N_9868);
nor U10903 (N_10903,N_9327,N_9560);
nand U10904 (N_10904,N_9790,N_9079);
nor U10905 (N_10905,N_9881,N_9590);
or U10906 (N_10906,N_9593,N_9483);
xor U10907 (N_10907,N_9772,N_9757);
xor U10908 (N_10908,N_9206,N_9020);
or U10909 (N_10909,N_9629,N_9450);
nand U10910 (N_10910,N_9543,N_9084);
xor U10911 (N_10911,N_9172,N_9280);
and U10912 (N_10912,N_9673,N_9819);
xnor U10913 (N_10913,N_9759,N_9501);
nand U10914 (N_10914,N_9203,N_9305);
and U10915 (N_10915,N_9166,N_9545);
nand U10916 (N_10916,N_9930,N_9556);
nor U10917 (N_10917,N_9648,N_9306);
nor U10918 (N_10918,N_9685,N_9400);
xnor U10919 (N_10919,N_9799,N_9652);
and U10920 (N_10920,N_9084,N_9196);
nand U10921 (N_10921,N_9276,N_9936);
or U10922 (N_10922,N_9423,N_9612);
or U10923 (N_10923,N_9532,N_9204);
xnor U10924 (N_10924,N_9453,N_9900);
xnor U10925 (N_10925,N_9978,N_9272);
nor U10926 (N_10926,N_9277,N_9084);
nand U10927 (N_10927,N_9668,N_9275);
xor U10928 (N_10928,N_9166,N_9167);
or U10929 (N_10929,N_9453,N_9376);
or U10930 (N_10930,N_9356,N_9086);
or U10931 (N_10931,N_9330,N_9588);
or U10932 (N_10932,N_9823,N_9411);
nor U10933 (N_10933,N_9451,N_9418);
nand U10934 (N_10934,N_9534,N_9409);
and U10935 (N_10935,N_9903,N_9335);
or U10936 (N_10936,N_9724,N_9517);
and U10937 (N_10937,N_9760,N_9615);
nor U10938 (N_10938,N_9415,N_9074);
xnor U10939 (N_10939,N_9972,N_9939);
or U10940 (N_10940,N_9513,N_9879);
nand U10941 (N_10941,N_9692,N_9713);
nor U10942 (N_10942,N_9598,N_9160);
or U10943 (N_10943,N_9505,N_9670);
nand U10944 (N_10944,N_9685,N_9964);
nand U10945 (N_10945,N_9668,N_9395);
xor U10946 (N_10946,N_9045,N_9219);
and U10947 (N_10947,N_9448,N_9186);
nor U10948 (N_10948,N_9126,N_9972);
nor U10949 (N_10949,N_9581,N_9863);
or U10950 (N_10950,N_9285,N_9886);
or U10951 (N_10951,N_9404,N_9499);
nor U10952 (N_10952,N_9670,N_9196);
nor U10953 (N_10953,N_9142,N_9300);
nor U10954 (N_10954,N_9239,N_9683);
or U10955 (N_10955,N_9986,N_9880);
or U10956 (N_10956,N_9870,N_9114);
nor U10957 (N_10957,N_9195,N_9411);
and U10958 (N_10958,N_9638,N_9462);
and U10959 (N_10959,N_9136,N_9655);
and U10960 (N_10960,N_9909,N_9328);
or U10961 (N_10961,N_9097,N_9028);
nand U10962 (N_10962,N_9997,N_9483);
nand U10963 (N_10963,N_9696,N_9360);
and U10964 (N_10964,N_9149,N_9745);
nand U10965 (N_10965,N_9473,N_9332);
and U10966 (N_10966,N_9849,N_9730);
nand U10967 (N_10967,N_9002,N_9520);
nor U10968 (N_10968,N_9203,N_9516);
nor U10969 (N_10969,N_9574,N_9418);
or U10970 (N_10970,N_9683,N_9221);
nand U10971 (N_10971,N_9584,N_9312);
nand U10972 (N_10972,N_9024,N_9970);
nand U10973 (N_10973,N_9469,N_9704);
nor U10974 (N_10974,N_9696,N_9547);
nand U10975 (N_10975,N_9522,N_9715);
and U10976 (N_10976,N_9005,N_9709);
and U10977 (N_10977,N_9755,N_9207);
nor U10978 (N_10978,N_9877,N_9868);
or U10979 (N_10979,N_9130,N_9801);
nand U10980 (N_10980,N_9228,N_9723);
or U10981 (N_10981,N_9643,N_9532);
and U10982 (N_10982,N_9489,N_9684);
or U10983 (N_10983,N_9069,N_9142);
or U10984 (N_10984,N_9760,N_9304);
and U10985 (N_10985,N_9230,N_9109);
and U10986 (N_10986,N_9243,N_9518);
nand U10987 (N_10987,N_9691,N_9726);
or U10988 (N_10988,N_9242,N_9193);
and U10989 (N_10989,N_9908,N_9059);
nor U10990 (N_10990,N_9207,N_9620);
xnor U10991 (N_10991,N_9787,N_9432);
nand U10992 (N_10992,N_9341,N_9042);
or U10993 (N_10993,N_9008,N_9979);
nor U10994 (N_10994,N_9106,N_9596);
nand U10995 (N_10995,N_9186,N_9512);
nand U10996 (N_10996,N_9083,N_9452);
and U10997 (N_10997,N_9690,N_9056);
or U10998 (N_10998,N_9780,N_9289);
or U10999 (N_10999,N_9265,N_9842);
nor U11000 (N_11000,N_10996,N_10641);
nor U11001 (N_11001,N_10630,N_10416);
nand U11002 (N_11002,N_10004,N_10895);
nor U11003 (N_11003,N_10749,N_10619);
and U11004 (N_11004,N_10794,N_10428);
nor U11005 (N_11005,N_10847,N_10675);
xnor U11006 (N_11006,N_10534,N_10068);
xor U11007 (N_11007,N_10928,N_10627);
and U11008 (N_11008,N_10560,N_10899);
xor U11009 (N_11009,N_10244,N_10500);
and U11010 (N_11010,N_10870,N_10857);
nand U11011 (N_11011,N_10883,N_10310);
nor U11012 (N_11012,N_10320,N_10540);
nand U11013 (N_11013,N_10229,N_10580);
and U11014 (N_11014,N_10280,N_10113);
nand U11015 (N_11015,N_10406,N_10232);
xor U11016 (N_11016,N_10678,N_10803);
nor U11017 (N_11017,N_10139,N_10112);
or U11018 (N_11018,N_10102,N_10818);
xor U11019 (N_11019,N_10839,N_10833);
nand U11020 (N_11020,N_10546,N_10699);
nand U11021 (N_11021,N_10849,N_10062);
nand U11022 (N_11022,N_10153,N_10172);
or U11023 (N_11023,N_10090,N_10369);
and U11024 (N_11024,N_10159,N_10567);
nor U11025 (N_11025,N_10765,N_10910);
nand U11026 (N_11026,N_10027,N_10659);
or U11027 (N_11027,N_10029,N_10798);
or U11028 (N_11028,N_10271,N_10418);
or U11029 (N_11029,N_10167,N_10423);
nor U11030 (N_11030,N_10609,N_10755);
nand U11031 (N_11031,N_10439,N_10242);
or U11032 (N_11032,N_10478,N_10510);
and U11033 (N_11033,N_10703,N_10264);
or U11034 (N_11034,N_10597,N_10115);
nor U11035 (N_11035,N_10254,N_10867);
or U11036 (N_11036,N_10421,N_10760);
and U11037 (N_11037,N_10484,N_10083);
nor U11038 (N_11038,N_10455,N_10824);
nand U11039 (N_11039,N_10807,N_10188);
and U11040 (N_11040,N_10862,N_10373);
and U11041 (N_11041,N_10983,N_10008);
and U11042 (N_11042,N_10555,N_10941);
nor U11043 (N_11043,N_10956,N_10997);
nand U11044 (N_11044,N_10639,N_10492);
nand U11045 (N_11045,N_10353,N_10668);
xor U11046 (N_11046,N_10537,N_10448);
and U11047 (N_11047,N_10776,N_10123);
nor U11048 (N_11048,N_10992,N_10786);
nand U11049 (N_11049,N_10907,N_10969);
nand U11050 (N_11050,N_10042,N_10177);
or U11051 (N_11051,N_10838,N_10038);
nor U11052 (N_11052,N_10122,N_10213);
nor U11053 (N_11053,N_10007,N_10359);
and U11054 (N_11054,N_10502,N_10579);
or U11055 (N_11055,N_10957,N_10735);
nor U11056 (N_11056,N_10340,N_10712);
xor U11057 (N_11057,N_10916,N_10160);
and U11058 (N_11058,N_10044,N_10162);
xor U11059 (N_11059,N_10987,N_10601);
or U11060 (N_11060,N_10544,N_10877);
nand U11061 (N_11061,N_10911,N_10660);
or U11062 (N_11062,N_10125,N_10391);
xnor U11063 (N_11063,N_10404,N_10001);
xor U11064 (N_11064,N_10479,N_10780);
nor U11065 (N_11065,N_10679,N_10816);
and U11066 (N_11066,N_10485,N_10058);
nor U11067 (N_11067,N_10135,N_10727);
nand U11068 (N_11068,N_10021,N_10566);
or U11069 (N_11069,N_10395,N_10813);
nor U11070 (N_11070,N_10563,N_10236);
nor U11071 (N_11071,N_10164,N_10684);
xnor U11072 (N_11072,N_10696,N_10051);
xnor U11073 (N_11073,N_10517,N_10345);
nand U11074 (N_11074,N_10014,N_10884);
or U11075 (N_11075,N_10393,N_10300);
nor U11076 (N_11076,N_10430,N_10010);
nor U11077 (N_11077,N_10783,N_10046);
and U11078 (N_11078,N_10318,N_10193);
nor U11079 (N_11079,N_10405,N_10772);
xor U11080 (N_11080,N_10901,N_10497);
nand U11081 (N_11081,N_10142,N_10531);
and U11082 (N_11082,N_10460,N_10770);
nor U11083 (N_11083,N_10635,N_10097);
nor U11084 (N_11084,N_10821,N_10955);
nor U11085 (N_11085,N_10671,N_10575);
nor U11086 (N_11086,N_10933,N_10876);
and U11087 (N_11087,N_10388,N_10127);
and U11088 (N_11088,N_10495,N_10401);
and U11089 (N_11089,N_10819,N_10032);
and U11090 (N_11090,N_10331,N_10033);
or U11091 (N_11091,N_10767,N_10194);
and U11092 (N_11092,N_10722,N_10055);
nor U11093 (N_11093,N_10469,N_10729);
nor U11094 (N_11094,N_10754,N_10269);
and U11095 (N_11095,N_10644,N_10514);
xor U11096 (N_11096,N_10191,N_10267);
or U11097 (N_11097,N_10185,N_10399);
or U11098 (N_11098,N_10995,N_10059);
nand U11099 (N_11099,N_10964,N_10349);
nor U11100 (N_11100,N_10572,N_10060);
and U11101 (N_11101,N_10268,N_10990);
and U11102 (N_11102,N_10384,N_10801);
nand U11103 (N_11103,N_10315,N_10912);
nor U11104 (N_11104,N_10614,N_10666);
nor U11105 (N_11105,N_10364,N_10530);
nor U11106 (N_11106,N_10578,N_10805);
xnor U11107 (N_11107,N_10480,N_10545);
nand U11108 (N_11108,N_10716,N_10473);
nand U11109 (N_11109,N_10207,N_10661);
nor U11110 (N_11110,N_10440,N_10812);
nor U11111 (N_11111,N_10230,N_10169);
or U11112 (N_11112,N_10974,N_10622);
nand U11113 (N_11113,N_10085,N_10978);
and U11114 (N_11114,N_10950,N_10157);
nor U11115 (N_11115,N_10192,N_10790);
or U11116 (N_11116,N_10312,N_10730);
and U11117 (N_11117,N_10588,N_10855);
and U11118 (N_11118,N_10685,N_10149);
nand U11119 (N_11119,N_10420,N_10952);
and U11120 (N_11120,N_10251,N_10132);
nor U11121 (N_11121,N_10472,N_10773);
nor U11122 (N_11122,N_10657,N_10586);
nor U11123 (N_11123,N_10282,N_10830);
nand U11124 (N_11124,N_10494,N_10348);
or U11125 (N_11125,N_10652,N_10605);
xnor U11126 (N_11126,N_10832,N_10926);
and U11127 (N_11127,N_10260,N_10713);
or U11128 (N_11128,N_10152,N_10189);
or U11129 (N_11129,N_10902,N_10319);
nand U11130 (N_11130,N_10233,N_10810);
and U11131 (N_11131,N_10284,N_10719);
or U11132 (N_11132,N_10827,N_10625);
or U11133 (N_11133,N_10371,N_10356);
and U11134 (N_11134,N_10690,N_10809);
or U11135 (N_11135,N_10934,N_10250);
or U11136 (N_11136,N_10589,N_10873);
and U11137 (N_11137,N_10991,N_10844);
nor U11138 (N_11138,N_10746,N_10413);
nor U11139 (N_11139,N_10715,N_10655);
and U11140 (N_11140,N_10882,N_10664);
or U11141 (N_11141,N_10370,N_10930);
and U11142 (N_11142,N_10561,N_10209);
or U11143 (N_11143,N_10092,N_10170);
nand U11144 (N_11144,N_10972,N_10931);
and U11145 (N_11145,N_10266,N_10527);
nor U11146 (N_11146,N_10327,N_10487);
or U11147 (N_11147,N_10144,N_10342);
and U11148 (N_11148,N_10680,N_10724);
xor U11149 (N_11149,N_10082,N_10071);
xor U11150 (N_11150,N_10925,N_10012);
xnor U11151 (N_11151,N_10878,N_10938);
nor U11152 (N_11152,N_10651,N_10670);
nand U11153 (N_11153,N_10378,N_10241);
nor U11154 (N_11154,N_10116,N_10415);
xnor U11155 (N_11155,N_10292,N_10442);
nor U11156 (N_11156,N_10204,N_10898);
or U11157 (N_11157,N_10299,N_10493);
or U11158 (N_11158,N_10409,N_10396);
or U11159 (N_11159,N_10748,N_10171);
nor U11160 (N_11160,N_10023,N_10459);
and U11161 (N_11161,N_10020,N_10261);
nor U11162 (N_11162,N_10103,N_10272);
nand U11163 (N_11163,N_10604,N_10558);
nand U11164 (N_11164,N_10620,N_10278);
and U11165 (N_11165,N_10757,N_10141);
and U11166 (N_11166,N_10146,N_10505);
and U11167 (N_11167,N_10326,N_10096);
xor U11168 (N_11168,N_10017,N_10520);
nand U11169 (N_11169,N_10887,N_10245);
nand U11170 (N_11170,N_10199,N_10221);
or U11171 (N_11171,N_10000,N_10206);
nand U11172 (N_11172,N_10360,N_10994);
or U11173 (N_11173,N_10297,N_10638);
xor U11174 (N_11174,N_10425,N_10585);
nand U11175 (N_11175,N_10403,N_10959);
nand U11176 (N_11176,N_10550,N_10362);
and U11177 (N_11177,N_10653,N_10771);
or U11178 (N_11178,N_10564,N_10165);
and U11179 (N_11179,N_10147,N_10195);
or U11180 (N_11180,N_10337,N_10202);
and U11181 (N_11181,N_10306,N_10329);
nand U11182 (N_11182,N_10547,N_10759);
xor U11183 (N_11183,N_10307,N_10408);
nand U11184 (N_11184,N_10960,N_10845);
nand U11185 (N_11185,N_10491,N_10971);
and U11186 (N_11186,N_10441,N_10640);
nand U11187 (N_11187,N_10443,N_10488);
or U11188 (N_11188,N_10450,N_10366);
nor U11189 (N_11189,N_10205,N_10909);
or U11190 (N_11190,N_10741,N_10596);
nand U11191 (N_11191,N_10768,N_10054);
or U11192 (N_11192,N_10259,N_10341);
nand U11193 (N_11193,N_10196,N_10045);
nand U11194 (N_11194,N_10277,N_10865);
nor U11195 (N_11195,N_10982,N_10467);
or U11196 (N_11196,N_10281,N_10357);
nand U11197 (N_11197,N_10607,N_10247);
nor U11198 (N_11198,N_10963,N_10052);
or U11199 (N_11199,N_10894,N_10304);
nand U11200 (N_11200,N_10049,N_10183);
and U11201 (N_11201,N_10673,N_10394);
nor U11202 (N_11202,N_10101,N_10943);
xnor U11203 (N_11203,N_10654,N_10829);
nor U11204 (N_11204,N_10466,N_10940);
and U11205 (N_11205,N_10035,N_10015);
or U11206 (N_11206,N_10677,N_10968);
or U11207 (N_11207,N_10066,N_10521);
nor U11208 (N_11208,N_10904,N_10501);
nor U11209 (N_11209,N_10100,N_10180);
nand U11210 (N_11210,N_10584,N_10201);
nand U11211 (N_11211,N_10248,N_10915);
or U11212 (N_11212,N_10662,N_10255);
and U11213 (N_11213,N_10869,N_10778);
and U11214 (N_11214,N_10782,N_10513);
nand U11215 (N_11215,N_10752,N_10186);
and U11216 (N_11216,N_10293,N_10444);
and U11217 (N_11217,N_10802,N_10559);
nor U11218 (N_11218,N_10470,N_10649);
nor U11219 (N_11219,N_10246,N_10842);
nand U11220 (N_11220,N_10223,N_10458);
or U11221 (N_11221,N_10063,N_10321);
nor U11222 (N_11222,N_10217,N_10150);
or U11223 (N_11223,N_10892,N_10775);
nor U11224 (N_11224,N_10064,N_10900);
or U11225 (N_11225,N_10412,N_10515);
xnor U11226 (N_11226,N_10462,N_10507);
and U11227 (N_11227,N_10238,N_10235);
and U11228 (N_11228,N_10476,N_10379);
and U11229 (N_11229,N_10872,N_10815);
and U11230 (N_11230,N_10031,N_10463);
and U11231 (N_11231,N_10411,N_10128);
or U11232 (N_11232,N_10006,N_10851);
or U11233 (N_11233,N_10541,N_10875);
nor U11234 (N_11234,N_10942,N_10323);
nand U11235 (N_11235,N_10253,N_10881);
nor U11236 (N_11236,N_10322,N_10538);
nor U11237 (N_11237,N_10287,N_10854);
and U11238 (N_11238,N_10486,N_10067);
and U11239 (N_11239,N_10524,N_10731);
nand U11240 (N_11240,N_10539,N_10927);
nand U11241 (N_11241,N_10707,N_10228);
or U11242 (N_11242,N_10407,N_10612);
and U11243 (N_11243,N_10710,N_10908);
nor U11244 (N_11244,N_10945,N_10693);
nor U11245 (N_11245,N_10951,N_10993);
nand U11246 (N_11246,N_10240,N_10929);
or U11247 (N_11247,N_10350,N_10826);
nand U11248 (N_11248,N_10890,N_10435);
nand U11249 (N_11249,N_10610,N_10222);
nand U11250 (N_11250,N_10758,N_10871);
xor U11251 (N_11251,N_10795,N_10631);
and U11252 (N_11252,N_10275,N_10156);
or U11253 (N_11253,N_10094,N_10747);
nand U11254 (N_11254,N_10701,N_10903);
or U11255 (N_11255,N_10283,N_10744);
nand U11256 (N_11256,N_10108,N_10363);
nand U11257 (N_11257,N_10828,N_10069);
or U11258 (N_11258,N_10543,N_10037);
or U11259 (N_11259,N_10896,N_10973);
nor U11260 (N_11260,N_10295,N_10294);
nand U11261 (N_11261,N_10026,N_10099);
nor U11262 (N_11262,N_10846,N_10243);
nor U11263 (N_11263,N_10129,N_10637);
or U11264 (N_11264,N_10075,N_10120);
or U11265 (N_11265,N_10397,N_10708);
and U11266 (N_11266,N_10858,N_10114);
and U11267 (N_11267,N_10823,N_10965);
or U11268 (N_11268,N_10118,N_10779);
or U11269 (N_11269,N_10107,N_10019);
and U11270 (N_11270,N_10988,N_10548);
or U11271 (N_11271,N_10769,N_10499);
xnor U11272 (N_11272,N_10856,N_10398);
nor U11273 (N_11273,N_10695,N_10065);
nor U11274 (N_11274,N_10325,N_10553);
and U11275 (N_11275,N_10457,N_10745);
nand U11276 (N_11276,N_10452,N_10984);
nand U11277 (N_11277,N_10726,N_10226);
nand U11278 (N_11278,N_10667,N_10674);
xnor U11279 (N_11279,N_10848,N_10714);
or U11280 (N_11280,N_10874,N_10840);
or U11281 (N_11281,N_10665,N_10117);
nor U11282 (N_11282,N_10806,N_10985);
and U11283 (N_11283,N_10656,N_10098);
or U11284 (N_11284,N_10796,N_10650);
nor U11285 (N_11285,N_10317,N_10104);
and U11286 (N_11286,N_10562,N_10239);
or U11287 (N_11287,N_10225,N_10628);
xor U11288 (N_11288,N_10289,N_10743);
and U11289 (N_11289,N_10750,N_10864);
nor U11290 (N_11290,N_10569,N_10753);
or U11291 (N_11291,N_10863,N_10937);
or U11292 (N_11292,N_10518,N_10291);
or U11293 (N_11293,N_10590,N_10134);
xor U11294 (N_11294,N_10953,N_10338);
nand U11295 (N_11295,N_10332,N_10600);
xor U11296 (N_11296,N_10346,N_10257);
nor U11297 (N_11297,N_10800,N_10718);
and U11298 (N_11298,N_10761,N_10962);
nor U11299 (N_11299,N_10088,N_10148);
and U11300 (N_11300,N_10918,N_10265);
xnor U11301 (N_11301,N_10616,N_10372);
nor U11302 (N_11302,N_10961,N_10451);
xor U11303 (N_11303,N_10498,N_10924);
and U11304 (N_11304,N_10227,N_10948);
or U11305 (N_11305,N_10121,N_10390);
nor U11306 (N_11306,N_10136,N_10302);
or U11307 (N_11307,N_10554,N_10025);
nand U11308 (N_11308,N_10935,N_10793);
xnor U11309 (N_11309,N_10009,N_10595);
nor U11310 (N_11310,N_10742,N_10050);
nor U11311 (N_11311,N_10119,N_10419);
nand U11312 (N_11312,N_10036,N_10445);
or U11313 (N_11313,N_10914,N_10005);
nor U11314 (N_11314,N_10155,N_10301);
nand U11315 (N_11315,N_10781,N_10468);
and U11316 (N_11316,N_10946,N_10621);
nand U11317 (N_11317,N_10296,N_10424);
nand U11318 (N_11318,N_10697,N_10138);
nand U11319 (N_11319,N_10519,N_10509);
xnor U11320 (N_11320,N_10137,N_10556);
xor U11321 (N_11321,N_10262,N_10324);
or U11322 (N_11322,N_10822,N_10290);
xnor U11323 (N_11323,N_10133,N_10154);
nor U11324 (N_11324,N_10885,N_10110);
nor U11325 (N_11325,N_10532,N_10219);
xor U11326 (N_11326,N_10879,N_10905);
or U11327 (N_11327,N_10181,N_10581);
and U11328 (N_11328,N_10681,N_10273);
nand U11329 (N_11329,N_10535,N_10512);
nand U11330 (N_11330,N_10161,N_10429);
nor U11331 (N_11331,N_10151,N_10013);
or U11332 (N_11332,N_10756,N_10936);
and U11333 (N_11333,N_10016,N_10347);
xnor U11334 (N_11334,N_10218,N_10076);
or U11335 (N_11335,N_10920,N_10740);
or U11336 (N_11336,N_10565,N_10105);
or U11337 (N_11337,N_10377,N_10529);
and U11338 (N_11338,N_10056,N_10788);
or U11339 (N_11339,N_10906,N_10400);
and U11340 (N_11340,N_10465,N_10024);
nor U11341 (N_11341,N_10568,N_10176);
nor U11342 (N_11342,N_10095,N_10888);
and U11343 (N_11343,N_10763,N_10891);
xor U11344 (N_11344,N_10453,N_10339);
nor U11345 (N_11345,N_10426,N_10328);
and U11346 (N_11346,N_10179,N_10184);
nor U11347 (N_11347,N_10613,N_10808);
xor U11348 (N_11348,N_10456,N_10410);
and U11349 (N_11349,N_10922,N_10041);
and U11350 (N_11350,N_10316,N_10536);
and U11351 (N_11351,N_10837,N_10592);
nor U11352 (N_11352,N_10367,N_10078);
nand U11353 (N_11353,N_10506,N_10286);
nor U11354 (N_11354,N_10886,N_10949);
nand U11355 (N_11355,N_10481,N_10311);
and U11356 (N_11356,N_10003,N_10214);
and U11357 (N_11357,N_10522,N_10070);
xor U11358 (N_11358,N_10704,N_10970);
or U11359 (N_11359,N_10721,N_10599);
nor U11360 (N_11360,N_10669,N_10976);
xor U11361 (N_11361,N_10437,N_10389);
and U11362 (N_11362,N_10381,N_10921);
and U11363 (N_11363,N_10427,N_10417);
and U11364 (N_11364,N_10576,N_10002);
xnor U11365 (N_11365,N_10725,N_10799);
and U11366 (N_11366,N_10077,N_10190);
xor U11367 (N_11367,N_10689,N_10158);
and U11368 (N_11368,N_10496,N_10618);
nand U11369 (N_11369,N_10999,N_10593);
or U11370 (N_11370,N_10843,N_10431);
nand U11371 (N_11371,N_10224,N_10081);
and U11372 (N_11372,N_10089,N_10571);
or U11373 (N_11373,N_10836,N_10923);
and U11374 (N_11374,N_10617,N_10361);
nor U11375 (N_11375,N_10525,N_10633);
nand U11376 (N_11376,N_10355,N_10061);
nand U11377 (N_11377,N_10594,N_10860);
nand U11378 (N_11378,N_10954,N_10454);
nor U11379 (N_11379,N_10804,N_10611);
nor U11380 (N_11380,N_10608,N_10237);
nor U11381 (N_11381,N_10958,N_10392);
nor U11382 (N_11382,N_10087,N_10841);
or U11383 (N_11383,N_10475,N_10314);
or U11384 (N_11384,N_10057,N_10814);
and U11385 (N_11385,N_10197,N_10382);
or U11386 (N_11386,N_10643,N_10734);
and U11387 (N_11387,N_10040,N_10508);
nor U11388 (N_11388,N_10706,N_10034);
nand U11389 (N_11389,N_10698,N_10091);
nand U11390 (N_11390,N_10380,N_10022);
and U11391 (N_11391,N_10709,N_10642);
nor U11392 (N_11392,N_10549,N_10376);
and U11393 (N_11393,N_10447,N_10252);
nor U11394 (N_11394,N_10489,N_10820);
nor U11395 (N_11395,N_10817,N_10705);
nand U11396 (N_11396,N_10676,N_10130);
nand U11397 (N_11397,N_10072,N_10503);
and U11398 (N_11398,N_10028,N_10811);
xor U11399 (N_11399,N_10720,N_10220);
nor U11400 (N_11400,N_10374,N_10335);
and U11401 (N_11401,N_10048,N_10182);
or U11402 (N_11402,N_10831,N_10145);
or U11403 (N_11403,N_10975,N_10889);
nor U11404 (N_11404,N_10163,N_10648);
nor U11405 (N_11405,N_10691,N_10079);
nor U11406 (N_11406,N_10762,N_10368);
nor U11407 (N_11407,N_10629,N_10850);
nor U11408 (N_11408,N_10511,N_10490);
nor U11409 (N_11409,N_10672,N_10789);
nor U11410 (N_11410,N_10603,N_10852);
or U11411 (N_11411,N_10215,N_10203);
or U11412 (N_11412,N_10835,N_10234);
and U11413 (N_11413,N_10692,N_10106);
or U11414 (N_11414,N_10624,N_10047);
or U11415 (N_11415,N_10623,N_10212);
and U11416 (N_11416,N_10687,N_10343);
xnor U11417 (N_11417,N_10305,N_10168);
and U11418 (N_11418,N_10777,N_10577);
nand U11419 (N_11419,N_10626,N_10615);
and U11420 (N_11420,N_10231,N_10387);
nor U11421 (N_11421,N_10274,N_10533);
or U11422 (N_11422,N_10483,N_10979);
or U11423 (N_11423,N_10737,N_10313);
nand U11424 (N_11424,N_10279,N_10258);
or U11425 (N_11425,N_10732,N_10433);
nor U11426 (N_11426,N_10111,N_10528);
and U11427 (N_11427,N_10939,N_10256);
nor U11428 (N_11428,N_10330,N_10043);
or U11429 (N_11429,N_10682,N_10140);
nand U11430 (N_11430,N_10998,N_10504);
and U11431 (N_11431,N_10591,N_10733);
nor U11432 (N_11432,N_10298,N_10053);
or U11433 (N_11433,N_10344,N_10124);
or U11434 (N_11434,N_10583,N_10986);
nand U11435 (N_11435,N_10526,N_10173);
and U11436 (N_11436,N_10825,N_10523);
and U11437 (N_11437,N_10717,N_10178);
nand U11438 (N_11438,N_10552,N_10967);
xor U11439 (N_11439,N_10977,N_10434);
nor U11440 (N_11440,N_10216,N_10602);
or U11441 (N_11441,N_10309,N_10200);
and U11442 (N_11442,N_10474,N_10436);
nand U11443 (N_11443,N_10919,N_10471);
and U11444 (N_11444,N_10482,N_10438);
or U11445 (N_11445,N_10868,N_10308);
xnor U11446 (N_11446,N_10574,N_10785);
xnor U11447 (N_11447,N_10573,N_10385);
and U11448 (N_11448,N_10166,N_10636);
and U11449 (N_11449,N_10913,N_10386);
nor U11450 (N_11450,N_10866,N_10551);
xnor U11451 (N_11451,N_10093,N_10736);
or U11452 (N_11452,N_10333,N_10880);
and U11453 (N_11453,N_10646,N_10477);
or U11454 (N_11454,N_10688,N_10792);
nor U11455 (N_11455,N_10861,N_10989);
nand U11456 (N_11456,N_10764,N_10375);
nand U11457 (N_11457,N_10446,N_10131);
and U11458 (N_11458,N_10039,N_10011);
and U11459 (N_11459,N_10352,N_10634);
and U11460 (N_11460,N_10542,N_10109);
nand U11461 (N_11461,N_10658,N_10464);
nor U11462 (N_11462,N_10738,N_10084);
and U11463 (N_11463,N_10126,N_10187);
and U11464 (N_11464,N_10694,N_10080);
nor U11465 (N_11465,N_10947,N_10647);
nor U11466 (N_11466,N_10897,N_10211);
nand U11467 (N_11467,N_10351,N_10645);
nand U11468 (N_11468,N_10587,N_10336);
nand U11469 (N_11469,N_10784,N_10570);
or U11470 (N_11470,N_10285,N_10739);
nor U11471 (N_11471,N_10893,N_10365);
or U11472 (N_11472,N_10174,N_10751);
nor U11473 (N_11473,N_10700,N_10663);
and U11474 (N_11474,N_10422,N_10288);
nand U11475 (N_11475,N_10598,N_10711);
and U11476 (N_11476,N_10516,N_10632);
and U11477 (N_11477,N_10175,N_10774);
nor U11478 (N_11478,N_10198,N_10834);
nor U11479 (N_11479,N_10917,N_10853);
or U11480 (N_11480,N_10074,N_10334);
nand U11481 (N_11481,N_10030,N_10944);
nor U11482 (N_11482,N_10728,N_10073);
nand U11483 (N_11483,N_10263,N_10981);
nor U11484 (N_11484,N_10787,N_10208);
xor U11485 (N_11485,N_10766,N_10210);
nor U11486 (N_11486,N_10354,N_10932);
or U11487 (N_11487,N_10723,N_10303);
or U11488 (N_11488,N_10686,N_10270);
nand U11489 (N_11489,N_10383,N_10432);
or U11490 (N_11490,N_10086,N_10859);
nand U11491 (N_11491,N_10402,N_10557);
or U11492 (N_11492,N_10966,N_10797);
nand U11493 (N_11493,N_10606,N_10702);
nand U11494 (N_11494,N_10582,N_10683);
nand U11495 (N_11495,N_10358,N_10791);
and U11496 (N_11496,N_10249,N_10414);
nor U11497 (N_11497,N_10018,N_10449);
and U11498 (N_11498,N_10143,N_10276);
and U11499 (N_11499,N_10980,N_10461);
nor U11500 (N_11500,N_10004,N_10801);
or U11501 (N_11501,N_10609,N_10754);
nor U11502 (N_11502,N_10470,N_10915);
nor U11503 (N_11503,N_10578,N_10218);
nand U11504 (N_11504,N_10136,N_10082);
and U11505 (N_11505,N_10079,N_10591);
and U11506 (N_11506,N_10602,N_10441);
or U11507 (N_11507,N_10373,N_10049);
and U11508 (N_11508,N_10118,N_10228);
or U11509 (N_11509,N_10294,N_10299);
and U11510 (N_11510,N_10211,N_10988);
nand U11511 (N_11511,N_10876,N_10645);
or U11512 (N_11512,N_10829,N_10842);
and U11513 (N_11513,N_10683,N_10484);
nand U11514 (N_11514,N_10308,N_10853);
and U11515 (N_11515,N_10093,N_10448);
nand U11516 (N_11516,N_10640,N_10140);
and U11517 (N_11517,N_10991,N_10412);
and U11518 (N_11518,N_10283,N_10626);
xnor U11519 (N_11519,N_10774,N_10381);
xor U11520 (N_11520,N_10734,N_10377);
nand U11521 (N_11521,N_10789,N_10997);
and U11522 (N_11522,N_10086,N_10516);
nand U11523 (N_11523,N_10495,N_10675);
and U11524 (N_11524,N_10318,N_10591);
or U11525 (N_11525,N_10925,N_10485);
and U11526 (N_11526,N_10341,N_10176);
and U11527 (N_11527,N_10898,N_10551);
xor U11528 (N_11528,N_10251,N_10734);
and U11529 (N_11529,N_10581,N_10676);
and U11530 (N_11530,N_10600,N_10918);
nand U11531 (N_11531,N_10277,N_10793);
and U11532 (N_11532,N_10108,N_10937);
nand U11533 (N_11533,N_10015,N_10920);
and U11534 (N_11534,N_10903,N_10904);
and U11535 (N_11535,N_10227,N_10310);
or U11536 (N_11536,N_10446,N_10112);
nand U11537 (N_11537,N_10393,N_10491);
nand U11538 (N_11538,N_10841,N_10737);
xor U11539 (N_11539,N_10719,N_10225);
xor U11540 (N_11540,N_10611,N_10502);
nand U11541 (N_11541,N_10140,N_10041);
nand U11542 (N_11542,N_10957,N_10550);
nand U11543 (N_11543,N_10963,N_10662);
nand U11544 (N_11544,N_10044,N_10314);
and U11545 (N_11545,N_10923,N_10370);
and U11546 (N_11546,N_10962,N_10767);
and U11547 (N_11547,N_10373,N_10313);
nand U11548 (N_11548,N_10027,N_10573);
xnor U11549 (N_11549,N_10997,N_10302);
or U11550 (N_11550,N_10053,N_10490);
or U11551 (N_11551,N_10659,N_10839);
and U11552 (N_11552,N_10593,N_10586);
nor U11553 (N_11553,N_10828,N_10665);
nor U11554 (N_11554,N_10688,N_10458);
xnor U11555 (N_11555,N_10697,N_10334);
nor U11556 (N_11556,N_10888,N_10660);
nor U11557 (N_11557,N_10597,N_10555);
or U11558 (N_11558,N_10732,N_10022);
nand U11559 (N_11559,N_10114,N_10449);
or U11560 (N_11560,N_10152,N_10257);
nand U11561 (N_11561,N_10656,N_10499);
nand U11562 (N_11562,N_10816,N_10446);
or U11563 (N_11563,N_10017,N_10313);
and U11564 (N_11564,N_10743,N_10453);
and U11565 (N_11565,N_10420,N_10037);
nor U11566 (N_11566,N_10648,N_10553);
and U11567 (N_11567,N_10189,N_10767);
nor U11568 (N_11568,N_10466,N_10857);
or U11569 (N_11569,N_10776,N_10960);
or U11570 (N_11570,N_10450,N_10529);
and U11571 (N_11571,N_10588,N_10834);
and U11572 (N_11572,N_10860,N_10626);
nor U11573 (N_11573,N_10145,N_10965);
nor U11574 (N_11574,N_10921,N_10882);
and U11575 (N_11575,N_10122,N_10129);
or U11576 (N_11576,N_10793,N_10392);
nand U11577 (N_11577,N_10286,N_10872);
or U11578 (N_11578,N_10211,N_10569);
or U11579 (N_11579,N_10014,N_10320);
nor U11580 (N_11580,N_10113,N_10548);
or U11581 (N_11581,N_10401,N_10500);
nand U11582 (N_11582,N_10232,N_10353);
xor U11583 (N_11583,N_10520,N_10754);
or U11584 (N_11584,N_10232,N_10963);
or U11585 (N_11585,N_10447,N_10777);
and U11586 (N_11586,N_10529,N_10671);
and U11587 (N_11587,N_10591,N_10224);
and U11588 (N_11588,N_10316,N_10915);
or U11589 (N_11589,N_10408,N_10991);
nor U11590 (N_11590,N_10688,N_10270);
nor U11591 (N_11591,N_10284,N_10879);
xor U11592 (N_11592,N_10993,N_10029);
nor U11593 (N_11593,N_10903,N_10463);
nor U11594 (N_11594,N_10234,N_10490);
nand U11595 (N_11595,N_10842,N_10980);
and U11596 (N_11596,N_10599,N_10127);
nor U11597 (N_11597,N_10114,N_10739);
nand U11598 (N_11598,N_10949,N_10364);
and U11599 (N_11599,N_10823,N_10025);
nand U11600 (N_11600,N_10424,N_10263);
nand U11601 (N_11601,N_10541,N_10953);
xor U11602 (N_11602,N_10792,N_10179);
nand U11603 (N_11603,N_10917,N_10933);
nand U11604 (N_11604,N_10692,N_10191);
nand U11605 (N_11605,N_10678,N_10771);
nand U11606 (N_11606,N_10829,N_10099);
xnor U11607 (N_11607,N_10538,N_10992);
and U11608 (N_11608,N_10701,N_10289);
nand U11609 (N_11609,N_10817,N_10655);
nor U11610 (N_11610,N_10135,N_10624);
and U11611 (N_11611,N_10073,N_10352);
xnor U11612 (N_11612,N_10370,N_10990);
nor U11613 (N_11613,N_10711,N_10181);
or U11614 (N_11614,N_10174,N_10046);
nand U11615 (N_11615,N_10749,N_10583);
nand U11616 (N_11616,N_10705,N_10921);
nand U11617 (N_11617,N_10204,N_10846);
nand U11618 (N_11618,N_10023,N_10572);
nor U11619 (N_11619,N_10159,N_10120);
nor U11620 (N_11620,N_10919,N_10682);
nand U11621 (N_11621,N_10150,N_10438);
or U11622 (N_11622,N_10635,N_10123);
nand U11623 (N_11623,N_10450,N_10267);
and U11624 (N_11624,N_10351,N_10152);
or U11625 (N_11625,N_10096,N_10567);
nor U11626 (N_11626,N_10413,N_10624);
and U11627 (N_11627,N_10539,N_10412);
and U11628 (N_11628,N_10180,N_10748);
or U11629 (N_11629,N_10806,N_10369);
or U11630 (N_11630,N_10502,N_10358);
xnor U11631 (N_11631,N_10167,N_10458);
nor U11632 (N_11632,N_10129,N_10081);
or U11633 (N_11633,N_10735,N_10637);
nand U11634 (N_11634,N_10319,N_10652);
nor U11635 (N_11635,N_10797,N_10667);
nand U11636 (N_11636,N_10909,N_10459);
xor U11637 (N_11637,N_10174,N_10018);
or U11638 (N_11638,N_10673,N_10921);
xor U11639 (N_11639,N_10567,N_10154);
nand U11640 (N_11640,N_10192,N_10252);
and U11641 (N_11641,N_10171,N_10646);
xor U11642 (N_11642,N_10682,N_10524);
and U11643 (N_11643,N_10907,N_10867);
nor U11644 (N_11644,N_10712,N_10987);
nand U11645 (N_11645,N_10012,N_10081);
xnor U11646 (N_11646,N_10763,N_10363);
nor U11647 (N_11647,N_10363,N_10758);
nor U11648 (N_11648,N_10204,N_10859);
or U11649 (N_11649,N_10374,N_10072);
and U11650 (N_11650,N_10296,N_10149);
and U11651 (N_11651,N_10916,N_10278);
nor U11652 (N_11652,N_10800,N_10821);
and U11653 (N_11653,N_10019,N_10170);
or U11654 (N_11654,N_10538,N_10334);
nor U11655 (N_11655,N_10554,N_10147);
and U11656 (N_11656,N_10330,N_10498);
xnor U11657 (N_11657,N_10957,N_10729);
and U11658 (N_11658,N_10489,N_10673);
or U11659 (N_11659,N_10566,N_10134);
nor U11660 (N_11660,N_10775,N_10588);
and U11661 (N_11661,N_10748,N_10348);
nor U11662 (N_11662,N_10804,N_10071);
or U11663 (N_11663,N_10431,N_10815);
or U11664 (N_11664,N_10966,N_10504);
or U11665 (N_11665,N_10747,N_10386);
xnor U11666 (N_11666,N_10395,N_10159);
nor U11667 (N_11667,N_10048,N_10859);
or U11668 (N_11668,N_10878,N_10676);
or U11669 (N_11669,N_10342,N_10873);
nor U11670 (N_11670,N_10695,N_10393);
xor U11671 (N_11671,N_10432,N_10625);
nand U11672 (N_11672,N_10045,N_10208);
nor U11673 (N_11673,N_10579,N_10429);
nor U11674 (N_11674,N_10627,N_10099);
nor U11675 (N_11675,N_10990,N_10510);
nand U11676 (N_11676,N_10735,N_10482);
and U11677 (N_11677,N_10250,N_10946);
nand U11678 (N_11678,N_10937,N_10401);
nor U11679 (N_11679,N_10643,N_10823);
nor U11680 (N_11680,N_10780,N_10071);
nor U11681 (N_11681,N_10649,N_10167);
or U11682 (N_11682,N_10786,N_10030);
or U11683 (N_11683,N_10387,N_10653);
nand U11684 (N_11684,N_10635,N_10880);
and U11685 (N_11685,N_10299,N_10723);
or U11686 (N_11686,N_10991,N_10125);
or U11687 (N_11687,N_10820,N_10211);
xor U11688 (N_11688,N_10594,N_10893);
xor U11689 (N_11689,N_10420,N_10374);
and U11690 (N_11690,N_10907,N_10026);
and U11691 (N_11691,N_10134,N_10257);
nand U11692 (N_11692,N_10113,N_10337);
and U11693 (N_11693,N_10363,N_10442);
nor U11694 (N_11694,N_10715,N_10380);
nand U11695 (N_11695,N_10078,N_10176);
or U11696 (N_11696,N_10766,N_10645);
or U11697 (N_11697,N_10692,N_10451);
or U11698 (N_11698,N_10583,N_10215);
nor U11699 (N_11699,N_10898,N_10957);
and U11700 (N_11700,N_10074,N_10066);
nand U11701 (N_11701,N_10703,N_10764);
nand U11702 (N_11702,N_10001,N_10606);
or U11703 (N_11703,N_10723,N_10162);
or U11704 (N_11704,N_10814,N_10577);
nand U11705 (N_11705,N_10326,N_10169);
or U11706 (N_11706,N_10697,N_10007);
or U11707 (N_11707,N_10698,N_10836);
and U11708 (N_11708,N_10994,N_10516);
nor U11709 (N_11709,N_10659,N_10230);
nand U11710 (N_11710,N_10281,N_10767);
nand U11711 (N_11711,N_10702,N_10481);
and U11712 (N_11712,N_10360,N_10677);
nor U11713 (N_11713,N_10536,N_10569);
nand U11714 (N_11714,N_10794,N_10101);
nor U11715 (N_11715,N_10573,N_10356);
xnor U11716 (N_11716,N_10397,N_10289);
or U11717 (N_11717,N_10688,N_10249);
or U11718 (N_11718,N_10091,N_10930);
nor U11719 (N_11719,N_10506,N_10130);
or U11720 (N_11720,N_10952,N_10776);
xor U11721 (N_11721,N_10013,N_10311);
nor U11722 (N_11722,N_10670,N_10541);
nand U11723 (N_11723,N_10741,N_10803);
or U11724 (N_11724,N_10490,N_10607);
nor U11725 (N_11725,N_10492,N_10985);
or U11726 (N_11726,N_10197,N_10661);
and U11727 (N_11727,N_10963,N_10438);
nor U11728 (N_11728,N_10563,N_10089);
and U11729 (N_11729,N_10267,N_10868);
nand U11730 (N_11730,N_10744,N_10854);
nor U11731 (N_11731,N_10959,N_10184);
nor U11732 (N_11732,N_10012,N_10057);
or U11733 (N_11733,N_10108,N_10042);
or U11734 (N_11734,N_10205,N_10397);
nand U11735 (N_11735,N_10404,N_10059);
xor U11736 (N_11736,N_10644,N_10538);
and U11737 (N_11737,N_10470,N_10164);
and U11738 (N_11738,N_10777,N_10477);
nand U11739 (N_11739,N_10180,N_10281);
nor U11740 (N_11740,N_10675,N_10551);
or U11741 (N_11741,N_10149,N_10151);
or U11742 (N_11742,N_10002,N_10108);
xor U11743 (N_11743,N_10832,N_10861);
nor U11744 (N_11744,N_10185,N_10827);
and U11745 (N_11745,N_10359,N_10406);
nor U11746 (N_11746,N_10850,N_10973);
and U11747 (N_11747,N_10351,N_10414);
or U11748 (N_11748,N_10172,N_10253);
or U11749 (N_11749,N_10178,N_10877);
nand U11750 (N_11750,N_10995,N_10308);
and U11751 (N_11751,N_10173,N_10971);
xnor U11752 (N_11752,N_10319,N_10351);
nor U11753 (N_11753,N_10713,N_10618);
or U11754 (N_11754,N_10597,N_10152);
nand U11755 (N_11755,N_10710,N_10453);
nor U11756 (N_11756,N_10293,N_10116);
or U11757 (N_11757,N_10552,N_10573);
xnor U11758 (N_11758,N_10082,N_10172);
nor U11759 (N_11759,N_10870,N_10768);
or U11760 (N_11760,N_10845,N_10532);
and U11761 (N_11761,N_10661,N_10179);
nand U11762 (N_11762,N_10412,N_10811);
nand U11763 (N_11763,N_10938,N_10598);
or U11764 (N_11764,N_10386,N_10207);
nand U11765 (N_11765,N_10602,N_10104);
xor U11766 (N_11766,N_10508,N_10031);
or U11767 (N_11767,N_10013,N_10659);
nor U11768 (N_11768,N_10738,N_10833);
and U11769 (N_11769,N_10461,N_10886);
nand U11770 (N_11770,N_10671,N_10730);
nor U11771 (N_11771,N_10014,N_10556);
nor U11772 (N_11772,N_10535,N_10523);
or U11773 (N_11773,N_10269,N_10313);
nand U11774 (N_11774,N_10836,N_10835);
or U11775 (N_11775,N_10291,N_10472);
xor U11776 (N_11776,N_10167,N_10281);
or U11777 (N_11777,N_10113,N_10355);
nor U11778 (N_11778,N_10613,N_10799);
nand U11779 (N_11779,N_10329,N_10046);
nand U11780 (N_11780,N_10877,N_10690);
nor U11781 (N_11781,N_10850,N_10020);
nand U11782 (N_11782,N_10456,N_10583);
nand U11783 (N_11783,N_10832,N_10325);
nor U11784 (N_11784,N_10701,N_10913);
xor U11785 (N_11785,N_10310,N_10466);
or U11786 (N_11786,N_10622,N_10409);
nor U11787 (N_11787,N_10346,N_10874);
or U11788 (N_11788,N_10162,N_10151);
nor U11789 (N_11789,N_10528,N_10164);
nand U11790 (N_11790,N_10278,N_10664);
xor U11791 (N_11791,N_10524,N_10944);
nor U11792 (N_11792,N_10019,N_10061);
and U11793 (N_11793,N_10678,N_10286);
nand U11794 (N_11794,N_10347,N_10792);
nor U11795 (N_11795,N_10857,N_10064);
nand U11796 (N_11796,N_10077,N_10181);
and U11797 (N_11797,N_10211,N_10168);
nand U11798 (N_11798,N_10336,N_10062);
or U11799 (N_11799,N_10864,N_10294);
nor U11800 (N_11800,N_10276,N_10046);
nand U11801 (N_11801,N_10725,N_10280);
nand U11802 (N_11802,N_10991,N_10458);
nor U11803 (N_11803,N_10209,N_10935);
nand U11804 (N_11804,N_10092,N_10067);
and U11805 (N_11805,N_10108,N_10729);
nand U11806 (N_11806,N_10166,N_10924);
nand U11807 (N_11807,N_10814,N_10361);
nand U11808 (N_11808,N_10676,N_10517);
or U11809 (N_11809,N_10619,N_10804);
xor U11810 (N_11810,N_10553,N_10481);
nor U11811 (N_11811,N_10764,N_10131);
or U11812 (N_11812,N_10023,N_10298);
or U11813 (N_11813,N_10971,N_10773);
nand U11814 (N_11814,N_10668,N_10293);
and U11815 (N_11815,N_10593,N_10971);
nor U11816 (N_11816,N_10243,N_10295);
or U11817 (N_11817,N_10024,N_10279);
nand U11818 (N_11818,N_10793,N_10235);
or U11819 (N_11819,N_10567,N_10819);
xor U11820 (N_11820,N_10561,N_10627);
nor U11821 (N_11821,N_10900,N_10925);
or U11822 (N_11822,N_10048,N_10782);
and U11823 (N_11823,N_10336,N_10145);
and U11824 (N_11824,N_10668,N_10817);
nand U11825 (N_11825,N_10305,N_10659);
and U11826 (N_11826,N_10681,N_10623);
nand U11827 (N_11827,N_10874,N_10407);
or U11828 (N_11828,N_10462,N_10752);
xor U11829 (N_11829,N_10464,N_10314);
xor U11830 (N_11830,N_10794,N_10061);
or U11831 (N_11831,N_10482,N_10901);
and U11832 (N_11832,N_10614,N_10615);
or U11833 (N_11833,N_10702,N_10076);
or U11834 (N_11834,N_10058,N_10117);
nor U11835 (N_11835,N_10899,N_10784);
nor U11836 (N_11836,N_10099,N_10214);
nand U11837 (N_11837,N_10093,N_10271);
and U11838 (N_11838,N_10313,N_10736);
nand U11839 (N_11839,N_10979,N_10725);
nand U11840 (N_11840,N_10980,N_10552);
nand U11841 (N_11841,N_10439,N_10610);
nor U11842 (N_11842,N_10651,N_10175);
nand U11843 (N_11843,N_10595,N_10273);
nand U11844 (N_11844,N_10853,N_10960);
nor U11845 (N_11845,N_10052,N_10955);
and U11846 (N_11846,N_10911,N_10481);
nand U11847 (N_11847,N_10859,N_10581);
or U11848 (N_11848,N_10377,N_10888);
or U11849 (N_11849,N_10202,N_10583);
nor U11850 (N_11850,N_10969,N_10785);
nor U11851 (N_11851,N_10882,N_10052);
and U11852 (N_11852,N_10750,N_10333);
nand U11853 (N_11853,N_10654,N_10932);
and U11854 (N_11854,N_10349,N_10285);
nor U11855 (N_11855,N_10613,N_10894);
or U11856 (N_11856,N_10902,N_10190);
xor U11857 (N_11857,N_10636,N_10526);
and U11858 (N_11858,N_10591,N_10095);
nor U11859 (N_11859,N_10604,N_10239);
nor U11860 (N_11860,N_10984,N_10312);
nor U11861 (N_11861,N_10181,N_10566);
or U11862 (N_11862,N_10625,N_10445);
xor U11863 (N_11863,N_10663,N_10569);
or U11864 (N_11864,N_10975,N_10858);
or U11865 (N_11865,N_10714,N_10374);
xor U11866 (N_11866,N_10440,N_10089);
nand U11867 (N_11867,N_10440,N_10706);
or U11868 (N_11868,N_10437,N_10905);
and U11869 (N_11869,N_10919,N_10320);
nor U11870 (N_11870,N_10022,N_10728);
and U11871 (N_11871,N_10617,N_10074);
and U11872 (N_11872,N_10642,N_10126);
or U11873 (N_11873,N_10927,N_10222);
and U11874 (N_11874,N_10864,N_10621);
nor U11875 (N_11875,N_10064,N_10458);
and U11876 (N_11876,N_10517,N_10935);
nor U11877 (N_11877,N_10946,N_10025);
nor U11878 (N_11878,N_10379,N_10085);
or U11879 (N_11879,N_10944,N_10519);
or U11880 (N_11880,N_10757,N_10229);
nand U11881 (N_11881,N_10026,N_10877);
or U11882 (N_11882,N_10583,N_10764);
nor U11883 (N_11883,N_10105,N_10529);
nand U11884 (N_11884,N_10896,N_10665);
nand U11885 (N_11885,N_10611,N_10643);
nand U11886 (N_11886,N_10594,N_10271);
and U11887 (N_11887,N_10754,N_10407);
and U11888 (N_11888,N_10196,N_10953);
and U11889 (N_11889,N_10681,N_10661);
nand U11890 (N_11890,N_10784,N_10472);
and U11891 (N_11891,N_10591,N_10979);
or U11892 (N_11892,N_10665,N_10418);
nand U11893 (N_11893,N_10544,N_10092);
or U11894 (N_11894,N_10141,N_10207);
nor U11895 (N_11895,N_10367,N_10086);
nor U11896 (N_11896,N_10233,N_10131);
or U11897 (N_11897,N_10773,N_10045);
nand U11898 (N_11898,N_10761,N_10950);
or U11899 (N_11899,N_10133,N_10459);
or U11900 (N_11900,N_10253,N_10742);
or U11901 (N_11901,N_10533,N_10424);
or U11902 (N_11902,N_10457,N_10438);
nand U11903 (N_11903,N_10188,N_10789);
nor U11904 (N_11904,N_10962,N_10571);
xnor U11905 (N_11905,N_10302,N_10999);
xnor U11906 (N_11906,N_10243,N_10386);
nand U11907 (N_11907,N_10694,N_10266);
nor U11908 (N_11908,N_10167,N_10706);
or U11909 (N_11909,N_10232,N_10091);
and U11910 (N_11910,N_10049,N_10022);
or U11911 (N_11911,N_10102,N_10580);
and U11912 (N_11912,N_10677,N_10905);
or U11913 (N_11913,N_10865,N_10135);
and U11914 (N_11914,N_10934,N_10147);
or U11915 (N_11915,N_10192,N_10414);
and U11916 (N_11916,N_10551,N_10925);
nor U11917 (N_11917,N_10971,N_10595);
nor U11918 (N_11918,N_10124,N_10707);
nor U11919 (N_11919,N_10443,N_10835);
xor U11920 (N_11920,N_10534,N_10240);
nor U11921 (N_11921,N_10641,N_10463);
or U11922 (N_11922,N_10082,N_10878);
nand U11923 (N_11923,N_10654,N_10476);
or U11924 (N_11924,N_10967,N_10670);
and U11925 (N_11925,N_10622,N_10786);
nand U11926 (N_11926,N_10460,N_10931);
nor U11927 (N_11927,N_10936,N_10975);
nand U11928 (N_11928,N_10920,N_10130);
and U11929 (N_11929,N_10539,N_10883);
nor U11930 (N_11930,N_10573,N_10442);
xnor U11931 (N_11931,N_10967,N_10436);
nand U11932 (N_11932,N_10567,N_10412);
xnor U11933 (N_11933,N_10090,N_10362);
nor U11934 (N_11934,N_10307,N_10527);
xnor U11935 (N_11935,N_10557,N_10226);
and U11936 (N_11936,N_10137,N_10655);
and U11937 (N_11937,N_10227,N_10241);
nor U11938 (N_11938,N_10178,N_10451);
nand U11939 (N_11939,N_10254,N_10524);
nand U11940 (N_11940,N_10976,N_10468);
and U11941 (N_11941,N_10012,N_10002);
nand U11942 (N_11942,N_10608,N_10399);
nor U11943 (N_11943,N_10313,N_10152);
nor U11944 (N_11944,N_10673,N_10072);
nand U11945 (N_11945,N_10588,N_10809);
nand U11946 (N_11946,N_10093,N_10836);
nor U11947 (N_11947,N_10289,N_10945);
or U11948 (N_11948,N_10631,N_10659);
and U11949 (N_11949,N_10392,N_10957);
and U11950 (N_11950,N_10122,N_10901);
nand U11951 (N_11951,N_10529,N_10066);
and U11952 (N_11952,N_10137,N_10778);
nand U11953 (N_11953,N_10400,N_10966);
nor U11954 (N_11954,N_10390,N_10812);
and U11955 (N_11955,N_10585,N_10650);
nand U11956 (N_11956,N_10878,N_10444);
or U11957 (N_11957,N_10104,N_10898);
and U11958 (N_11958,N_10589,N_10122);
nor U11959 (N_11959,N_10193,N_10816);
xor U11960 (N_11960,N_10082,N_10650);
and U11961 (N_11961,N_10392,N_10696);
and U11962 (N_11962,N_10358,N_10610);
and U11963 (N_11963,N_10293,N_10808);
and U11964 (N_11964,N_10670,N_10232);
nor U11965 (N_11965,N_10053,N_10941);
or U11966 (N_11966,N_10760,N_10766);
nand U11967 (N_11967,N_10217,N_10487);
nand U11968 (N_11968,N_10570,N_10705);
and U11969 (N_11969,N_10434,N_10425);
and U11970 (N_11970,N_10928,N_10226);
nor U11971 (N_11971,N_10571,N_10149);
xnor U11972 (N_11972,N_10397,N_10623);
or U11973 (N_11973,N_10360,N_10911);
or U11974 (N_11974,N_10978,N_10586);
nand U11975 (N_11975,N_10665,N_10724);
nand U11976 (N_11976,N_10107,N_10135);
nor U11977 (N_11977,N_10685,N_10448);
xor U11978 (N_11978,N_10166,N_10450);
nand U11979 (N_11979,N_10464,N_10691);
and U11980 (N_11980,N_10972,N_10477);
nor U11981 (N_11981,N_10829,N_10154);
or U11982 (N_11982,N_10557,N_10941);
or U11983 (N_11983,N_10862,N_10155);
and U11984 (N_11984,N_10913,N_10408);
nor U11985 (N_11985,N_10915,N_10451);
xor U11986 (N_11986,N_10370,N_10006);
nor U11987 (N_11987,N_10871,N_10765);
nor U11988 (N_11988,N_10173,N_10668);
nor U11989 (N_11989,N_10710,N_10985);
nand U11990 (N_11990,N_10225,N_10073);
nor U11991 (N_11991,N_10807,N_10786);
nor U11992 (N_11992,N_10466,N_10285);
xnor U11993 (N_11993,N_10266,N_10442);
or U11994 (N_11994,N_10627,N_10076);
or U11995 (N_11995,N_10030,N_10129);
nand U11996 (N_11996,N_10168,N_10378);
nor U11997 (N_11997,N_10118,N_10679);
nor U11998 (N_11998,N_10176,N_10102);
nand U11999 (N_11999,N_10158,N_10657);
nor U12000 (N_12000,N_11135,N_11571);
or U12001 (N_12001,N_11228,N_11494);
nand U12002 (N_12002,N_11021,N_11885);
or U12003 (N_12003,N_11102,N_11967);
xor U12004 (N_12004,N_11321,N_11703);
nor U12005 (N_12005,N_11841,N_11618);
nor U12006 (N_12006,N_11659,N_11392);
nand U12007 (N_12007,N_11338,N_11906);
or U12008 (N_12008,N_11755,N_11534);
and U12009 (N_12009,N_11472,N_11501);
nand U12010 (N_12010,N_11203,N_11638);
nand U12011 (N_12011,N_11700,N_11038);
nand U12012 (N_12012,N_11729,N_11304);
nor U12013 (N_12013,N_11427,N_11836);
xor U12014 (N_12014,N_11145,N_11679);
and U12015 (N_12015,N_11759,N_11599);
xnor U12016 (N_12016,N_11593,N_11281);
and U12017 (N_12017,N_11344,N_11044);
and U12018 (N_12018,N_11452,N_11006);
and U12019 (N_12019,N_11750,N_11416);
and U12020 (N_12020,N_11737,N_11847);
nor U12021 (N_12021,N_11129,N_11968);
or U12022 (N_12022,N_11943,N_11349);
nand U12023 (N_12023,N_11456,N_11610);
and U12024 (N_12024,N_11993,N_11916);
or U12025 (N_12025,N_11589,N_11517);
or U12026 (N_12026,N_11300,N_11326);
nand U12027 (N_12027,N_11185,N_11165);
and U12028 (N_12028,N_11786,N_11744);
nor U12029 (N_12029,N_11592,N_11940);
or U12030 (N_12030,N_11341,N_11290);
nor U12031 (N_12031,N_11495,N_11143);
nor U12032 (N_12032,N_11381,N_11560);
or U12033 (N_12033,N_11011,N_11698);
xor U12034 (N_12034,N_11407,N_11773);
and U12035 (N_12035,N_11628,N_11696);
or U12036 (N_12036,N_11106,N_11764);
or U12037 (N_12037,N_11997,N_11117);
nor U12038 (N_12038,N_11438,N_11709);
nor U12039 (N_12039,N_11607,N_11119);
and U12040 (N_12040,N_11098,N_11911);
or U12041 (N_12041,N_11633,N_11950);
and U12042 (N_12042,N_11431,N_11666);
nand U12043 (N_12043,N_11842,N_11315);
and U12044 (N_12044,N_11749,N_11463);
xor U12045 (N_12045,N_11374,N_11208);
or U12046 (N_12046,N_11367,N_11311);
and U12047 (N_12047,N_11704,N_11382);
nor U12048 (N_12048,N_11273,N_11234);
or U12049 (N_12049,N_11296,N_11695);
and U12050 (N_12050,N_11733,N_11664);
and U12051 (N_12051,N_11174,N_11964);
xnor U12052 (N_12052,N_11553,N_11516);
nand U12053 (N_12053,N_11752,N_11858);
and U12054 (N_12054,N_11319,N_11863);
and U12055 (N_12055,N_11913,N_11909);
nand U12056 (N_12056,N_11265,N_11678);
nor U12057 (N_12057,N_11897,N_11433);
nand U12058 (N_12058,N_11107,N_11739);
or U12059 (N_12059,N_11328,N_11160);
nand U12060 (N_12060,N_11167,N_11423);
and U12061 (N_12061,N_11757,N_11142);
and U12062 (N_12062,N_11201,N_11039);
and U12063 (N_12063,N_11364,N_11820);
nand U12064 (N_12064,N_11153,N_11450);
xnor U12065 (N_12065,N_11988,N_11594);
or U12066 (N_12066,N_11653,N_11198);
and U12067 (N_12067,N_11444,N_11280);
nand U12068 (N_12068,N_11957,N_11779);
nand U12069 (N_12069,N_11715,N_11510);
and U12070 (N_12070,N_11697,N_11683);
or U12071 (N_12071,N_11730,N_11164);
and U12072 (N_12072,N_11978,N_11914);
or U12073 (N_12073,N_11542,N_11806);
nor U12074 (N_12074,N_11958,N_11190);
nor U12075 (N_12075,N_11413,N_11702);
nor U12076 (N_12076,N_11356,N_11357);
and U12077 (N_12077,N_11802,N_11561);
nor U12078 (N_12078,N_11071,N_11948);
and U12079 (N_12079,N_11229,N_11788);
or U12080 (N_12080,N_11034,N_11708);
xor U12081 (N_12081,N_11713,N_11591);
nor U12082 (N_12082,N_11566,N_11912);
xnor U12083 (N_12083,N_11101,N_11742);
and U12084 (N_12084,N_11987,N_11536);
and U12085 (N_12085,N_11838,N_11782);
and U12086 (N_12086,N_11794,N_11166);
nor U12087 (N_12087,N_11324,N_11586);
or U12088 (N_12088,N_11353,N_11279);
xor U12089 (N_12089,N_11045,N_11617);
and U12090 (N_12090,N_11230,N_11099);
nand U12091 (N_12091,N_11146,N_11642);
nor U12092 (N_12092,N_11677,N_11161);
xnor U12093 (N_12093,N_11078,N_11148);
and U12094 (N_12094,N_11524,N_11616);
xnor U12095 (N_12095,N_11743,N_11317);
nand U12096 (N_12096,N_11938,N_11065);
nor U12097 (N_12097,N_11196,N_11475);
and U12098 (N_12098,N_11012,N_11956);
or U12099 (N_12099,N_11687,N_11865);
nand U12100 (N_12100,N_11226,N_11428);
nor U12101 (N_12101,N_11981,N_11640);
nor U12102 (N_12102,N_11636,N_11086);
nor U12103 (N_12103,N_11037,N_11422);
nor U12104 (N_12104,N_11798,N_11067);
nand U12105 (N_12105,N_11665,N_11725);
or U12106 (N_12106,N_11758,N_11881);
and U12107 (N_12107,N_11077,N_11796);
xor U12108 (N_12108,N_11396,N_11545);
nor U12109 (N_12109,N_11057,N_11890);
and U12110 (N_12110,N_11900,N_11479);
nand U12111 (N_12111,N_11249,N_11803);
nand U12112 (N_12112,N_11685,N_11974);
xnor U12113 (N_12113,N_11060,N_11630);
nand U12114 (N_12114,N_11309,N_11676);
nand U12115 (N_12115,N_11944,N_11351);
nor U12116 (N_12116,N_11492,N_11980);
and U12117 (N_12117,N_11046,N_11136);
nand U12118 (N_12118,N_11606,N_11214);
nand U12119 (N_12119,N_11140,N_11110);
and U12120 (N_12120,N_11929,N_11888);
and U12121 (N_12121,N_11476,N_11787);
and U12122 (N_12122,N_11503,N_11092);
or U12123 (N_12123,N_11031,N_11986);
and U12124 (N_12124,N_11923,N_11732);
nor U12125 (N_12125,N_11932,N_11043);
and U12126 (N_12126,N_11570,N_11850);
nor U12127 (N_12127,N_11483,N_11731);
nand U12128 (N_12128,N_11118,N_11019);
and U12129 (N_12129,N_11445,N_11761);
and U12130 (N_12130,N_11042,N_11216);
or U12131 (N_12131,N_11139,N_11651);
or U12132 (N_12132,N_11939,N_11079);
or U12133 (N_12133,N_11626,N_11849);
nand U12134 (N_12134,N_11096,N_11833);
nand U12135 (N_12135,N_11669,N_11104);
nor U12136 (N_12136,N_11578,N_11706);
or U12137 (N_12137,N_11276,N_11920);
or U12138 (N_12138,N_11998,N_11083);
nand U12139 (N_12139,N_11644,N_11791);
or U12140 (N_12140,N_11500,N_11574);
nand U12141 (N_12141,N_11675,N_11984);
and U12142 (N_12142,N_11391,N_11657);
nor U12143 (N_12143,N_11686,N_11152);
nand U12144 (N_12144,N_11793,N_11267);
or U12145 (N_12145,N_11187,N_11063);
or U12146 (N_12146,N_11587,N_11222);
and U12147 (N_12147,N_11223,N_11648);
nor U12148 (N_12148,N_11903,N_11816);
nand U12149 (N_12149,N_11023,N_11255);
and U12150 (N_12150,N_11360,N_11851);
and U12151 (N_12151,N_11013,N_11514);
nor U12152 (N_12152,N_11458,N_11859);
nor U12153 (N_12153,N_11499,N_11236);
nand U12154 (N_12154,N_11585,N_11085);
nor U12155 (N_12155,N_11928,N_11639);
and U12156 (N_12156,N_11699,N_11384);
nor U12157 (N_12157,N_11965,N_11840);
nand U12158 (N_12158,N_11496,N_11723);
nand U12159 (N_12159,N_11466,N_11380);
nand U12160 (N_12160,N_11470,N_11763);
nand U12161 (N_12161,N_11959,N_11128);
nand U12162 (N_12162,N_11537,N_11507);
nor U12163 (N_12163,N_11263,N_11745);
xor U12164 (N_12164,N_11058,N_11896);
or U12165 (N_12165,N_11783,N_11398);
nor U12166 (N_12166,N_11995,N_11753);
nor U12167 (N_12167,N_11760,N_11894);
and U12168 (N_12168,N_11949,N_11855);
nor U12169 (N_12169,N_11435,N_11714);
nand U12170 (N_12170,N_11432,N_11935);
nand U12171 (N_12171,N_11907,N_11918);
or U12172 (N_12172,N_11688,N_11168);
or U12173 (N_12173,N_11875,N_11989);
and U12174 (N_12174,N_11689,N_11778);
or U12175 (N_12175,N_11879,N_11401);
and U12176 (N_12176,N_11191,N_11970);
nor U12177 (N_12177,N_11632,N_11523);
and U12178 (N_12178,N_11557,N_11634);
nand U12179 (N_12179,N_11133,N_11370);
and U12180 (N_12180,N_11905,N_11212);
and U12181 (N_12181,N_11355,N_11769);
nand U12182 (N_12182,N_11818,N_11768);
nand U12183 (N_12183,N_11443,N_11286);
nor U12184 (N_12184,N_11717,N_11183);
nand U12185 (N_12185,N_11721,N_11658);
nand U12186 (N_12186,N_11204,N_11154);
and U12187 (N_12187,N_11990,N_11527);
and U12188 (N_12188,N_11804,N_11792);
nand U12189 (N_12189,N_11813,N_11623);
or U12190 (N_12190,N_11805,N_11565);
nor U12191 (N_12191,N_11608,N_11766);
nor U12192 (N_12192,N_11221,N_11017);
xnor U12193 (N_12193,N_11091,N_11141);
or U12194 (N_12194,N_11720,N_11457);
or U12195 (N_12195,N_11654,N_11854);
or U12196 (N_12196,N_11138,N_11245);
and U12197 (N_12197,N_11218,N_11027);
nand U12198 (N_12198,N_11330,N_11904);
nand U12199 (N_12199,N_11576,N_11460);
nor U12200 (N_12200,N_11213,N_11403);
nor U12201 (N_12201,N_11268,N_11983);
nor U12202 (N_12202,N_11022,N_11826);
and U12203 (N_12203,N_11182,N_11252);
nor U12204 (N_12204,N_11868,N_11404);
nor U12205 (N_12205,N_11246,N_11643);
or U12206 (N_12206,N_11335,N_11856);
nor U12207 (N_12207,N_11175,N_11811);
and U12208 (N_12208,N_11004,N_11238);
and U12209 (N_12209,N_11559,N_11785);
nand U12210 (N_12210,N_11740,N_11810);
nor U12211 (N_12211,N_11600,N_11188);
nor U12212 (N_12212,N_11332,N_11960);
and U12213 (N_12213,N_11348,N_11872);
nand U12214 (N_12214,N_11346,N_11624);
xor U12215 (N_12215,N_11105,N_11192);
and U12216 (N_12216,N_11162,N_11055);
nor U12217 (N_12217,N_11070,N_11969);
and U12218 (N_12218,N_11926,N_11240);
or U12219 (N_12219,N_11756,N_11358);
nand U12220 (N_12220,N_11605,N_11490);
and U12221 (N_12221,N_11054,N_11320);
nor U12222 (N_12222,N_11886,N_11925);
and U12223 (N_12223,N_11746,N_11439);
and U12224 (N_12224,N_11159,N_11899);
or U12225 (N_12225,N_11541,N_11126);
or U12226 (N_12226,N_11227,N_11048);
nand U12227 (N_12227,N_11340,N_11331);
xnor U12228 (N_12228,N_11303,N_11951);
nand U12229 (N_12229,N_11464,N_11409);
or U12230 (N_12230,N_11113,N_11436);
nor U12231 (N_12231,N_11829,N_11784);
xor U12232 (N_12232,N_11563,N_11525);
nand U12233 (N_12233,N_11917,N_11962);
and U12234 (N_12234,N_11845,N_11482);
xnor U12235 (N_12235,N_11082,N_11402);
or U12236 (N_12236,N_11365,N_11971);
nand U12237 (N_12237,N_11163,N_11692);
nand U12238 (N_12238,N_11269,N_11947);
xnor U12239 (N_12239,N_11954,N_11088);
and U12240 (N_12240,N_11548,N_11277);
nand U12241 (N_12241,N_11220,N_11502);
nor U12242 (N_12242,N_11184,N_11846);
and U12243 (N_12243,N_11857,N_11511);
nand U12244 (N_12244,N_11646,N_11519);
or U12245 (N_12245,N_11861,N_11361);
nand U12246 (N_12246,N_11284,N_11933);
nand U12247 (N_12247,N_11376,N_11233);
xnor U12248 (N_12248,N_11362,N_11690);
and U12249 (N_12249,N_11059,N_11109);
and U12250 (N_12250,N_11069,N_11674);
nor U12251 (N_12251,N_11497,N_11274);
nor U12252 (N_12252,N_11823,N_11211);
nand U12253 (N_12253,N_11812,N_11941);
or U12254 (N_12254,N_11555,N_11285);
nand U12255 (N_12255,N_11531,N_11822);
nor U12256 (N_12256,N_11197,N_11075);
nand U12257 (N_12257,N_11478,N_11972);
nor U12258 (N_12258,N_11506,N_11459);
and U12259 (N_12259,N_11580,N_11535);
nor U12260 (N_12260,N_11420,N_11345);
and U12261 (N_12261,N_11097,N_11880);
nor U12262 (N_12262,N_11915,N_11572);
nor U12263 (N_12263,N_11232,N_11144);
nand U12264 (N_12264,N_11707,N_11405);
nor U12265 (N_12265,N_11830,N_11001);
or U12266 (N_12266,N_11489,N_11125);
nand U12267 (N_12267,N_11189,N_11339);
and U12268 (N_12268,N_11526,N_11976);
xor U12269 (N_12269,N_11588,N_11000);
nor U12270 (N_12270,N_11532,N_11074);
nor U12271 (N_12271,N_11115,N_11831);
and U12272 (N_12272,N_11295,N_11081);
and U12273 (N_12273,N_11417,N_11884);
or U12274 (N_12274,N_11620,N_11751);
nand U12275 (N_12275,N_11799,N_11350);
or U12276 (N_12276,N_11372,N_11064);
or U12277 (N_12277,N_11538,N_11352);
and U12278 (N_12278,N_11461,N_11299);
nor U12279 (N_12279,N_11235,N_11641);
and U12280 (N_12280,N_11275,N_11441);
nor U12281 (N_12281,N_11655,N_11780);
or U12282 (N_12282,N_11415,N_11862);
nand U12283 (N_12283,N_11771,N_11029);
and U12284 (N_12284,N_11518,N_11596);
or U12285 (N_12285,N_11512,N_11515);
nor U12286 (N_12286,N_11584,N_11016);
nand U12287 (N_12287,N_11181,N_11611);
or U12288 (N_12288,N_11206,N_11522);
and U12289 (N_12289,N_11602,N_11504);
or U12290 (N_12290,N_11663,N_11480);
xnor U12291 (N_12291,N_11193,N_11336);
and U12292 (N_12292,N_11656,N_11824);
or U12293 (N_12293,N_11177,N_11852);
nand U12294 (N_12294,N_11051,N_11807);
nor U12295 (N_12295,N_11789,N_11754);
nand U12296 (N_12296,N_11712,N_11934);
and U12297 (N_12297,N_11672,N_11323);
and U12298 (N_12298,N_11597,N_11041);
and U12299 (N_12299,N_11910,N_11217);
nand U12300 (N_12300,N_11781,N_11258);
xor U12301 (N_12301,N_11305,N_11251);
and U12302 (N_12302,N_11334,N_11395);
or U12303 (N_12303,N_11030,N_11414);
or U12304 (N_12304,N_11325,N_11224);
nor U12305 (N_12305,N_11327,N_11891);
and U12306 (N_12306,N_11631,N_11400);
and U12307 (N_12307,N_11953,N_11772);
xnor U12308 (N_12308,N_11619,N_11738);
nand U12309 (N_12309,N_11992,N_11024);
nand U12310 (N_12310,N_11601,N_11150);
or U12311 (N_12311,N_11869,N_11681);
and U12312 (N_12312,N_11484,N_11289);
and U12313 (N_12313,N_11622,N_11134);
nor U12314 (N_12314,N_11449,N_11260);
and U12315 (N_12315,N_11018,N_11394);
xor U12316 (N_12316,N_11540,N_11363);
or U12317 (N_12317,N_11178,N_11662);
nor U12318 (N_12318,N_11343,N_11583);
or U12319 (N_12319,N_11388,N_11108);
or U12320 (N_12320,N_11378,N_11080);
or U12321 (N_12321,N_11200,N_11765);
or U12322 (N_12322,N_11529,N_11577);
nor U12323 (N_12323,N_11825,N_11329);
and U12324 (N_12324,N_11169,N_11726);
nand U12325 (N_12325,N_11158,N_11293);
or U12326 (N_12326,N_11945,N_11288);
nand U12327 (N_12327,N_11581,N_11895);
nand U12328 (N_12328,N_11467,N_11015);
nand U12329 (N_12329,N_11710,N_11387);
and U12330 (N_12330,N_11005,N_11377);
and U12331 (N_12331,N_11313,N_11173);
and U12332 (N_12332,N_11547,N_11114);
and U12333 (N_12333,N_11292,N_11421);
nor U12334 (N_12334,N_11930,N_11615);
and U12335 (N_12335,N_11477,N_11982);
or U12336 (N_12336,N_11835,N_11179);
or U12337 (N_12337,N_11966,N_11207);
nor U12338 (N_12338,N_11287,N_11454);
nor U12339 (N_12339,N_11877,N_11076);
nor U12340 (N_12340,N_11660,N_11123);
or U12341 (N_12341,N_11775,N_11199);
nor U12342 (N_12342,N_11243,N_11734);
and U12343 (N_12343,N_11567,N_11471);
xnor U12344 (N_12344,N_11952,N_11544);
nor U12345 (N_12345,N_11008,N_11375);
or U12346 (N_12346,N_11131,N_11368);
nand U12347 (N_12347,N_11385,N_11429);
and U12348 (N_12348,N_11468,N_11493);
nor U12349 (N_12349,N_11487,N_11568);
xor U12350 (N_12350,N_11393,N_11533);
or U12351 (N_12351,N_11558,N_11294);
or U12352 (N_12352,N_11007,N_11670);
and U12353 (N_12353,N_11942,N_11171);
and U12354 (N_12354,N_11727,N_11047);
nand U12355 (N_12355,N_11337,N_11736);
or U12356 (N_12356,N_11864,N_11090);
nor U12357 (N_12357,N_11264,N_11121);
nor U12358 (N_12358,N_11298,N_11735);
or U12359 (N_12359,N_11595,N_11546);
xnor U12360 (N_12360,N_11072,N_11882);
or U12361 (N_12361,N_11225,N_11874);
nor U12362 (N_12362,N_11116,N_11157);
nor U12363 (N_12363,N_11955,N_11866);
or U12364 (N_12364,N_11440,N_11575);
or U12365 (N_12365,N_11867,N_11383);
xor U12366 (N_12366,N_11087,N_11722);
or U12367 (N_12367,N_11564,N_11270);
and U12368 (N_12368,N_11342,N_11680);
and U12369 (N_12369,N_11815,N_11112);
nand U12370 (N_12370,N_11176,N_11120);
nor U12371 (N_12371,N_11552,N_11333);
nor U12372 (N_12372,N_11020,N_11465);
nand U12373 (N_12373,N_11817,N_11062);
nor U12374 (N_12374,N_11261,N_11156);
nand U12375 (N_12375,N_11963,N_11770);
nor U12376 (N_12376,N_11025,N_11718);
xor U12377 (N_12377,N_11627,N_11111);
and U12378 (N_12378,N_11301,N_11050);
nand U12379 (N_12379,N_11386,N_11776);
and U12380 (N_12380,N_11979,N_11996);
xor U12381 (N_12381,N_11239,N_11127);
or U12382 (N_12382,N_11569,N_11425);
and U12383 (N_12383,N_11314,N_11652);
xor U12384 (N_12384,N_11266,N_11604);
nand U12385 (N_12385,N_11447,N_11579);
nor U12386 (N_12386,N_11562,N_11219);
and U12387 (N_12387,N_11889,N_11549);
xnor U12388 (N_12388,N_11250,N_11035);
nand U12389 (N_12389,N_11132,N_11318);
xnor U12390 (N_12390,N_11486,N_11418);
and U12391 (N_12391,N_11210,N_11590);
xor U12392 (N_12392,N_11056,N_11582);
nor U12393 (N_12393,N_11053,N_11919);
nand U12394 (N_12394,N_11612,N_11257);
nand U12395 (N_12395,N_11508,N_11613);
or U12396 (N_12396,N_11209,N_11271);
nand U12397 (N_12397,N_11625,N_11924);
and U12398 (N_12398,N_11282,N_11180);
nand U12399 (N_12399,N_11248,N_11808);
nand U12400 (N_12400,N_11898,N_11767);
nand U12401 (N_12401,N_11728,N_11262);
nand U12402 (N_12402,N_11312,N_11014);
or U12403 (N_12403,N_11366,N_11446);
and U12404 (N_12404,N_11936,N_11237);
nor U12405 (N_12405,N_11094,N_11379);
or U12406 (N_12406,N_11434,N_11556);
and U12407 (N_12407,N_11650,N_11195);
xor U12408 (N_12408,N_11844,N_11701);
nor U12409 (N_12409,N_11040,N_11661);
nor U12410 (N_12410,N_11991,N_11322);
xor U12411 (N_12411,N_11902,N_11748);
and U12412 (N_12412,N_11927,N_11253);
or U12413 (N_12413,N_11921,N_11800);
and U12414 (N_12414,N_11066,N_11052);
xnor U12415 (N_12415,N_11481,N_11084);
nand U12416 (N_12416,N_11172,N_11424);
xor U12417 (N_12417,N_11272,N_11419);
nand U12418 (N_12418,N_11870,N_11241);
nor U12419 (N_12419,N_11186,N_11774);
nand U12420 (N_12420,N_11975,N_11887);
and U12421 (N_12421,N_11839,N_11278);
or U12422 (N_12422,N_11716,N_11883);
and U12423 (N_12423,N_11242,N_11521);
or U12424 (N_12424,N_11853,N_11999);
and U12425 (N_12425,N_11819,N_11977);
nand U12426 (N_12426,N_11033,N_11124);
xnor U12427 (N_12427,N_11860,N_11509);
nand U12428 (N_12428,N_11247,N_11347);
and U12429 (N_12429,N_11554,N_11520);
and U12430 (N_12430,N_11310,N_11821);
xor U12431 (N_12431,N_11621,N_11684);
nor U12432 (N_12432,N_11389,N_11194);
and U12433 (N_12433,N_11649,N_11061);
nor U12434 (N_12434,N_11307,N_11316);
nor U12435 (N_12435,N_11406,N_11306);
or U12436 (N_12436,N_11871,N_11103);
nand U12437 (N_12437,N_11892,N_11691);
nand U12438 (N_12438,N_11485,N_11068);
nand U12439 (N_12439,N_11922,N_11291);
nor U12440 (N_12440,N_11550,N_11371);
nor U12441 (N_12441,N_11410,N_11283);
xnor U12442 (N_12442,N_11151,N_11297);
nor U12443 (N_12443,N_11215,N_11551);
nor U12444 (N_12444,N_11451,N_11032);
nor U12445 (N_12445,N_11667,N_11801);
nand U12446 (N_12446,N_11876,N_11430);
xnor U12447 (N_12447,N_11645,N_11901);
or U12448 (N_12448,N_11878,N_11149);
and U12449 (N_12449,N_11513,N_11469);
or U12450 (N_12450,N_11827,N_11946);
and U12451 (N_12451,N_11530,N_11724);
nor U12452 (N_12452,N_11426,N_11937);
or U12453 (N_12453,N_11637,N_11834);
nand U12454 (N_12454,N_11028,N_11448);
nand U12455 (N_12455,N_11647,N_11437);
or U12456 (N_12456,N_11009,N_11036);
nand U12457 (N_12457,N_11003,N_11100);
nor U12458 (N_12458,N_11488,N_11155);
or U12459 (N_12459,N_11244,N_11412);
xnor U12460 (N_12460,N_11961,N_11762);
and U12461 (N_12461,N_11673,N_11994);
or U12462 (N_12462,N_11049,N_11302);
xor U12463 (N_12463,N_11543,N_11843);
nor U12464 (N_12464,N_11373,N_11719);
nor U12465 (N_12465,N_11973,N_11442);
nor U12466 (N_12466,N_11453,N_11397);
nor U12467 (N_12467,N_11491,N_11010);
nor U12468 (N_12468,N_11828,N_11893);
nor U12469 (N_12469,N_11908,N_11832);
nor U12470 (N_12470,N_11668,N_11694);
nor U12471 (N_12471,N_11795,N_11693);
or U12472 (N_12472,N_11254,N_11256);
nand U12473 (N_12473,N_11026,N_11259);
nor U12474 (N_12474,N_11705,N_11848);
nand U12475 (N_12475,N_11505,N_11137);
or U12476 (N_12476,N_11814,N_11359);
xor U12477 (N_12477,N_11473,N_11629);
nand U12478 (N_12478,N_11399,N_11231);
xnor U12479 (N_12479,N_11809,N_11170);
or U12480 (N_12480,N_11682,N_11462);
and U12481 (N_12481,N_11777,N_11603);
nand U12482 (N_12482,N_11408,N_11837);
and U12483 (N_12483,N_11202,N_11095);
or U12484 (N_12484,N_11390,N_11093);
nor U12485 (N_12485,N_11455,N_11002);
and U12486 (N_12486,N_11797,N_11539);
xnor U12487 (N_12487,N_11130,N_11790);
and U12488 (N_12488,N_11671,N_11089);
nor U12489 (N_12489,N_11985,N_11598);
and U12490 (N_12490,N_11711,N_11354);
nor U12491 (N_12491,N_11122,N_11573);
nand U12492 (N_12492,N_11498,N_11205);
nand U12493 (N_12493,N_11308,N_11609);
xor U12494 (N_12494,N_11073,N_11931);
or U12495 (N_12495,N_11411,N_11741);
and U12496 (N_12496,N_11614,N_11747);
or U12497 (N_12497,N_11369,N_11474);
xor U12498 (N_12498,N_11147,N_11528);
xnor U12499 (N_12499,N_11635,N_11873);
or U12500 (N_12500,N_11328,N_11432);
xor U12501 (N_12501,N_11022,N_11166);
and U12502 (N_12502,N_11436,N_11545);
nor U12503 (N_12503,N_11765,N_11370);
nand U12504 (N_12504,N_11973,N_11928);
or U12505 (N_12505,N_11169,N_11897);
and U12506 (N_12506,N_11661,N_11976);
nand U12507 (N_12507,N_11454,N_11486);
and U12508 (N_12508,N_11725,N_11496);
and U12509 (N_12509,N_11490,N_11055);
nor U12510 (N_12510,N_11443,N_11717);
or U12511 (N_12511,N_11446,N_11991);
and U12512 (N_12512,N_11838,N_11506);
xor U12513 (N_12513,N_11716,N_11176);
or U12514 (N_12514,N_11088,N_11390);
nand U12515 (N_12515,N_11862,N_11866);
nand U12516 (N_12516,N_11508,N_11964);
xor U12517 (N_12517,N_11126,N_11625);
nor U12518 (N_12518,N_11068,N_11512);
and U12519 (N_12519,N_11491,N_11780);
nor U12520 (N_12520,N_11968,N_11367);
and U12521 (N_12521,N_11921,N_11670);
nor U12522 (N_12522,N_11263,N_11068);
nand U12523 (N_12523,N_11508,N_11621);
nand U12524 (N_12524,N_11212,N_11839);
and U12525 (N_12525,N_11405,N_11480);
nor U12526 (N_12526,N_11074,N_11681);
or U12527 (N_12527,N_11400,N_11467);
and U12528 (N_12528,N_11200,N_11564);
nand U12529 (N_12529,N_11767,N_11279);
or U12530 (N_12530,N_11180,N_11709);
and U12531 (N_12531,N_11467,N_11391);
xor U12532 (N_12532,N_11209,N_11453);
nor U12533 (N_12533,N_11800,N_11841);
nor U12534 (N_12534,N_11103,N_11235);
nand U12535 (N_12535,N_11586,N_11743);
nor U12536 (N_12536,N_11261,N_11160);
or U12537 (N_12537,N_11571,N_11780);
nand U12538 (N_12538,N_11205,N_11837);
and U12539 (N_12539,N_11992,N_11343);
and U12540 (N_12540,N_11909,N_11262);
nand U12541 (N_12541,N_11722,N_11014);
xnor U12542 (N_12542,N_11199,N_11933);
nor U12543 (N_12543,N_11091,N_11062);
or U12544 (N_12544,N_11856,N_11799);
or U12545 (N_12545,N_11332,N_11304);
or U12546 (N_12546,N_11616,N_11413);
nand U12547 (N_12547,N_11864,N_11619);
and U12548 (N_12548,N_11445,N_11497);
nand U12549 (N_12549,N_11359,N_11336);
and U12550 (N_12550,N_11517,N_11884);
xnor U12551 (N_12551,N_11311,N_11727);
nor U12552 (N_12552,N_11721,N_11668);
nor U12553 (N_12553,N_11698,N_11426);
and U12554 (N_12554,N_11152,N_11928);
nor U12555 (N_12555,N_11099,N_11041);
nand U12556 (N_12556,N_11624,N_11229);
nor U12557 (N_12557,N_11651,N_11677);
nor U12558 (N_12558,N_11621,N_11712);
and U12559 (N_12559,N_11109,N_11214);
nand U12560 (N_12560,N_11065,N_11963);
nor U12561 (N_12561,N_11762,N_11717);
nand U12562 (N_12562,N_11391,N_11776);
nor U12563 (N_12563,N_11513,N_11534);
nor U12564 (N_12564,N_11228,N_11706);
or U12565 (N_12565,N_11532,N_11298);
nand U12566 (N_12566,N_11148,N_11457);
nand U12567 (N_12567,N_11651,N_11065);
and U12568 (N_12568,N_11484,N_11291);
and U12569 (N_12569,N_11689,N_11773);
xor U12570 (N_12570,N_11964,N_11918);
xor U12571 (N_12571,N_11257,N_11034);
and U12572 (N_12572,N_11671,N_11839);
and U12573 (N_12573,N_11922,N_11404);
nor U12574 (N_12574,N_11806,N_11322);
nor U12575 (N_12575,N_11008,N_11701);
and U12576 (N_12576,N_11455,N_11464);
nand U12577 (N_12577,N_11714,N_11345);
or U12578 (N_12578,N_11083,N_11875);
or U12579 (N_12579,N_11686,N_11728);
nand U12580 (N_12580,N_11196,N_11467);
or U12581 (N_12581,N_11875,N_11689);
and U12582 (N_12582,N_11330,N_11924);
or U12583 (N_12583,N_11981,N_11996);
or U12584 (N_12584,N_11387,N_11224);
nand U12585 (N_12585,N_11007,N_11360);
and U12586 (N_12586,N_11183,N_11874);
xor U12587 (N_12587,N_11144,N_11989);
nor U12588 (N_12588,N_11948,N_11593);
nor U12589 (N_12589,N_11987,N_11937);
nand U12590 (N_12590,N_11194,N_11957);
nor U12591 (N_12591,N_11953,N_11179);
and U12592 (N_12592,N_11592,N_11298);
nand U12593 (N_12593,N_11132,N_11171);
nand U12594 (N_12594,N_11754,N_11363);
or U12595 (N_12595,N_11520,N_11038);
xor U12596 (N_12596,N_11455,N_11063);
nand U12597 (N_12597,N_11197,N_11474);
nor U12598 (N_12598,N_11807,N_11213);
nor U12599 (N_12599,N_11386,N_11251);
or U12600 (N_12600,N_11395,N_11336);
nand U12601 (N_12601,N_11525,N_11546);
xor U12602 (N_12602,N_11178,N_11276);
and U12603 (N_12603,N_11898,N_11780);
xnor U12604 (N_12604,N_11850,N_11514);
and U12605 (N_12605,N_11358,N_11474);
and U12606 (N_12606,N_11495,N_11427);
nor U12607 (N_12607,N_11419,N_11102);
xor U12608 (N_12608,N_11457,N_11192);
nor U12609 (N_12609,N_11256,N_11414);
or U12610 (N_12610,N_11781,N_11283);
or U12611 (N_12611,N_11862,N_11815);
and U12612 (N_12612,N_11342,N_11869);
nor U12613 (N_12613,N_11657,N_11813);
and U12614 (N_12614,N_11837,N_11276);
and U12615 (N_12615,N_11461,N_11667);
nor U12616 (N_12616,N_11786,N_11136);
nand U12617 (N_12617,N_11471,N_11670);
or U12618 (N_12618,N_11956,N_11500);
or U12619 (N_12619,N_11163,N_11966);
nand U12620 (N_12620,N_11977,N_11774);
nor U12621 (N_12621,N_11050,N_11078);
and U12622 (N_12622,N_11645,N_11580);
nor U12623 (N_12623,N_11194,N_11229);
or U12624 (N_12624,N_11974,N_11006);
nand U12625 (N_12625,N_11731,N_11681);
nand U12626 (N_12626,N_11157,N_11742);
and U12627 (N_12627,N_11815,N_11901);
nor U12628 (N_12628,N_11588,N_11745);
or U12629 (N_12629,N_11125,N_11036);
and U12630 (N_12630,N_11077,N_11017);
nor U12631 (N_12631,N_11398,N_11282);
nand U12632 (N_12632,N_11129,N_11125);
and U12633 (N_12633,N_11336,N_11053);
nor U12634 (N_12634,N_11568,N_11596);
and U12635 (N_12635,N_11654,N_11448);
and U12636 (N_12636,N_11746,N_11938);
xor U12637 (N_12637,N_11859,N_11740);
or U12638 (N_12638,N_11895,N_11430);
and U12639 (N_12639,N_11337,N_11687);
and U12640 (N_12640,N_11171,N_11621);
and U12641 (N_12641,N_11354,N_11034);
and U12642 (N_12642,N_11430,N_11281);
or U12643 (N_12643,N_11505,N_11924);
xnor U12644 (N_12644,N_11358,N_11179);
xor U12645 (N_12645,N_11945,N_11368);
nand U12646 (N_12646,N_11290,N_11050);
nand U12647 (N_12647,N_11577,N_11616);
xor U12648 (N_12648,N_11215,N_11155);
and U12649 (N_12649,N_11124,N_11561);
nand U12650 (N_12650,N_11218,N_11535);
and U12651 (N_12651,N_11278,N_11844);
nand U12652 (N_12652,N_11349,N_11551);
or U12653 (N_12653,N_11389,N_11000);
or U12654 (N_12654,N_11856,N_11939);
nand U12655 (N_12655,N_11042,N_11461);
or U12656 (N_12656,N_11486,N_11737);
and U12657 (N_12657,N_11869,N_11742);
nor U12658 (N_12658,N_11107,N_11975);
and U12659 (N_12659,N_11098,N_11745);
or U12660 (N_12660,N_11404,N_11394);
xnor U12661 (N_12661,N_11855,N_11973);
or U12662 (N_12662,N_11092,N_11790);
nand U12663 (N_12663,N_11971,N_11405);
and U12664 (N_12664,N_11596,N_11769);
nand U12665 (N_12665,N_11645,N_11158);
nor U12666 (N_12666,N_11336,N_11943);
nand U12667 (N_12667,N_11740,N_11785);
nand U12668 (N_12668,N_11557,N_11652);
nor U12669 (N_12669,N_11243,N_11736);
nand U12670 (N_12670,N_11909,N_11445);
or U12671 (N_12671,N_11109,N_11647);
and U12672 (N_12672,N_11579,N_11914);
or U12673 (N_12673,N_11977,N_11658);
nor U12674 (N_12674,N_11731,N_11615);
nand U12675 (N_12675,N_11048,N_11443);
or U12676 (N_12676,N_11951,N_11341);
nor U12677 (N_12677,N_11641,N_11229);
nor U12678 (N_12678,N_11793,N_11395);
nand U12679 (N_12679,N_11096,N_11968);
or U12680 (N_12680,N_11769,N_11038);
nor U12681 (N_12681,N_11534,N_11697);
nor U12682 (N_12682,N_11761,N_11002);
nand U12683 (N_12683,N_11513,N_11141);
nor U12684 (N_12684,N_11532,N_11104);
or U12685 (N_12685,N_11922,N_11672);
nand U12686 (N_12686,N_11941,N_11612);
or U12687 (N_12687,N_11554,N_11738);
nand U12688 (N_12688,N_11643,N_11269);
and U12689 (N_12689,N_11406,N_11832);
and U12690 (N_12690,N_11432,N_11533);
and U12691 (N_12691,N_11412,N_11712);
nor U12692 (N_12692,N_11735,N_11812);
nor U12693 (N_12693,N_11118,N_11712);
nor U12694 (N_12694,N_11898,N_11069);
nand U12695 (N_12695,N_11523,N_11842);
and U12696 (N_12696,N_11087,N_11434);
nor U12697 (N_12697,N_11915,N_11475);
nand U12698 (N_12698,N_11341,N_11744);
and U12699 (N_12699,N_11433,N_11929);
and U12700 (N_12700,N_11245,N_11284);
and U12701 (N_12701,N_11725,N_11569);
nand U12702 (N_12702,N_11416,N_11985);
nand U12703 (N_12703,N_11877,N_11595);
xnor U12704 (N_12704,N_11861,N_11603);
and U12705 (N_12705,N_11716,N_11038);
nand U12706 (N_12706,N_11188,N_11102);
or U12707 (N_12707,N_11370,N_11524);
nor U12708 (N_12708,N_11180,N_11465);
nand U12709 (N_12709,N_11581,N_11619);
nor U12710 (N_12710,N_11794,N_11961);
and U12711 (N_12711,N_11298,N_11438);
nor U12712 (N_12712,N_11552,N_11555);
nor U12713 (N_12713,N_11514,N_11309);
and U12714 (N_12714,N_11296,N_11672);
or U12715 (N_12715,N_11521,N_11060);
or U12716 (N_12716,N_11169,N_11758);
nand U12717 (N_12717,N_11416,N_11885);
and U12718 (N_12718,N_11258,N_11157);
or U12719 (N_12719,N_11193,N_11921);
xnor U12720 (N_12720,N_11901,N_11464);
nor U12721 (N_12721,N_11891,N_11237);
nor U12722 (N_12722,N_11060,N_11971);
nand U12723 (N_12723,N_11703,N_11209);
nor U12724 (N_12724,N_11080,N_11257);
or U12725 (N_12725,N_11665,N_11433);
or U12726 (N_12726,N_11780,N_11619);
nand U12727 (N_12727,N_11393,N_11439);
nand U12728 (N_12728,N_11565,N_11680);
nand U12729 (N_12729,N_11487,N_11114);
nor U12730 (N_12730,N_11598,N_11852);
nand U12731 (N_12731,N_11248,N_11757);
nor U12732 (N_12732,N_11573,N_11915);
nand U12733 (N_12733,N_11401,N_11073);
nand U12734 (N_12734,N_11279,N_11993);
or U12735 (N_12735,N_11556,N_11091);
or U12736 (N_12736,N_11738,N_11140);
nand U12737 (N_12737,N_11840,N_11867);
xor U12738 (N_12738,N_11411,N_11719);
nand U12739 (N_12739,N_11611,N_11103);
or U12740 (N_12740,N_11464,N_11952);
xor U12741 (N_12741,N_11359,N_11160);
and U12742 (N_12742,N_11843,N_11777);
or U12743 (N_12743,N_11338,N_11031);
xor U12744 (N_12744,N_11917,N_11696);
nand U12745 (N_12745,N_11714,N_11579);
nand U12746 (N_12746,N_11898,N_11282);
and U12747 (N_12747,N_11217,N_11352);
nand U12748 (N_12748,N_11217,N_11825);
nor U12749 (N_12749,N_11031,N_11766);
and U12750 (N_12750,N_11882,N_11421);
or U12751 (N_12751,N_11549,N_11105);
nand U12752 (N_12752,N_11130,N_11642);
and U12753 (N_12753,N_11073,N_11995);
nor U12754 (N_12754,N_11261,N_11590);
and U12755 (N_12755,N_11948,N_11136);
or U12756 (N_12756,N_11326,N_11290);
nor U12757 (N_12757,N_11885,N_11791);
and U12758 (N_12758,N_11552,N_11348);
nor U12759 (N_12759,N_11709,N_11812);
or U12760 (N_12760,N_11606,N_11691);
xnor U12761 (N_12761,N_11244,N_11460);
xor U12762 (N_12762,N_11989,N_11011);
xor U12763 (N_12763,N_11828,N_11722);
nand U12764 (N_12764,N_11261,N_11492);
and U12765 (N_12765,N_11742,N_11437);
and U12766 (N_12766,N_11096,N_11065);
and U12767 (N_12767,N_11406,N_11642);
nor U12768 (N_12768,N_11861,N_11310);
nor U12769 (N_12769,N_11240,N_11401);
nor U12770 (N_12770,N_11721,N_11526);
or U12771 (N_12771,N_11527,N_11209);
nor U12772 (N_12772,N_11616,N_11661);
nor U12773 (N_12773,N_11314,N_11690);
nand U12774 (N_12774,N_11554,N_11591);
nor U12775 (N_12775,N_11679,N_11820);
xnor U12776 (N_12776,N_11557,N_11350);
nand U12777 (N_12777,N_11515,N_11144);
nand U12778 (N_12778,N_11020,N_11564);
and U12779 (N_12779,N_11197,N_11780);
and U12780 (N_12780,N_11185,N_11255);
xor U12781 (N_12781,N_11521,N_11078);
or U12782 (N_12782,N_11368,N_11482);
nor U12783 (N_12783,N_11673,N_11524);
or U12784 (N_12784,N_11500,N_11232);
and U12785 (N_12785,N_11901,N_11484);
or U12786 (N_12786,N_11373,N_11063);
nand U12787 (N_12787,N_11008,N_11725);
nor U12788 (N_12788,N_11406,N_11078);
nand U12789 (N_12789,N_11796,N_11793);
xnor U12790 (N_12790,N_11738,N_11055);
or U12791 (N_12791,N_11656,N_11937);
or U12792 (N_12792,N_11751,N_11984);
nand U12793 (N_12793,N_11611,N_11579);
nor U12794 (N_12794,N_11892,N_11718);
or U12795 (N_12795,N_11372,N_11425);
and U12796 (N_12796,N_11614,N_11511);
and U12797 (N_12797,N_11199,N_11124);
and U12798 (N_12798,N_11744,N_11322);
or U12799 (N_12799,N_11649,N_11431);
nand U12800 (N_12800,N_11292,N_11321);
nor U12801 (N_12801,N_11683,N_11785);
nor U12802 (N_12802,N_11111,N_11701);
and U12803 (N_12803,N_11330,N_11376);
and U12804 (N_12804,N_11918,N_11861);
and U12805 (N_12805,N_11189,N_11067);
nand U12806 (N_12806,N_11807,N_11619);
nand U12807 (N_12807,N_11921,N_11314);
nor U12808 (N_12808,N_11947,N_11827);
and U12809 (N_12809,N_11425,N_11206);
nand U12810 (N_12810,N_11004,N_11378);
nand U12811 (N_12811,N_11120,N_11575);
or U12812 (N_12812,N_11197,N_11657);
xor U12813 (N_12813,N_11430,N_11072);
nand U12814 (N_12814,N_11670,N_11510);
or U12815 (N_12815,N_11994,N_11040);
nor U12816 (N_12816,N_11744,N_11791);
xor U12817 (N_12817,N_11177,N_11897);
nand U12818 (N_12818,N_11577,N_11796);
nor U12819 (N_12819,N_11145,N_11314);
and U12820 (N_12820,N_11725,N_11301);
nor U12821 (N_12821,N_11630,N_11161);
and U12822 (N_12822,N_11106,N_11509);
nor U12823 (N_12823,N_11825,N_11787);
or U12824 (N_12824,N_11106,N_11645);
nor U12825 (N_12825,N_11311,N_11107);
xnor U12826 (N_12826,N_11623,N_11298);
or U12827 (N_12827,N_11773,N_11190);
nand U12828 (N_12828,N_11430,N_11752);
or U12829 (N_12829,N_11579,N_11565);
nand U12830 (N_12830,N_11393,N_11099);
xor U12831 (N_12831,N_11662,N_11981);
xor U12832 (N_12832,N_11490,N_11337);
nor U12833 (N_12833,N_11245,N_11730);
xor U12834 (N_12834,N_11193,N_11792);
or U12835 (N_12835,N_11619,N_11134);
nand U12836 (N_12836,N_11902,N_11736);
nor U12837 (N_12837,N_11530,N_11467);
or U12838 (N_12838,N_11633,N_11300);
xnor U12839 (N_12839,N_11330,N_11772);
nand U12840 (N_12840,N_11405,N_11177);
nor U12841 (N_12841,N_11592,N_11561);
nand U12842 (N_12842,N_11782,N_11182);
nor U12843 (N_12843,N_11984,N_11076);
nor U12844 (N_12844,N_11623,N_11340);
and U12845 (N_12845,N_11781,N_11065);
nor U12846 (N_12846,N_11969,N_11501);
xnor U12847 (N_12847,N_11467,N_11117);
and U12848 (N_12848,N_11637,N_11822);
nor U12849 (N_12849,N_11885,N_11902);
nand U12850 (N_12850,N_11412,N_11037);
or U12851 (N_12851,N_11895,N_11125);
nand U12852 (N_12852,N_11166,N_11002);
nor U12853 (N_12853,N_11504,N_11120);
and U12854 (N_12854,N_11669,N_11606);
nor U12855 (N_12855,N_11027,N_11607);
xnor U12856 (N_12856,N_11233,N_11513);
nand U12857 (N_12857,N_11366,N_11404);
and U12858 (N_12858,N_11232,N_11123);
xnor U12859 (N_12859,N_11212,N_11677);
nor U12860 (N_12860,N_11050,N_11592);
xor U12861 (N_12861,N_11740,N_11776);
nor U12862 (N_12862,N_11562,N_11660);
xnor U12863 (N_12863,N_11156,N_11972);
xnor U12864 (N_12864,N_11660,N_11623);
xnor U12865 (N_12865,N_11199,N_11383);
nand U12866 (N_12866,N_11856,N_11398);
and U12867 (N_12867,N_11017,N_11693);
nor U12868 (N_12868,N_11284,N_11319);
and U12869 (N_12869,N_11153,N_11726);
or U12870 (N_12870,N_11660,N_11200);
or U12871 (N_12871,N_11484,N_11153);
and U12872 (N_12872,N_11723,N_11849);
nor U12873 (N_12873,N_11819,N_11473);
and U12874 (N_12874,N_11277,N_11375);
nand U12875 (N_12875,N_11743,N_11665);
and U12876 (N_12876,N_11541,N_11527);
xor U12877 (N_12877,N_11845,N_11189);
and U12878 (N_12878,N_11857,N_11293);
and U12879 (N_12879,N_11707,N_11135);
nand U12880 (N_12880,N_11149,N_11786);
or U12881 (N_12881,N_11970,N_11119);
nor U12882 (N_12882,N_11100,N_11308);
nand U12883 (N_12883,N_11500,N_11420);
xnor U12884 (N_12884,N_11967,N_11751);
nor U12885 (N_12885,N_11706,N_11171);
and U12886 (N_12886,N_11278,N_11773);
or U12887 (N_12887,N_11262,N_11379);
nand U12888 (N_12888,N_11869,N_11985);
nor U12889 (N_12889,N_11779,N_11867);
nor U12890 (N_12890,N_11821,N_11852);
or U12891 (N_12891,N_11776,N_11384);
and U12892 (N_12892,N_11959,N_11935);
or U12893 (N_12893,N_11184,N_11384);
or U12894 (N_12894,N_11024,N_11440);
nor U12895 (N_12895,N_11429,N_11986);
or U12896 (N_12896,N_11203,N_11049);
nor U12897 (N_12897,N_11535,N_11304);
nand U12898 (N_12898,N_11186,N_11503);
xor U12899 (N_12899,N_11802,N_11252);
nand U12900 (N_12900,N_11729,N_11625);
or U12901 (N_12901,N_11852,N_11288);
nor U12902 (N_12902,N_11059,N_11100);
nor U12903 (N_12903,N_11830,N_11715);
nand U12904 (N_12904,N_11336,N_11674);
nor U12905 (N_12905,N_11534,N_11337);
and U12906 (N_12906,N_11574,N_11314);
nand U12907 (N_12907,N_11425,N_11843);
nor U12908 (N_12908,N_11846,N_11296);
nor U12909 (N_12909,N_11185,N_11863);
and U12910 (N_12910,N_11351,N_11223);
xnor U12911 (N_12911,N_11003,N_11539);
or U12912 (N_12912,N_11854,N_11999);
nand U12913 (N_12913,N_11482,N_11013);
nor U12914 (N_12914,N_11410,N_11704);
nor U12915 (N_12915,N_11528,N_11234);
or U12916 (N_12916,N_11812,N_11518);
nand U12917 (N_12917,N_11024,N_11035);
and U12918 (N_12918,N_11296,N_11824);
nand U12919 (N_12919,N_11557,N_11254);
nor U12920 (N_12920,N_11448,N_11173);
or U12921 (N_12921,N_11142,N_11648);
nor U12922 (N_12922,N_11634,N_11119);
nand U12923 (N_12923,N_11249,N_11118);
or U12924 (N_12924,N_11011,N_11288);
nand U12925 (N_12925,N_11838,N_11981);
nor U12926 (N_12926,N_11122,N_11548);
nor U12927 (N_12927,N_11858,N_11183);
or U12928 (N_12928,N_11199,N_11558);
and U12929 (N_12929,N_11392,N_11907);
nor U12930 (N_12930,N_11485,N_11182);
nand U12931 (N_12931,N_11252,N_11953);
nand U12932 (N_12932,N_11596,N_11088);
nand U12933 (N_12933,N_11764,N_11671);
nor U12934 (N_12934,N_11010,N_11246);
or U12935 (N_12935,N_11248,N_11582);
or U12936 (N_12936,N_11800,N_11553);
xor U12937 (N_12937,N_11816,N_11840);
nand U12938 (N_12938,N_11102,N_11479);
and U12939 (N_12939,N_11013,N_11336);
or U12940 (N_12940,N_11012,N_11248);
or U12941 (N_12941,N_11708,N_11238);
or U12942 (N_12942,N_11432,N_11825);
or U12943 (N_12943,N_11285,N_11953);
nand U12944 (N_12944,N_11287,N_11055);
xnor U12945 (N_12945,N_11987,N_11944);
nand U12946 (N_12946,N_11475,N_11854);
xor U12947 (N_12947,N_11622,N_11938);
nor U12948 (N_12948,N_11006,N_11900);
xor U12949 (N_12949,N_11030,N_11840);
nor U12950 (N_12950,N_11376,N_11268);
nand U12951 (N_12951,N_11867,N_11196);
and U12952 (N_12952,N_11734,N_11101);
xnor U12953 (N_12953,N_11535,N_11233);
or U12954 (N_12954,N_11443,N_11588);
and U12955 (N_12955,N_11746,N_11971);
nand U12956 (N_12956,N_11206,N_11000);
and U12957 (N_12957,N_11986,N_11825);
nand U12958 (N_12958,N_11677,N_11295);
nand U12959 (N_12959,N_11377,N_11594);
nor U12960 (N_12960,N_11094,N_11906);
or U12961 (N_12961,N_11347,N_11586);
nor U12962 (N_12962,N_11424,N_11597);
or U12963 (N_12963,N_11879,N_11257);
nand U12964 (N_12964,N_11232,N_11825);
and U12965 (N_12965,N_11612,N_11697);
and U12966 (N_12966,N_11205,N_11576);
nand U12967 (N_12967,N_11837,N_11285);
nor U12968 (N_12968,N_11036,N_11568);
nor U12969 (N_12969,N_11855,N_11444);
nand U12970 (N_12970,N_11325,N_11721);
nand U12971 (N_12971,N_11772,N_11970);
and U12972 (N_12972,N_11251,N_11215);
and U12973 (N_12973,N_11442,N_11287);
nand U12974 (N_12974,N_11578,N_11067);
nor U12975 (N_12975,N_11487,N_11387);
nand U12976 (N_12976,N_11331,N_11079);
nor U12977 (N_12977,N_11696,N_11262);
or U12978 (N_12978,N_11159,N_11452);
xor U12979 (N_12979,N_11790,N_11996);
xnor U12980 (N_12980,N_11937,N_11497);
or U12981 (N_12981,N_11529,N_11475);
xor U12982 (N_12982,N_11059,N_11377);
and U12983 (N_12983,N_11628,N_11928);
or U12984 (N_12984,N_11831,N_11246);
nor U12985 (N_12985,N_11548,N_11533);
or U12986 (N_12986,N_11385,N_11492);
nor U12987 (N_12987,N_11303,N_11185);
and U12988 (N_12988,N_11758,N_11088);
or U12989 (N_12989,N_11965,N_11747);
nor U12990 (N_12990,N_11520,N_11477);
or U12991 (N_12991,N_11861,N_11175);
and U12992 (N_12992,N_11014,N_11345);
nor U12993 (N_12993,N_11822,N_11426);
and U12994 (N_12994,N_11614,N_11510);
or U12995 (N_12995,N_11954,N_11992);
nor U12996 (N_12996,N_11920,N_11047);
or U12997 (N_12997,N_11787,N_11589);
or U12998 (N_12998,N_11831,N_11451);
xnor U12999 (N_12999,N_11670,N_11831);
nor U13000 (N_13000,N_12569,N_12775);
nor U13001 (N_13001,N_12605,N_12714);
nor U13002 (N_13002,N_12794,N_12607);
nand U13003 (N_13003,N_12183,N_12863);
or U13004 (N_13004,N_12987,N_12222);
and U13005 (N_13005,N_12464,N_12325);
nand U13006 (N_13006,N_12049,N_12213);
or U13007 (N_13007,N_12483,N_12187);
nand U13008 (N_13008,N_12473,N_12395);
and U13009 (N_13009,N_12503,N_12564);
nor U13010 (N_13010,N_12414,N_12783);
xor U13011 (N_13011,N_12955,N_12740);
nand U13012 (N_13012,N_12695,N_12170);
and U13013 (N_13013,N_12590,N_12001);
or U13014 (N_13014,N_12883,N_12957);
and U13015 (N_13015,N_12120,N_12494);
or U13016 (N_13016,N_12710,N_12484);
nor U13017 (N_13017,N_12412,N_12941);
xnor U13018 (N_13018,N_12108,N_12920);
and U13019 (N_13019,N_12531,N_12450);
nand U13020 (N_13020,N_12602,N_12432);
and U13021 (N_13021,N_12877,N_12057);
nand U13022 (N_13022,N_12834,N_12547);
nor U13023 (N_13023,N_12096,N_12565);
or U13024 (N_13024,N_12596,N_12479);
or U13025 (N_13025,N_12995,N_12211);
and U13026 (N_13026,N_12106,N_12840);
xnor U13027 (N_13027,N_12302,N_12337);
nor U13028 (N_13028,N_12345,N_12760);
nor U13029 (N_13029,N_12850,N_12028);
nor U13030 (N_13030,N_12053,N_12280);
nand U13031 (N_13031,N_12196,N_12192);
or U13032 (N_13032,N_12027,N_12301);
nand U13033 (N_13033,N_12698,N_12693);
and U13034 (N_13034,N_12146,N_12438);
xor U13035 (N_13035,N_12133,N_12919);
nand U13036 (N_13036,N_12772,N_12523);
nor U13037 (N_13037,N_12066,N_12952);
nor U13038 (N_13038,N_12386,N_12847);
nand U13039 (N_13039,N_12906,N_12765);
or U13040 (N_13040,N_12989,N_12220);
nor U13041 (N_13041,N_12421,N_12499);
and U13042 (N_13042,N_12713,N_12258);
and U13043 (N_13043,N_12029,N_12524);
and U13044 (N_13044,N_12022,N_12176);
and U13045 (N_13045,N_12809,N_12384);
or U13046 (N_13046,N_12927,N_12568);
and U13047 (N_13047,N_12836,N_12904);
nor U13048 (N_13048,N_12428,N_12401);
xor U13049 (N_13049,N_12510,N_12154);
or U13050 (N_13050,N_12604,N_12411);
and U13051 (N_13051,N_12744,N_12977);
or U13052 (N_13052,N_12806,N_12289);
nor U13053 (N_13053,N_12673,N_12459);
or U13054 (N_13054,N_12086,N_12805);
xnor U13055 (N_13055,N_12762,N_12758);
or U13056 (N_13056,N_12644,N_12374);
and U13057 (N_13057,N_12777,N_12145);
xnor U13058 (N_13058,N_12467,N_12773);
and U13059 (N_13059,N_12160,N_12686);
nor U13060 (N_13060,N_12320,N_12574);
xor U13061 (N_13061,N_12480,N_12191);
nor U13062 (N_13062,N_12413,N_12925);
and U13063 (N_13063,N_12930,N_12255);
nand U13064 (N_13064,N_12439,N_12129);
nor U13065 (N_13065,N_12288,N_12718);
nor U13066 (N_13066,N_12333,N_12383);
nand U13067 (N_13067,N_12167,N_12313);
or U13068 (N_13068,N_12814,N_12425);
or U13069 (N_13069,N_12729,N_12983);
nand U13070 (N_13070,N_12733,N_12627);
or U13071 (N_13071,N_12190,N_12339);
xor U13072 (N_13072,N_12463,N_12529);
xnor U13073 (N_13073,N_12406,N_12228);
or U13074 (N_13074,N_12330,N_12680);
nand U13075 (N_13075,N_12918,N_12371);
and U13076 (N_13076,N_12197,N_12731);
xnor U13077 (N_13077,N_12709,N_12298);
nor U13078 (N_13078,N_12079,N_12246);
or U13079 (N_13079,N_12748,N_12984);
nor U13080 (N_13080,N_12243,N_12442);
nor U13081 (N_13081,N_12198,N_12894);
and U13082 (N_13082,N_12005,N_12789);
nand U13083 (N_13083,N_12914,N_12727);
and U13084 (N_13084,N_12575,N_12263);
nor U13085 (N_13085,N_12964,N_12618);
nand U13086 (N_13086,N_12861,N_12282);
and U13087 (N_13087,N_12236,N_12248);
or U13088 (N_13088,N_12553,N_12141);
nor U13089 (N_13089,N_12515,N_12763);
nor U13090 (N_13090,N_12309,N_12471);
nand U13091 (N_13091,N_12430,N_12436);
or U13092 (N_13092,N_12972,N_12804);
or U13093 (N_13093,N_12490,N_12550);
nor U13094 (N_13094,N_12181,N_12291);
nor U13095 (N_13095,N_12101,N_12098);
and U13096 (N_13096,N_12707,N_12849);
nor U13097 (N_13097,N_12712,N_12455);
and U13098 (N_13098,N_12589,N_12319);
and U13099 (N_13099,N_12461,N_12277);
nor U13100 (N_13100,N_12268,N_12629);
nor U13101 (N_13101,N_12084,N_12979);
nor U13102 (N_13102,N_12722,N_12570);
and U13103 (N_13103,N_12265,N_12328);
xor U13104 (N_13104,N_12105,N_12721);
or U13105 (N_13105,N_12481,N_12324);
and U13106 (N_13106,N_12766,N_12224);
nand U13107 (N_13107,N_12612,N_12089);
nor U13108 (N_13108,N_12993,N_12162);
xnor U13109 (N_13109,N_12125,N_12608);
nor U13110 (N_13110,N_12715,N_12951);
nor U13111 (N_13111,N_12953,N_12530);
nand U13112 (N_13112,N_12936,N_12491);
nor U13113 (N_13113,N_12054,N_12254);
nor U13114 (N_13114,N_12915,N_12965);
nand U13115 (N_13115,N_12980,N_12071);
nand U13116 (N_13116,N_12825,N_12905);
or U13117 (N_13117,N_12420,N_12034);
xor U13118 (N_13118,N_12819,N_12387);
and U13119 (N_13119,N_12394,N_12683);
nand U13120 (N_13120,N_12950,N_12601);
or U13121 (N_13121,N_12099,N_12303);
xor U13122 (N_13122,N_12356,N_12283);
xnor U13123 (N_13123,N_12080,N_12373);
nand U13124 (N_13124,N_12020,N_12381);
and U13125 (N_13125,N_12485,N_12469);
nor U13126 (N_13126,N_12179,N_12642);
and U13127 (N_13127,N_12889,N_12043);
nor U13128 (N_13128,N_12663,N_12150);
nor U13129 (N_13129,N_12315,N_12127);
xnor U13130 (N_13130,N_12634,N_12451);
nor U13131 (N_13131,N_12357,N_12078);
xor U13132 (N_13132,N_12175,N_12841);
nor U13133 (N_13133,N_12716,N_12492);
xnor U13134 (N_13134,N_12975,N_12045);
nor U13135 (N_13135,N_12063,N_12546);
nor U13136 (N_13136,N_12507,N_12286);
nand U13137 (N_13137,N_12219,N_12854);
nand U13138 (N_13138,N_12363,N_12512);
nor U13139 (N_13139,N_12747,N_12177);
nand U13140 (N_13140,N_12932,N_12545);
nand U13141 (N_13141,N_12542,N_12314);
and U13142 (N_13142,N_12441,N_12521);
nand U13143 (N_13143,N_12842,N_12871);
nor U13144 (N_13144,N_12824,N_12617);
and U13145 (N_13145,N_12233,N_12583);
nor U13146 (N_13146,N_12046,N_12784);
and U13147 (N_13147,N_12923,N_12435);
nor U13148 (N_13148,N_12959,N_12974);
or U13149 (N_13149,N_12639,N_12408);
and U13150 (N_13150,N_12402,N_12422);
or U13151 (N_13151,N_12807,N_12573);
nor U13152 (N_13152,N_12505,N_12969);
nor U13153 (N_13153,N_12872,N_12667);
or U13154 (N_13154,N_12234,N_12083);
and U13155 (N_13155,N_12278,N_12584);
xnor U13156 (N_13156,N_12603,N_12225);
xnor U13157 (N_13157,N_12161,N_12067);
or U13158 (N_13158,N_12931,N_12717);
nor U13159 (N_13159,N_12555,N_12973);
nor U13160 (N_13160,N_12743,N_12788);
or U13161 (N_13161,N_12831,N_12600);
and U13162 (N_13162,N_12535,N_12229);
nor U13163 (N_13163,N_12012,N_12454);
and U13164 (N_13164,N_12377,N_12645);
or U13165 (N_13165,N_12866,N_12937);
and U13166 (N_13166,N_12870,N_12221);
nor U13167 (N_13167,N_12830,N_12676);
and U13168 (N_13168,N_12929,N_12011);
nand U13169 (N_13169,N_12654,N_12398);
nor U13170 (N_13170,N_12749,N_12403);
nand U13171 (N_13171,N_12694,N_12567);
or U13172 (N_13172,N_12802,N_12540);
nor U13173 (N_13173,N_12554,N_12041);
or U13174 (N_13174,N_12334,N_12679);
nand U13175 (N_13175,N_12657,N_12085);
nand U13176 (N_13176,N_12040,N_12780);
or U13177 (N_13177,N_12934,N_12818);
and U13178 (N_13178,N_12399,N_12251);
xnor U13179 (N_13179,N_12134,N_12201);
xor U13180 (N_13180,N_12292,N_12878);
nor U13181 (N_13181,N_12227,N_12130);
nor U13182 (N_13182,N_12856,N_12658);
nor U13183 (N_13183,N_12536,N_12050);
nand U13184 (N_13184,N_12072,N_12405);
nand U13185 (N_13185,N_12826,N_12967);
nor U13186 (N_13186,N_12660,N_12591);
nor U13187 (N_13187,N_12666,N_12588);
and U13188 (N_13188,N_12578,N_12582);
nor U13189 (N_13189,N_12862,N_12400);
xor U13190 (N_13190,N_12606,N_12256);
or U13191 (N_13191,N_12349,N_12166);
and U13192 (N_13192,N_12882,N_12981);
or U13193 (N_13193,N_12264,N_12552);
nand U13194 (N_13194,N_12791,N_12104);
or U13195 (N_13195,N_12711,N_12558);
nor U13196 (N_13196,N_12344,N_12477);
xor U13197 (N_13197,N_12586,N_12138);
and U13198 (N_13198,N_12643,N_12646);
or U13199 (N_13199,N_12655,N_12396);
or U13200 (N_13200,N_12839,N_12092);
nand U13201 (N_13201,N_12688,N_12311);
nor U13202 (N_13202,N_12128,N_12456);
nor U13203 (N_13203,N_12656,N_12126);
or U13204 (N_13204,N_12297,N_12902);
nor U13205 (N_13205,N_12185,N_12622);
nor U13206 (N_13206,N_12538,N_12235);
and U13207 (N_13207,N_12155,N_12188);
and U13208 (N_13208,N_12390,N_12734);
xnor U13209 (N_13209,N_12482,N_12453);
xnor U13210 (N_13210,N_12633,N_12719);
or U13211 (N_13211,N_12991,N_12241);
nor U13212 (N_13212,N_12094,N_12835);
nor U13213 (N_13213,N_12039,N_12184);
nand U13214 (N_13214,N_12052,N_12911);
xor U13215 (N_13215,N_12010,N_12061);
nand U13216 (N_13216,N_12811,N_12323);
or U13217 (N_13217,N_12764,N_12290);
xor U13218 (N_13218,N_12116,N_12230);
and U13219 (N_13219,N_12924,N_12385);
or U13220 (N_13220,N_12468,N_12091);
nor U13221 (N_13221,N_12843,N_12174);
and U13222 (N_13222,N_12901,N_12443);
nor U13223 (N_13223,N_12368,N_12100);
or U13224 (N_13224,N_12427,N_12738);
nand U13225 (N_13225,N_12090,N_12912);
nand U13226 (N_13226,N_12599,N_12647);
or U13227 (N_13227,N_12369,N_12496);
or U13228 (N_13228,N_12753,N_12501);
nor U13229 (N_13229,N_12495,N_12142);
xor U13230 (N_13230,N_12682,N_12677);
nand U13231 (N_13231,N_12994,N_12609);
or U13232 (N_13232,N_12416,N_12947);
nand U13233 (N_13233,N_12095,N_12284);
nand U13234 (N_13234,N_12940,N_12070);
nand U13235 (N_13235,N_12628,N_12869);
nand U13236 (N_13236,N_12648,N_12409);
or U13237 (N_13237,N_12511,N_12075);
and U13238 (N_13238,N_12522,N_12316);
or U13239 (N_13239,N_12685,N_12779);
nand U13240 (N_13240,N_12561,N_12017);
nor U13241 (N_13241,N_12064,N_12741);
nor U13242 (N_13242,N_12532,N_12702);
or U13243 (N_13243,N_12030,N_12876);
and U13244 (N_13244,N_12305,N_12308);
nor U13245 (N_13245,N_12757,N_12853);
and U13246 (N_13246,N_12509,N_12486);
and U13247 (N_13247,N_12475,N_12004);
nor U13248 (N_13248,N_12110,N_12525);
nor U13249 (N_13249,N_12124,N_12641);
and U13250 (N_13250,N_12121,N_12770);
or U13251 (N_13251,N_12304,N_12347);
nor U13252 (N_13252,N_12418,N_12415);
nor U13253 (N_13253,N_12055,N_12956);
nor U13254 (N_13254,N_12332,N_12670);
and U13255 (N_13255,N_12434,N_12331);
and U13256 (N_13256,N_12855,N_12426);
nor U13257 (N_13257,N_12037,N_12759);
or U13258 (N_13258,N_12990,N_12787);
nand U13259 (N_13259,N_12489,N_12244);
or U13260 (N_13260,N_12771,N_12173);
xor U13261 (N_13261,N_12820,N_12706);
and U13262 (N_13262,N_12335,N_12792);
nand U13263 (N_13263,N_12838,N_12382);
nand U13264 (N_13264,N_12294,N_12502);
nor U13265 (N_13265,N_12899,N_12886);
nand U13266 (N_13266,N_12452,N_12518);
and U13267 (N_13267,N_12527,N_12370);
nor U13268 (N_13268,N_12214,N_12295);
or U13269 (N_13269,N_12595,N_12253);
and U13270 (N_13270,N_12659,N_12218);
xor U13271 (N_13271,N_12031,N_12143);
xor U13272 (N_13272,N_12058,N_12164);
nor U13273 (N_13273,N_12487,N_12392);
xnor U13274 (N_13274,N_12970,N_12497);
or U13275 (N_13275,N_12249,N_12287);
nor U13276 (N_13276,N_12252,N_12921);
nor U13277 (N_13277,N_12204,N_12135);
or U13278 (N_13278,N_12571,N_12354);
nand U13279 (N_13279,N_12514,N_12585);
nand U13280 (N_13280,N_12739,N_12625);
or U13281 (N_13281,N_12708,N_12216);
nor U13282 (N_13282,N_12781,N_12472);
nor U13283 (N_13283,N_12868,N_12267);
nor U13284 (N_13284,N_12864,N_12423);
xnor U13285 (N_13285,N_12665,N_12375);
nand U13286 (N_13286,N_12704,N_12730);
and U13287 (N_13287,N_12465,N_12163);
nand U13288 (N_13288,N_12500,N_12897);
and U13289 (N_13289,N_12598,N_12036);
or U13290 (N_13290,N_12581,N_12774);
and U13291 (N_13291,N_12113,N_12768);
or U13292 (N_13292,N_12960,N_12881);
nor U13293 (N_13293,N_12798,N_12611);
and U13294 (N_13294,N_12449,N_12945);
nand U13295 (N_13295,N_12752,N_12378);
nand U13296 (N_13296,N_12372,N_12242);
nor U13297 (N_13297,N_12391,N_12720);
nand U13298 (N_13298,N_12669,N_12801);
or U13299 (N_13299,N_12207,N_12816);
nor U13300 (N_13300,N_12107,N_12274);
nor U13301 (N_13301,N_12488,N_12351);
nand U13302 (N_13302,N_12821,N_12103);
nand U13303 (N_13303,N_12988,N_12796);
nand U13304 (N_13304,N_12913,N_12732);
or U13305 (N_13305,N_12151,N_12273);
or U13306 (N_13306,N_12786,N_12437);
nor U13307 (N_13307,N_12696,N_12885);
and U13308 (N_13308,N_12875,N_12329);
nand U13309 (N_13309,N_12879,N_12671);
and U13310 (N_13310,N_12093,N_12038);
nor U13311 (N_13311,N_12701,N_12365);
or U13312 (N_13312,N_12968,N_12827);
nand U13313 (N_13313,N_12458,N_12194);
nor U13314 (N_13314,N_12534,N_12350);
and U13315 (N_13315,N_12285,N_12828);
or U13316 (N_13316,N_12587,N_12322);
and U13317 (N_13317,N_12448,N_12852);
xor U13318 (N_13318,N_12003,N_12903);
nor U13319 (N_13319,N_12577,N_12009);
xnor U13320 (N_13320,N_12065,N_12082);
or U13321 (N_13321,N_12736,N_12232);
or U13322 (N_13322,N_12238,N_12355);
nand U13323 (N_13323,N_12942,N_12541);
or U13324 (N_13324,N_12636,N_12884);
or U13325 (N_13325,N_12006,N_12735);
nand U13326 (N_13326,N_12858,N_12069);
and U13327 (N_13327,N_12528,N_12132);
nand U13328 (N_13328,N_12678,N_12812);
and U13329 (N_13329,N_12563,N_12446);
and U13330 (N_13330,N_12767,N_12195);
nand U13331 (N_13331,N_12362,N_12189);
nand U13332 (N_13332,N_12478,N_12014);
or U13333 (N_13333,N_12896,N_12650);
and U13334 (N_13334,N_12353,N_12986);
nor U13335 (N_13335,N_12844,N_12470);
and U13336 (N_13336,N_12306,N_12597);
nand U13337 (N_13337,N_12703,N_12073);
xnor U13338 (N_13338,N_12019,N_12312);
or U13339 (N_13339,N_12444,N_12358);
nand U13340 (N_13340,N_12321,N_12180);
and U13341 (N_13341,N_12149,N_12074);
and U13342 (N_13342,N_12240,N_12815);
and U13343 (N_13343,N_12662,N_12077);
and U13344 (N_13344,N_12388,N_12380);
nor U13345 (N_13345,N_12122,N_12631);
and U13346 (N_13346,N_12266,N_12572);
nand U13347 (N_13347,N_12200,N_12144);
or U13348 (N_13348,N_12136,N_12217);
or U13349 (N_13349,N_12307,N_12907);
and U13350 (N_13350,N_12954,N_12171);
xnor U13351 (N_13351,N_12193,N_12750);
or U13352 (N_13352,N_12649,N_12076);
nand U13353 (N_13353,N_12048,N_12700);
xnor U13354 (N_13354,N_12737,N_12999);
nand U13355 (N_13355,N_12359,N_12250);
or U13356 (N_13356,N_12140,N_12998);
nand U13357 (N_13357,N_12621,N_12326);
or U13358 (N_13358,N_12393,N_12336);
nor U13359 (N_13359,N_12111,N_12664);
nand U13360 (N_13360,N_12205,N_12087);
nor U13361 (N_13361,N_12559,N_12837);
nand U13362 (N_13362,N_12165,N_12462);
and U13363 (N_13363,N_12259,N_12520);
or U13364 (N_13364,N_12551,N_12203);
nand U13365 (N_13365,N_12756,N_12630);
or U13366 (N_13366,N_12948,N_12044);
xor U13367 (N_13367,N_12626,N_12209);
nor U13368 (N_13368,N_12576,N_12042);
nand U13369 (N_13369,N_12687,N_12429);
xor U13370 (N_13370,N_12047,N_12544);
or U13371 (N_13371,N_12724,N_12318);
nand U13372 (N_13372,N_12892,N_12691);
xor U13373 (N_13373,N_12675,N_12966);
or U13374 (N_13374,N_12379,N_12909);
nand U13375 (N_13375,N_12247,N_12342);
or U13376 (N_13376,N_12300,N_12874);
nor U13377 (N_13377,N_12799,N_12109);
nor U13378 (N_13378,N_12615,N_12493);
or U13379 (N_13379,N_12971,N_12156);
or U13380 (N_13380,N_12212,N_12661);
or U13381 (N_13381,N_12389,N_12526);
and U13382 (N_13382,N_12513,N_12033);
nand U13383 (N_13383,N_12845,N_12088);
or U13384 (N_13384,N_12404,N_12653);
and U13385 (N_13385,N_12186,N_12440);
or U13386 (N_13386,N_12352,N_12900);
or U13387 (N_13387,N_12566,N_12958);
nor U13388 (N_13388,N_12982,N_12865);
nand U13389 (N_13389,N_12782,N_12118);
nand U13390 (N_13390,N_12797,N_12257);
nor U13391 (N_13391,N_12823,N_12310);
nor U13392 (N_13392,N_12560,N_12279);
or U13393 (N_13393,N_12725,N_12916);
and U13394 (N_13394,N_12476,N_12832);
nor U13395 (N_13395,N_12623,N_12025);
nand U13396 (N_13396,N_12846,N_12051);
or U13397 (N_13397,N_12466,N_12963);
and U13398 (N_13398,N_12260,N_12857);
xnor U13399 (N_13399,N_12202,N_12018);
xor U13400 (N_13400,N_12119,N_12364);
or U13401 (N_13401,N_12624,N_12343);
nor U13402 (N_13402,N_12115,N_12299);
or U13403 (N_13403,N_12272,N_12593);
xnor U13404 (N_13404,N_12651,N_12504);
or U13405 (N_13405,N_12457,N_12159);
or U13406 (N_13406,N_12056,N_12594);
xnor U13407 (N_13407,N_12873,N_12460);
and U13408 (N_13408,N_12638,N_12275);
and U13409 (N_13409,N_12008,N_12007);
and U13410 (N_13410,N_12237,N_12206);
and U13411 (N_13411,N_12726,N_12158);
and U13412 (N_13412,N_12139,N_12778);
and U13413 (N_13413,N_12992,N_12580);
or U13414 (N_13414,N_12153,N_12813);
nand U13415 (N_13415,N_12859,N_12944);
or U13416 (N_13416,N_12293,N_12997);
and U13417 (N_13417,N_12117,N_12338);
or U13418 (N_13418,N_12208,N_12985);
nand U13419 (N_13419,N_12013,N_12271);
and U13420 (N_13420,N_12182,N_12178);
and U13421 (N_13421,N_12681,N_12269);
and U13422 (N_13422,N_12557,N_12754);
and U13423 (N_13423,N_12032,N_12172);
xnor U13424 (N_13424,N_12539,N_12949);
nand U13425 (N_13425,N_12785,N_12376);
or U13426 (N_13426,N_12592,N_12935);
or U13427 (N_13427,N_12431,N_12867);
or U13428 (N_13428,N_12062,N_12692);
xnor U13429 (N_13429,N_12674,N_12537);
nand U13430 (N_13430,N_12829,N_12723);
nand U13431 (N_13431,N_12668,N_12933);
or U13432 (N_13432,N_12168,N_12517);
and U13433 (N_13433,N_12616,N_12776);
nand U13434 (N_13434,N_12407,N_12728);
or U13435 (N_13435,N_12498,N_12346);
nor U13436 (N_13436,N_12637,N_12516);
nand U13437 (N_13437,N_12943,N_12632);
and U13438 (N_13438,N_12474,N_12548);
nand U13439 (N_13439,N_12231,N_12223);
nand U13440 (N_13440,N_12652,N_12926);
and U13441 (N_13441,N_12397,N_12131);
or U13442 (N_13442,N_12361,N_12833);
or U13443 (N_13443,N_12917,N_12635);
nand U13444 (N_13444,N_12790,N_12035);
or U13445 (N_13445,N_12508,N_12147);
nor U13446 (N_13446,N_12579,N_12543);
xor U13447 (N_13447,N_12137,N_12619);
or U13448 (N_13448,N_12000,N_12097);
nor U13449 (N_13449,N_12939,N_12023);
or U13450 (N_13450,N_12016,N_12152);
nand U13451 (N_13451,N_12002,N_12803);
xor U13452 (N_13452,N_12114,N_12068);
and U13453 (N_13453,N_12976,N_12697);
or U13454 (N_13454,N_12021,N_12751);
nor U13455 (N_13455,N_12961,N_12793);
nand U13456 (N_13456,N_12690,N_12417);
and U13457 (N_13457,N_12360,N_12742);
and U13458 (N_13458,N_12898,N_12059);
or U13459 (N_13459,N_12112,N_12340);
or U13460 (N_13460,N_12506,N_12245);
xor U13461 (N_13461,N_12102,N_12795);
nand U13462 (N_13462,N_12808,N_12199);
nand U13463 (N_13463,N_12239,N_12946);
or U13464 (N_13464,N_12746,N_12519);
or U13465 (N_13465,N_12928,N_12445);
or U13466 (N_13466,N_12769,N_12887);
nor U13467 (N_13467,N_12419,N_12060);
nor U13468 (N_13468,N_12556,N_12367);
and U13469 (N_13469,N_12978,N_12433);
xor U13470 (N_13470,N_12123,N_12015);
xnor U13471 (N_13471,N_12341,N_12893);
xor U13472 (N_13472,N_12908,N_12169);
or U13473 (N_13473,N_12962,N_12755);
nor U13474 (N_13474,N_12689,N_12890);
nand U13475 (N_13475,N_12888,N_12296);
nor U13476 (N_13476,N_12891,N_12822);
xor U13477 (N_13477,N_12613,N_12317);
and U13478 (N_13478,N_12880,N_12424);
and U13479 (N_13479,N_12148,N_12447);
and U13480 (N_13480,N_12410,N_12761);
or U13481 (N_13481,N_12276,N_12705);
nor U13482 (N_13482,N_12215,N_12549);
nor U13483 (N_13483,N_12684,N_12081);
or U13484 (N_13484,N_12281,N_12910);
or U13485 (N_13485,N_12938,N_12327);
xor U13486 (N_13486,N_12562,N_12672);
or U13487 (N_13487,N_12614,N_12810);
nand U13488 (N_13488,N_12800,N_12366);
nor U13489 (N_13489,N_12817,N_12895);
and U13490 (N_13490,N_12024,N_12533);
or U13491 (N_13491,N_12745,N_12026);
and U13492 (N_13492,N_12620,N_12848);
xor U13493 (N_13493,N_12860,N_12851);
or U13494 (N_13494,N_12922,N_12261);
xor U13495 (N_13495,N_12157,N_12640);
and U13496 (N_13496,N_12996,N_12699);
nor U13497 (N_13497,N_12226,N_12210);
and U13498 (N_13498,N_12348,N_12270);
and U13499 (N_13499,N_12262,N_12610);
or U13500 (N_13500,N_12918,N_12806);
and U13501 (N_13501,N_12015,N_12571);
nand U13502 (N_13502,N_12561,N_12866);
nand U13503 (N_13503,N_12335,N_12692);
nand U13504 (N_13504,N_12334,N_12898);
or U13505 (N_13505,N_12096,N_12897);
and U13506 (N_13506,N_12309,N_12255);
nand U13507 (N_13507,N_12845,N_12757);
or U13508 (N_13508,N_12921,N_12974);
or U13509 (N_13509,N_12922,N_12422);
nand U13510 (N_13510,N_12001,N_12363);
xor U13511 (N_13511,N_12496,N_12300);
or U13512 (N_13512,N_12534,N_12687);
nor U13513 (N_13513,N_12423,N_12377);
and U13514 (N_13514,N_12436,N_12359);
or U13515 (N_13515,N_12046,N_12210);
and U13516 (N_13516,N_12673,N_12371);
xnor U13517 (N_13517,N_12441,N_12563);
nor U13518 (N_13518,N_12440,N_12304);
or U13519 (N_13519,N_12070,N_12463);
or U13520 (N_13520,N_12265,N_12800);
nand U13521 (N_13521,N_12470,N_12261);
or U13522 (N_13522,N_12229,N_12435);
and U13523 (N_13523,N_12098,N_12996);
xor U13524 (N_13524,N_12864,N_12458);
and U13525 (N_13525,N_12593,N_12633);
nand U13526 (N_13526,N_12947,N_12041);
nor U13527 (N_13527,N_12015,N_12028);
or U13528 (N_13528,N_12033,N_12629);
nor U13529 (N_13529,N_12044,N_12932);
or U13530 (N_13530,N_12744,N_12420);
nor U13531 (N_13531,N_12046,N_12231);
nor U13532 (N_13532,N_12772,N_12487);
or U13533 (N_13533,N_12145,N_12377);
and U13534 (N_13534,N_12838,N_12858);
nand U13535 (N_13535,N_12546,N_12753);
and U13536 (N_13536,N_12003,N_12275);
and U13537 (N_13537,N_12212,N_12143);
nand U13538 (N_13538,N_12154,N_12451);
nor U13539 (N_13539,N_12285,N_12450);
and U13540 (N_13540,N_12708,N_12337);
xnor U13541 (N_13541,N_12067,N_12950);
nand U13542 (N_13542,N_12690,N_12002);
and U13543 (N_13543,N_12862,N_12308);
nand U13544 (N_13544,N_12229,N_12886);
or U13545 (N_13545,N_12612,N_12794);
and U13546 (N_13546,N_12905,N_12655);
or U13547 (N_13547,N_12500,N_12975);
nand U13548 (N_13548,N_12177,N_12504);
nand U13549 (N_13549,N_12477,N_12001);
and U13550 (N_13550,N_12331,N_12689);
xnor U13551 (N_13551,N_12839,N_12751);
and U13552 (N_13552,N_12443,N_12838);
xnor U13553 (N_13553,N_12411,N_12333);
nor U13554 (N_13554,N_12032,N_12026);
nand U13555 (N_13555,N_12582,N_12364);
nor U13556 (N_13556,N_12907,N_12273);
nand U13557 (N_13557,N_12818,N_12632);
or U13558 (N_13558,N_12947,N_12344);
nand U13559 (N_13559,N_12015,N_12493);
and U13560 (N_13560,N_12146,N_12154);
nor U13561 (N_13561,N_12127,N_12742);
and U13562 (N_13562,N_12951,N_12847);
xnor U13563 (N_13563,N_12332,N_12393);
and U13564 (N_13564,N_12509,N_12566);
or U13565 (N_13565,N_12029,N_12179);
nor U13566 (N_13566,N_12761,N_12962);
or U13567 (N_13567,N_12849,N_12400);
or U13568 (N_13568,N_12700,N_12339);
nor U13569 (N_13569,N_12319,N_12427);
nor U13570 (N_13570,N_12208,N_12261);
or U13571 (N_13571,N_12641,N_12928);
or U13572 (N_13572,N_12710,N_12108);
or U13573 (N_13573,N_12403,N_12443);
nor U13574 (N_13574,N_12693,N_12935);
xnor U13575 (N_13575,N_12707,N_12604);
nand U13576 (N_13576,N_12934,N_12641);
or U13577 (N_13577,N_12748,N_12526);
and U13578 (N_13578,N_12454,N_12661);
nand U13579 (N_13579,N_12102,N_12605);
xor U13580 (N_13580,N_12250,N_12242);
or U13581 (N_13581,N_12238,N_12734);
nand U13582 (N_13582,N_12166,N_12302);
nand U13583 (N_13583,N_12906,N_12670);
or U13584 (N_13584,N_12013,N_12402);
and U13585 (N_13585,N_12697,N_12919);
nand U13586 (N_13586,N_12701,N_12180);
nor U13587 (N_13587,N_12377,N_12999);
and U13588 (N_13588,N_12723,N_12487);
and U13589 (N_13589,N_12713,N_12276);
xor U13590 (N_13590,N_12635,N_12308);
and U13591 (N_13591,N_12629,N_12880);
nor U13592 (N_13592,N_12903,N_12024);
nor U13593 (N_13593,N_12550,N_12258);
nor U13594 (N_13594,N_12669,N_12005);
or U13595 (N_13595,N_12197,N_12097);
nor U13596 (N_13596,N_12657,N_12314);
or U13597 (N_13597,N_12800,N_12781);
or U13598 (N_13598,N_12478,N_12129);
or U13599 (N_13599,N_12017,N_12303);
nand U13600 (N_13600,N_12791,N_12645);
nor U13601 (N_13601,N_12543,N_12254);
or U13602 (N_13602,N_12645,N_12232);
nand U13603 (N_13603,N_12212,N_12163);
nor U13604 (N_13604,N_12258,N_12950);
or U13605 (N_13605,N_12749,N_12303);
or U13606 (N_13606,N_12465,N_12407);
and U13607 (N_13607,N_12238,N_12925);
nor U13608 (N_13608,N_12620,N_12805);
and U13609 (N_13609,N_12523,N_12229);
and U13610 (N_13610,N_12346,N_12333);
nand U13611 (N_13611,N_12529,N_12689);
and U13612 (N_13612,N_12647,N_12684);
or U13613 (N_13613,N_12429,N_12843);
nand U13614 (N_13614,N_12715,N_12263);
nand U13615 (N_13615,N_12926,N_12840);
nor U13616 (N_13616,N_12680,N_12394);
or U13617 (N_13617,N_12891,N_12711);
or U13618 (N_13618,N_12075,N_12570);
xnor U13619 (N_13619,N_12353,N_12442);
and U13620 (N_13620,N_12403,N_12742);
or U13621 (N_13621,N_12795,N_12370);
nand U13622 (N_13622,N_12294,N_12877);
and U13623 (N_13623,N_12674,N_12761);
and U13624 (N_13624,N_12993,N_12034);
xor U13625 (N_13625,N_12506,N_12381);
nand U13626 (N_13626,N_12215,N_12452);
and U13627 (N_13627,N_12511,N_12587);
and U13628 (N_13628,N_12194,N_12955);
xnor U13629 (N_13629,N_12438,N_12511);
nand U13630 (N_13630,N_12720,N_12560);
nand U13631 (N_13631,N_12049,N_12131);
and U13632 (N_13632,N_12554,N_12315);
nand U13633 (N_13633,N_12984,N_12512);
nor U13634 (N_13634,N_12219,N_12464);
and U13635 (N_13635,N_12466,N_12390);
or U13636 (N_13636,N_12815,N_12968);
and U13637 (N_13637,N_12168,N_12355);
nor U13638 (N_13638,N_12945,N_12631);
nand U13639 (N_13639,N_12860,N_12327);
or U13640 (N_13640,N_12954,N_12603);
xor U13641 (N_13641,N_12074,N_12433);
xor U13642 (N_13642,N_12353,N_12296);
or U13643 (N_13643,N_12222,N_12986);
and U13644 (N_13644,N_12186,N_12227);
and U13645 (N_13645,N_12967,N_12662);
xnor U13646 (N_13646,N_12947,N_12866);
and U13647 (N_13647,N_12669,N_12835);
nor U13648 (N_13648,N_12750,N_12843);
nand U13649 (N_13649,N_12979,N_12512);
xor U13650 (N_13650,N_12507,N_12605);
and U13651 (N_13651,N_12109,N_12995);
or U13652 (N_13652,N_12957,N_12489);
or U13653 (N_13653,N_12786,N_12003);
nand U13654 (N_13654,N_12018,N_12960);
xnor U13655 (N_13655,N_12502,N_12681);
and U13656 (N_13656,N_12838,N_12228);
or U13657 (N_13657,N_12368,N_12041);
or U13658 (N_13658,N_12533,N_12062);
or U13659 (N_13659,N_12240,N_12646);
nand U13660 (N_13660,N_12755,N_12297);
nand U13661 (N_13661,N_12789,N_12218);
nor U13662 (N_13662,N_12535,N_12757);
nor U13663 (N_13663,N_12030,N_12148);
and U13664 (N_13664,N_12278,N_12972);
nor U13665 (N_13665,N_12732,N_12084);
or U13666 (N_13666,N_12275,N_12447);
nand U13667 (N_13667,N_12117,N_12701);
nor U13668 (N_13668,N_12035,N_12497);
nor U13669 (N_13669,N_12690,N_12243);
or U13670 (N_13670,N_12434,N_12344);
xnor U13671 (N_13671,N_12711,N_12974);
xor U13672 (N_13672,N_12388,N_12018);
nand U13673 (N_13673,N_12521,N_12911);
or U13674 (N_13674,N_12480,N_12331);
xor U13675 (N_13675,N_12533,N_12359);
and U13676 (N_13676,N_12216,N_12078);
or U13677 (N_13677,N_12443,N_12200);
and U13678 (N_13678,N_12225,N_12579);
or U13679 (N_13679,N_12954,N_12987);
and U13680 (N_13680,N_12314,N_12765);
or U13681 (N_13681,N_12746,N_12301);
nand U13682 (N_13682,N_12560,N_12325);
or U13683 (N_13683,N_12900,N_12045);
xor U13684 (N_13684,N_12909,N_12468);
or U13685 (N_13685,N_12114,N_12709);
nand U13686 (N_13686,N_12891,N_12498);
or U13687 (N_13687,N_12928,N_12870);
nand U13688 (N_13688,N_12533,N_12397);
or U13689 (N_13689,N_12157,N_12130);
nand U13690 (N_13690,N_12255,N_12032);
nand U13691 (N_13691,N_12737,N_12179);
nand U13692 (N_13692,N_12736,N_12949);
or U13693 (N_13693,N_12411,N_12769);
nor U13694 (N_13694,N_12248,N_12819);
nand U13695 (N_13695,N_12118,N_12506);
xnor U13696 (N_13696,N_12549,N_12771);
nand U13697 (N_13697,N_12000,N_12219);
nand U13698 (N_13698,N_12074,N_12796);
nand U13699 (N_13699,N_12778,N_12614);
nor U13700 (N_13700,N_12717,N_12163);
nor U13701 (N_13701,N_12205,N_12363);
nand U13702 (N_13702,N_12253,N_12506);
and U13703 (N_13703,N_12446,N_12791);
nor U13704 (N_13704,N_12864,N_12155);
or U13705 (N_13705,N_12523,N_12099);
nand U13706 (N_13706,N_12375,N_12908);
or U13707 (N_13707,N_12953,N_12769);
and U13708 (N_13708,N_12863,N_12145);
or U13709 (N_13709,N_12096,N_12208);
or U13710 (N_13710,N_12019,N_12135);
nand U13711 (N_13711,N_12809,N_12727);
nand U13712 (N_13712,N_12136,N_12265);
nor U13713 (N_13713,N_12050,N_12695);
or U13714 (N_13714,N_12844,N_12971);
nand U13715 (N_13715,N_12800,N_12395);
and U13716 (N_13716,N_12059,N_12949);
nand U13717 (N_13717,N_12942,N_12463);
or U13718 (N_13718,N_12070,N_12447);
nand U13719 (N_13719,N_12126,N_12826);
and U13720 (N_13720,N_12752,N_12978);
nand U13721 (N_13721,N_12468,N_12792);
nor U13722 (N_13722,N_12202,N_12096);
xnor U13723 (N_13723,N_12922,N_12446);
nand U13724 (N_13724,N_12387,N_12033);
or U13725 (N_13725,N_12827,N_12945);
nand U13726 (N_13726,N_12487,N_12663);
and U13727 (N_13727,N_12702,N_12075);
nor U13728 (N_13728,N_12966,N_12140);
and U13729 (N_13729,N_12141,N_12273);
or U13730 (N_13730,N_12368,N_12917);
xnor U13731 (N_13731,N_12987,N_12274);
or U13732 (N_13732,N_12769,N_12789);
nor U13733 (N_13733,N_12365,N_12757);
nand U13734 (N_13734,N_12773,N_12759);
or U13735 (N_13735,N_12520,N_12830);
nand U13736 (N_13736,N_12875,N_12596);
xnor U13737 (N_13737,N_12093,N_12328);
and U13738 (N_13738,N_12982,N_12574);
and U13739 (N_13739,N_12456,N_12191);
nor U13740 (N_13740,N_12392,N_12928);
xnor U13741 (N_13741,N_12977,N_12870);
xnor U13742 (N_13742,N_12778,N_12564);
and U13743 (N_13743,N_12044,N_12591);
nand U13744 (N_13744,N_12145,N_12641);
nand U13745 (N_13745,N_12971,N_12000);
nor U13746 (N_13746,N_12463,N_12321);
nand U13747 (N_13747,N_12373,N_12535);
nand U13748 (N_13748,N_12417,N_12014);
nor U13749 (N_13749,N_12102,N_12293);
or U13750 (N_13750,N_12746,N_12558);
nor U13751 (N_13751,N_12683,N_12842);
and U13752 (N_13752,N_12666,N_12480);
nor U13753 (N_13753,N_12750,N_12459);
xor U13754 (N_13754,N_12562,N_12208);
nor U13755 (N_13755,N_12208,N_12186);
and U13756 (N_13756,N_12389,N_12902);
and U13757 (N_13757,N_12194,N_12444);
nor U13758 (N_13758,N_12477,N_12046);
and U13759 (N_13759,N_12650,N_12491);
xnor U13760 (N_13760,N_12429,N_12572);
nand U13761 (N_13761,N_12610,N_12066);
and U13762 (N_13762,N_12732,N_12516);
nand U13763 (N_13763,N_12077,N_12104);
nand U13764 (N_13764,N_12064,N_12971);
or U13765 (N_13765,N_12185,N_12469);
or U13766 (N_13766,N_12677,N_12296);
and U13767 (N_13767,N_12667,N_12433);
or U13768 (N_13768,N_12000,N_12164);
or U13769 (N_13769,N_12433,N_12465);
nor U13770 (N_13770,N_12913,N_12764);
nor U13771 (N_13771,N_12723,N_12009);
and U13772 (N_13772,N_12882,N_12516);
and U13773 (N_13773,N_12190,N_12180);
or U13774 (N_13774,N_12249,N_12988);
nand U13775 (N_13775,N_12635,N_12100);
nor U13776 (N_13776,N_12380,N_12072);
or U13777 (N_13777,N_12452,N_12691);
nand U13778 (N_13778,N_12982,N_12213);
nand U13779 (N_13779,N_12605,N_12865);
nand U13780 (N_13780,N_12448,N_12889);
xor U13781 (N_13781,N_12757,N_12740);
and U13782 (N_13782,N_12066,N_12925);
or U13783 (N_13783,N_12282,N_12816);
and U13784 (N_13784,N_12468,N_12778);
or U13785 (N_13785,N_12256,N_12976);
nor U13786 (N_13786,N_12958,N_12107);
nor U13787 (N_13787,N_12278,N_12087);
or U13788 (N_13788,N_12471,N_12742);
or U13789 (N_13789,N_12794,N_12675);
nor U13790 (N_13790,N_12233,N_12079);
or U13791 (N_13791,N_12240,N_12493);
nor U13792 (N_13792,N_12332,N_12723);
xnor U13793 (N_13793,N_12346,N_12541);
nand U13794 (N_13794,N_12777,N_12221);
and U13795 (N_13795,N_12430,N_12096);
and U13796 (N_13796,N_12707,N_12869);
nor U13797 (N_13797,N_12942,N_12932);
or U13798 (N_13798,N_12055,N_12983);
nand U13799 (N_13799,N_12246,N_12559);
nor U13800 (N_13800,N_12693,N_12213);
and U13801 (N_13801,N_12482,N_12594);
or U13802 (N_13802,N_12907,N_12720);
or U13803 (N_13803,N_12494,N_12674);
or U13804 (N_13804,N_12970,N_12922);
or U13805 (N_13805,N_12964,N_12183);
and U13806 (N_13806,N_12369,N_12347);
nor U13807 (N_13807,N_12056,N_12385);
and U13808 (N_13808,N_12088,N_12313);
nor U13809 (N_13809,N_12648,N_12238);
nor U13810 (N_13810,N_12569,N_12872);
nand U13811 (N_13811,N_12099,N_12386);
and U13812 (N_13812,N_12862,N_12209);
or U13813 (N_13813,N_12849,N_12059);
nand U13814 (N_13814,N_12855,N_12427);
nand U13815 (N_13815,N_12096,N_12674);
nor U13816 (N_13816,N_12025,N_12425);
and U13817 (N_13817,N_12299,N_12380);
nor U13818 (N_13818,N_12165,N_12229);
and U13819 (N_13819,N_12280,N_12480);
or U13820 (N_13820,N_12289,N_12734);
nand U13821 (N_13821,N_12204,N_12819);
nor U13822 (N_13822,N_12283,N_12686);
and U13823 (N_13823,N_12353,N_12399);
and U13824 (N_13824,N_12345,N_12600);
or U13825 (N_13825,N_12453,N_12312);
nor U13826 (N_13826,N_12197,N_12722);
or U13827 (N_13827,N_12072,N_12558);
nor U13828 (N_13828,N_12361,N_12865);
or U13829 (N_13829,N_12442,N_12199);
and U13830 (N_13830,N_12766,N_12901);
nor U13831 (N_13831,N_12372,N_12741);
or U13832 (N_13832,N_12185,N_12671);
and U13833 (N_13833,N_12048,N_12744);
and U13834 (N_13834,N_12498,N_12363);
nand U13835 (N_13835,N_12782,N_12142);
nor U13836 (N_13836,N_12767,N_12402);
or U13837 (N_13837,N_12042,N_12557);
nor U13838 (N_13838,N_12001,N_12275);
nand U13839 (N_13839,N_12362,N_12382);
nor U13840 (N_13840,N_12642,N_12603);
nor U13841 (N_13841,N_12017,N_12004);
or U13842 (N_13842,N_12971,N_12238);
or U13843 (N_13843,N_12414,N_12175);
and U13844 (N_13844,N_12287,N_12491);
or U13845 (N_13845,N_12176,N_12336);
nand U13846 (N_13846,N_12097,N_12521);
nand U13847 (N_13847,N_12801,N_12374);
nor U13848 (N_13848,N_12569,N_12318);
and U13849 (N_13849,N_12630,N_12974);
nand U13850 (N_13850,N_12355,N_12034);
xnor U13851 (N_13851,N_12098,N_12932);
or U13852 (N_13852,N_12452,N_12813);
and U13853 (N_13853,N_12359,N_12430);
xor U13854 (N_13854,N_12255,N_12490);
nor U13855 (N_13855,N_12214,N_12227);
xnor U13856 (N_13856,N_12456,N_12292);
or U13857 (N_13857,N_12150,N_12670);
and U13858 (N_13858,N_12984,N_12094);
or U13859 (N_13859,N_12869,N_12422);
and U13860 (N_13860,N_12002,N_12726);
and U13861 (N_13861,N_12996,N_12781);
xnor U13862 (N_13862,N_12856,N_12174);
nand U13863 (N_13863,N_12311,N_12963);
nor U13864 (N_13864,N_12878,N_12489);
and U13865 (N_13865,N_12898,N_12740);
nor U13866 (N_13866,N_12092,N_12222);
nand U13867 (N_13867,N_12188,N_12341);
or U13868 (N_13868,N_12284,N_12778);
and U13869 (N_13869,N_12353,N_12492);
nand U13870 (N_13870,N_12770,N_12937);
nor U13871 (N_13871,N_12792,N_12413);
and U13872 (N_13872,N_12465,N_12860);
or U13873 (N_13873,N_12038,N_12347);
nor U13874 (N_13874,N_12162,N_12920);
nand U13875 (N_13875,N_12879,N_12356);
nand U13876 (N_13876,N_12011,N_12436);
xnor U13877 (N_13877,N_12574,N_12568);
or U13878 (N_13878,N_12354,N_12889);
nand U13879 (N_13879,N_12797,N_12617);
nand U13880 (N_13880,N_12539,N_12351);
and U13881 (N_13881,N_12251,N_12190);
or U13882 (N_13882,N_12552,N_12053);
nand U13883 (N_13883,N_12071,N_12874);
or U13884 (N_13884,N_12968,N_12154);
xor U13885 (N_13885,N_12686,N_12867);
nor U13886 (N_13886,N_12862,N_12353);
or U13887 (N_13887,N_12773,N_12553);
nand U13888 (N_13888,N_12110,N_12569);
and U13889 (N_13889,N_12583,N_12771);
nand U13890 (N_13890,N_12386,N_12013);
nand U13891 (N_13891,N_12749,N_12660);
and U13892 (N_13892,N_12782,N_12840);
xor U13893 (N_13893,N_12228,N_12250);
and U13894 (N_13894,N_12534,N_12885);
nand U13895 (N_13895,N_12299,N_12873);
nand U13896 (N_13896,N_12420,N_12927);
and U13897 (N_13897,N_12922,N_12279);
and U13898 (N_13898,N_12961,N_12604);
or U13899 (N_13899,N_12069,N_12011);
nor U13900 (N_13900,N_12976,N_12705);
and U13901 (N_13901,N_12434,N_12913);
nor U13902 (N_13902,N_12228,N_12553);
or U13903 (N_13903,N_12342,N_12626);
and U13904 (N_13904,N_12270,N_12941);
nand U13905 (N_13905,N_12123,N_12240);
nor U13906 (N_13906,N_12684,N_12532);
nor U13907 (N_13907,N_12676,N_12892);
nor U13908 (N_13908,N_12216,N_12033);
nand U13909 (N_13909,N_12068,N_12764);
nand U13910 (N_13910,N_12471,N_12317);
or U13911 (N_13911,N_12752,N_12805);
or U13912 (N_13912,N_12029,N_12501);
xor U13913 (N_13913,N_12125,N_12555);
or U13914 (N_13914,N_12150,N_12494);
or U13915 (N_13915,N_12929,N_12760);
nor U13916 (N_13916,N_12993,N_12423);
nand U13917 (N_13917,N_12693,N_12277);
nand U13918 (N_13918,N_12258,N_12367);
and U13919 (N_13919,N_12330,N_12959);
xor U13920 (N_13920,N_12185,N_12204);
xor U13921 (N_13921,N_12771,N_12777);
and U13922 (N_13922,N_12722,N_12644);
and U13923 (N_13923,N_12271,N_12088);
nand U13924 (N_13924,N_12413,N_12016);
nand U13925 (N_13925,N_12830,N_12835);
or U13926 (N_13926,N_12019,N_12023);
and U13927 (N_13927,N_12665,N_12363);
and U13928 (N_13928,N_12563,N_12517);
nor U13929 (N_13929,N_12940,N_12474);
nand U13930 (N_13930,N_12615,N_12334);
xnor U13931 (N_13931,N_12780,N_12675);
xnor U13932 (N_13932,N_12767,N_12879);
xnor U13933 (N_13933,N_12964,N_12988);
or U13934 (N_13934,N_12103,N_12774);
nor U13935 (N_13935,N_12868,N_12913);
or U13936 (N_13936,N_12549,N_12171);
nor U13937 (N_13937,N_12356,N_12167);
and U13938 (N_13938,N_12501,N_12649);
and U13939 (N_13939,N_12278,N_12962);
and U13940 (N_13940,N_12114,N_12688);
and U13941 (N_13941,N_12557,N_12039);
nor U13942 (N_13942,N_12553,N_12267);
and U13943 (N_13943,N_12136,N_12079);
nand U13944 (N_13944,N_12517,N_12834);
nand U13945 (N_13945,N_12278,N_12296);
nor U13946 (N_13946,N_12498,N_12274);
or U13947 (N_13947,N_12916,N_12390);
xor U13948 (N_13948,N_12722,N_12519);
and U13949 (N_13949,N_12112,N_12870);
and U13950 (N_13950,N_12254,N_12397);
or U13951 (N_13951,N_12026,N_12471);
nand U13952 (N_13952,N_12651,N_12360);
and U13953 (N_13953,N_12180,N_12514);
and U13954 (N_13954,N_12596,N_12952);
xnor U13955 (N_13955,N_12965,N_12380);
and U13956 (N_13956,N_12819,N_12429);
nor U13957 (N_13957,N_12534,N_12498);
and U13958 (N_13958,N_12767,N_12162);
and U13959 (N_13959,N_12193,N_12012);
nor U13960 (N_13960,N_12545,N_12843);
and U13961 (N_13961,N_12552,N_12444);
and U13962 (N_13962,N_12206,N_12371);
nor U13963 (N_13963,N_12855,N_12344);
nor U13964 (N_13964,N_12564,N_12237);
nor U13965 (N_13965,N_12581,N_12783);
or U13966 (N_13966,N_12107,N_12899);
nand U13967 (N_13967,N_12482,N_12457);
and U13968 (N_13968,N_12978,N_12972);
nand U13969 (N_13969,N_12824,N_12727);
or U13970 (N_13970,N_12639,N_12189);
nand U13971 (N_13971,N_12788,N_12007);
nor U13972 (N_13972,N_12991,N_12692);
nand U13973 (N_13973,N_12487,N_12108);
and U13974 (N_13974,N_12538,N_12280);
and U13975 (N_13975,N_12513,N_12184);
or U13976 (N_13976,N_12809,N_12507);
and U13977 (N_13977,N_12314,N_12907);
nor U13978 (N_13978,N_12665,N_12173);
nor U13979 (N_13979,N_12845,N_12984);
or U13980 (N_13980,N_12638,N_12214);
nor U13981 (N_13981,N_12925,N_12193);
or U13982 (N_13982,N_12266,N_12593);
or U13983 (N_13983,N_12799,N_12551);
or U13984 (N_13984,N_12468,N_12855);
nor U13985 (N_13985,N_12763,N_12579);
or U13986 (N_13986,N_12404,N_12046);
nor U13987 (N_13987,N_12106,N_12415);
nand U13988 (N_13988,N_12394,N_12365);
or U13989 (N_13989,N_12225,N_12045);
or U13990 (N_13990,N_12150,N_12823);
nand U13991 (N_13991,N_12135,N_12304);
nand U13992 (N_13992,N_12803,N_12625);
nand U13993 (N_13993,N_12949,N_12578);
xnor U13994 (N_13994,N_12621,N_12724);
nand U13995 (N_13995,N_12353,N_12594);
nand U13996 (N_13996,N_12606,N_12772);
xor U13997 (N_13997,N_12513,N_12113);
or U13998 (N_13998,N_12009,N_12734);
nor U13999 (N_13999,N_12766,N_12909);
nand U14000 (N_14000,N_13303,N_13545);
or U14001 (N_14001,N_13081,N_13880);
nand U14002 (N_14002,N_13171,N_13702);
nor U14003 (N_14003,N_13480,N_13247);
nand U14004 (N_14004,N_13503,N_13540);
nand U14005 (N_14005,N_13878,N_13906);
or U14006 (N_14006,N_13309,N_13846);
and U14007 (N_14007,N_13167,N_13570);
or U14008 (N_14008,N_13196,N_13583);
xnor U14009 (N_14009,N_13618,N_13689);
nor U14010 (N_14010,N_13682,N_13304);
and U14011 (N_14011,N_13924,N_13329);
xnor U14012 (N_14012,N_13378,N_13202);
and U14013 (N_14013,N_13027,N_13705);
and U14014 (N_14014,N_13730,N_13148);
nor U14015 (N_14015,N_13987,N_13893);
nor U14016 (N_14016,N_13512,N_13157);
and U14017 (N_14017,N_13007,N_13984);
or U14018 (N_14018,N_13737,N_13700);
or U14019 (N_14019,N_13429,N_13733);
nand U14020 (N_14020,N_13346,N_13975);
xnor U14021 (N_14021,N_13103,N_13745);
nand U14022 (N_14022,N_13079,N_13129);
or U14023 (N_14023,N_13375,N_13664);
nor U14024 (N_14024,N_13798,N_13553);
nand U14025 (N_14025,N_13248,N_13711);
or U14026 (N_14026,N_13505,N_13881);
nand U14027 (N_14027,N_13960,N_13038);
or U14028 (N_14028,N_13147,N_13900);
and U14029 (N_14029,N_13504,N_13067);
or U14030 (N_14030,N_13982,N_13001);
nor U14031 (N_14031,N_13190,N_13670);
nand U14032 (N_14032,N_13181,N_13322);
nand U14033 (N_14033,N_13811,N_13792);
and U14034 (N_14034,N_13245,N_13986);
nand U14035 (N_14035,N_13568,N_13166);
nor U14036 (N_14036,N_13841,N_13518);
and U14037 (N_14037,N_13966,N_13735);
and U14038 (N_14038,N_13951,N_13337);
and U14039 (N_14039,N_13845,N_13954);
or U14040 (N_14040,N_13649,N_13617);
nand U14041 (N_14041,N_13660,N_13866);
nor U14042 (N_14042,N_13569,N_13615);
nand U14043 (N_14043,N_13541,N_13361);
nor U14044 (N_14044,N_13099,N_13921);
or U14045 (N_14045,N_13952,N_13176);
nand U14046 (N_14046,N_13392,N_13738);
and U14047 (N_14047,N_13749,N_13755);
nor U14048 (N_14048,N_13348,N_13474);
and U14049 (N_14049,N_13154,N_13944);
xor U14050 (N_14050,N_13035,N_13150);
nor U14051 (N_14051,N_13650,N_13973);
nand U14052 (N_14052,N_13642,N_13253);
and U14053 (N_14053,N_13076,N_13736);
nand U14054 (N_14054,N_13370,N_13580);
nor U14055 (N_14055,N_13529,N_13948);
nand U14056 (N_14056,N_13972,N_13255);
or U14057 (N_14057,N_13808,N_13544);
nor U14058 (N_14058,N_13832,N_13399);
or U14059 (N_14059,N_13108,N_13827);
or U14060 (N_14060,N_13719,N_13352);
nor U14061 (N_14061,N_13523,N_13968);
xnor U14062 (N_14062,N_13587,N_13913);
nor U14063 (N_14063,N_13121,N_13620);
nor U14064 (N_14064,N_13416,N_13830);
and U14065 (N_14065,N_13115,N_13863);
nor U14066 (N_14066,N_13117,N_13957);
nand U14067 (N_14067,N_13934,N_13872);
nand U14068 (N_14068,N_13596,N_13419);
xnor U14069 (N_14069,N_13888,N_13442);
and U14070 (N_14070,N_13050,N_13272);
and U14071 (N_14071,N_13669,N_13712);
nand U14072 (N_14072,N_13155,N_13858);
and U14073 (N_14073,N_13572,N_13242);
nand U14074 (N_14074,N_13661,N_13233);
nand U14075 (N_14075,N_13856,N_13410);
nand U14076 (N_14076,N_13066,N_13211);
or U14077 (N_14077,N_13899,N_13327);
xnor U14078 (N_14078,N_13078,N_13110);
and U14079 (N_14079,N_13034,N_13377);
xnor U14080 (N_14080,N_13360,N_13292);
and U14081 (N_14081,N_13051,N_13964);
or U14082 (N_14082,N_13491,N_13865);
nand U14083 (N_14083,N_13404,N_13720);
and U14084 (N_14084,N_13767,N_13376);
and U14085 (N_14085,N_13867,N_13036);
or U14086 (N_14086,N_13500,N_13374);
nor U14087 (N_14087,N_13631,N_13422);
and U14088 (N_14088,N_13042,N_13123);
and U14089 (N_14089,N_13852,N_13462);
or U14090 (N_14090,N_13588,N_13601);
or U14091 (N_14091,N_13552,N_13160);
or U14092 (N_14092,N_13603,N_13930);
and U14093 (N_14093,N_13903,N_13291);
xnor U14094 (N_14094,N_13581,N_13164);
nand U14095 (N_14095,N_13061,N_13116);
or U14096 (N_14096,N_13482,N_13560);
and U14097 (N_14097,N_13006,N_13487);
nor U14098 (N_14098,N_13198,N_13688);
nor U14099 (N_14099,N_13473,N_13916);
or U14100 (N_14100,N_13046,N_13999);
and U14101 (N_14101,N_13842,N_13988);
or U14102 (N_14102,N_13490,N_13470);
or U14103 (N_14103,N_13056,N_13464);
nand U14104 (N_14104,N_13140,N_13862);
nor U14105 (N_14105,N_13223,N_13850);
or U14106 (N_14106,N_13188,N_13525);
and U14107 (N_14107,N_13831,N_13119);
or U14108 (N_14108,N_13182,N_13721);
nand U14109 (N_14109,N_13316,N_13278);
and U14110 (N_14110,N_13232,N_13911);
xnor U14111 (N_14111,N_13195,N_13270);
or U14112 (N_14112,N_13695,N_13691);
xor U14113 (N_14113,N_13187,N_13648);
or U14114 (N_14114,N_13288,N_13917);
and U14115 (N_14115,N_13566,N_13633);
and U14116 (N_14116,N_13716,N_13991);
nor U14117 (N_14117,N_13124,N_13112);
nand U14118 (N_14118,N_13969,N_13571);
and U14119 (N_14119,N_13282,N_13179);
nand U14120 (N_14120,N_13443,N_13795);
or U14121 (N_14121,N_13889,N_13380);
nand U14122 (N_14122,N_13997,N_13373);
or U14123 (N_14123,N_13463,N_13345);
nor U14124 (N_14124,N_13747,N_13275);
nor U14125 (N_14125,N_13130,N_13848);
xnor U14126 (N_14126,N_13885,N_13684);
nand U14127 (N_14127,N_13237,N_13871);
or U14128 (N_14128,N_13981,N_13467);
and U14129 (N_14129,N_13174,N_13090);
xnor U14130 (N_14130,N_13805,N_13979);
or U14131 (N_14131,N_13853,N_13213);
and U14132 (N_14132,N_13200,N_13877);
xnor U14133 (N_14133,N_13135,N_13466);
xnor U14134 (N_14134,N_13479,N_13677);
nor U14135 (N_14135,N_13353,N_13168);
or U14136 (N_14136,N_13502,N_13536);
or U14137 (N_14137,N_13004,N_13744);
or U14138 (N_14138,N_13976,N_13388);
xnor U14139 (N_14139,N_13514,N_13980);
and U14140 (N_14140,N_13883,N_13335);
xnor U14141 (N_14141,N_13136,N_13595);
or U14142 (N_14142,N_13229,N_13221);
or U14143 (N_14143,N_13177,N_13073);
nand U14144 (N_14144,N_13095,N_13000);
and U14145 (N_14145,N_13647,N_13781);
or U14146 (N_14146,N_13582,N_13923);
or U14147 (N_14147,N_13936,N_13801);
xnor U14148 (N_14148,N_13494,N_13797);
nor U14149 (N_14149,N_13059,N_13778);
xor U14150 (N_14150,N_13608,N_13817);
and U14151 (N_14151,N_13891,N_13683);
nand U14152 (N_14152,N_13365,N_13325);
or U14153 (N_14153,N_13089,N_13996);
or U14154 (N_14154,N_13145,N_13731);
and U14155 (N_14155,N_13412,N_13816);
nor U14156 (N_14156,N_13704,N_13803);
or U14157 (N_14157,N_13457,N_13426);
and U14158 (N_14158,N_13625,N_13561);
nor U14159 (N_14159,N_13896,N_13387);
and U14160 (N_14160,N_13113,N_13486);
and U14161 (N_14161,N_13768,N_13409);
nand U14162 (N_14162,N_13098,N_13860);
nor U14163 (N_14163,N_13125,N_13630);
and U14164 (N_14164,N_13501,N_13144);
and U14165 (N_14165,N_13926,N_13932);
and U14166 (N_14166,N_13260,N_13092);
or U14167 (N_14167,N_13937,N_13591);
or U14168 (N_14168,N_13551,N_13105);
nor U14169 (N_14169,N_13621,N_13268);
or U14170 (N_14170,N_13657,N_13938);
xnor U14171 (N_14171,N_13658,N_13756);
nor U14172 (N_14172,N_13386,N_13524);
nor U14173 (N_14173,N_13610,N_13029);
or U14174 (N_14174,N_13822,N_13623);
xor U14175 (N_14175,N_13220,N_13793);
nor U14176 (N_14176,N_13199,N_13653);
or U14177 (N_14177,N_13989,N_13627);
and U14178 (N_14178,N_13879,N_13192);
or U14179 (N_14179,N_13077,N_13334);
nand U14180 (N_14180,N_13602,N_13687);
and U14181 (N_14181,N_13363,N_13895);
nor U14182 (N_14182,N_13306,N_13507);
nor U14183 (N_14183,N_13718,N_13611);
nand U14184 (N_14184,N_13577,N_13598);
nor U14185 (N_14185,N_13537,N_13178);
and U14186 (N_14186,N_13428,N_13481);
or U14187 (N_14187,N_13834,N_13234);
xnor U14188 (N_14188,N_13813,N_13590);
nand U14189 (N_14189,N_13604,N_13405);
nor U14190 (N_14190,N_13764,N_13641);
or U14191 (N_14191,N_13654,N_13946);
or U14192 (N_14192,N_13472,N_13851);
or U14193 (N_14193,N_13806,N_13918);
nand U14194 (N_14194,N_13025,N_13120);
nor U14195 (N_14195,N_13939,N_13681);
and U14196 (N_14196,N_13209,N_13995);
nand U14197 (N_14197,N_13673,N_13859);
xor U14198 (N_14198,N_13478,N_13638);
xor U14199 (N_14199,N_13364,N_13186);
and U14200 (N_14200,N_13301,N_13729);
nand U14201 (N_14201,N_13499,N_13096);
and U14202 (N_14202,N_13037,N_13520);
nor U14203 (N_14203,N_13751,N_13961);
nand U14204 (N_14204,N_13055,N_13983);
or U14205 (N_14205,N_13314,N_13297);
and U14206 (N_14206,N_13875,N_13323);
nor U14207 (N_14207,N_13236,N_13897);
and U14208 (N_14208,N_13715,N_13384);
nor U14209 (N_14209,N_13251,N_13597);
or U14210 (N_14210,N_13840,N_13224);
xor U14211 (N_14211,N_13819,N_13488);
nor U14212 (N_14212,N_13743,N_13626);
or U14213 (N_14213,N_13773,N_13243);
nor U14214 (N_14214,N_13857,N_13225);
nand U14215 (N_14215,N_13100,N_13599);
or U14216 (N_14216,N_13958,N_13530);
nor U14217 (N_14217,N_13635,N_13458);
nor U14218 (N_14218,N_13414,N_13726);
nand U14219 (N_14219,N_13444,N_13172);
xnor U14220 (N_14220,N_13040,N_13210);
xnor U14221 (N_14221,N_13252,N_13927);
or U14222 (N_14222,N_13855,N_13022);
nand U14223 (N_14223,N_13293,N_13612);
or U14224 (N_14224,N_13928,N_13065);
nand U14225 (N_14225,N_13261,N_13894);
xnor U14226 (N_14226,N_13655,N_13594);
nor U14227 (N_14227,N_13132,N_13344);
and U14228 (N_14228,N_13723,N_13156);
and U14229 (N_14229,N_13315,N_13519);
and U14230 (N_14230,N_13777,N_13060);
nand U14231 (N_14231,N_13824,N_13455);
and U14232 (N_14232,N_13393,N_13699);
nor U14233 (N_14233,N_13139,N_13593);
nor U14234 (N_14234,N_13692,N_13659);
or U14235 (N_14235,N_13047,N_13672);
nor U14236 (N_14236,N_13403,N_13212);
nor U14237 (N_14237,N_13489,N_13531);
xnor U14238 (N_14238,N_13574,N_13727);
nand U14239 (N_14239,N_13411,N_13671);
or U14240 (N_14240,N_13041,N_13904);
nor U14241 (N_14241,N_13662,N_13576);
nor U14242 (N_14242,N_13397,N_13362);
nor U14243 (N_14243,N_13656,N_13667);
and U14244 (N_14244,N_13907,N_13732);
nand U14245 (N_14245,N_13026,N_13356);
and U14246 (N_14246,N_13821,N_13133);
or U14247 (N_14247,N_13943,N_13039);
and U14248 (N_14248,N_13543,N_13249);
and U14249 (N_14249,N_13319,N_13350);
nand U14250 (N_14250,N_13963,N_13475);
nor U14251 (N_14251,N_13790,N_13789);
and U14252 (N_14252,N_13636,N_13367);
nand U14253 (N_14253,N_13250,N_13624);
or U14254 (N_14254,N_13456,N_13369);
nand U14255 (N_14255,N_13146,N_13263);
and U14256 (N_14256,N_13746,N_13535);
and U14257 (N_14257,N_13030,N_13754);
nor U14258 (N_14258,N_13031,N_13508);
xnor U14259 (N_14259,N_13759,N_13575);
nor U14260 (N_14260,N_13750,N_13521);
and U14261 (N_14261,N_13064,N_13045);
and U14262 (N_14262,N_13358,N_13945);
xnor U14263 (N_14263,N_13436,N_13433);
and U14264 (N_14264,N_13740,N_13246);
and U14265 (N_14265,N_13728,N_13752);
and U14266 (N_14266,N_13407,N_13547);
or U14267 (N_14267,N_13804,N_13506);
nor U14268 (N_14268,N_13940,N_13493);
or U14269 (N_14269,N_13516,N_13843);
and U14270 (N_14270,N_13269,N_13153);
or U14271 (N_14271,N_13548,N_13775);
nand U14272 (N_14272,N_13629,N_13418);
nor U14273 (N_14273,N_13435,N_13573);
xor U14274 (N_14274,N_13787,N_13083);
nand U14275 (N_14275,N_13628,N_13469);
or U14276 (N_14276,N_13734,N_13998);
and U14277 (N_14277,N_13640,N_13425);
nand U14278 (N_14278,N_13043,N_13835);
nand U14279 (N_14279,N_13258,N_13698);
or U14280 (N_14280,N_13554,N_13368);
and U14281 (N_14281,N_13665,N_13977);
nor U14282 (N_14282,N_13185,N_13949);
nand U14283 (N_14283,N_13825,N_13231);
and U14284 (N_14284,N_13194,N_13956);
and U14285 (N_14285,N_13854,N_13622);
nor U14286 (N_14286,N_13613,N_13564);
or U14287 (N_14287,N_13710,N_13351);
and U14288 (N_14288,N_13703,N_13605);
nor U14289 (N_14289,N_13336,N_13460);
nor U14290 (N_14290,N_13158,N_13317);
or U14291 (N_14291,N_13757,N_13401);
xnor U14292 (N_14292,N_13522,N_13607);
nand U14293 (N_14293,N_13539,N_13389);
nand U14294 (N_14294,N_13244,N_13550);
nor U14295 (N_14295,N_13873,N_13484);
or U14296 (N_14296,N_13264,N_13072);
or U14297 (N_14297,N_13033,N_13398);
nand U14298 (N_14298,N_13011,N_13406);
nand U14299 (N_14299,N_13791,N_13289);
and U14300 (N_14300,N_13024,N_13953);
xor U14301 (N_14301,N_13826,N_13302);
or U14302 (N_14302,N_13241,N_13218);
xor U14303 (N_14303,N_13111,N_13510);
xor U14304 (N_14304,N_13277,N_13708);
nand U14305 (N_14305,N_13391,N_13417);
xor U14306 (N_14306,N_13257,N_13465);
xor U14307 (N_14307,N_13562,N_13839);
nand U14308 (N_14308,N_13205,N_13844);
nand U14309 (N_14309,N_13634,N_13328);
nand U14310 (N_14310,N_13044,N_13062);
nand U14311 (N_14311,N_13676,N_13382);
nand U14312 (N_14312,N_13696,N_13651);
or U14313 (N_14313,N_13955,N_13584);
and U14314 (N_14314,N_13320,N_13163);
nor U14315 (N_14315,N_13993,N_13935);
nand U14316 (N_14316,N_13057,N_13886);
and U14317 (N_14317,N_13152,N_13300);
nand U14318 (N_14318,N_13606,N_13343);
or U14319 (N_14319,N_13197,N_13355);
nand U14320 (N_14320,N_13912,N_13170);
or U14321 (N_14321,N_13141,N_13015);
or U14322 (N_14322,N_13020,N_13459);
and U14323 (N_14323,N_13632,N_13331);
nor U14324 (N_14324,N_13400,N_13592);
nand U14325 (N_14325,N_13772,N_13093);
nor U14326 (N_14326,N_13215,N_13742);
xor U14327 (N_14327,N_13274,N_13347);
and U14328 (N_14328,N_13219,N_13052);
nand U14329 (N_14329,N_13313,N_13714);
nand U14330 (N_14330,N_13922,N_13214);
nand U14331 (N_14331,N_13183,N_13204);
xnor U14332 (N_14332,N_13513,N_13496);
nor U14333 (N_14333,N_13441,N_13019);
nand U14334 (N_14334,N_13118,N_13637);
and U14335 (N_14335,N_13546,N_13697);
nor U14336 (N_14336,N_13396,N_13271);
xnor U14337 (N_14337,N_13449,N_13450);
and U14338 (N_14338,N_13138,N_13833);
and U14339 (N_14339,N_13498,N_13295);
and U14340 (N_14340,N_13495,N_13959);
nor U14341 (N_14341,N_13162,N_13238);
nor U14342 (N_14342,N_13947,N_13330);
nor U14343 (N_14343,N_13189,N_13201);
or U14344 (N_14344,N_13965,N_13909);
nor U14345 (N_14345,N_13794,N_13070);
or U14346 (N_14346,N_13383,N_13701);
and U14347 (N_14347,N_13780,N_13137);
and U14348 (N_14348,N_13305,N_13771);
nor U14349 (N_14349,N_13942,N_13685);
and U14350 (N_14350,N_13381,N_13101);
nor U14351 (N_14351,N_13785,N_13799);
or U14352 (N_14352,N_13753,N_13408);
nand U14353 (N_14353,N_13901,N_13748);
and U14354 (N_14354,N_13003,N_13276);
and U14355 (N_14355,N_13849,N_13925);
xnor U14356 (N_14356,N_13663,N_13437);
nor U14357 (N_14357,N_13675,N_13193);
nor U14358 (N_14358,N_13892,N_13774);
and U14359 (N_14359,N_13461,N_13340);
nor U14360 (N_14360,N_13049,N_13971);
nor U14361 (N_14361,N_13281,N_13517);
nand U14362 (N_14362,N_13818,N_13788);
and U14363 (N_14363,N_13807,N_13102);
and U14364 (N_14364,N_13010,N_13016);
xnor U14365 (N_14365,N_13287,N_13762);
nand U14366 (N_14366,N_13814,N_13332);
and U14367 (N_14367,N_13898,N_13173);
or U14368 (N_14368,N_13294,N_13431);
and U14369 (N_14369,N_13532,N_13578);
and U14370 (N_14370,N_13815,N_13706);
or U14371 (N_14371,N_13349,N_13962);
or U14372 (N_14372,N_13549,N_13165);
and U14373 (N_14373,N_13616,N_13679);
and U14374 (N_14374,N_13161,N_13453);
and U14375 (N_14375,N_13446,N_13829);
or U14376 (N_14376,N_13870,N_13882);
nand U14377 (N_14377,N_13021,N_13722);
and U14378 (N_14378,N_13134,N_13652);
nor U14379 (N_14379,N_13765,N_13589);
or U14380 (N_14380,N_13018,N_13782);
nor U14381 (N_14381,N_13823,N_13142);
and U14382 (N_14382,N_13143,N_13690);
and U14383 (N_14383,N_13283,N_13087);
nor U14384 (N_14384,N_13239,N_13985);
or U14385 (N_14385,N_13739,N_13326);
nor U14386 (N_14386,N_13254,N_13312);
and U14387 (N_14387,N_13311,N_13256);
and U14388 (N_14388,N_13216,N_13267);
and U14389 (N_14389,N_13694,N_13128);
nand U14390 (N_14390,N_13424,N_13088);
nand U14391 (N_14391,N_13837,N_13228);
nand U14392 (N_14392,N_13678,N_13071);
nand U14393 (N_14393,N_13509,N_13008);
nand U14394 (N_14394,N_13600,N_13126);
nand U14395 (N_14395,N_13763,N_13206);
nand U14396 (N_14396,N_13032,N_13299);
or U14397 (N_14397,N_13929,N_13438);
nor U14398 (N_14398,N_13674,N_13371);
or U14399 (N_14399,N_13222,N_13127);
nor U14400 (N_14400,N_13920,N_13014);
nand U14401 (N_14401,N_13235,N_13884);
and U14402 (N_14402,N_13448,N_13796);
or U14403 (N_14403,N_13741,N_13447);
nand U14404 (N_14404,N_13009,N_13800);
or U14405 (N_14405,N_13420,N_13868);
and U14406 (N_14406,N_13054,N_13151);
xor U14407 (N_14407,N_13555,N_13203);
or U14408 (N_14408,N_13810,N_13874);
or U14409 (N_14409,N_13109,N_13012);
nand U14410 (N_14410,N_13324,N_13802);
nand U14411 (N_14411,N_13556,N_13869);
and U14412 (N_14412,N_13230,N_13533);
nor U14413 (N_14413,N_13421,N_13339);
and U14414 (N_14414,N_13227,N_13887);
nand U14415 (N_14415,N_13614,N_13298);
xnor U14416 (N_14416,N_13082,N_13058);
or U14417 (N_14417,N_13013,N_13492);
xnor U14418 (N_14418,N_13342,N_13864);
nor U14419 (N_14419,N_13511,N_13526);
nor U14420 (N_14420,N_13713,N_13318);
nand U14421 (N_14421,N_13760,N_13075);
nand U14422 (N_14422,N_13717,N_13028);
xor U14423 (N_14423,N_13776,N_13266);
and U14424 (N_14424,N_13693,N_13159);
and U14425 (N_14425,N_13766,N_13538);
nor U14426 (N_14426,N_13415,N_13341);
xor U14427 (N_14427,N_13668,N_13114);
nor U14428 (N_14428,N_13497,N_13941);
nor U14429 (N_14429,N_13445,N_13828);
or U14430 (N_14430,N_13586,N_13709);
or U14431 (N_14431,N_13812,N_13104);
nor U14432 (N_14432,N_13423,N_13908);
nor U14433 (N_14433,N_13184,N_13786);
nor U14434 (N_14434,N_13534,N_13847);
nor U14435 (N_14435,N_13567,N_13273);
or U14436 (N_14436,N_13413,N_13515);
or U14437 (N_14437,N_13175,N_13558);
and U14438 (N_14438,N_13053,N_13069);
and U14439 (N_14439,N_13565,N_13149);
and U14440 (N_14440,N_13394,N_13820);
nor U14441 (N_14441,N_13372,N_13779);
and U14442 (N_14442,N_13131,N_13310);
or U14443 (N_14443,N_13085,N_13191);
nand U14444 (N_14444,N_13080,N_13023);
and U14445 (N_14445,N_13307,N_13468);
nor U14446 (N_14446,N_13094,N_13333);
xnor U14447 (N_14447,N_13645,N_13666);
nand U14448 (N_14448,N_13528,N_13485);
or U14449 (N_14449,N_13974,N_13395);
xor U14450 (N_14450,N_13914,N_13402);
nor U14451 (N_14451,N_13861,N_13440);
or U14452 (N_14452,N_13097,N_13296);
xnor U14453 (N_14453,N_13385,N_13279);
and U14454 (N_14454,N_13207,N_13290);
nor U14455 (N_14455,N_13876,N_13579);
xor U14456 (N_14456,N_13454,N_13905);
nand U14457 (N_14457,N_13262,N_13240);
and U14458 (N_14458,N_13770,N_13619);
nand U14459 (N_14459,N_13265,N_13427);
xor U14460 (N_14460,N_13338,N_13559);
and U14461 (N_14461,N_13005,N_13725);
or U14462 (N_14462,N_13563,N_13259);
and U14463 (N_14463,N_13122,N_13091);
nand U14464 (N_14464,N_13542,N_13086);
or U14465 (N_14465,N_13308,N_13068);
nand U14466 (N_14466,N_13180,N_13390);
nor U14467 (N_14467,N_13919,N_13439);
nand U14468 (N_14468,N_13724,N_13285);
or U14469 (N_14469,N_13769,N_13838);
xor U14470 (N_14470,N_13107,N_13048);
nand U14471 (N_14471,N_13451,N_13002);
or U14472 (N_14472,N_13017,N_13284);
nand U14473 (N_14473,N_13217,N_13483);
and U14474 (N_14474,N_13471,N_13950);
nor U14475 (N_14475,N_13992,N_13910);
or U14476 (N_14476,N_13477,N_13761);
xnor U14477 (N_14477,N_13783,N_13585);
nor U14478 (N_14478,N_13639,N_13434);
nand U14479 (N_14479,N_13784,N_13933);
nand U14480 (N_14480,N_13354,N_13379);
or U14481 (N_14481,N_13644,N_13990);
nand U14482 (N_14482,N_13967,N_13359);
nand U14483 (N_14483,N_13890,N_13432);
and U14484 (N_14484,N_13994,N_13452);
nand U14485 (N_14485,N_13280,N_13646);
nand U14486 (N_14486,N_13836,N_13809);
or U14487 (N_14487,N_13430,N_13931);
or U14488 (N_14488,N_13226,N_13978);
and U14489 (N_14489,N_13758,N_13970);
and U14490 (N_14490,N_13902,N_13084);
nand U14491 (N_14491,N_13643,N_13321);
and U14492 (N_14492,N_13707,N_13063);
nor U14493 (N_14493,N_13208,N_13609);
or U14494 (N_14494,N_13680,N_13686);
nor U14495 (N_14495,N_13286,N_13476);
and U14496 (N_14496,N_13169,N_13915);
and U14497 (N_14497,N_13074,N_13106);
or U14498 (N_14498,N_13366,N_13527);
nor U14499 (N_14499,N_13357,N_13557);
nand U14500 (N_14500,N_13735,N_13250);
and U14501 (N_14501,N_13668,N_13157);
nor U14502 (N_14502,N_13780,N_13581);
nand U14503 (N_14503,N_13667,N_13949);
nor U14504 (N_14504,N_13968,N_13536);
nand U14505 (N_14505,N_13160,N_13122);
nand U14506 (N_14506,N_13317,N_13857);
nor U14507 (N_14507,N_13814,N_13712);
and U14508 (N_14508,N_13497,N_13364);
and U14509 (N_14509,N_13590,N_13343);
nor U14510 (N_14510,N_13040,N_13104);
nor U14511 (N_14511,N_13850,N_13969);
nor U14512 (N_14512,N_13591,N_13121);
nor U14513 (N_14513,N_13596,N_13593);
or U14514 (N_14514,N_13830,N_13612);
nand U14515 (N_14515,N_13442,N_13082);
or U14516 (N_14516,N_13728,N_13057);
nand U14517 (N_14517,N_13792,N_13711);
nand U14518 (N_14518,N_13287,N_13885);
xnor U14519 (N_14519,N_13888,N_13495);
and U14520 (N_14520,N_13938,N_13500);
and U14521 (N_14521,N_13476,N_13255);
nor U14522 (N_14522,N_13559,N_13764);
nor U14523 (N_14523,N_13334,N_13833);
or U14524 (N_14524,N_13817,N_13827);
nand U14525 (N_14525,N_13488,N_13383);
or U14526 (N_14526,N_13120,N_13692);
and U14527 (N_14527,N_13535,N_13334);
or U14528 (N_14528,N_13365,N_13113);
or U14529 (N_14529,N_13442,N_13131);
xor U14530 (N_14530,N_13885,N_13972);
nand U14531 (N_14531,N_13720,N_13032);
or U14532 (N_14532,N_13539,N_13725);
nand U14533 (N_14533,N_13586,N_13885);
or U14534 (N_14534,N_13387,N_13681);
and U14535 (N_14535,N_13532,N_13778);
nand U14536 (N_14536,N_13554,N_13922);
nor U14537 (N_14537,N_13907,N_13948);
xnor U14538 (N_14538,N_13458,N_13228);
or U14539 (N_14539,N_13388,N_13212);
nand U14540 (N_14540,N_13937,N_13115);
nand U14541 (N_14541,N_13721,N_13154);
and U14542 (N_14542,N_13829,N_13802);
or U14543 (N_14543,N_13305,N_13006);
and U14544 (N_14544,N_13481,N_13641);
nor U14545 (N_14545,N_13552,N_13774);
and U14546 (N_14546,N_13624,N_13582);
nand U14547 (N_14547,N_13379,N_13784);
nand U14548 (N_14548,N_13613,N_13995);
xor U14549 (N_14549,N_13548,N_13063);
and U14550 (N_14550,N_13720,N_13163);
nand U14551 (N_14551,N_13226,N_13801);
nand U14552 (N_14552,N_13343,N_13454);
nand U14553 (N_14553,N_13418,N_13176);
nor U14554 (N_14554,N_13808,N_13640);
nor U14555 (N_14555,N_13966,N_13911);
or U14556 (N_14556,N_13200,N_13454);
nor U14557 (N_14557,N_13178,N_13105);
nor U14558 (N_14558,N_13695,N_13619);
or U14559 (N_14559,N_13691,N_13994);
nand U14560 (N_14560,N_13036,N_13930);
nand U14561 (N_14561,N_13672,N_13923);
nor U14562 (N_14562,N_13962,N_13805);
nor U14563 (N_14563,N_13002,N_13895);
or U14564 (N_14564,N_13582,N_13869);
and U14565 (N_14565,N_13506,N_13980);
nand U14566 (N_14566,N_13740,N_13800);
or U14567 (N_14567,N_13570,N_13812);
or U14568 (N_14568,N_13929,N_13974);
or U14569 (N_14569,N_13538,N_13649);
nand U14570 (N_14570,N_13948,N_13511);
and U14571 (N_14571,N_13208,N_13916);
xor U14572 (N_14572,N_13713,N_13861);
nor U14573 (N_14573,N_13329,N_13896);
or U14574 (N_14574,N_13045,N_13489);
xnor U14575 (N_14575,N_13855,N_13846);
nor U14576 (N_14576,N_13694,N_13925);
nand U14577 (N_14577,N_13249,N_13521);
nor U14578 (N_14578,N_13291,N_13584);
nand U14579 (N_14579,N_13254,N_13936);
or U14580 (N_14580,N_13656,N_13417);
or U14581 (N_14581,N_13761,N_13185);
and U14582 (N_14582,N_13722,N_13408);
nor U14583 (N_14583,N_13501,N_13606);
nand U14584 (N_14584,N_13579,N_13263);
nand U14585 (N_14585,N_13533,N_13786);
or U14586 (N_14586,N_13289,N_13954);
or U14587 (N_14587,N_13272,N_13818);
or U14588 (N_14588,N_13414,N_13482);
nand U14589 (N_14589,N_13537,N_13179);
or U14590 (N_14590,N_13761,N_13942);
and U14591 (N_14591,N_13673,N_13327);
or U14592 (N_14592,N_13606,N_13926);
nor U14593 (N_14593,N_13250,N_13233);
and U14594 (N_14594,N_13703,N_13568);
or U14595 (N_14595,N_13447,N_13788);
and U14596 (N_14596,N_13205,N_13964);
nor U14597 (N_14597,N_13657,N_13790);
nor U14598 (N_14598,N_13139,N_13511);
nor U14599 (N_14599,N_13546,N_13884);
and U14600 (N_14600,N_13780,N_13363);
nor U14601 (N_14601,N_13475,N_13075);
or U14602 (N_14602,N_13928,N_13238);
nand U14603 (N_14603,N_13468,N_13973);
xnor U14604 (N_14604,N_13436,N_13518);
nor U14605 (N_14605,N_13413,N_13334);
and U14606 (N_14606,N_13054,N_13724);
or U14607 (N_14607,N_13168,N_13857);
or U14608 (N_14608,N_13250,N_13709);
xor U14609 (N_14609,N_13262,N_13487);
nand U14610 (N_14610,N_13207,N_13137);
xnor U14611 (N_14611,N_13208,N_13743);
nor U14612 (N_14612,N_13800,N_13266);
nand U14613 (N_14613,N_13015,N_13265);
or U14614 (N_14614,N_13995,N_13121);
nor U14615 (N_14615,N_13909,N_13822);
and U14616 (N_14616,N_13548,N_13204);
nor U14617 (N_14617,N_13159,N_13177);
nor U14618 (N_14618,N_13450,N_13182);
nor U14619 (N_14619,N_13471,N_13899);
xor U14620 (N_14620,N_13273,N_13071);
nor U14621 (N_14621,N_13297,N_13700);
nor U14622 (N_14622,N_13241,N_13433);
xnor U14623 (N_14623,N_13214,N_13640);
or U14624 (N_14624,N_13601,N_13272);
and U14625 (N_14625,N_13530,N_13589);
and U14626 (N_14626,N_13072,N_13842);
or U14627 (N_14627,N_13424,N_13236);
and U14628 (N_14628,N_13768,N_13733);
nand U14629 (N_14629,N_13620,N_13575);
nand U14630 (N_14630,N_13316,N_13068);
nor U14631 (N_14631,N_13796,N_13592);
or U14632 (N_14632,N_13848,N_13317);
xor U14633 (N_14633,N_13473,N_13841);
nand U14634 (N_14634,N_13943,N_13025);
nor U14635 (N_14635,N_13027,N_13171);
xnor U14636 (N_14636,N_13238,N_13686);
xnor U14637 (N_14637,N_13668,N_13244);
or U14638 (N_14638,N_13446,N_13417);
xor U14639 (N_14639,N_13617,N_13588);
nand U14640 (N_14640,N_13897,N_13935);
or U14641 (N_14641,N_13314,N_13033);
xnor U14642 (N_14642,N_13049,N_13956);
and U14643 (N_14643,N_13476,N_13549);
nand U14644 (N_14644,N_13202,N_13655);
nor U14645 (N_14645,N_13629,N_13416);
or U14646 (N_14646,N_13520,N_13263);
and U14647 (N_14647,N_13884,N_13028);
nand U14648 (N_14648,N_13103,N_13918);
nor U14649 (N_14649,N_13593,N_13617);
and U14650 (N_14650,N_13797,N_13725);
nor U14651 (N_14651,N_13038,N_13276);
and U14652 (N_14652,N_13880,N_13927);
nor U14653 (N_14653,N_13852,N_13099);
or U14654 (N_14654,N_13673,N_13433);
and U14655 (N_14655,N_13639,N_13320);
nand U14656 (N_14656,N_13800,N_13581);
and U14657 (N_14657,N_13550,N_13293);
nand U14658 (N_14658,N_13647,N_13139);
and U14659 (N_14659,N_13571,N_13019);
or U14660 (N_14660,N_13748,N_13946);
and U14661 (N_14661,N_13025,N_13380);
nor U14662 (N_14662,N_13058,N_13556);
nor U14663 (N_14663,N_13222,N_13729);
nand U14664 (N_14664,N_13098,N_13553);
nor U14665 (N_14665,N_13373,N_13555);
nor U14666 (N_14666,N_13336,N_13975);
xnor U14667 (N_14667,N_13945,N_13368);
or U14668 (N_14668,N_13292,N_13043);
xor U14669 (N_14669,N_13262,N_13219);
or U14670 (N_14670,N_13984,N_13655);
xor U14671 (N_14671,N_13997,N_13506);
and U14672 (N_14672,N_13523,N_13167);
nand U14673 (N_14673,N_13143,N_13221);
nor U14674 (N_14674,N_13631,N_13293);
xnor U14675 (N_14675,N_13420,N_13628);
nor U14676 (N_14676,N_13918,N_13552);
and U14677 (N_14677,N_13881,N_13730);
nand U14678 (N_14678,N_13217,N_13745);
and U14679 (N_14679,N_13541,N_13798);
nor U14680 (N_14680,N_13630,N_13806);
nor U14681 (N_14681,N_13114,N_13947);
or U14682 (N_14682,N_13824,N_13109);
and U14683 (N_14683,N_13772,N_13840);
or U14684 (N_14684,N_13490,N_13760);
and U14685 (N_14685,N_13400,N_13150);
xor U14686 (N_14686,N_13423,N_13564);
and U14687 (N_14687,N_13169,N_13832);
nor U14688 (N_14688,N_13795,N_13734);
and U14689 (N_14689,N_13440,N_13018);
and U14690 (N_14690,N_13789,N_13650);
or U14691 (N_14691,N_13778,N_13479);
nor U14692 (N_14692,N_13671,N_13787);
or U14693 (N_14693,N_13762,N_13405);
and U14694 (N_14694,N_13382,N_13690);
or U14695 (N_14695,N_13756,N_13759);
nor U14696 (N_14696,N_13663,N_13673);
nand U14697 (N_14697,N_13172,N_13813);
and U14698 (N_14698,N_13090,N_13544);
nand U14699 (N_14699,N_13365,N_13289);
nand U14700 (N_14700,N_13101,N_13994);
or U14701 (N_14701,N_13557,N_13492);
nand U14702 (N_14702,N_13378,N_13854);
xnor U14703 (N_14703,N_13651,N_13788);
xnor U14704 (N_14704,N_13965,N_13406);
nand U14705 (N_14705,N_13254,N_13835);
nor U14706 (N_14706,N_13492,N_13269);
and U14707 (N_14707,N_13925,N_13269);
nor U14708 (N_14708,N_13379,N_13713);
or U14709 (N_14709,N_13131,N_13708);
and U14710 (N_14710,N_13855,N_13505);
nand U14711 (N_14711,N_13431,N_13821);
and U14712 (N_14712,N_13024,N_13439);
nor U14713 (N_14713,N_13806,N_13438);
nor U14714 (N_14714,N_13046,N_13593);
and U14715 (N_14715,N_13992,N_13489);
nor U14716 (N_14716,N_13428,N_13767);
and U14717 (N_14717,N_13142,N_13890);
nand U14718 (N_14718,N_13383,N_13726);
nor U14719 (N_14719,N_13582,N_13065);
nand U14720 (N_14720,N_13848,N_13168);
xor U14721 (N_14721,N_13579,N_13808);
or U14722 (N_14722,N_13645,N_13298);
nand U14723 (N_14723,N_13447,N_13023);
xnor U14724 (N_14724,N_13344,N_13455);
or U14725 (N_14725,N_13203,N_13977);
or U14726 (N_14726,N_13003,N_13876);
or U14727 (N_14727,N_13871,N_13083);
nor U14728 (N_14728,N_13137,N_13227);
and U14729 (N_14729,N_13734,N_13181);
or U14730 (N_14730,N_13415,N_13401);
and U14731 (N_14731,N_13115,N_13552);
xnor U14732 (N_14732,N_13088,N_13399);
nor U14733 (N_14733,N_13582,N_13448);
nor U14734 (N_14734,N_13554,N_13267);
nor U14735 (N_14735,N_13171,N_13256);
xnor U14736 (N_14736,N_13259,N_13093);
and U14737 (N_14737,N_13804,N_13310);
and U14738 (N_14738,N_13985,N_13643);
or U14739 (N_14739,N_13628,N_13408);
or U14740 (N_14740,N_13704,N_13485);
or U14741 (N_14741,N_13930,N_13342);
and U14742 (N_14742,N_13966,N_13755);
nor U14743 (N_14743,N_13299,N_13428);
and U14744 (N_14744,N_13966,N_13370);
nor U14745 (N_14745,N_13544,N_13183);
nand U14746 (N_14746,N_13921,N_13103);
nand U14747 (N_14747,N_13672,N_13194);
and U14748 (N_14748,N_13776,N_13098);
nand U14749 (N_14749,N_13382,N_13464);
nand U14750 (N_14750,N_13988,N_13389);
nand U14751 (N_14751,N_13102,N_13028);
nor U14752 (N_14752,N_13385,N_13564);
and U14753 (N_14753,N_13561,N_13498);
or U14754 (N_14754,N_13478,N_13521);
xnor U14755 (N_14755,N_13767,N_13336);
and U14756 (N_14756,N_13517,N_13258);
nand U14757 (N_14757,N_13663,N_13953);
nor U14758 (N_14758,N_13173,N_13505);
nand U14759 (N_14759,N_13401,N_13782);
xor U14760 (N_14760,N_13773,N_13607);
nor U14761 (N_14761,N_13635,N_13320);
or U14762 (N_14762,N_13074,N_13566);
xnor U14763 (N_14763,N_13337,N_13884);
or U14764 (N_14764,N_13351,N_13751);
nand U14765 (N_14765,N_13164,N_13458);
nor U14766 (N_14766,N_13133,N_13810);
nand U14767 (N_14767,N_13877,N_13655);
or U14768 (N_14768,N_13064,N_13083);
xnor U14769 (N_14769,N_13968,N_13207);
nor U14770 (N_14770,N_13798,N_13468);
nor U14771 (N_14771,N_13457,N_13152);
or U14772 (N_14772,N_13215,N_13812);
nand U14773 (N_14773,N_13419,N_13977);
nand U14774 (N_14774,N_13269,N_13329);
and U14775 (N_14775,N_13246,N_13675);
nand U14776 (N_14776,N_13889,N_13985);
xor U14777 (N_14777,N_13142,N_13161);
or U14778 (N_14778,N_13952,N_13642);
and U14779 (N_14779,N_13231,N_13060);
xor U14780 (N_14780,N_13824,N_13831);
nand U14781 (N_14781,N_13420,N_13545);
and U14782 (N_14782,N_13477,N_13486);
nor U14783 (N_14783,N_13374,N_13020);
nand U14784 (N_14784,N_13637,N_13064);
or U14785 (N_14785,N_13854,N_13549);
and U14786 (N_14786,N_13537,N_13612);
nor U14787 (N_14787,N_13928,N_13891);
or U14788 (N_14788,N_13889,N_13860);
or U14789 (N_14789,N_13024,N_13484);
and U14790 (N_14790,N_13982,N_13019);
nand U14791 (N_14791,N_13674,N_13421);
or U14792 (N_14792,N_13705,N_13649);
or U14793 (N_14793,N_13793,N_13588);
and U14794 (N_14794,N_13349,N_13156);
nand U14795 (N_14795,N_13428,N_13199);
nand U14796 (N_14796,N_13209,N_13235);
nor U14797 (N_14797,N_13001,N_13627);
nand U14798 (N_14798,N_13657,N_13564);
xnor U14799 (N_14799,N_13673,N_13627);
nor U14800 (N_14800,N_13674,N_13048);
or U14801 (N_14801,N_13428,N_13156);
nand U14802 (N_14802,N_13825,N_13614);
nand U14803 (N_14803,N_13915,N_13694);
nand U14804 (N_14804,N_13893,N_13226);
nor U14805 (N_14805,N_13675,N_13336);
or U14806 (N_14806,N_13091,N_13931);
and U14807 (N_14807,N_13043,N_13093);
and U14808 (N_14808,N_13682,N_13468);
and U14809 (N_14809,N_13783,N_13995);
nand U14810 (N_14810,N_13852,N_13311);
nand U14811 (N_14811,N_13614,N_13666);
or U14812 (N_14812,N_13612,N_13369);
nand U14813 (N_14813,N_13586,N_13684);
nor U14814 (N_14814,N_13853,N_13454);
xor U14815 (N_14815,N_13111,N_13693);
nand U14816 (N_14816,N_13920,N_13098);
nand U14817 (N_14817,N_13922,N_13358);
and U14818 (N_14818,N_13273,N_13405);
nand U14819 (N_14819,N_13105,N_13499);
or U14820 (N_14820,N_13735,N_13337);
or U14821 (N_14821,N_13273,N_13641);
nand U14822 (N_14822,N_13552,N_13169);
nand U14823 (N_14823,N_13329,N_13142);
xnor U14824 (N_14824,N_13718,N_13198);
and U14825 (N_14825,N_13493,N_13634);
and U14826 (N_14826,N_13768,N_13694);
or U14827 (N_14827,N_13661,N_13501);
nand U14828 (N_14828,N_13233,N_13790);
nor U14829 (N_14829,N_13673,N_13405);
or U14830 (N_14830,N_13364,N_13357);
nand U14831 (N_14831,N_13670,N_13507);
and U14832 (N_14832,N_13921,N_13430);
and U14833 (N_14833,N_13439,N_13492);
and U14834 (N_14834,N_13943,N_13638);
nor U14835 (N_14835,N_13484,N_13154);
xor U14836 (N_14836,N_13936,N_13339);
nand U14837 (N_14837,N_13510,N_13051);
nand U14838 (N_14838,N_13532,N_13305);
and U14839 (N_14839,N_13504,N_13675);
nor U14840 (N_14840,N_13640,N_13873);
nand U14841 (N_14841,N_13682,N_13454);
and U14842 (N_14842,N_13639,N_13240);
nor U14843 (N_14843,N_13231,N_13011);
or U14844 (N_14844,N_13425,N_13482);
xor U14845 (N_14845,N_13170,N_13794);
or U14846 (N_14846,N_13046,N_13451);
nor U14847 (N_14847,N_13967,N_13740);
nor U14848 (N_14848,N_13331,N_13184);
and U14849 (N_14849,N_13392,N_13359);
or U14850 (N_14850,N_13057,N_13260);
xor U14851 (N_14851,N_13089,N_13060);
nand U14852 (N_14852,N_13181,N_13715);
or U14853 (N_14853,N_13285,N_13233);
or U14854 (N_14854,N_13395,N_13056);
nand U14855 (N_14855,N_13581,N_13240);
and U14856 (N_14856,N_13624,N_13845);
nand U14857 (N_14857,N_13608,N_13324);
or U14858 (N_14858,N_13193,N_13399);
and U14859 (N_14859,N_13542,N_13381);
nand U14860 (N_14860,N_13134,N_13080);
or U14861 (N_14861,N_13346,N_13771);
xor U14862 (N_14862,N_13307,N_13050);
and U14863 (N_14863,N_13582,N_13922);
xor U14864 (N_14864,N_13169,N_13831);
and U14865 (N_14865,N_13671,N_13094);
and U14866 (N_14866,N_13690,N_13679);
or U14867 (N_14867,N_13177,N_13179);
nand U14868 (N_14868,N_13387,N_13135);
or U14869 (N_14869,N_13910,N_13007);
or U14870 (N_14870,N_13583,N_13169);
or U14871 (N_14871,N_13481,N_13111);
or U14872 (N_14872,N_13380,N_13857);
nor U14873 (N_14873,N_13655,N_13875);
nand U14874 (N_14874,N_13432,N_13701);
or U14875 (N_14875,N_13790,N_13807);
nor U14876 (N_14876,N_13625,N_13000);
and U14877 (N_14877,N_13771,N_13307);
xnor U14878 (N_14878,N_13071,N_13574);
nor U14879 (N_14879,N_13867,N_13479);
nor U14880 (N_14880,N_13612,N_13506);
nor U14881 (N_14881,N_13334,N_13554);
nor U14882 (N_14882,N_13729,N_13337);
nand U14883 (N_14883,N_13844,N_13228);
nor U14884 (N_14884,N_13947,N_13829);
xnor U14885 (N_14885,N_13567,N_13271);
nor U14886 (N_14886,N_13741,N_13759);
nor U14887 (N_14887,N_13455,N_13152);
nand U14888 (N_14888,N_13213,N_13636);
or U14889 (N_14889,N_13102,N_13465);
and U14890 (N_14890,N_13826,N_13259);
or U14891 (N_14891,N_13101,N_13366);
nand U14892 (N_14892,N_13949,N_13009);
or U14893 (N_14893,N_13034,N_13641);
nor U14894 (N_14894,N_13634,N_13196);
or U14895 (N_14895,N_13835,N_13045);
nor U14896 (N_14896,N_13132,N_13898);
and U14897 (N_14897,N_13612,N_13349);
and U14898 (N_14898,N_13711,N_13543);
nor U14899 (N_14899,N_13786,N_13991);
or U14900 (N_14900,N_13553,N_13419);
nor U14901 (N_14901,N_13264,N_13268);
or U14902 (N_14902,N_13567,N_13391);
xor U14903 (N_14903,N_13711,N_13934);
nor U14904 (N_14904,N_13523,N_13531);
and U14905 (N_14905,N_13688,N_13059);
nand U14906 (N_14906,N_13438,N_13783);
nand U14907 (N_14907,N_13134,N_13122);
or U14908 (N_14908,N_13671,N_13298);
nand U14909 (N_14909,N_13311,N_13134);
nor U14910 (N_14910,N_13604,N_13863);
or U14911 (N_14911,N_13725,N_13165);
or U14912 (N_14912,N_13708,N_13539);
nand U14913 (N_14913,N_13681,N_13511);
and U14914 (N_14914,N_13699,N_13480);
or U14915 (N_14915,N_13034,N_13317);
nand U14916 (N_14916,N_13813,N_13360);
xor U14917 (N_14917,N_13139,N_13900);
or U14918 (N_14918,N_13033,N_13189);
or U14919 (N_14919,N_13522,N_13507);
xnor U14920 (N_14920,N_13277,N_13659);
or U14921 (N_14921,N_13817,N_13639);
nand U14922 (N_14922,N_13324,N_13988);
and U14923 (N_14923,N_13845,N_13927);
or U14924 (N_14924,N_13401,N_13709);
xor U14925 (N_14925,N_13244,N_13782);
and U14926 (N_14926,N_13624,N_13730);
and U14927 (N_14927,N_13186,N_13324);
xnor U14928 (N_14928,N_13768,N_13854);
or U14929 (N_14929,N_13524,N_13713);
nor U14930 (N_14930,N_13024,N_13588);
nor U14931 (N_14931,N_13526,N_13638);
nor U14932 (N_14932,N_13234,N_13273);
nor U14933 (N_14933,N_13059,N_13947);
nand U14934 (N_14934,N_13923,N_13329);
or U14935 (N_14935,N_13719,N_13294);
or U14936 (N_14936,N_13783,N_13947);
nand U14937 (N_14937,N_13713,N_13290);
nor U14938 (N_14938,N_13331,N_13550);
and U14939 (N_14939,N_13542,N_13663);
nand U14940 (N_14940,N_13349,N_13241);
or U14941 (N_14941,N_13789,N_13316);
nor U14942 (N_14942,N_13682,N_13501);
or U14943 (N_14943,N_13493,N_13975);
nor U14944 (N_14944,N_13427,N_13703);
or U14945 (N_14945,N_13238,N_13327);
nor U14946 (N_14946,N_13333,N_13233);
nor U14947 (N_14947,N_13283,N_13263);
nand U14948 (N_14948,N_13037,N_13364);
nand U14949 (N_14949,N_13339,N_13193);
and U14950 (N_14950,N_13037,N_13545);
and U14951 (N_14951,N_13015,N_13130);
and U14952 (N_14952,N_13081,N_13726);
nor U14953 (N_14953,N_13329,N_13451);
nand U14954 (N_14954,N_13374,N_13611);
xor U14955 (N_14955,N_13762,N_13269);
nor U14956 (N_14956,N_13106,N_13888);
or U14957 (N_14957,N_13284,N_13945);
or U14958 (N_14958,N_13812,N_13713);
and U14959 (N_14959,N_13474,N_13180);
and U14960 (N_14960,N_13751,N_13962);
and U14961 (N_14961,N_13931,N_13503);
xnor U14962 (N_14962,N_13048,N_13207);
nor U14963 (N_14963,N_13000,N_13534);
and U14964 (N_14964,N_13985,N_13684);
nor U14965 (N_14965,N_13910,N_13213);
nor U14966 (N_14966,N_13355,N_13901);
or U14967 (N_14967,N_13893,N_13840);
xnor U14968 (N_14968,N_13939,N_13908);
or U14969 (N_14969,N_13373,N_13372);
and U14970 (N_14970,N_13932,N_13685);
or U14971 (N_14971,N_13738,N_13511);
and U14972 (N_14972,N_13834,N_13528);
or U14973 (N_14973,N_13930,N_13179);
and U14974 (N_14974,N_13750,N_13952);
nor U14975 (N_14975,N_13663,N_13397);
or U14976 (N_14976,N_13010,N_13357);
and U14977 (N_14977,N_13922,N_13766);
nor U14978 (N_14978,N_13502,N_13820);
nand U14979 (N_14979,N_13674,N_13360);
and U14980 (N_14980,N_13961,N_13858);
nand U14981 (N_14981,N_13037,N_13060);
xnor U14982 (N_14982,N_13559,N_13717);
and U14983 (N_14983,N_13236,N_13912);
nand U14984 (N_14984,N_13573,N_13519);
or U14985 (N_14985,N_13980,N_13800);
or U14986 (N_14986,N_13531,N_13679);
or U14987 (N_14987,N_13750,N_13254);
nor U14988 (N_14988,N_13910,N_13870);
or U14989 (N_14989,N_13825,N_13441);
xnor U14990 (N_14990,N_13451,N_13842);
or U14991 (N_14991,N_13867,N_13459);
xor U14992 (N_14992,N_13950,N_13172);
nor U14993 (N_14993,N_13057,N_13062);
and U14994 (N_14994,N_13675,N_13313);
and U14995 (N_14995,N_13094,N_13844);
and U14996 (N_14996,N_13159,N_13421);
nand U14997 (N_14997,N_13212,N_13895);
and U14998 (N_14998,N_13081,N_13907);
and U14999 (N_14999,N_13285,N_13730);
or UO_0 (O_0,N_14188,N_14485);
xor UO_1 (O_1,N_14289,N_14488);
nor UO_2 (O_2,N_14463,N_14554);
and UO_3 (O_3,N_14281,N_14231);
or UO_4 (O_4,N_14001,N_14148);
and UO_5 (O_5,N_14610,N_14564);
or UO_6 (O_6,N_14867,N_14410);
xor UO_7 (O_7,N_14614,N_14743);
or UO_8 (O_8,N_14484,N_14780);
nand UO_9 (O_9,N_14057,N_14389);
and UO_10 (O_10,N_14322,N_14073);
and UO_11 (O_11,N_14327,N_14159);
nand UO_12 (O_12,N_14816,N_14293);
nor UO_13 (O_13,N_14225,N_14184);
nand UO_14 (O_14,N_14285,N_14502);
nor UO_15 (O_15,N_14622,N_14070);
nand UO_16 (O_16,N_14600,N_14124);
nand UO_17 (O_17,N_14556,N_14744);
nand UO_18 (O_18,N_14457,N_14911);
nor UO_19 (O_19,N_14863,N_14045);
nor UO_20 (O_20,N_14336,N_14062);
xnor UO_21 (O_21,N_14925,N_14658);
nand UO_22 (O_22,N_14015,N_14724);
and UO_23 (O_23,N_14802,N_14870);
and UO_24 (O_24,N_14982,N_14102);
and UO_25 (O_25,N_14803,N_14357);
or UO_26 (O_26,N_14604,N_14306);
nand UO_27 (O_27,N_14352,N_14694);
or UO_28 (O_28,N_14751,N_14790);
nand UO_29 (O_29,N_14893,N_14248);
nand UO_30 (O_30,N_14137,N_14493);
nor UO_31 (O_31,N_14123,N_14421);
xor UO_32 (O_32,N_14771,N_14512);
nor UO_33 (O_33,N_14508,N_14473);
nor UO_34 (O_34,N_14047,N_14196);
or UO_35 (O_35,N_14118,N_14858);
nand UO_36 (O_36,N_14317,N_14535);
xor UO_37 (O_37,N_14239,N_14301);
nand UO_38 (O_38,N_14179,N_14416);
and UO_39 (O_39,N_14194,N_14745);
nand UO_40 (O_40,N_14048,N_14868);
and UO_41 (O_41,N_14601,N_14243);
xor UO_42 (O_42,N_14752,N_14534);
and UO_43 (O_43,N_14789,N_14006);
nand UO_44 (O_44,N_14002,N_14312);
nor UO_45 (O_45,N_14656,N_14873);
nor UO_46 (O_46,N_14869,N_14795);
xnor UO_47 (O_47,N_14424,N_14400);
and UO_48 (O_48,N_14612,N_14326);
or UO_49 (O_49,N_14072,N_14517);
nand UO_50 (O_50,N_14447,N_14445);
or UO_51 (O_51,N_14372,N_14263);
nor UO_52 (O_52,N_14418,N_14584);
or UO_53 (O_53,N_14677,N_14081);
nor UO_54 (O_54,N_14528,N_14419);
and UO_55 (O_55,N_14334,N_14271);
xor UO_56 (O_56,N_14806,N_14230);
nand UO_57 (O_57,N_14210,N_14452);
and UO_58 (O_58,N_14609,N_14283);
xor UO_59 (O_59,N_14580,N_14432);
nor UO_60 (O_60,N_14759,N_14200);
and UO_61 (O_61,N_14232,N_14250);
nand UO_62 (O_62,N_14350,N_14822);
or UO_63 (O_63,N_14278,N_14178);
nor UO_64 (O_64,N_14549,N_14593);
xor UO_65 (O_65,N_14847,N_14059);
nand UO_66 (O_66,N_14020,N_14567);
xor UO_67 (O_67,N_14687,N_14074);
or UO_68 (O_68,N_14246,N_14937);
and UO_69 (O_69,N_14097,N_14638);
nand UO_70 (O_70,N_14646,N_14272);
or UO_71 (O_71,N_14568,N_14189);
nor UO_72 (O_72,N_14674,N_14037);
and UO_73 (O_73,N_14036,N_14799);
and UO_74 (O_74,N_14437,N_14163);
xor UO_75 (O_75,N_14865,N_14125);
or UO_76 (O_76,N_14122,N_14695);
nand UO_77 (O_77,N_14499,N_14726);
nor UO_78 (O_78,N_14224,N_14040);
nor UO_79 (O_79,N_14819,N_14676);
and UO_80 (O_80,N_14725,N_14960);
nor UO_81 (O_81,N_14815,N_14533);
nor UO_82 (O_82,N_14460,N_14854);
or UO_83 (O_83,N_14434,N_14689);
and UO_84 (O_84,N_14112,N_14891);
nor UO_85 (O_85,N_14089,N_14343);
and UO_86 (O_86,N_14041,N_14288);
and UO_87 (O_87,N_14558,N_14409);
xnor UO_88 (O_88,N_14441,N_14427);
nand UO_89 (O_89,N_14019,N_14055);
and UO_90 (O_90,N_14722,N_14207);
or UO_91 (O_91,N_14510,N_14860);
or UO_92 (O_92,N_14295,N_14141);
nand UO_93 (O_93,N_14364,N_14487);
nor UO_94 (O_94,N_14913,N_14561);
nor UO_95 (O_95,N_14856,N_14160);
nand UO_96 (O_96,N_14862,N_14618);
and UO_97 (O_97,N_14637,N_14536);
xnor UO_98 (O_98,N_14866,N_14713);
and UO_99 (O_99,N_14111,N_14500);
nor UO_100 (O_100,N_14165,N_14109);
or UO_101 (O_101,N_14589,N_14791);
and UO_102 (O_102,N_14634,N_14025);
nor UO_103 (O_103,N_14008,N_14588);
xnor UO_104 (O_104,N_14537,N_14208);
and UO_105 (O_105,N_14299,N_14974);
nand UO_106 (O_106,N_14607,N_14947);
xor UO_107 (O_107,N_14665,N_14261);
or UO_108 (O_108,N_14956,N_14628);
or UO_109 (O_109,N_14135,N_14832);
or UO_110 (O_110,N_14579,N_14693);
nor UO_111 (O_111,N_14023,N_14086);
nor UO_112 (O_112,N_14572,N_14716);
nand UO_113 (O_113,N_14879,N_14910);
or UO_114 (O_114,N_14117,N_14814);
nor UO_115 (O_115,N_14472,N_14895);
xor UO_116 (O_116,N_14375,N_14669);
and UO_117 (O_117,N_14800,N_14942);
xor UO_118 (O_118,N_14605,N_14335);
or UO_119 (O_119,N_14099,N_14912);
and UO_120 (O_120,N_14852,N_14798);
nand UO_121 (O_121,N_14769,N_14620);
xor UO_122 (O_122,N_14007,N_14110);
nor UO_123 (O_123,N_14642,N_14311);
or UO_124 (O_124,N_14741,N_14773);
or UO_125 (O_125,N_14162,N_14240);
nor UO_126 (O_126,N_14578,N_14962);
xnor UO_127 (O_127,N_14169,N_14010);
and UO_128 (O_128,N_14813,N_14943);
nor UO_129 (O_129,N_14843,N_14082);
nand UO_130 (O_130,N_14241,N_14191);
nand UO_131 (O_131,N_14166,N_14763);
nand UO_132 (O_132,N_14206,N_14571);
and UO_133 (O_133,N_14918,N_14906);
and UO_134 (O_134,N_14292,N_14919);
nand UO_135 (O_135,N_14058,N_14595);
and UO_136 (O_136,N_14318,N_14548);
nand UO_137 (O_137,N_14946,N_14202);
nor UO_138 (O_138,N_14654,N_14221);
xnor UO_139 (O_139,N_14147,N_14168);
or UO_140 (O_140,N_14750,N_14325);
nand UO_141 (O_141,N_14353,N_14466);
nand UO_142 (O_142,N_14399,N_14965);
nand UO_143 (O_143,N_14114,N_14126);
and UO_144 (O_144,N_14670,N_14190);
nor UO_145 (O_145,N_14371,N_14192);
nor UO_146 (O_146,N_14603,N_14107);
and UO_147 (O_147,N_14955,N_14778);
and UO_148 (O_148,N_14043,N_14762);
nor UO_149 (O_149,N_14249,N_14054);
or UO_150 (O_150,N_14345,N_14987);
nand UO_151 (O_151,N_14429,N_14131);
nor UO_152 (O_152,N_14155,N_14258);
xnor UO_153 (O_153,N_14134,N_14924);
nand UO_154 (O_154,N_14841,N_14018);
and UO_155 (O_155,N_14539,N_14707);
xor UO_156 (O_156,N_14631,N_14067);
xnor UO_157 (O_157,N_14753,N_14875);
or UO_158 (O_158,N_14804,N_14455);
xor UO_159 (O_159,N_14507,N_14296);
nand UO_160 (O_160,N_14935,N_14754);
nand UO_161 (O_161,N_14986,N_14775);
xor UO_162 (O_162,N_14187,N_14864);
nand UO_163 (O_163,N_14412,N_14063);
nand UO_164 (O_164,N_14586,N_14739);
and UO_165 (O_165,N_14084,N_14524);
or UO_166 (O_166,N_14254,N_14598);
nand UO_167 (O_167,N_14204,N_14997);
nand UO_168 (O_168,N_14384,N_14645);
nand UO_169 (O_169,N_14222,N_14801);
or UO_170 (O_170,N_14826,N_14330);
and UO_171 (O_171,N_14808,N_14520);
nand UO_172 (O_172,N_14308,N_14358);
nand UO_173 (O_173,N_14423,N_14228);
nor UO_174 (O_174,N_14276,N_14747);
nand UO_175 (O_175,N_14393,N_14303);
and UO_176 (O_176,N_14993,N_14104);
nor UO_177 (O_177,N_14378,N_14476);
xnor UO_178 (O_178,N_14181,N_14356);
nor UO_179 (O_179,N_14951,N_14321);
and UO_180 (O_180,N_14220,N_14142);
xor UO_181 (O_181,N_14623,N_14619);
and UO_182 (O_182,N_14782,N_14596);
nand UO_183 (O_183,N_14483,N_14590);
nor UO_184 (O_184,N_14274,N_14717);
and UO_185 (O_185,N_14602,N_14459);
nand UO_186 (O_186,N_14735,N_14643);
nand UO_187 (O_187,N_14840,N_14850);
or UO_188 (O_188,N_14709,N_14538);
xor UO_189 (O_189,N_14933,N_14736);
and UO_190 (O_190,N_14105,N_14298);
or UO_191 (O_191,N_14923,N_14662);
nor UO_192 (O_192,N_14329,N_14161);
and UO_193 (O_193,N_14121,N_14821);
or UO_194 (O_194,N_14103,N_14098);
or UO_195 (O_195,N_14839,N_14708);
and UO_196 (O_196,N_14733,N_14038);
and UO_197 (O_197,N_14650,N_14518);
or UO_198 (O_198,N_14738,N_14881);
nor UO_199 (O_199,N_14742,N_14851);
or UO_200 (O_200,N_14907,N_14899);
or UO_201 (O_201,N_14992,N_14000);
and UO_202 (O_202,N_14053,N_14252);
and UO_203 (O_203,N_14390,N_14562);
or UO_204 (O_204,N_14414,N_14932);
or UO_205 (O_205,N_14976,N_14448);
and UO_206 (O_206,N_14217,N_14316);
xnor UO_207 (O_207,N_14758,N_14044);
nor UO_208 (O_208,N_14730,N_14969);
or UO_209 (O_209,N_14836,N_14146);
nor UO_210 (O_210,N_14787,N_14201);
and UO_211 (O_211,N_14545,N_14442);
or UO_212 (O_212,N_14017,N_14376);
nor UO_213 (O_213,N_14282,N_14158);
or UO_214 (O_214,N_14226,N_14973);
or UO_215 (O_215,N_14195,N_14908);
nand UO_216 (O_216,N_14127,N_14715);
or UO_217 (O_217,N_14952,N_14964);
and UO_218 (O_218,N_14939,N_14757);
or UO_219 (O_219,N_14917,N_14264);
or UO_220 (O_220,N_14324,N_14233);
and UO_221 (O_221,N_14209,N_14591);
nand UO_222 (O_222,N_14404,N_14692);
and UO_223 (O_223,N_14016,N_14894);
nor UO_224 (O_224,N_14766,N_14003);
nor UO_225 (O_225,N_14031,N_14422);
or UO_226 (O_226,N_14544,N_14765);
nor UO_227 (O_227,N_14632,N_14608);
nor UO_228 (O_228,N_14234,N_14411);
nand UO_229 (O_229,N_14185,N_14443);
or UO_230 (O_230,N_14990,N_14838);
and UO_231 (O_231,N_14830,N_14113);
nor UO_232 (O_232,N_14844,N_14344);
and UO_233 (O_233,N_14855,N_14461);
or UO_234 (O_234,N_14262,N_14706);
xor UO_235 (O_235,N_14033,N_14013);
nand UO_236 (O_236,N_14648,N_14872);
and UO_237 (O_237,N_14468,N_14898);
and UO_238 (O_238,N_14582,N_14565);
xor UO_239 (O_239,N_14647,N_14085);
and UO_240 (O_240,N_14480,N_14398);
and UO_241 (O_241,N_14164,N_14705);
nand UO_242 (O_242,N_14700,N_14569);
or UO_243 (O_243,N_14391,N_14383);
nor UO_244 (O_244,N_14996,N_14630);
nand UO_245 (O_245,N_14551,N_14878);
or UO_246 (O_246,N_14408,N_14106);
and UO_247 (O_247,N_14433,N_14767);
or UO_248 (O_248,N_14219,N_14402);
nor UO_249 (O_249,N_14686,N_14810);
nand UO_250 (O_250,N_14711,N_14088);
or UO_251 (O_251,N_14489,N_14080);
or UO_252 (O_252,N_14175,N_14892);
and UO_253 (O_253,N_14351,N_14474);
or UO_254 (O_254,N_14368,N_14774);
or UO_255 (O_255,N_14890,N_14138);
and UO_256 (O_256,N_14842,N_14144);
nand UO_257 (O_257,N_14557,N_14347);
or UO_258 (O_258,N_14186,N_14024);
nor UO_259 (O_259,N_14959,N_14833);
nand UO_260 (O_260,N_14180,N_14145);
xor UO_261 (O_261,N_14575,N_14793);
or UO_262 (O_262,N_14256,N_14245);
nor UO_263 (O_263,N_14691,N_14363);
nand UO_264 (O_264,N_14022,N_14011);
nand UO_265 (O_265,N_14922,N_14928);
nor UO_266 (O_266,N_14837,N_14994);
nor UO_267 (O_267,N_14170,N_14749);
or UO_268 (O_268,N_14305,N_14269);
nand UO_269 (O_269,N_14215,N_14218);
nand UO_270 (O_270,N_14497,N_14673);
xor UO_271 (O_271,N_14672,N_14587);
xor UO_272 (O_272,N_14685,N_14555);
and UO_273 (O_273,N_14783,N_14119);
nor UO_274 (O_274,N_14541,N_14889);
xor UO_275 (O_275,N_14639,N_14005);
or UO_276 (O_276,N_14611,N_14482);
nor UO_277 (O_277,N_14259,N_14794);
nor UO_278 (O_278,N_14491,N_14966);
or UO_279 (O_279,N_14475,N_14511);
and UO_280 (O_280,N_14060,N_14133);
xor UO_281 (O_281,N_14174,N_14069);
xor UO_282 (O_282,N_14392,N_14236);
nor UO_283 (O_283,N_14379,N_14214);
nor UO_284 (O_284,N_14247,N_14129);
nor UO_285 (O_285,N_14989,N_14313);
xnor UO_286 (O_286,N_14576,N_14944);
and UO_287 (O_287,N_14167,N_14823);
xor UO_288 (O_288,N_14012,N_14380);
or UO_289 (O_289,N_14506,N_14941);
or UO_290 (O_290,N_14636,N_14359);
nor UO_291 (O_291,N_14300,N_14728);
nand UO_292 (O_292,N_14029,N_14065);
and UO_293 (O_293,N_14199,N_14051);
nand UO_294 (O_294,N_14177,N_14406);
nand UO_295 (O_295,N_14405,N_14828);
or UO_296 (O_296,N_14616,N_14690);
nand UO_297 (O_297,N_14504,N_14776);
nand UO_298 (O_298,N_14337,N_14035);
nor UO_299 (O_299,N_14958,N_14294);
and UO_300 (O_300,N_14042,N_14710);
nand UO_301 (O_301,N_14615,N_14286);
xor UO_302 (O_302,N_14530,N_14428);
nor UO_303 (O_303,N_14902,N_14915);
nand UO_304 (O_304,N_14513,N_14644);
nand UO_305 (O_305,N_14640,N_14394);
or UO_306 (O_306,N_14501,N_14831);
or UO_307 (O_307,N_14349,N_14339);
and UO_308 (O_308,N_14755,N_14370);
nor UO_309 (O_309,N_14523,N_14027);
xor UO_310 (O_310,N_14760,N_14087);
nor UO_311 (O_311,N_14157,N_14515);
nor UO_312 (O_312,N_14154,N_14213);
xnor UO_313 (O_313,N_14028,N_14546);
nor UO_314 (O_314,N_14657,N_14302);
nor UO_315 (O_315,N_14718,N_14101);
nand UO_316 (O_316,N_14279,N_14046);
nand UO_317 (O_317,N_14792,N_14980);
nand UO_318 (O_318,N_14521,N_14328);
or UO_319 (O_319,N_14439,N_14514);
or UO_320 (O_320,N_14066,N_14784);
and UO_321 (O_321,N_14977,N_14469);
or UO_322 (O_322,N_14857,N_14998);
or UO_323 (O_323,N_14205,N_14624);
or UO_324 (O_324,N_14663,N_14203);
nor UO_325 (O_325,N_14467,N_14477);
nor UO_326 (O_326,N_14516,N_14307);
or UO_327 (O_327,N_14212,N_14887);
nor UO_328 (O_328,N_14679,N_14756);
and UO_329 (O_329,N_14785,N_14449);
and UO_330 (O_330,N_14734,N_14635);
xnor UO_331 (O_331,N_14583,N_14094);
nor UO_332 (O_332,N_14934,N_14348);
or UO_333 (O_333,N_14874,N_14182);
nor UO_334 (O_334,N_14342,N_14291);
nand UO_335 (O_335,N_14978,N_14970);
nor UO_336 (O_336,N_14540,N_14988);
nor UO_337 (O_337,N_14267,N_14824);
nand UO_338 (O_338,N_14573,N_14975);
xor UO_339 (O_339,N_14967,N_14809);
nand UO_340 (O_340,N_14495,N_14304);
and UO_341 (O_341,N_14396,N_14323);
and UO_342 (O_342,N_14369,N_14438);
nor UO_343 (O_343,N_14426,N_14825);
nand UO_344 (O_344,N_14667,N_14971);
nand UO_345 (O_345,N_14255,N_14772);
xor UO_346 (O_346,N_14770,N_14340);
or UO_347 (O_347,N_14139,N_14446);
or UO_348 (O_348,N_14812,N_14381);
or UO_349 (O_349,N_14731,N_14309);
xor UO_350 (O_350,N_14963,N_14366);
nor UO_351 (O_351,N_14173,N_14004);
nand UO_352 (O_352,N_14211,N_14697);
nand UO_353 (O_353,N_14197,N_14244);
nor UO_354 (O_354,N_14542,N_14968);
or UO_355 (O_355,N_14021,N_14931);
xnor UO_356 (O_356,N_14039,N_14559);
and UO_357 (O_357,N_14786,N_14130);
xor UO_358 (O_358,N_14817,N_14712);
nand UO_359 (O_359,N_14574,N_14684);
and UO_360 (O_360,N_14362,N_14076);
nor UO_361 (O_361,N_14532,N_14140);
or UO_362 (O_362,N_14310,N_14949);
or UO_363 (O_363,N_14714,N_14617);
and UO_364 (O_364,N_14257,N_14268);
nor UO_365 (O_365,N_14183,N_14884);
nand UO_366 (O_366,N_14284,N_14985);
or UO_367 (O_367,N_14599,N_14355);
and UO_368 (O_368,N_14651,N_14275);
and UO_369 (O_369,N_14664,N_14503);
nor UO_370 (O_370,N_14655,N_14885);
and UO_371 (O_371,N_14277,N_14095);
nor UO_372 (O_372,N_14176,N_14732);
and UO_373 (O_373,N_14903,N_14699);
and UO_374 (O_374,N_14083,N_14827);
nand UO_375 (O_375,N_14904,N_14120);
or UO_376 (O_376,N_14314,N_14888);
or UO_377 (O_377,N_14216,N_14387);
nand UO_378 (O_378,N_14068,N_14936);
and UO_379 (O_379,N_14818,N_14957);
nand UO_380 (O_380,N_14064,N_14981);
or UO_381 (O_381,N_14811,N_14729);
xnor UO_382 (O_382,N_14519,N_14242);
or UO_383 (O_383,N_14481,N_14435);
and UO_384 (O_384,N_14365,N_14382);
nand UO_385 (O_385,N_14845,N_14633);
nand UO_386 (O_386,N_14566,N_14346);
and UO_387 (O_387,N_14149,N_14153);
xor UO_388 (O_388,N_14338,N_14577);
nor UO_389 (O_389,N_14652,N_14462);
or UO_390 (O_390,N_14543,N_14471);
and UO_391 (O_391,N_14594,N_14407);
and UO_392 (O_392,N_14075,N_14625);
nor UO_393 (O_393,N_14172,N_14032);
nor UO_394 (O_394,N_14152,N_14675);
or UO_395 (O_395,N_14505,N_14496);
nor UO_396 (O_396,N_14876,N_14397);
nor UO_397 (O_397,N_14198,N_14265);
and UO_398 (O_398,N_14948,N_14108);
nand UO_399 (O_399,N_14034,N_14287);
or UO_400 (O_400,N_14882,N_14090);
nand UO_401 (O_401,N_14470,N_14420);
nand UO_402 (O_402,N_14796,N_14401);
nand UO_403 (O_403,N_14367,N_14229);
and UO_404 (O_404,N_14266,N_14629);
nor UO_405 (O_405,N_14659,N_14115);
and UO_406 (O_406,N_14683,N_14227);
nor UO_407 (O_407,N_14509,N_14374);
and UO_408 (O_408,N_14768,N_14954);
or UO_409 (O_409,N_14486,N_14553);
and UO_410 (O_410,N_14388,N_14078);
xnor UO_411 (O_411,N_14332,N_14171);
nand UO_412 (O_412,N_14193,N_14896);
and UO_413 (O_413,N_14999,N_14525);
and UO_414 (O_414,N_14585,N_14280);
nor UO_415 (O_415,N_14143,N_14333);
xor UO_416 (O_416,N_14661,N_14490);
and UO_417 (O_417,N_14748,N_14597);
and UO_418 (O_418,N_14492,N_14498);
and UO_419 (O_419,N_14260,N_14270);
nand UO_420 (O_420,N_14052,N_14829);
or UO_421 (O_421,N_14315,N_14805);
and UO_422 (O_422,N_14440,N_14720);
or UO_423 (O_423,N_14849,N_14871);
nor UO_424 (O_424,N_14238,N_14395);
and UO_425 (O_425,N_14253,N_14853);
nand UO_426 (O_426,N_14660,N_14938);
nand UO_427 (O_427,N_14386,N_14702);
or UO_428 (O_428,N_14071,N_14235);
and UO_429 (O_429,N_14444,N_14682);
and UO_430 (O_430,N_14050,N_14450);
and UO_431 (O_431,N_14251,N_14746);
and UO_432 (O_432,N_14927,N_14547);
or UO_433 (O_433,N_14570,N_14914);
nor UO_434 (O_434,N_14764,N_14136);
nand UO_435 (O_435,N_14464,N_14984);
nand UO_436 (O_436,N_14385,N_14897);
or UO_437 (O_437,N_14678,N_14413);
and UO_438 (O_438,N_14649,N_14861);
xor UO_439 (O_439,N_14417,N_14454);
and UO_440 (O_440,N_14688,N_14527);
and UO_441 (O_441,N_14877,N_14696);
or UO_442 (O_442,N_14560,N_14737);
nand UO_443 (O_443,N_14727,N_14883);
nor UO_444 (O_444,N_14950,N_14009);
nand UO_445 (O_445,N_14132,N_14671);
xor UO_446 (O_446,N_14431,N_14797);
or UO_447 (O_447,N_14983,N_14848);
nand UO_448 (O_448,N_14719,N_14100);
nor UO_449 (O_449,N_14613,N_14320);
or UO_450 (O_450,N_14930,N_14479);
and UO_451 (O_451,N_14953,N_14704);
nor UO_452 (O_452,N_14451,N_14621);
nand UO_453 (O_453,N_14526,N_14698);
and UO_454 (O_454,N_14297,N_14550);
nor UO_455 (O_455,N_14237,N_14092);
nand UO_456 (O_456,N_14360,N_14781);
nor UO_457 (O_457,N_14331,N_14151);
and UO_458 (O_458,N_14886,N_14835);
nor UO_459 (O_459,N_14606,N_14079);
xnor UO_460 (O_460,N_14478,N_14415);
or UO_461 (O_461,N_14995,N_14156);
and UO_462 (O_462,N_14723,N_14880);
and UO_463 (O_463,N_14453,N_14425);
and UO_464 (O_464,N_14859,N_14056);
or UO_465 (O_465,N_14680,N_14093);
and UO_466 (O_466,N_14456,N_14740);
nand UO_467 (O_467,N_14701,N_14552);
nand UO_468 (O_468,N_14779,N_14014);
and UO_469 (O_469,N_14026,N_14721);
nand UO_470 (O_470,N_14049,N_14077);
nor UO_471 (O_471,N_14091,N_14531);
or UO_472 (O_472,N_14436,N_14929);
or UO_473 (O_473,N_14581,N_14666);
nor UO_474 (O_474,N_14529,N_14592);
and UO_475 (O_475,N_14223,N_14373);
and UO_476 (O_476,N_14909,N_14641);
or UO_477 (O_477,N_14150,N_14920);
and UO_478 (O_478,N_14627,N_14777);
nor UO_479 (O_479,N_14653,N_14458);
nand UO_480 (O_480,N_14945,N_14403);
or UO_481 (O_481,N_14926,N_14061);
nand UO_482 (O_482,N_14626,N_14377);
nand UO_483 (O_483,N_14921,N_14494);
nand UO_484 (O_484,N_14681,N_14788);
nand UO_485 (O_485,N_14807,N_14991);
and UO_486 (O_486,N_14761,N_14834);
or UO_487 (O_487,N_14128,N_14273);
nor UO_488 (O_488,N_14940,N_14905);
and UO_489 (O_489,N_14703,N_14979);
and UO_490 (O_490,N_14972,N_14901);
xor UO_491 (O_491,N_14961,N_14341);
and UO_492 (O_492,N_14030,N_14430);
and UO_493 (O_493,N_14465,N_14361);
or UO_494 (O_494,N_14522,N_14096);
and UO_495 (O_495,N_14668,N_14820);
nor UO_496 (O_496,N_14290,N_14846);
nor UO_497 (O_497,N_14354,N_14916);
xor UO_498 (O_498,N_14563,N_14900);
nor UO_499 (O_499,N_14116,N_14319);
nor UO_500 (O_500,N_14577,N_14432);
nor UO_501 (O_501,N_14923,N_14888);
or UO_502 (O_502,N_14024,N_14068);
and UO_503 (O_503,N_14990,N_14517);
and UO_504 (O_504,N_14657,N_14168);
and UO_505 (O_505,N_14268,N_14653);
or UO_506 (O_506,N_14231,N_14705);
xnor UO_507 (O_507,N_14229,N_14141);
or UO_508 (O_508,N_14716,N_14374);
nor UO_509 (O_509,N_14718,N_14154);
nand UO_510 (O_510,N_14559,N_14131);
nor UO_511 (O_511,N_14379,N_14182);
and UO_512 (O_512,N_14019,N_14160);
nor UO_513 (O_513,N_14167,N_14602);
and UO_514 (O_514,N_14781,N_14994);
nor UO_515 (O_515,N_14941,N_14257);
or UO_516 (O_516,N_14105,N_14627);
nor UO_517 (O_517,N_14633,N_14812);
nor UO_518 (O_518,N_14984,N_14923);
and UO_519 (O_519,N_14830,N_14945);
and UO_520 (O_520,N_14377,N_14050);
or UO_521 (O_521,N_14677,N_14781);
xnor UO_522 (O_522,N_14389,N_14136);
xor UO_523 (O_523,N_14815,N_14192);
or UO_524 (O_524,N_14379,N_14645);
nor UO_525 (O_525,N_14913,N_14355);
nand UO_526 (O_526,N_14803,N_14861);
and UO_527 (O_527,N_14362,N_14574);
and UO_528 (O_528,N_14717,N_14791);
nand UO_529 (O_529,N_14456,N_14402);
and UO_530 (O_530,N_14583,N_14782);
nor UO_531 (O_531,N_14311,N_14926);
nand UO_532 (O_532,N_14103,N_14449);
xor UO_533 (O_533,N_14236,N_14038);
nor UO_534 (O_534,N_14909,N_14348);
nand UO_535 (O_535,N_14849,N_14416);
and UO_536 (O_536,N_14903,N_14416);
xor UO_537 (O_537,N_14566,N_14109);
and UO_538 (O_538,N_14468,N_14710);
or UO_539 (O_539,N_14562,N_14998);
nand UO_540 (O_540,N_14476,N_14978);
and UO_541 (O_541,N_14722,N_14533);
and UO_542 (O_542,N_14870,N_14893);
or UO_543 (O_543,N_14335,N_14867);
or UO_544 (O_544,N_14838,N_14806);
or UO_545 (O_545,N_14835,N_14583);
or UO_546 (O_546,N_14479,N_14967);
nand UO_547 (O_547,N_14825,N_14161);
nand UO_548 (O_548,N_14976,N_14650);
or UO_549 (O_549,N_14047,N_14106);
nand UO_550 (O_550,N_14582,N_14986);
and UO_551 (O_551,N_14029,N_14090);
nor UO_552 (O_552,N_14248,N_14797);
and UO_553 (O_553,N_14961,N_14044);
nand UO_554 (O_554,N_14823,N_14944);
and UO_555 (O_555,N_14652,N_14724);
nand UO_556 (O_556,N_14302,N_14901);
and UO_557 (O_557,N_14041,N_14268);
or UO_558 (O_558,N_14043,N_14401);
or UO_559 (O_559,N_14677,N_14760);
nor UO_560 (O_560,N_14722,N_14284);
and UO_561 (O_561,N_14435,N_14404);
xnor UO_562 (O_562,N_14423,N_14763);
xor UO_563 (O_563,N_14725,N_14601);
nand UO_564 (O_564,N_14122,N_14262);
and UO_565 (O_565,N_14904,N_14040);
or UO_566 (O_566,N_14412,N_14489);
or UO_567 (O_567,N_14135,N_14355);
nand UO_568 (O_568,N_14928,N_14033);
and UO_569 (O_569,N_14360,N_14975);
nor UO_570 (O_570,N_14841,N_14399);
nor UO_571 (O_571,N_14188,N_14469);
or UO_572 (O_572,N_14930,N_14465);
nand UO_573 (O_573,N_14833,N_14885);
xor UO_574 (O_574,N_14956,N_14974);
or UO_575 (O_575,N_14758,N_14309);
nor UO_576 (O_576,N_14325,N_14475);
nand UO_577 (O_577,N_14836,N_14305);
nand UO_578 (O_578,N_14401,N_14682);
xor UO_579 (O_579,N_14668,N_14773);
nand UO_580 (O_580,N_14611,N_14322);
or UO_581 (O_581,N_14413,N_14786);
and UO_582 (O_582,N_14550,N_14236);
nand UO_583 (O_583,N_14576,N_14152);
and UO_584 (O_584,N_14232,N_14580);
xnor UO_585 (O_585,N_14101,N_14421);
nand UO_586 (O_586,N_14948,N_14087);
and UO_587 (O_587,N_14651,N_14328);
xor UO_588 (O_588,N_14769,N_14167);
or UO_589 (O_589,N_14620,N_14578);
nand UO_590 (O_590,N_14894,N_14994);
or UO_591 (O_591,N_14253,N_14611);
or UO_592 (O_592,N_14259,N_14927);
xnor UO_593 (O_593,N_14338,N_14238);
nand UO_594 (O_594,N_14578,N_14386);
and UO_595 (O_595,N_14448,N_14614);
xnor UO_596 (O_596,N_14939,N_14698);
xor UO_597 (O_597,N_14741,N_14364);
xnor UO_598 (O_598,N_14644,N_14279);
nand UO_599 (O_599,N_14596,N_14389);
and UO_600 (O_600,N_14820,N_14930);
nand UO_601 (O_601,N_14559,N_14602);
or UO_602 (O_602,N_14410,N_14291);
and UO_603 (O_603,N_14634,N_14846);
nor UO_604 (O_604,N_14802,N_14954);
nor UO_605 (O_605,N_14018,N_14809);
nor UO_606 (O_606,N_14982,N_14033);
and UO_607 (O_607,N_14764,N_14896);
or UO_608 (O_608,N_14183,N_14727);
or UO_609 (O_609,N_14048,N_14217);
nand UO_610 (O_610,N_14404,N_14554);
nand UO_611 (O_611,N_14636,N_14429);
nor UO_612 (O_612,N_14317,N_14834);
nand UO_613 (O_613,N_14273,N_14884);
nand UO_614 (O_614,N_14115,N_14475);
and UO_615 (O_615,N_14320,N_14191);
nor UO_616 (O_616,N_14369,N_14373);
nand UO_617 (O_617,N_14573,N_14742);
xor UO_618 (O_618,N_14110,N_14244);
and UO_619 (O_619,N_14277,N_14876);
or UO_620 (O_620,N_14275,N_14599);
or UO_621 (O_621,N_14106,N_14962);
or UO_622 (O_622,N_14719,N_14043);
and UO_623 (O_623,N_14905,N_14080);
nor UO_624 (O_624,N_14890,N_14233);
and UO_625 (O_625,N_14409,N_14090);
nor UO_626 (O_626,N_14715,N_14233);
nand UO_627 (O_627,N_14254,N_14287);
nand UO_628 (O_628,N_14217,N_14448);
or UO_629 (O_629,N_14196,N_14401);
nor UO_630 (O_630,N_14751,N_14632);
or UO_631 (O_631,N_14989,N_14150);
or UO_632 (O_632,N_14059,N_14781);
nor UO_633 (O_633,N_14332,N_14818);
and UO_634 (O_634,N_14968,N_14002);
or UO_635 (O_635,N_14175,N_14252);
nor UO_636 (O_636,N_14316,N_14080);
nand UO_637 (O_637,N_14363,N_14419);
nor UO_638 (O_638,N_14081,N_14378);
nor UO_639 (O_639,N_14270,N_14859);
nand UO_640 (O_640,N_14026,N_14032);
xor UO_641 (O_641,N_14428,N_14274);
or UO_642 (O_642,N_14762,N_14115);
nor UO_643 (O_643,N_14900,N_14019);
and UO_644 (O_644,N_14113,N_14597);
and UO_645 (O_645,N_14944,N_14443);
or UO_646 (O_646,N_14975,N_14033);
nand UO_647 (O_647,N_14178,N_14645);
nand UO_648 (O_648,N_14208,N_14412);
or UO_649 (O_649,N_14232,N_14944);
and UO_650 (O_650,N_14886,N_14126);
nand UO_651 (O_651,N_14196,N_14353);
xnor UO_652 (O_652,N_14604,N_14014);
and UO_653 (O_653,N_14615,N_14551);
nand UO_654 (O_654,N_14847,N_14619);
nand UO_655 (O_655,N_14747,N_14436);
nor UO_656 (O_656,N_14910,N_14794);
xor UO_657 (O_657,N_14968,N_14108);
xnor UO_658 (O_658,N_14559,N_14458);
or UO_659 (O_659,N_14463,N_14515);
nor UO_660 (O_660,N_14182,N_14895);
nor UO_661 (O_661,N_14026,N_14010);
nor UO_662 (O_662,N_14121,N_14966);
or UO_663 (O_663,N_14680,N_14157);
nor UO_664 (O_664,N_14780,N_14071);
xnor UO_665 (O_665,N_14835,N_14049);
or UO_666 (O_666,N_14310,N_14551);
nor UO_667 (O_667,N_14051,N_14097);
or UO_668 (O_668,N_14082,N_14756);
nor UO_669 (O_669,N_14588,N_14340);
xor UO_670 (O_670,N_14119,N_14160);
nand UO_671 (O_671,N_14448,N_14638);
or UO_672 (O_672,N_14584,N_14083);
xnor UO_673 (O_673,N_14059,N_14658);
xor UO_674 (O_674,N_14163,N_14400);
and UO_675 (O_675,N_14144,N_14832);
nand UO_676 (O_676,N_14043,N_14874);
or UO_677 (O_677,N_14955,N_14630);
and UO_678 (O_678,N_14440,N_14675);
xor UO_679 (O_679,N_14889,N_14574);
and UO_680 (O_680,N_14372,N_14317);
and UO_681 (O_681,N_14473,N_14526);
nand UO_682 (O_682,N_14170,N_14309);
nand UO_683 (O_683,N_14967,N_14368);
and UO_684 (O_684,N_14621,N_14244);
and UO_685 (O_685,N_14439,N_14254);
and UO_686 (O_686,N_14304,N_14411);
nor UO_687 (O_687,N_14695,N_14768);
or UO_688 (O_688,N_14432,N_14635);
or UO_689 (O_689,N_14354,N_14052);
nor UO_690 (O_690,N_14590,N_14024);
and UO_691 (O_691,N_14221,N_14894);
nor UO_692 (O_692,N_14464,N_14524);
or UO_693 (O_693,N_14727,N_14327);
and UO_694 (O_694,N_14372,N_14347);
nand UO_695 (O_695,N_14861,N_14348);
nor UO_696 (O_696,N_14822,N_14123);
and UO_697 (O_697,N_14593,N_14883);
and UO_698 (O_698,N_14439,N_14923);
nor UO_699 (O_699,N_14080,N_14601);
and UO_700 (O_700,N_14083,N_14911);
and UO_701 (O_701,N_14235,N_14026);
nor UO_702 (O_702,N_14494,N_14255);
and UO_703 (O_703,N_14490,N_14298);
nor UO_704 (O_704,N_14222,N_14427);
and UO_705 (O_705,N_14985,N_14719);
and UO_706 (O_706,N_14657,N_14054);
or UO_707 (O_707,N_14332,N_14704);
and UO_708 (O_708,N_14040,N_14612);
and UO_709 (O_709,N_14944,N_14855);
and UO_710 (O_710,N_14773,N_14757);
nand UO_711 (O_711,N_14083,N_14327);
nor UO_712 (O_712,N_14738,N_14426);
nor UO_713 (O_713,N_14695,N_14216);
nand UO_714 (O_714,N_14818,N_14780);
or UO_715 (O_715,N_14750,N_14308);
and UO_716 (O_716,N_14348,N_14807);
nor UO_717 (O_717,N_14164,N_14994);
or UO_718 (O_718,N_14142,N_14017);
nand UO_719 (O_719,N_14492,N_14572);
xnor UO_720 (O_720,N_14676,N_14807);
nor UO_721 (O_721,N_14690,N_14685);
nand UO_722 (O_722,N_14662,N_14515);
nor UO_723 (O_723,N_14096,N_14821);
nand UO_724 (O_724,N_14391,N_14673);
and UO_725 (O_725,N_14799,N_14181);
or UO_726 (O_726,N_14355,N_14021);
nor UO_727 (O_727,N_14926,N_14485);
or UO_728 (O_728,N_14976,N_14614);
or UO_729 (O_729,N_14773,N_14402);
nand UO_730 (O_730,N_14945,N_14710);
xnor UO_731 (O_731,N_14508,N_14061);
or UO_732 (O_732,N_14018,N_14693);
xor UO_733 (O_733,N_14506,N_14545);
nand UO_734 (O_734,N_14969,N_14799);
nand UO_735 (O_735,N_14742,N_14891);
xor UO_736 (O_736,N_14925,N_14991);
nor UO_737 (O_737,N_14561,N_14315);
or UO_738 (O_738,N_14575,N_14239);
and UO_739 (O_739,N_14576,N_14733);
and UO_740 (O_740,N_14259,N_14659);
nor UO_741 (O_741,N_14480,N_14374);
or UO_742 (O_742,N_14992,N_14362);
nor UO_743 (O_743,N_14114,N_14043);
or UO_744 (O_744,N_14253,N_14617);
nand UO_745 (O_745,N_14939,N_14213);
and UO_746 (O_746,N_14377,N_14152);
nand UO_747 (O_747,N_14415,N_14286);
nor UO_748 (O_748,N_14668,N_14771);
nand UO_749 (O_749,N_14080,N_14197);
nor UO_750 (O_750,N_14980,N_14465);
and UO_751 (O_751,N_14582,N_14812);
nand UO_752 (O_752,N_14803,N_14128);
and UO_753 (O_753,N_14946,N_14655);
xnor UO_754 (O_754,N_14230,N_14665);
and UO_755 (O_755,N_14016,N_14606);
nor UO_756 (O_756,N_14648,N_14843);
nor UO_757 (O_757,N_14159,N_14146);
xnor UO_758 (O_758,N_14799,N_14877);
and UO_759 (O_759,N_14980,N_14550);
nor UO_760 (O_760,N_14691,N_14561);
nor UO_761 (O_761,N_14048,N_14179);
nand UO_762 (O_762,N_14806,N_14599);
nand UO_763 (O_763,N_14018,N_14878);
or UO_764 (O_764,N_14568,N_14056);
nor UO_765 (O_765,N_14447,N_14443);
or UO_766 (O_766,N_14446,N_14902);
or UO_767 (O_767,N_14051,N_14670);
nand UO_768 (O_768,N_14424,N_14463);
and UO_769 (O_769,N_14311,N_14110);
and UO_770 (O_770,N_14069,N_14619);
and UO_771 (O_771,N_14464,N_14958);
nand UO_772 (O_772,N_14097,N_14171);
nand UO_773 (O_773,N_14407,N_14785);
nand UO_774 (O_774,N_14173,N_14035);
nor UO_775 (O_775,N_14818,N_14966);
and UO_776 (O_776,N_14617,N_14277);
nor UO_777 (O_777,N_14134,N_14732);
or UO_778 (O_778,N_14309,N_14133);
and UO_779 (O_779,N_14058,N_14800);
and UO_780 (O_780,N_14602,N_14223);
nor UO_781 (O_781,N_14490,N_14043);
or UO_782 (O_782,N_14348,N_14541);
nand UO_783 (O_783,N_14218,N_14295);
nor UO_784 (O_784,N_14691,N_14744);
and UO_785 (O_785,N_14937,N_14605);
nor UO_786 (O_786,N_14106,N_14246);
nand UO_787 (O_787,N_14428,N_14810);
nand UO_788 (O_788,N_14412,N_14580);
nand UO_789 (O_789,N_14329,N_14847);
and UO_790 (O_790,N_14048,N_14663);
and UO_791 (O_791,N_14787,N_14673);
nand UO_792 (O_792,N_14540,N_14602);
nor UO_793 (O_793,N_14749,N_14340);
and UO_794 (O_794,N_14272,N_14170);
xnor UO_795 (O_795,N_14286,N_14896);
nor UO_796 (O_796,N_14178,N_14173);
nor UO_797 (O_797,N_14561,N_14082);
and UO_798 (O_798,N_14465,N_14756);
nor UO_799 (O_799,N_14353,N_14773);
nand UO_800 (O_800,N_14427,N_14595);
nand UO_801 (O_801,N_14563,N_14390);
nor UO_802 (O_802,N_14425,N_14011);
xor UO_803 (O_803,N_14234,N_14603);
nor UO_804 (O_804,N_14192,N_14200);
nor UO_805 (O_805,N_14845,N_14866);
nand UO_806 (O_806,N_14760,N_14804);
or UO_807 (O_807,N_14751,N_14062);
nor UO_808 (O_808,N_14107,N_14691);
nor UO_809 (O_809,N_14582,N_14789);
and UO_810 (O_810,N_14412,N_14374);
or UO_811 (O_811,N_14293,N_14907);
nand UO_812 (O_812,N_14661,N_14778);
nand UO_813 (O_813,N_14501,N_14880);
nor UO_814 (O_814,N_14538,N_14738);
and UO_815 (O_815,N_14849,N_14012);
or UO_816 (O_816,N_14297,N_14116);
and UO_817 (O_817,N_14905,N_14748);
or UO_818 (O_818,N_14137,N_14696);
nand UO_819 (O_819,N_14140,N_14344);
or UO_820 (O_820,N_14578,N_14429);
nand UO_821 (O_821,N_14538,N_14596);
or UO_822 (O_822,N_14795,N_14344);
and UO_823 (O_823,N_14431,N_14172);
and UO_824 (O_824,N_14980,N_14304);
xnor UO_825 (O_825,N_14472,N_14570);
nand UO_826 (O_826,N_14841,N_14393);
and UO_827 (O_827,N_14955,N_14425);
or UO_828 (O_828,N_14081,N_14355);
nand UO_829 (O_829,N_14280,N_14323);
and UO_830 (O_830,N_14529,N_14215);
nor UO_831 (O_831,N_14791,N_14491);
or UO_832 (O_832,N_14506,N_14516);
xor UO_833 (O_833,N_14602,N_14677);
or UO_834 (O_834,N_14655,N_14217);
or UO_835 (O_835,N_14240,N_14582);
nand UO_836 (O_836,N_14252,N_14096);
or UO_837 (O_837,N_14534,N_14887);
and UO_838 (O_838,N_14996,N_14093);
nor UO_839 (O_839,N_14504,N_14016);
nor UO_840 (O_840,N_14381,N_14239);
xor UO_841 (O_841,N_14840,N_14340);
and UO_842 (O_842,N_14760,N_14868);
nand UO_843 (O_843,N_14302,N_14289);
nand UO_844 (O_844,N_14505,N_14039);
nor UO_845 (O_845,N_14240,N_14170);
nand UO_846 (O_846,N_14227,N_14257);
nand UO_847 (O_847,N_14276,N_14380);
or UO_848 (O_848,N_14454,N_14182);
xnor UO_849 (O_849,N_14307,N_14440);
nor UO_850 (O_850,N_14556,N_14673);
nand UO_851 (O_851,N_14392,N_14707);
nand UO_852 (O_852,N_14845,N_14640);
or UO_853 (O_853,N_14350,N_14739);
nand UO_854 (O_854,N_14233,N_14520);
nand UO_855 (O_855,N_14689,N_14955);
nand UO_856 (O_856,N_14235,N_14369);
xor UO_857 (O_857,N_14955,N_14319);
or UO_858 (O_858,N_14356,N_14211);
or UO_859 (O_859,N_14214,N_14253);
and UO_860 (O_860,N_14193,N_14926);
or UO_861 (O_861,N_14493,N_14679);
xor UO_862 (O_862,N_14596,N_14453);
xor UO_863 (O_863,N_14346,N_14432);
and UO_864 (O_864,N_14067,N_14194);
nand UO_865 (O_865,N_14042,N_14865);
and UO_866 (O_866,N_14503,N_14403);
nand UO_867 (O_867,N_14189,N_14049);
and UO_868 (O_868,N_14675,N_14749);
nand UO_869 (O_869,N_14561,N_14593);
or UO_870 (O_870,N_14524,N_14818);
xor UO_871 (O_871,N_14578,N_14400);
or UO_872 (O_872,N_14729,N_14227);
and UO_873 (O_873,N_14424,N_14818);
nor UO_874 (O_874,N_14855,N_14008);
nor UO_875 (O_875,N_14716,N_14189);
or UO_876 (O_876,N_14952,N_14096);
or UO_877 (O_877,N_14021,N_14944);
nor UO_878 (O_878,N_14455,N_14387);
or UO_879 (O_879,N_14086,N_14750);
nand UO_880 (O_880,N_14298,N_14169);
or UO_881 (O_881,N_14735,N_14032);
nor UO_882 (O_882,N_14361,N_14059);
nor UO_883 (O_883,N_14627,N_14662);
nor UO_884 (O_884,N_14603,N_14192);
or UO_885 (O_885,N_14796,N_14239);
nor UO_886 (O_886,N_14756,N_14416);
and UO_887 (O_887,N_14487,N_14322);
or UO_888 (O_888,N_14672,N_14004);
xnor UO_889 (O_889,N_14133,N_14172);
nor UO_890 (O_890,N_14187,N_14545);
nand UO_891 (O_891,N_14048,N_14746);
or UO_892 (O_892,N_14725,N_14714);
nor UO_893 (O_893,N_14218,N_14153);
nor UO_894 (O_894,N_14602,N_14646);
xnor UO_895 (O_895,N_14152,N_14663);
or UO_896 (O_896,N_14428,N_14500);
or UO_897 (O_897,N_14966,N_14679);
nor UO_898 (O_898,N_14517,N_14322);
and UO_899 (O_899,N_14691,N_14846);
or UO_900 (O_900,N_14961,N_14893);
or UO_901 (O_901,N_14614,N_14517);
or UO_902 (O_902,N_14135,N_14091);
nand UO_903 (O_903,N_14730,N_14344);
and UO_904 (O_904,N_14295,N_14758);
nand UO_905 (O_905,N_14827,N_14389);
or UO_906 (O_906,N_14942,N_14559);
nor UO_907 (O_907,N_14459,N_14187);
or UO_908 (O_908,N_14782,N_14806);
nor UO_909 (O_909,N_14207,N_14083);
and UO_910 (O_910,N_14630,N_14336);
nor UO_911 (O_911,N_14760,N_14628);
and UO_912 (O_912,N_14800,N_14420);
nor UO_913 (O_913,N_14333,N_14927);
nor UO_914 (O_914,N_14562,N_14169);
nor UO_915 (O_915,N_14953,N_14991);
nor UO_916 (O_916,N_14942,N_14490);
and UO_917 (O_917,N_14250,N_14341);
or UO_918 (O_918,N_14865,N_14964);
nand UO_919 (O_919,N_14004,N_14308);
and UO_920 (O_920,N_14203,N_14830);
nor UO_921 (O_921,N_14158,N_14504);
nor UO_922 (O_922,N_14256,N_14234);
or UO_923 (O_923,N_14037,N_14694);
nor UO_924 (O_924,N_14230,N_14590);
nor UO_925 (O_925,N_14725,N_14177);
or UO_926 (O_926,N_14253,N_14505);
or UO_927 (O_927,N_14303,N_14235);
or UO_928 (O_928,N_14195,N_14574);
and UO_929 (O_929,N_14937,N_14614);
and UO_930 (O_930,N_14032,N_14751);
nor UO_931 (O_931,N_14247,N_14490);
and UO_932 (O_932,N_14264,N_14929);
and UO_933 (O_933,N_14016,N_14896);
nand UO_934 (O_934,N_14497,N_14821);
and UO_935 (O_935,N_14206,N_14234);
and UO_936 (O_936,N_14503,N_14278);
nor UO_937 (O_937,N_14043,N_14788);
and UO_938 (O_938,N_14522,N_14573);
or UO_939 (O_939,N_14980,N_14166);
nand UO_940 (O_940,N_14302,N_14644);
or UO_941 (O_941,N_14629,N_14093);
or UO_942 (O_942,N_14499,N_14476);
or UO_943 (O_943,N_14829,N_14137);
or UO_944 (O_944,N_14754,N_14316);
and UO_945 (O_945,N_14467,N_14921);
and UO_946 (O_946,N_14252,N_14904);
and UO_947 (O_947,N_14177,N_14450);
xnor UO_948 (O_948,N_14350,N_14633);
or UO_949 (O_949,N_14527,N_14691);
nand UO_950 (O_950,N_14557,N_14822);
and UO_951 (O_951,N_14589,N_14179);
and UO_952 (O_952,N_14727,N_14470);
or UO_953 (O_953,N_14737,N_14644);
and UO_954 (O_954,N_14071,N_14339);
and UO_955 (O_955,N_14638,N_14252);
or UO_956 (O_956,N_14645,N_14561);
nor UO_957 (O_957,N_14386,N_14676);
nand UO_958 (O_958,N_14509,N_14015);
or UO_959 (O_959,N_14531,N_14757);
nor UO_960 (O_960,N_14859,N_14022);
nand UO_961 (O_961,N_14139,N_14362);
or UO_962 (O_962,N_14980,N_14612);
nor UO_963 (O_963,N_14481,N_14492);
and UO_964 (O_964,N_14157,N_14698);
or UO_965 (O_965,N_14217,N_14452);
nand UO_966 (O_966,N_14106,N_14982);
or UO_967 (O_967,N_14044,N_14294);
xnor UO_968 (O_968,N_14623,N_14157);
and UO_969 (O_969,N_14152,N_14939);
or UO_970 (O_970,N_14871,N_14391);
or UO_971 (O_971,N_14962,N_14453);
xor UO_972 (O_972,N_14029,N_14354);
nand UO_973 (O_973,N_14338,N_14098);
nor UO_974 (O_974,N_14731,N_14082);
nor UO_975 (O_975,N_14980,N_14250);
nor UO_976 (O_976,N_14654,N_14943);
xor UO_977 (O_977,N_14895,N_14752);
xor UO_978 (O_978,N_14258,N_14014);
nand UO_979 (O_979,N_14951,N_14778);
and UO_980 (O_980,N_14908,N_14939);
nor UO_981 (O_981,N_14522,N_14798);
and UO_982 (O_982,N_14209,N_14235);
nand UO_983 (O_983,N_14512,N_14946);
nand UO_984 (O_984,N_14095,N_14480);
or UO_985 (O_985,N_14283,N_14491);
or UO_986 (O_986,N_14564,N_14752);
or UO_987 (O_987,N_14317,N_14376);
or UO_988 (O_988,N_14740,N_14566);
xor UO_989 (O_989,N_14756,N_14202);
and UO_990 (O_990,N_14116,N_14163);
nand UO_991 (O_991,N_14224,N_14340);
or UO_992 (O_992,N_14133,N_14664);
and UO_993 (O_993,N_14928,N_14337);
and UO_994 (O_994,N_14013,N_14130);
and UO_995 (O_995,N_14467,N_14918);
nand UO_996 (O_996,N_14630,N_14750);
or UO_997 (O_997,N_14464,N_14255);
xnor UO_998 (O_998,N_14283,N_14592);
or UO_999 (O_999,N_14243,N_14810);
nand UO_1000 (O_1000,N_14638,N_14224);
or UO_1001 (O_1001,N_14339,N_14520);
xor UO_1002 (O_1002,N_14481,N_14731);
xnor UO_1003 (O_1003,N_14754,N_14508);
nor UO_1004 (O_1004,N_14409,N_14337);
nand UO_1005 (O_1005,N_14219,N_14966);
nor UO_1006 (O_1006,N_14068,N_14373);
nand UO_1007 (O_1007,N_14034,N_14187);
or UO_1008 (O_1008,N_14362,N_14689);
nor UO_1009 (O_1009,N_14767,N_14357);
and UO_1010 (O_1010,N_14676,N_14613);
nor UO_1011 (O_1011,N_14305,N_14915);
or UO_1012 (O_1012,N_14535,N_14507);
nand UO_1013 (O_1013,N_14689,N_14718);
nand UO_1014 (O_1014,N_14127,N_14392);
nand UO_1015 (O_1015,N_14916,N_14306);
and UO_1016 (O_1016,N_14021,N_14357);
and UO_1017 (O_1017,N_14152,N_14534);
or UO_1018 (O_1018,N_14688,N_14746);
nand UO_1019 (O_1019,N_14786,N_14004);
or UO_1020 (O_1020,N_14698,N_14142);
or UO_1021 (O_1021,N_14982,N_14230);
nand UO_1022 (O_1022,N_14150,N_14915);
nand UO_1023 (O_1023,N_14499,N_14897);
nand UO_1024 (O_1024,N_14408,N_14739);
nor UO_1025 (O_1025,N_14791,N_14129);
nand UO_1026 (O_1026,N_14125,N_14475);
nor UO_1027 (O_1027,N_14671,N_14944);
nand UO_1028 (O_1028,N_14566,N_14269);
nor UO_1029 (O_1029,N_14805,N_14244);
or UO_1030 (O_1030,N_14349,N_14933);
nand UO_1031 (O_1031,N_14870,N_14170);
nor UO_1032 (O_1032,N_14511,N_14150);
nand UO_1033 (O_1033,N_14108,N_14701);
nand UO_1034 (O_1034,N_14467,N_14393);
xnor UO_1035 (O_1035,N_14712,N_14979);
nor UO_1036 (O_1036,N_14923,N_14530);
nor UO_1037 (O_1037,N_14408,N_14098);
or UO_1038 (O_1038,N_14283,N_14424);
nand UO_1039 (O_1039,N_14753,N_14218);
nor UO_1040 (O_1040,N_14752,N_14504);
xor UO_1041 (O_1041,N_14852,N_14609);
nand UO_1042 (O_1042,N_14103,N_14495);
nand UO_1043 (O_1043,N_14881,N_14687);
and UO_1044 (O_1044,N_14879,N_14061);
or UO_1045 (O_1045,N_14879,N_14213);
nor UO_1046 (O_1046,N_14244,N_14489);
or UO_1047 (O_1047,N_14536,N_14005);
or UO_1048 (O_1048,N_14536,N_14643);
nor UO_1049 (O_1049,N_14283,N_14299);
and UO_1050 (O_1050,N_14117,N_14412);
and UO_1051 (O_1051,N_14896,N_14418);
nor UO_1052 (O_1052,N_14534,N_14289);
or UO_1053 (O_1053,N_14674,N_14366);
nor UO_1054 (O_1054,N_14086,N_14709);
nor UO_1055 (O_1055,N_14376,N_14299);
nand UO_1056 (O_1056,N_14210,N_14480);
nand UO_1057 (O_1057,N_14729,N_14221);
and UO_1058 (O_1058,N_14451,N_14917);
and UO_1059 (O_1059,N_14753,N_14565);
or UO_1060 (O_1060,N_14566,N_14963);
or UO_1061 (O_1061,N_14702,N_14115);
nand UO_1062 (O_1062,N_14168,N_14776);
and UO_1063 (O_1063,N_14041,N_14461);
xnor UO_1064 (O_1064,N_14035,N_14540);
xor UO_1065 (O_1065,N_14661,N_14726);
and UO_1066 (O_1066,N_14293,N_14446);
xor UO_1067 (O_1067,N_14565,N_14646);
nor UO_1068 (O_1068,N_14958,N_14363);
nor UO_1069 (O_1069,N_14710,N_14454);
and UO_1070 (O_1070,N_14464,N_14587);
nand UO_1071 (O_1071,N_14495,N_14362);
or UO_1072 (O_1072,N_14846,N_14355);
or UO_1073 (O_1073,N_14905,N_14344);
nor UO_1074 (O_1074,N_14541,N_14229);
and UO_1075 (O_1075,N_14844,N_14783);
or UO_1076 (O_1076,N_14415,N_14324);
and UO_1077 (O_1077,N_14428,N_14738);
nand UO_1078 (O_1078,N_14949,N_14626);
and UO_1079 (O_1079,N_14918,N_14322);
nor UO_1080 (O_1080,N_14861,N_14334);
nand UO_1081 (O_1081,N_14555,N_14947);
and UO_1082 (O_1082,N_14209,N_14983);
nand UO_1083 (O_1083,N_14477,N_14960);
and UO_1084 (O_1084,N_14923,N_14910);
nor UO_1085 (O_1085,N_14884,N_14558);
nor UO_1086 (O_1086,N_14373,N_14334);
and UO_1087 (O_1087,N_14719,N_14702);
nor UO_1088 (O_1088,N_14406,N_14380);
nand UO_1089 (O_1089,N_14920,N_14697);
xnor UO_1090 (O_1090,N_14197,N_14100);
or UO_1091 (O_1091,N_14096,N_14966);
nor UO_1092 (O_1092,N_14885,N_14323);
nor UO_1093 (O_1093,N_14451,N_14295);
or UO_1094 (O_1094,N_14310,N_14169);
or UO_1095 (O_1095,N_14682,N_14761);
or UO_1096 (O_1096,N_14968,N_14008);
or UO_1097 (O_1097,N_14457,N_14170);
and UO_1098 (O_1098,N_14121,N_14979);
nor UO_1099 (O_1099,N_14511,N_14711);
or UO_1100 (O_1100,N_14537,N_14412);
and UO_1101 (O_1101,N_14930,N_14642);
or UO_1102 (O_1102,N_14454,N_14452);
and UO_1103 (O_1103,N_14799,N_14892);
or UO_1104 (O_1104,N_14706,N_14732);
nor UO_1105 (O_1105,N_14379,N_14262);
or UO_1106 (O_1106,N_14966,N_14456);
and UO_1107 (O_1107,N_14966,N_14710);
or UO_1108 (O_1108,N_14529,N_14422);
nand UO_1109 (O_1109,N_14261,N_14385);
and UO_1110 (O_1110,N_14127,N_14135);
nor UO_1111 (O_1111,N_14903,N_14295);
or UO_1112 (O_1112,N_14767,N_14652);
nand UO_1113 (O_1113,N_14624,N_14130);
nand UO_1114 (O_1114,N_14327,N_14268);
xnor UO_1115 (O_1115,N_14809,N_14411);
nand UO_1116 (O_1116,N_14491,N_14853);
and UO_1117 (O_1117,N_14536,N_14811);
or UO_1118 (O_1118,N_14230,N_14221);
or UO_1119 (O_1119,N_14596,N_14941);
nor UO_1120 (O_1120,N_14325,N_14247);
and UO_1121 (O_1121,N_14095,N_14979);
xor UO_1122 (O_1122,N_14055,N_14525);
or UO_1123 (O_1123,N_14396,N_14516);
nor UO_1124 (O_1124,N_14323,N_14423);
or UO_1125 (O_1125,N_14360,N_14248);
and UO_1126 (O_1126,N_14674,N_14730);
or UO_1127 (O_1127,N_14958,N_14635);
nor UO_1128 (O_1128,N_14586,N_14079);
nand UO_1129 (O_1129,N_14361,N_14328);
nand UO_1130 (O_1130,N_14945,N_14749);
and UO_1131 (O_1131,N_14276,N_14255);
nand UO_1132 (O_1132,N_14685,N_14416);
xnor UO_1133 (O_1133,N_14219,N_14496);
nand UO_1134 (O_1134,N_14600,N_14742);
and UO_1135 (O_1135,N_14278,N_14392);
nor UO_1136 (O_1136,N_14658,N_14688);
or UO_1137 (O_1137,N_14353,N_14048);
and UO_1138 (O_1138,N_14610,N_14669);
and UO_1139 (O_1139,N_14613,N_14102);
nor UO_1140 (O_1140,N_14790,N_14687);
xor UO_1141 (O_1141,N_14875,N_14561);
nand UO_1142 (O_1142,N_14619,N_14881);
nor UO_1143 (O_1143,N_14589,N_14919);
nand UO_1144 (O_1144,N_14902,N_14296);
nand UO_1145 (O_1145,N_14069,N_14207);
or UO_1146 (O_1146,N_14992,N_14043);
nand UO_1147 (O_1147,N_14394,N_14197);
nor UO_1148 (O_1148,N_14869,N_14633);
nand UO_1149 (O_1149,N_14873,N_14821);
nand UO_1150 (O_1150,N_14407,N_14576);
nor UO_1151 (O_1151,N_14824,N_14488);
and UO_1152 (O_1152,N_14040,N_14937);
and UO_1153 (O_1153,N_14758,N_14372);
or UO_1154 (O_1154,N_14870,N_14733);
nor UO_1155 (O_1155,N_14682,N_14216);
xor UO_1156 (O_1156,N_14768,N_14654);
and UO_1157 (O_1157,N_14279,N_14291);
nor UO_1158 (O_1158,N_14486,N_14795);
and UO_1159 (O_1159,N_14879,N_14918);
nand UO_1160 (O_1160,N_14214,N_14070);
and UO_1161 (O_1161,N_14276,N_14830);
and UO_1162 (O_1162,N_14501,N_14533);
nor UO_1163 (O_1163,N_14904,N_14404);
and UO_1164 (O_1164,N_14004,N_14031);
xnor UO_1165 (O_1165,N_14449,N_14853);
and UO_1166 (O_1166,N_14518,N_14170);
nor UO_1167 (O_1167,N_14870,N_14403);
or UO_1168 (O_1168,N_14328,N_14915);
and UO_1169 (O_1169,N_14764,N_14278);
and UO_1170 (O_1170,N_14548,N_14992);
or UO_1171 (O_1171,N_14689,N_14628);
or UO_1172 (O_1172,N_14003,N_14602);
nand UO_1173 (O_1173,N_14984,N_14926);
and UO_1174 (O_1174,N_14404,N_14245);
nand UO_1175 (O_1175,N_14041,N_14031);
nor UO_1176 (O_1176,N_14413,N_14265);
nand UO_1177 (O_1177,N_14210,N_14643);
xor UO_1178 (O_1178,N_14178,N_14550);
nor UO_1179 (O_1179,N_14143,N_14036);
nor UO_1180 (O_1180,N_14662,N_14697);
nand UO_1181 (O_1181,N_14720,N_14288);
nor UO_1182 (O_1182,N_14824,N_14116);
nand UO_1183 (O_1183,N_14172,N_14489);
nor UO_1184 (O_1184,N_14314,N_14171);
nand UO_1185 (O_1185,N_14388,N_14334);
and UO_1186 (O_1186,N_14463,N_14410);
or UO_1187 (O_1187,N_14946,N_14230);
and UO_1188 (O_1188,N_14500,N_14185);
nor UO_1189 (O_1189,N_14101,N_14696);
xnor UO_1190 (O_1190,N_14319,N_14901);
nor UO_1191 (O_1191,N_14910,N_14216);
nand UO_1192 (O_1192,N_14957,N_14017);
and UO_1193 (O_1193,N_14380,N_14839);
and UO_1194 (O_1194,N_14006,N_14435);
or UO_1195 (O_1195,N_14955,N_14320);
and UO_1196 (O_1196,N_14682,N_14139);
or UO_1197 (O_1197,N_14880,N_14607);
xor UO_1198 (O_1198,N_14525,N_14449);
nand UO_1199 (O_1199,N_14770,N_14837);
xnor UO_1200 (O_1200,N_14622,N_14649);
nand UO_1201 (O_1201,N_14571,N_14647);
or UO_1202 (O_1202,N_14436,N_14785);
nand UO_1203 (O_1203,N_14864,N_14926);
xor UO_1204 (O_1204,N_14610,N_14684);
nand UO_1205 (O_1205,N_14098,N_14471);
xor UO_1206 (O_1206,N_14603,N_14469);
or UO_1207 (O_1207,N_14357,N_14667);
nor UO_1208 (O_1208,N_14465,N_14737);
and UO_1209 (O_1209,N_14213,N_14010);
nand UO_1210 (O_1210,N_14873,N_14295);
or UO_1211 (O_1211,N_14195,N_14734);
and UO_1212 (O_1212,N_14796,N_14691);
or UO_1213 (O_1213,N_14808,N_14860);
nor UO_1214 (O_1214,N_14739,N_14194);
or UO_1215 (O_1215,N_14140,N_14198);
xnor UO_1216 (O_1216,N_14393,N_14523);
and UO_1217 (O_1217,N_14574,N_14886);
and UO_1218 (O_1218,N_14165,N_14271);
nor UO_1219 (O_1219,N_14753,N_14665);
or UO_1220 (O_1220,N_14530,N_14319);
xnor UO_1221 (O_1221,N_14831,N_14631);
nand UO_1222 (O_1222,N_14163,N_14160);
nand UO_1223 (O_1223,N_14365,N_14066);
nand UO_1224 (O_1224,N_14199,N_14863);
xnor UO_1225 (O_1225,N_14054,N_14749);
nor UO_1226 (O_1226,N_14522,N_14156);
or UO_1227 (O_1227,N_14070,N_14511);
xor UO_1228 (O_1228,N_14768,N_14076);
and UO_1229 (O_1229,N_14739,N_14217);
nand UO_1230 (O_1230,N_14661,N_14520);
nand UO_1231 (O_1231,N_14619,N_14457);
and UO_1232 (O_1232,N_14743,N_14896);
xnor UO_1233 (O_1233,N_14414,N_14905);
nor UO_1234 (O_1234,N_14288,N_14110);
or UO_1235 (O_1235,N_14107,N_14466);
nand UO_1236 (O_1236,N_14051,N_14396);
or UO_1237 (O_1237,N_14447,N_14369);
or UO_1238 (O_1238,N_14929,N_14395);
xnor UO_1239 (O_1239,N_14590,N_14753);
nor UO_1240 (O_1240,N_14240,N_14522);
or UO_1241 (O_1241,N_14554,N_14025);
nand UO_1242 (O_1242,N_14708,N_14419);
nand UO_1243 (O_1243,N_14664,N_14900);
and UO_1244 (O_1244,N_14265,N_14087);
nand UO_1245 (O_1245,N_14503,N_14516);
and UO_1246 (O_1246,N_14803,N_14898);
and UO_1247 (O_1247,N_14684,N_14409);
nor UO_1248 (O_1248,N_14633,N_14374);
nor UO_1249 (O_1249,N_14766,N_14660);
nand UO_1250 (O_1250,N_14386,N_14525);
xnor UO_1251 (O_1251,N_14375,N_14659);
nand UO_1252 (O_1252,N_14112,N_14901);
nand UO_1253 (O_1253,N_14687,N_14871);
nand UO_1254 (O_1254,N_14489,N_14792);
nand UO_1255 (O_1255,N_14864,N_14821);
nand UO_1256 (O_1256,N_14176,N_14226);
xnor UO_1257 (O_1257,N_14693,N_14921);
xor UO_1258 (O_1258,N_14115,N_14024);
nor UO_1259 (O_1259,N_14921,N_14040);
xnor UO_1260 (O_1260,N_14807,N_14504);
nand UO_1261 (O_1261,N_14630,N_14405);
nand UO_1262 (O_1262,N_14739,N_14069);
or UO_1263 (O_1263,N_14432,N_14599);
or UO_1264 (O_1264,N_14252,N_14422);
or UO_1265 (O_1265,N_14026,N_14167);
nand UO_1266 (O_1266,N_14415,N_14338);
nor UO_1267 (O_1267,N_14899,N_14055);
or UO_1268 (O_1268,N_14828,N_14818);
nor UO_1269 (O_1269,N_14662,N_14122);
or UO_1270 (O_1270,N_14524,N_14394);
or UO_1271 (O_1271,N_14706,N_14962);
nor UO_1272 (O_1272,N_14186,N_14010);
nand UO_1273 (O_1273,N_14312,N_14195);
and UO_1274 (O_1274,N_14953,N_14596);
nor UO_1275 (O_1275,N_14787,N_14461);
nand UO_1276 (O_1276,N_14086,N_14857);
nand UO_1277 (O_1277,N_14157,N_14996);
or UO_1278 (O_1278,N_14753,N_14620);
or UO_1279 (O_1279,N_14484,N_14797);
nor UO_1280 (O_1280,N_14619,N_14915);
xor UO_1281 (O_1281,N_14165,N_14558);
or UO_1282 (O_1282,N_14077,N_14324);
nand UO_1283 (O_1283,N_14459,N_14305);
and UO_1284 (O_1284,N_14539,N_14234);
nand UO_1285 (O_1285,N_14785,N_14290);
nand UO_1286 (O_1286,N_14850,N_14004);
or UO_1287 (O_1287,N_14367,N_14250);
nand UO_1288 (O_1288,N_14276,N_14956);
xnor UO_1289 (O_1289,N_14307,N_14269);
and UO_1290 (O_1290,N_14261,N_14275);
and UO_1291 (O_1291,N_14241,N_14233);
or UO_1292 (O_1292,N_14477,N_14433);
nor UO_1293 (O_1293,N_14844,N_14853);
or UO_1294 (O_1294,N_14974,N_14479);
and UO_1295 (O_1295,N_14249,N_14371);
or UO_1296 (O_1296,N_14024,N_14032);
xor UO_1297 (O_1297,N_14963,N_14753);
and UO_1298 (O_1298,N_14120,N_14155);
and UO_1299 (O_1299,N_14707,N_14489);
nor UO_1300 (O_1300,N_14955,N_14642);
nand UO_1301 (O_1301,N_14065,N_14069);
nor UO_1302 (O_1302,N_14872,N_14215);
and UO_1303 (O_1303,N_14257,N_14730);
or UO_1304 (O_1304,N_14977,N_14978);
or UO_1305 (O_1305,N_14271,N_14333);
or UO_1306 (O_1306,N_14917,N_14888);
nand UO_1307 (O_1307,N_14613,N_14507);
and UO_1308 (O_1308,N_14598,N_14373);
nand UO_1309 (O_1309,N_14170,N_14331);
and UO_1310 (O_1310,N_14729,N_14020);
and UO_1311 (O_1311,N_14062,N_14023);
and UO_1312 (O_1312,N_14211,N_14941);
nand UO_1313 (O_1313,N_14722,N_14678);
nor UO_1314 (O_1314,N_14933,N_14745);
nor UO_1315 (O_1315,N_14195,N_14555);
nor UO_1316 (O_1316,N_14487,N_14662);
nor UO_1317 (O_1317,N_14295,N_14055);
nand UO_1318 (O_1318,N_14417,N_14743);
xnor UO_1319 (O_1319,N_14028,N_14353);
nor UO_1320 (O_1320,N_14196,N_14406);
nand UO_1321 (O_1321,N_14355,N_14806);
nor UO_1322 (O_1322,N_14257,N_14623);
xnor UO_1323 (O_1323,N_14087,N_14377);
nor UO_1324 (O_1324,N_14993,N_14786);
or UO_1325 (O_1325,N_14374,N_14000);
or UO_1326 (O_1326,N_14152,N_14002);
or UO_1327 (O_1327,N_14905,N_14983);
and UO_1328 (O_1328,N_14758,N_14172);
and UO_1329 (O_1329,N_14258,N_14248);
and UO_1330 (O_1330,N_14383,N_14891);
nand UO_1331 (O_1331,N_14546,N_14651);
and UO_1332 (O_1332,N_14394,N_14892);
and UO_1333 (O_1333,N_14877,N_14534);
or UO_1334 (O_1334,N_14172,N_14712);
nor UO_1335 (O_1335,N_14358,N_14236);
nor UO_1336 (O_1336,N_14623,N_14981);
nand UO_1337 (O_1337,N_14036,N_14127);
xnor UO_1338 (O_1338,N_14903,N_14743);
or UO_1339 (O_1339,N_14829,N_14899);
nor UO_1340 (O_1340,N_14982,N_14165);
nor UO_1341 (O_1341,N_14283,N_14525);
or UO_1342 (O_1342,N_14342,N_14523);
or UO_1343 (O_1343,N_14991,N_14970);
nor UO_1344 (O_1344,N_14292,N_14760);
nand UO_1345 (O_1345,N_14130,N_14334);
xor UO_1346 (O_1346,N_14853,N_14269);
nand UO_1347 (O_1347,N_14648,N_14538);
or UO_1348 (O_1348,N_14298,N_14349);
or UO_1349 (O_1349,N_14205,N_14371);
nand UO_1350 (O_1350,N_14282,N_14656);
nand UO_1351 (O_1351,N_14522,N_14905);
xnor UO_1352 (O_1352,N_14851,N_14391);
nand UO_1353 (O_1353,N_14478,N_14387);
xor UO_1354 (O_1354,N_14796,N_14255);
or UO_1355 (O_1355,N_14674,N_14962);
or UO_1356 (O_1356,N_14425,N_14726);
and UO_1357 (O_1357,N_14140,N_14537);
and UO_1358 (O_1358,N_14531,N_14605);
and UO_1359 (O_1359,N_14990,N_14853);
nor UO_1360 (O_1360,N_14965,N_14972);
or UO_1361 (O_1361,N_14906,N_14154);
or UO_1362 (O_1362,N_14381,N_14936);
nand UO_1363 (O_1363,N_14653,N_14574);
or UO_1364 (O_1364,N_14404,N_14263);
or UO_1365 (O_1365,N_14902,N_14440);
and UO_1366 (O_1366,N_14427,N_14179);
nor UO_1367 (O_1367,N_14101,N_14027);
nor UO_1368 (O_1368,N_14005,N_14924);
nor UO_1369 (O_1369,N_14665,N_14278);
nor UO_1370 (O_1370,N_14264,N_14525);
xnor UO_1371 (O_1371,N_14379,N_14674);
nand UO_1372 (O_1372,N_14003,N_14558);
and UO_1373 (O_1373,N_14269,N_14928);
and UO_1374 (O_1374,N_14705,N_14091);
or UO_1375 (O_1375,N_14442,N_14014);
nor UO_1376 (O_1376,N_14543,N_14764);
or UO_1377 (O_1377,N_14578,N_14024);
and UO_1378 (O_1378,N_14349,N_14691);
or UO_1379 (O_1379,N_14228,N_14120);
nor UO_1380 (O_1380,N_14552,N_14077);
or UO_1381 (O_1381,N_14830,N_14030);
nor UO_1382 (O_1382,N_14134,N_14057);
nor UO_1383 (O_1383,N_14059,N_14639);
or UO_1384 (O_1384,N_14987,N_14210);
and UO_1385 (O_1385,N_14197,N_14632);
or UO_1386 (O_1386,N_14535,N_14754);
nor UO_1387 (O_1387,N_14200,N_14717);
and UO_1388 (O_1388,N_14384,N_14514);
and UO_1389 (O_1389,N_14096,N_14665);
and UO_1390 (O_1390,N_14231,N_14558);
nor UO_1391 (O_1391,N_14726,N_14474);
or UO_1392 (O_1392,N_14810,N_14570);
or UO_1393 (O_1393,N_14576,N_14666);
nand UO_1394 (O_1394,N_14946,N_14146);
and UO_1395 (O_1395,N_14230,N_14432);
nand UO_1396 (O_1396,N_14817,N_14086);
nand UO_1397 (O_1397,N_14568,N_14344);
nor UO_1398 (O_1398,N_14775,N_14194);
or UO_1399 (O_1399,N_14069,N_14026);
nor UO_1400 (O_1400,N_14902,N_14143);
and UO_1401 (O_1401,N_14664,N_14813);
and UO_1402 (O_1402,N_14203,N_14515);
or UO_1403 (O_1403,N_14508,N_14391);
nor UO_1404 (O_1404,N_14308,N_14813);
or UO_1405 (O_1405,N_14955,N_14221);
or UO_1406 (O_1406,N_14579,N_14071);
xor UO_1407 (O_1407,N_14458,N_14657);
and UO_1408 (O_1408,N_14945,N_14153);
nand UO_1409 (O_1409,N_14915,N_14410);
nor UO_1410 (O_1410,N_14231,N_14979);
or UO_1411 (O_1411,N_14152,N_14233);
nor UO_1412 (O_1412,N_14137,N_14032);
nand UO_1413 (O_1413,N_14895,N_14038);
nor UO_1414 (O_1414,N_14732,N_14270);
and UO_1415 (O_1415,N_14010,N_14068);
nor UO_1416 (O_1416,N_14999,N_14511);
and UO_1417 (O_1417,N_14682,N_14203);
or UO_1418 (O_1418,N_14822,N_14931);
or UO_1419 (O_1419,N_14605,N_14165);
xnor UO_1420 (O_1420,N_14895,N_14386);
or UO_1421 (O_1421,N_14281,N_14645);
nor UO_1422 (O_1422,N_14309,N_14766);
or UO_1423 (O_1423,N_14506,N_14275);
xor UO_1424 (O_1424,N_14645,N_14661);
or UO_1425 (O_1425,N_14416,N_14749);
nor UO_1426 (O_1426,N_14029,N_14054);
nand UO_1427 (O_1427,N_14021,N_14708);
nor UO_1428 (O_1428,N_14411,N_14896);
nand UO_1429 (O_1429,N_14096,N_14710);
nor UO_1430 (O_1430,N_14769,N_14223);
nand UO_1431 (O_1431,N_14063,N_14093);
nand UO_1432 (O_1432,N_14852,N_14890);
nor UO_1433 (O_1433,N_14417,N_14613);
nor UO_1434 (O_1434,N_14429,N_14711);
xnor UO_1435 (O_1435,N_14852,N_14796);
nor UO_1436 (O_1436,N_14092,N_14725);
nor UO_1437 (O_1437,N_14116,N_14811);
or UO_1438 (O_1438,N_14846,N_14731);
nand UO_1439 (O_1439,N_14297,N_14750);
or UO_1440 (O_1440,N_14092,N_14297);
nor UO_1441 (O_1441,N_14200,N_14670);
nor UO_1442 (O_1442,N_14404,N_14807);
nand UO_1443 (O_1443,N_14647,N_14330);
or UO_1444 (O_1444,N_14701,N_14661);
nand UO_1445 (O_1445,N_14006,N_14677);
nand UO_1446 (O_1446,N_14520,N_14659);
or UO_1447 (O_1447,N_14474,N_14373);
or UO_1448 (O_1448,N_14860,N_14043);
nand UO_1449 (O_1449,N_14296,N_14949);
xnor UO_1450 (O_1450,N_14353,N_14291);
or UO_1451 (O_1451,N_14600,N_14282);
nor UO_1452 (O_1452,N_14678,N_14277);
nor UO_1453 (O_1453,N_14100,N_14706);
nor UO_1454 (O_1454,N_14389,N_14757);
nor UO_1455 (O_1455,N_14361,N_14814);
nand UO_1456 (O_1456,N_14841,N_14028);
xnor UO_1457 (O_1457,N_14151,N_14050);
or UO_1458 (O_1458,N_14609,N_14532);
or UO_1459 (O_1459,N_14354,N_14643);
nand UO_1460 (O_1460,N_14640,N_14411);
nand UO_1461 (O_1461,N_14859,N_14268);
and UO_1462 (O_1462,N_14261,N_14579);
xor UO_1463 (O_1463,N_14586,N_14607);
and UO_1464 (O_1464,N_14373,N_14239);
nand UO_1465 (O_1465,N_14983,N_14313);
nor UO_1466 (O_1466,N_14241,N_14224);
nor UO_1467 (O_1467,N_14920,N_14011);
nand UO_1468 (O_1468,N_14178,N_14616);
and UO_1469 (O_1469,N_14333,N_14179);
nand UO_1470 (O_1470,N_14791,N_14217);
and UO_1471 (O_1471,N_14554,N_14609);
or UO_1472 (O_1472,N_14136,N_14842);
or UO_1473 (O_1473,N_14590,N_14979);
xor UO_1474 (O_1474,N_14913,N_14642);
and UO_1475 (O_1475,N_14958,N_14888);
nor UO_1476 (O_1476,N_14101,N_14570);
or UO_1477 (O_1477,N_14615,N_14090);
xor UO_1478 (O_1478,N_14605,N_14736);
and UO_1479 (O_1479,N_14273,N_14709);
nor UO_1480 (O_1480,N_14068,N_14546);
nor UO_1481 (O_1481,N_14561,N_14651);
and UO_1482 (O_1482,N_14182,N_14516);
nor UO_1483 (O_1483,N_14074,N_14261);
and UO_1484 (O_1484,N_14070,N_14441);
nand UO_1485 (O_1485,N_14500,N_14002);
and UO_1486 (O_1486,N_14126,N_14427);
nand UO_1487 (O_1487,N_14986,N_14525);
xnor UO_1488 (O_1488,N_14495,N_14658);
nand UO_1489 (O_1489,N_14638,N_14679);
or UO_1490 (O_1490,N_14983,N_14150);
nand UO_1491 (O_1491,N_14080,N_14188);
nand UO_1492 (O_1492,N_14738,N_14288);
or UO_1493 (O_1493,N_14631,N_14530);
and UO_1494 (O_1494,N_14102,N_14231);
or UO_1495 (O_1495,N_14205,N_14609);
nor UO_1496 (O_1496,N_14337,N_14346);
and UO_1497 (O_1497,N_14861,N_14120);
nand UO_1498 (O_1498,N_14305,N_14376);
or UO_1499 (O_1499,N_14563,N_14807);
nor UO_1500 (O_1500,N_14060,N_14648);
nand UO_1501 (O_1501,N_14825,N_14853);
or UO_1502 (O_1502,N_14900,N_14402);
or UO_1503 (O_1503,N_14677,N_14916);
nand UO_1504 (O_1504,N_14178,N_14274);
xnor UO_1505 (O_1505,N_14330,N_14754);
nand UO_1506 (O_1506,N_14846,N_14262);
nor UO_1507 (O_1507,N_14263,N_14284);
and UO_1508 (O_1508,N_14475,N_14382);
nand UO_1509 (O_1509,N_14629,N_14661);
nand UO_1510 (O_1510,N_14558,N_14721);
xnor UO_1511 (O_1511,N_14543,N_14161);
nor UO_1512 (O_1512,N_14580,N_14347);
nor UO_1513 (O_1513,N_14169,N_14312);
nand UO_1514 (O_1514,N_14739,N_14879);
xor UO_1515 (O_1515,N_14010,N_14807);
or UO_1516 (O_1516,N_14437,N_14528);
nand UO_1517 (O_1517,N_14796,N_14841);
or UO_1518 (O_1518,N_14091,N_14494);
and UO_1519 (O_1519,N_14987,N_14855);
or UO_1520 (O_1520,N_14411,N_14349);
nand UO_1521 (O_1521,N_14518,N_14380);
nor UO_1522 (O_1522,N_14667,N_14917);
nor UO_1523 (O_1523,N_14247,N_14652);
or UO_1524 (O_1524,N_14980,N_14401);
nand UO_1525 (O_1525,N_14268,N_14031);
nor UO_1526 (O_1526,N_14135,N_14329);
or UO_1527 (O_1527,N_14746,N_14393);
nand UO_1528 (O_1528,N_14918,N_14151);
or UO_1529 (O_1529,N_14554,N_14177);
nor UO_1530 (O_1530,N_14421,N_14168);
nand UO_1531 (O_1531,N_14657,N_14630);
nor UO_1532 (O_1532,N_14085,N_14071);
nor UO_1533 (O_1533,N_14877,N_14876);
nor UO_1534 (O_1534,N_14747,N_14040);
or UO_1535 (O_1535,N_14575,N_14068);
and UO_1536 (O_1536,N_14414,N_14765);
or UO_1537 (O_1537,N_14205,N_14921);
and UO_1538 (O_1538,N_14305,N_14357);
xnor UO_1539 (O_1539,N_14356,N_14006);
xor UO_1540 (O_1540,N_14692,N_14174);
xnor UO_1541 (O_1541,N_14936,N_14220);
xnor UO_1542 (O_1542,N_14968,N_14434);
or UO_1543 (O_1543,N_14737,N_14397);
and UO_1544 (O_1544,N_14031,N_14264);
and UO_1545 (O_1545,N_14484,N_14631);
nor UO_1546 (O_1546,N_14059,N_14325);
and UO_1547 (O_1547,N_14149,N_14511);
xnor UO_1548 (O_1548,N_14582,N_14248);
nor UO_1549 (O_1549,N_14416,N_14034);
and UO_1550 (O_1550,N_14143,N_14469);
nor UO_1551 (O_1551,N_14401,N_14479);
and UO_1552 (O_1552,N_14898,N_14904);
xnor UO_1553 (O_1553,N_14812,N_14719);
nand UO_1554 (O_1554,N_14496,N_14440);
and UO_1555 (O_1555,N_14098,N_14979);
nand UO_1556 (O_1556,N_14025,N_14298);
nor UO_1557 (O_1557,N_14008,N_14027);
nand UO_1558 (O_1558,N_14286,N_14897);
and UO_1559 (O_1559,N_14549,N_14815);
or UO_1560 (O_1560,N_14341,N_14025);
xor UO_1561 (O_1561,N_14427,N_14960);
nor UO_1562 (O_1562,N_14749,N_14916);
nor UO_1563 (O_1563,N_14738,N_14981);
and UO_1564 (O_1564,N_14561,N_14620);
nand UO_1565 (O_1565,N_14623,N_14384);
nor UO_1566 (O_1566,N_14446,N_14665);
or UO_1567 (O_1567,N_14081,N_14406);
nand UO_1568 (O_1568,N_14542,N_14386);
xnor UO_1569 (O_1569,N_14540,N_14204);
nor UO_1570 (O_1570,N_14665,N_14597);
nor UO_1571 (O_1571,N_14904,N_14944);
nor UO_1572 (O_1572,N_14139,N_14241);
xor UO_1573 (O_1573,N_14812,N_14415);
nand UO_1574 (O_1574,N_14468,N_14675);
nor UO_1575 (O_1575,N_14086,N_14856);
and UO_1576 (O_1576,N_14950,N_14862);
nand UO_1577 (O_1577,N_14686,N_14616);
and UO_1578 (O_1578,N_14686,N_14723);
xnor UO_1579 (O_1579,N_14204,N_14334);
nor UO_1580 (O_1580,N_14023,N_14383);
or UO_1581 (O_1581,N_14752,N_14398);
nand UO_1582 (O_1582,N_14952,N_14787);
or UO_1583 (O_1583,N_14795,N_14034);
and UO_1584 (O_1584,N_14161,N_14933);
nand UO_1585 (O_1585,N_14814,N_14378);
nand UO_1586 (O_1586,N_14271,N_14420);
and UO_1587 (O_1587,N_14015,N_14983);
or UO_1588 (O_1588,N_14497,N_14378);
or UO_1589 (O_1589,N_14345,N_14518);
nor UO_1590 (O_1590,N_14216,N_14666);
nor UO_1591 (O_1591,N_14840,N_14285);
and UO_1592 (O_1592,N_14970,N_14225);
nor UO_1593 (O_1593,N_14549,N_14459);
nor UO_1594 (O_1594,N_14632,N_14791);
xor UO_1595 (O_1595,N_14531,N_14902);
and UO_1596 (O_1596,N_14667,N_14849);
nor UO_1597 (O_1597,N_14548,N_14003);
and UO_1598 (O_1598,N_14209,N_14701);
nand UO_1599 (O_1599,N_14707,N_14702);
or UO_1600 (O_1600,N_14883,N_14913);
nand UO_1601 (O_1601,N_14354,N_14775);
xnor UO_1602 (O_1602,N_14855,N_14026);
nand UO_1603 (O_1603,N_14094,N_14979);
or UO_1604 (O_1604,N_14094,N_14189);
nand UO_1605 (O_1605,N_14045,N_14069);
nor UO_1606 (O_1606,N_14492,N_14152);
xnor UO_1607 (O_1607,N_14224,N_14210);
xnor UO_1608 (O_1608,N_14666,N_14246);
nand UO_1609 (O_1609,N_14171,N_14600);
nand UO_1610 (O_1610,N_14113,N_14583);
or UO_1611 (O_1611,N_14239,N_14996);
and UO_1612 (O_1612,N_14024,N_14013);
and UO_1613 (O_1613,N_14380,N_14454);
nor UO_1614 (O_1614,N_14805,N_14630);
and UO_1615 (O_1615,N_14921,N_14089);
nand UO_1616 (O_1616,N_14290,N_14130);
nand UO_1617 (O_1617,N_14244,N_14629);
nand UO_1618 (O_1618,N_14706,N_14518);
nand UO_1619 (O_1619,N_14724,N_14916);
and UO_1620 (O_1620,N_14307,N_14719);
nor UO_1621 (O_1621,N_14731,N_14570);
and UO_1622 (O_1622,N_14939,N_14273);
or UO_1623 (O_1623,N_14087,N_14168);
and UO_1624 (O_1624,N_14370,N_14449);
xnor UO_1625 (O_1625,N_14212,N_14703);
and UO_1626 (O_1626,N_14549,N_14412);
xor UO_1627 (O_1627,N_14298,N_14975);
or UO_1628 (O_1628,N_14921,N_14970);
nand UO_1629 (O_1629,N_14082,N_14556);
xnor UO_1630 (O_1630,N_14787,N_14489);
or UO_1631 (O_1631,N_14993,N_14355);
nand UO_1632 (O_1632,N_14368,N_14111);
and UO_1633 (O_1633,N_14532,N_14968);
xor UO_1634 (O_1634,N_14744,N_14777);
or UO_1635 (O_1635,N_14509,N_14050);
xor UO_1636 (O_1636,N_14619,N_14269);
and UO_1637 (O_1637,N_14636,N_14720);
and UO_1638 (O_1638,N_14249,N_14481);
nand UO_1639 (O_1639,N_14947,N_14573);
and UO_1640 (O_1640,N_14508,N_14494);
and UO_1641 (O_1641,N_14103,N_14178);
nor UO_1642 (O_1642,N_14958,N_14568);
and UO_1643 (O_1643,N_14768,N_14483);
xnor UO_1644 (O_1644,N_14590,N_14931);
nand UO_1645 (O_1645,N_14528,N_14913);
or UO_1646 (O_1646,N_14673,N_14242);
nor UO_1647 (O_1647,N_14189,N_14615);
and UO_1648 (O_1648,N_14029,N_14694);
or UO_1649 (O_1649,N_14833,N_14825);
nor UO_1650 (O_1650,N_14805,N_14488);
nand UO_1651 (O_1651,N_14625,N_14521);
and UO_1652 (O_1652,N_14086,N_14969);
nor UO_1653 (O_1653,N_14184,N_14745);
or UO_1654 (O_1654,N_14331,N_14378);
nand UO_1655 (O_1655,N_14556,N_14451);
xor UO_1656 (O_1656,N_14459,N_14688);
xor UO_1657 (O_1657,N_14155,N_14188);
and UO_1658 (O_1658,N_14004,N_14118);
or UO_1659 (O_1659,N_14254,N_14748);
nand UO_1660 (O_1660,N_14742,N_14676);
and UO_1661 (O_1661,N_14010,N_14395);
xor UO_1662 (O_1662,N_14708,N_14458);
and UO_1663 (O_1663,N_14372,N_14354);
nand UO_1664 (O_1664,N_14349,N_14115);
and UO_1665 (O_1665,N_14430,N_14222);
or UO_1666 (O_1666,N_14880,N_14270);
nor UO_1667 (O_1667,N_14955,N_14293);
or UO_1668 (O_1668,N_14639,N_14586);
nand UO_1669 (O_1669,N_14565,N_14657);
nand UO_1670 (O_1670,N_14794,N_14605);
and UO_1671 (O_1671,N_14956,N_14371);
and UO_1672 (O_1672,N_14834,N_14924);
nand UO_1673 (O_1673,N_14562,N_14454);
and UO_1674 (O_1674,N_14162,N_14749);
nor UO_1675 (O_1675,N_14356,N_14567);
or UO_1676 (O_1676,N_14023,N_14156);
and UO_1677 (O_1677,N_14852,N_14703);
nor UO_1678 (O_1678,N_14957,N_14642);
xnor UO_1679 (O_1679,N_14332,N_14196);
xor UO_1680 (O_1680,N_14771,N_14179);
xnor UO_1681 (O_1681,N_14025,N_14129);
or UO_1682 (O_1682,N_14918,N_14882);
and UO_1683 (O_1683,N_14273,N_14170);
nand UO_1684 (O_1684,N_14972,N_14147);
nand UO_1685 (O_1685,N_14566,N_14557);
and UO_1686 (O_1686,N_14615,N_14390);
or UO_1687 (O_1687,N_14901,N_14007);
nand UO_1688 (O_1688,N_14856,N_14347);
nand UO_1689 (O_1689,N_14412,N_14052);
nor UO_1690 (O_1690,N_14350,N_14916);
and UO_1691 (O_1691,N_14451,N_14094);
or UO_1692 (O_1692,N_14776,N_14183);
and UO_1693 (O_1693,N_14448,N_14408);
and UO_1694 (O_1694,N_14554,N_14310);
xnor UO_1695 (O_1695,N_14565,N_14366);
or UO_1696 (O_1696,N_14722,N_14093);
nor UO_1697 (O_1697,N_14595,N_14864);
nor UO_1698 (O_1698,N_14154,N_14987);
xor UO_1699 (O_1699,N_14056,N_14781);
or UO_1700 (O_1700,N_14214,N_14303);
nand UO_1701 (O_1701,N_14534,N_14629);
or UO_1702 (O_1702,N_14953,N_14552);
nand UO_1703 (O_1703,N_14051,N_14466);
nand UO_1704 (O_1704,N_14582,N_14487);
and UO_1705 (O_1705,N_14279,N_14897);
and UO_1706 (O_1706,N_14491,N_14241);
or UO_1707 (O_1707,N_14617,N_14913);
nor UO_1708 (O_1708,N_14132,N_14305);
or UO_1709 (O_1709,N_14884,N_14847);
or UO_1710 (O_1710,N_14929,N_14447);
xnor UO_1711 (O_1711,N_14033,N_14843);
or UO_1712 (O_1712,N_14294,N_14505);
nand UO_1713 (O_1713,N_14762,N_14450);
or UO_1714 (O_1714,N_14741,N_14986);
nor UO_1715 (O_1715,N_14277,N_14629);
xor UO_1716 (O_1716,N_14881,N_14126);
nand UO_1717 (O_1717,N_14753,N_14716);
nor UO_1718 (O_1718,N_14124,N_14835);
and UO_1719 (O_1719,N_14810,N_14107);
and UO_1720 (O_1720,N_14364,N_14097);
and UO_1721 (O_1721,N_14989,N_14695);
nand UO_1722 (O_1722,N_14908,N_14535);
nor UO_1723 (O_1723,N_14550,N_14238);
or UO_1724 (O_1724,N_14446,N_14748);
nand UO_1725 (O_1725,N_14878,N_14606);
nor UO_1726 (O_1726,N_14158,N_14730);
nand UO_1727 (O_1727,N_14704,N_14222);
nand UO_1728 (O_1728,N_14909,N_14300);
and UO_1729 (O_1729,N_14166,N_14924);
xnor UO_1730 (O_1730,N_14812,N_14001);
or UO_1731 (O_1731,N_14511,N_14437);
nor UO_1732 (O_1732,N_14539,N_14782);
or UO_1733 (O_1733,N_14665,N_14911);
and UO_1734 (O_1734,N_14334,N_14122);
nor UO_1735 (O_1735,N_14646,N_14356);
nand UO_1736 (O_1736,N_14888,N_14901);
nand UO_1737 (O_1737,N_14198,N_14943);
nor UO_1738 (O_1738,N_14548,N_14702);
nand UO_1739 (O_1739,N_14096,N_14253);
or UO_1740 (O_1740,N_14323,N_14273);
or UO_1741 (O_1741,N_14899,N_14158);
and UO_1742 (O_1742,N_14368,N_14037);
or UO_1743 (O_1743,N_14328,N_14187);
and UO_1744 (O_1744,N_14366,N_14314);
and UO_1745 (O_1745,N_14281,N_14483);
nor UO_1746 (O_1746,N_14779,N_14356);
nor UO_1747 (O_1747,N_14115,N_14615);
xor UO_1748 (O_1748,N_14216,N_14863);
nand UO_1749 (O_1749,N_14205,N_14497);
nand UO_1750 (O_1750,N_14482,N_14636);
nor UO_1751 (O_1751,N_14610,N_14586);
nor UO_1752 (O_1752,N_14504,N_14167);
nor UO_1753 (O_1753,N_14565,N_14810);
or UO_1754 (O_1754,N_14550,N_14578);
and UO_1755 (O_1755,N_14799,N_14818);
nor UO_1756 (O_1756,N_14705,N_14810);
nor UO_1757 (O_1757,N_14916,N_14759);
or UO_1758 (O_1758,N_14741,N_14207);
and UO_1759 (O_1759,N_14907,N_14320);
and UO_1760 (O_1760,N_14359,N_14513);
and UO_1761 (O_1761,N_14056,N_14372);
and UO_1762 (O_1762,N_14051,N_14059);
and UO_1763 (O_1763,N_14056,N_14308);
or UO_1764 (O_1764,N_14176,N_14676);
nand UO_1765 (O_1765,N_14808,N_14358);
nand UO_1766 (O_1766,N_14831,N_14386);
nand UO_1767 (O_1767,N_14561,N_14301);
and UO_1768 (O_1768,N_14054,N_14802);
nand UO_1769 (O_1769,N_14210,N_14495);
and UO_1770 (O_1770,N_14683,N_14555);
nor UO_1771 (O_1771,N_14073,N_14944);
nor UO_1772 (O_1772,N_14599,N_14600);
nand UO_1773 (O_1773,N_14856,N_14673);
nor UO_1774 (O_1774,N_14034,N_14775);
nor UO_1775 (O_1775,N_14270,N_14690);
nand UO_1776 (O_1776,N_14152,N_14466);
nor UO_1777 (O_1777,N_14988,N_14260);
nand UO_1778 (O_1778,N_14033,N_14655);
nand UO_1779 (O_1779,N_14487,N_14173);
nor UO_1780 (O_1780,N_14944,N_14626);
nand UO_1781 (O_1781,N_14433,N_14834);
and UO_1782 (O_1782,N_14471,N_14768);
or UO_1783 (O_1783,N_14620,N_14402);
and UO_1784 (O_1784,N_14833,N_14864);
and UO_1785 (O_1785,N_14706,N_14949);
nor UO_1786 (O_1786,N_14605,N_14114);
and UO_1787 (O_1787,N_14471,N_14689);
nand UO_1788 (O_1788,N_14830,N_14313);
nand UO_1789 (O_1789,N_14094,N_14617);
xor UO_1790 (O_1790,N_14926,N_14117);
and UO_1791 (O_1791,N_14185,N_14432);
or UO_1792 (O_1792,N_14387,N_14234);
nor UO_1793 (O_1793,N_14523,N_14336);
nand UO_1794 (O_1794,N_14903,N_14014);
xor UO_1795 (O_1795,N_14182,N_14847);
nor UO_1796 (O_1796,N_14249,N_14639);
and UO_1797 (O_1797,N_14500,N_14706);
nand UO_1798 (O_1798,N_14784,N_14969);
or UO_1799 (O_1799,N_14510,N_14785);
nand UO_1800 (O_1800,N_14158,N_14499);
nand UO_1801 (O_1801,N_14791,N_14765);
nand UO_1802 (O_1802,N_14417,N_14054);
and UO_1803 (O_1803,N_14630,N_14210);
or UO_1804 (O_1804,N_14597,N_14508);
or UO_1805 (O_1805,N_14030,N_14073);
and UO_1806 (O_1806,N_14154,N_14692);
or UO_1807 (O_1807,N_14383,N_14740);
nand UO_1808 (O_1808,N_14760,N_14336);
and UO_1809 (O_1809,N_14422,N_14893);
nand UO_1810 (O_1810,N_14100,N_14777);
nor UO_1811 (O_1811,N_14976,N_14204);
nand UO_1812 (O_1812,N_14349,N_14462);
xnor UO_1813 (O_1813,N_14571,N_14633);
or UO_1814 (O_1814,N_14807,N_14000);
nand UO_1815 (O_1815,N_14710,N_14586);
and UO_1816 (O_1816,N_14580,N_14592);
or UO_1817 (O_1817,N_14962,N_14191);
or UO_1818 (O_1818,N_14653,N_14916);
and UO_1819 (O_1819,N_14652,N_14113);
or UO_1820 (O_1820,N_14087,N_14930);
nand UO_1821 (O_1821,N_14928,N_14318);
nor UO_1822 (O_1822,N_14935,N_14605);
nor UO_1823 (O_1823,N_14321,N_14031);
nand UO_1824 (O_1824,N_14853,N_14788);
and UO_1825 (O_1825,N_14375,N_14279);
or UO_1826 (O_1826,N_14834,N_14457);
or UO_1827 (O_1827,N_14753,N_14316);
nand UO_1828 (O_1828,N_14244,N_14112);
or UO_1829 (O_1829,N_14921,N_14166);
nand UO_1830 (O_1830,N_14513,N_14193);
and UO_1831 (O_1831,N_14084,N_14056);
xnor UO_1832 (O_1832,N_14124,N_14805);
nor UO_1833 (O_1833,N_14030,N_14544);
and UO_1834 (O_1834,N_14803,N_14941);
and UO_1835 (O_1835,N_14259,N_14666);
and UO_1836 (O_1836,N_14031,N_14637);
nor UO_1837 (O_1837,N_14565,N_14458);
or UO_1838 (O_1838,N_14786,N_14781);
nor UO_1839 (O_1839,N_14255,N_14226);
xnor UO_1840 (O_1840,N_14067,N_14817);
nand UO_1841 (O_1841,N_14625,N_14441);
nand UO_1842 (O_1842,N_14427,N_14752);
nor UO_1843 (O_1843,N_14649,N_14612);
or UO_1844 (O_1844,N_14800,N_14186);
xor UO_1845 (O_1845,N_14541,N_14651);
nand UO_1846 (O_1846,N_14167,N_14486);
or UO_1847 (O_1847,N_14583,N_14469);
and UO_1848 (O_1848,N_14270,N_14164);
nor UO_1849 (O_1849,N_14504,N_14563);
and UO_1850 (O_1850,N_14657,N_14031);
and UO_1851 (O_1851,N_14607,N_14716);
nand UO_1852 (O_1852,N_14440,N_14456);
or UO_1853 (O_1853,N_14704,N_14438);
or UO_1854 (O_1854,N_14172,N_14307);
xnor UO_1855 (O_1855,N_14421,N_14710);
or UO_1856 (O_1856,N_14359,N_14244);
or UO_1857 (O_1857,N_14193,N_14383);
and UO_1858 (O_1858,N_14153,N_14239);
nand UO_1859 (O_1859,N_14962,N_14777);
nor UO_1860 (O_1860,N_14178,N_14552);
and UO_1861 (O_1861,N_14737,N_14491);
nand UO_1862 (O_1862,N_14096,N_14339);
and UO_1863 (O_1863,N_14563,N_14058);
nor UO_1864 (O_1864,N_14774,N_14892);
or UO_1865 (O_1865,N_14997,N_14746);
xor UO_1866 (O_1866,N_14189,N_14778);
or UO_1867 (O_1867,N_14949,N_14514);
nand UO_1868 (O_1868,N_14215,N_14207);
and UO_1869 (O_1869,N_14940,N_14562);
or UO_1870 (O_1870,N_14493,N_14709);
or UO_1871 (O_1871,N_14202,N_14827);
xnor UO_1872 (O_1872,N_14077,N_14317);
nand UO_1873 (O_1873,N_14504,N_14438);
nand UO_1874 (O_1874,N_14908,N_14155);
nor UO_1875 (O_1875,N_14678,N_14457);
or UO_1876 (O_1876,N_14878,N_14264);
nand UO_1877 (O_1877,N_14289,N_14613);
or UO_1878 (O_1878,N_14348,N_14526);
nor UO_1879 (O_1879,N_14744,N_14116);
nand UO_1880 (O_1880,N_14808,N_14188);
and UO_1881 (O_1881,N_14105,N_14600);
or UO_1882 (O_1882,N_14300,N_14741);
and UO_1883 (O_1883,N_14792,N_14481);
nand UO_1884 (O_1884,N_14553,N_14623);
nor UO_1885 (O_1885,N_14343,N_14502);
and UO_1886 (O_1886,N_14312,N_14547);
and UO_1887 (O_1887,N_14004,N_14097);
nand UO_1888 (O_1888,N_14387,N_14153);
nor UO_1889 (O_1889,N_14710,N_14371);
or UO_1890 (O_1890,N_14293,N_14986);
nand UO_1891 (O_1891,N_14543,N_14659);
nand UO_1892 (O_1892,N_14175,N_14289);
nor UO_1893 (O_1893,N_14588,N_14416);
and UO_1894 (O_1894,N_14186,N_14866);
nor UO_1895 (O_1895,N_14820,N_14996);
nor UO_1896 (O_1896,N_14907,N_14911);
nand UO_1897 (O_1897,N_14063,N_14749);
or UO_1898 (O_1898,N_14334,N_14417);
and UO_1899 (O_1899,N_14932,N_14383);
nand UO_1900 (O_1900,N_14467,N_14184);
nor UO_1901 (O_1901,N_14847,N_14426);
or UO_1902 (O_1902,N_14310,N_14579);
or UO_1903 (O_1903,N_14170,N_14929);
nor UO_1904 (O_1904,N_14235,N_14078);
or UO_1905 (O_1905,N_14058,N_14426);
nor UO_1906 (O_1906,N_14420,N_14326);
nand UO_1907 (O_1907,N_14262,N_14860);
and UO_1908 (O_1908,N_14371,N_14688);
nor UO_1909 (O_1909,N_14613,N_14743);
nand UO_1910 (O_1910,N_14669,N_14963);
nand UO_1911 (O_1911,N_14358,N_14694);
or UO_1912 (O_1912,N_14367,N_14041);
nor UO_1913 (O_1913,N_14458,N_14374);
and UO_1914 (O_1914,N_14565,N_14538);
and UO_1915 (O_1915,N_14228,N_14376);
nand UO_1916 (O_1916,N_14658,N_14388);
and UO_1917 (O_1917,N_14577,N_14768);
nor UO_1918 (O_1918,N_14085,N_14966);
xor UO_1919 (O_1919,N_14955,N_14195);
nor UO_1920 (O_1920,N_14467,N_14923);
nor UO_1921 (O_1921,N_14018,N_14091);
or UO_1922 (O_1922,N_14799,N_14825);
xor UO_1923 (O_1923,N_14438,N_14267);
or UO_1924 (O_1924,N_14680,N_14955);
nor UO_1925 (O_1925,N_14851,N_14279);
and UO_1926 (O_1926,N_14515,N_14536);
or UO_1927 (O_1927,N_14634,N_14650);
and UO_1928 (O_1928,N_14817,N_14230);
or UO_1929 (O_1929,N_14943,N_14589);
or UO_1930 (O_1930,N_14703,N_14686);
nor UO_1931 (O_1931,N_14618,N_14497);
or UO_1932 (O_1932,N_14019,N_14133);
xnor UO_1933 (O_1933,N_14641,N_14482);
and UO_1934 (O_1934,N_14897,N_14099);
nor UO_1935 (O_1935,N_14136,N_14836);
nor UO_1936 (O_1936,N_14779,N_14080);
or UO_1937 (O_1937,N_14606,N_14597);
and UO_1938 (O_1938,N_14992,N_14009);
nor UO_1939 (O_1939,N_14436,N_14812);
nand UO_1940 (O_1940,N_14830,N_14449);
and UO_1941 (O_1941,N_14939,N_14409);
or UO_1942 (O_1942,N_14913,N_14621);
nor UO_1943 (O_1943,N_14383,N_14707);
nor UO_1944 (O_1944,N_14289,N_14120);
and UO_1945 (O_1945,N_14495,N_14562);
xnor UO_1946 (O_1946,N_14080,N_14475);
nand UO_1947 (O_1947,N_14808,N_14928);
or UO_1948 (O_1948,N_14210,N_14501);
nand UO_1949 (O_1949,N_14281,N_14813);
nand UO_1950 (O_1950,N_14351,N_14371);
xor UO_1951 (O_1951,N_14899,N_14298);
and UO_1952 (O_1952,N_14762,N_14914);
or UO_1953 (O_1953,N_14274,N_14956);
and UO_1954 (O_1954,N_14219,N_14628);
nand UO_1955 (O_1955,N_14014,N_14460);
nor UO_1956 (O_1956,N_14033,N_14569);
nand UO_1957 (O_1957,N_14585,N_14186);
and UO_1958 (O_1958,N_14144,N_14257);
nand UO_1959 (O_1959,N_14105,N_14046);
nand UO_1960 (O_1960,N_14370,N_14745);
and UO_1961 (O_1961,N_14044,N_14445);
nand UO_1962 (O_1962,N_14918,N_14428);
xnor UO_1963 (O_1963,N_14553,N_14088);
and UO_1964 (O_1964,N_14443,N_14862);
nand UO_1965 (O_1965,N_14054,N_14097);
nor UO_1966 (O_1966,N_14502,N_14242);
nor UO_1967 (O_1967,N_14389,N_14114);
nand UO_1968 (O_1968,N_14292,N_14753);
nand UO_1969 (O_1969,N_14416,N_14624);
and UO_1970 (O_1970,N_14855,N_14604);
or UO_1971 (O_1971,N_14490,N_14591);
nor UO_1972 (O_1972,N_14091,N_14787);
or UO_1973 (O_1973,N_14360,N_14356);
nand UO_1974 (O_1974,N_14299,N_14729);
or UO_1975 (O_1975,N_14475,N_14206);
and UO_1976 (O_1976,N_14757,N_14837);
nand UO_1977 (O_1977,N_14393,N_14179);
or UO_1978 (O_1978,N_14248,N_14490);
and UO_1979 (O_1979,N_14034,N_14172);
xor UO_1980 (O_1980,N_14701,N_14824);
or UO_1981 (O_1981,N_14363,N_14305);
or UO_1982 (O_1982,N_14499,N_14539);
or UO_1983 (O_1983,N_14792,N_14002);
and UO_1984 (O_1984,N_14109,N_14224);
nand UO_1985 (O_1985,N_14511,N_14450);
nor UO_1986 (O_1986,N_14616,N_14231);
nand UO_1987 (O_1987,N_14764,N_14343);
or UO_1988 (O_1988,N_14190,N_14530);
and UO_1989 (O_1989,N_14157,N_14368);
or UO_1990 (O_1990,N_14008,N_14705);
nor UO_1991 (O_1991,N_14141,N_14494);
nand UO_1992 (O_1992,N_14508,N_14994);
and UO_1993 (O_1993,N_14107,N_14574);
or UO_1994 (O_1994,N_14085,N_14089);
or UO_1995 (O_1995,N_14536,N_14091);
or UO_1996 (O_1996,N_14454,N_14738);
nand UO_1997 (O_1997,N_14495,N_14366);
xor UO_1998 (O_1998,N_14377,N_14362);
nand UO_1999 (O_1999,N_14898,N_14863);
endmodule