module basic_750_5000_1000_10_levels_2xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
nand U0 (N_0,In_23,In_715);
nand U1 (N_1,In_8,In_120);
nand U2 (N_2,In_636,In_360);
and U3 (N_3,In_585,In_702);
or U4 (N_4,In_233,In_41);
nand U5 (N_5,In_150,In_158);
and U6 (N_6,In_430,In_195);
and U7 (N_7,In_591,In_113);
or U8 (N_8,In_580,In_383);
nand U9 (N_9,In_24,In_109);
or U10 (N_10,In_644,In_535);
and U11 (N_11,In_296,In_9);
nor U12 (N_12,In_249,In_19);
nor U13 (N_13,In_440,In_499);
nand U14 (N_14,In_659,In_15);
and U15 (N_15,In_379,In_721);
nand U16 (N_16,In_122,In_123);
nor U17 (N_17,In_333,In_477);
and U18 (N_18,In_89,In_587);
nor U19 (N_19,In_205,In_688);
or U20 (N_20,In_457,In_394);
and U21 (N_21,In_505,In_625);
or U22 (N_22,In_471,In_298);
or U23 (N_23,In_260,In_98);
nand U24 (N_24,In_180,In_605);
or U25 (N_25,In_690,In_377);
nor U26 (N_26,In_447,In_621);
or U27 (N_27,In_281,In_689);
and U28 (N_28,In_337,In_594);
nand U29 (N_29,In_735,In_522);
nor U30 (N_30,In_575,In_431);
nand U31 (N_31,In_85,In_116);
or U32 (N_32,In_322,In_255);
nor U33 (N_33,In_581,In_395);
nor U34 (N_34,In_239,In_490);
or U35 (N_35,In_307,In_439);
nand U36 (N_36,In_536,In_194);
or U37 (N_37,In_677,In_501);
nand U38 (N_38,In_456,In_267);
nor U39 (N_39,In_583,In_172);
nor U40 (N_40,In_364,In_290);
or U41 (N_41,In_402,In_200);
or U42 (N_42,In_95,In_408);
nor U43 (N_43,In_468,In_48);
nand U44 (N_44,In_299,In_320);
nand U45 (N_45,In_17,In_243);
or U46 (N_46,In_616,In_230);
and U47 (N_47,In_657,In_295);
and U48 (N_48,In_227,In_97);
or U49 (N_49,In_466,In_592);
and U50 (N_50,In_486,In_665);
nand U51 (N_51,In_2,In_306);
xor U52 (N_52,In_598,In_265);
and U53 (N_53,In_642,In_429);
nor U54 (N_54,In_45,In_284);
nand U55 (N_55,In_71,In_404);
or U56 (N_56,In_669,In_631);
and U57 (N_57,In_280,In_484);
and U58 (N_58,In_272,In_606);
and U59 (N_59,In_99,In_115);
nor U60 (N_60,In_454,In_726);
or U61 (N_61,In_463,In_465);
or U62 (N_62,In_617,In_217);
nand U63 (N_63,In_413,In_170);
or U64 (N_64,In_332,In_136);
nor U65 (N_65,In_26,In_723);
and U66 (N_66,In_338,In_552);
nor U67 (N_67,In_528,In_668);
nor U68 (N_68,In_467,In_588);
nor U69 (N_69,In_571,In_162);
or U70 (N_70,In_237,In_341);
nor U71 (N_71,In_81,In_512);
nand U72 (N_72,In_32,In_179);
nor U73 (N_73,In_14,In_489);
or U74 (N_74,In_87,In_579);
nand U75 (N_75,In_736,In_40);
and U76 (N_76,In_416,In_185);
nand U77 (N_77,In_613,In_390);
or U78 (N_78,In_599,In_154);
nor U79 (N_79,In_112,In_167);
nand U80 (N_80,In_28,In_92);
or U81 (N_81,In_286,In_529);
or U82 (N_82,In_317,In_485);
nor U83 (N_83,In_472,In_421);
or U84 (N_84,In_737,In_168);
or U85 (N_85,In_70,In_662);
nor U86 (N_86,In_257,In_597);
nand U87 (N_87,In_746,In_334);
or U88 (N_88,In_258,In_564);
or U89 (N_89,In_343,In_107);
nor U90 (N_90,In_418,In_426);
and U91 (N_91,In_355,In_655);
nor U92 (N_92,In_69,In_254);
or U93 (N_93,In_119,In_104);
nand U94 (N_94,In_407,In_369);
or U95 (N_95,In_694,In_132);
nand U96 (N_96,In_7,In_156);
nand U97 (N_97,In_496,In_719);
and U98 (N_98,In_412,In_263);
and U99 (N_99,In_86,In_449);
nor U100 (N_100,In_716,In_483);
nand U101 (N_101,In_21,In_519);
nor U102 (N_102,In_538,In_387);
or U103 (N_103,In_91,In_503);
nor U104 (N_104,In_555,In_714);
nor U105 (N_105,In_600,In_675);
nor U106 (N_106,In_693,In_568);
or U107 (N_107,In_403,In_521);
or U108 (N_108,In_743,In_654);
and U109 (N_109,In_262,In_321);
and U110 (N_110,In_30,In_405);
and U111 (N_111,In_745,In_593);
nor U112 (N_112,In_370,In_530);
nand U113 (N_113,In_506,In_64);
xor U114 (N_114,In_221,In_209);
or U115 (N_115,In_228,In_31);
nor U116 (N_116,In_225,In_612);
and U117 (N_117,In_652,In_551);
nor U118 (N_118,In_352,In_685);
xnor U119 (N_119,In_208,In_229);
and U120 (N_120,In_663,In_549);
and U121 (N_121,In_201,In_684);
and U122 (N_122,In_118,In_410);
or U123 (N_123,In_121,In_645);
nor U124 (N_124,In_419,In_300);
and U125 (N_125,In_184,In_476);
and U126 (N_126,In_153,In_53);
nor U127 (N_127,In_371,In_117);
nand U128 (N_128,In_125,In_5);
and U129 (N_129,In_749,In_350);
xor U130 (N_130,In_103,In_683);
or U131 (N_131,In_135,In_482);
and U132 (N_132,In_713,In_703);
or U133 (N_133,In_311,In_247);
nor U134 (N_134,In_442,In_29);
and U135 (N_135,In_680,In_708);
and U136 (N_136,In_595,In_666);
or U137 (N_137,In_604,In_266);
nor U138 (N_138,In_141,In_236);
and U139 (N_139,In_65,In_459);
or U140 (N_140,In_565,In_546);
nor U141 (N_141,In_610,In_691);
nor U142 (N_142,In_640,In_509);
and U143 (N_143,In_562,In_314);
nor U144 (N_144,In_422,In_491);
nor U145 (N_145,In_312,In_537);
or U146 (N_146,In_382,In_235);
nand U147 (N_147,In_20,In_432);
nor U148 (N_148,In_176,In_169);
and U149 (N_149,In_58,In_560);
and U150 (N_150,In_363,In_539);
and U151 (N_151,In_508,In_473);
nand U152 (N_152,In_331,In_325);
and U153 (N_153,In_464,In_637);
nand U154 (N_154,In_687,In_740);
nor U155 (N_155,In_94,In_524);
nand U156 (N_156,In_189,In_618);
and U157 (N_157,In_202,In_301);
or U158 (N_158,In_705,In_566);
and U159 (N_159,In_603,In_544);
nand U160 (N_160,In_214,In_561);
xor U161 (N_161,In_177,In_542);
and U162 (N_162,In_540,In_651);
nor U163 (N_163,In_146,In_520);
nand U164 (N_164,In_61,In_10);
and U165 (N_165,In_347,In_151);
nand U166 (N_166,In_3,In_573);
or U167 (N_167,In_292,In_397);
nor U168 (N_168,In_191,In_149);
nand U169 (N_169,In_129,In_282);
or U170 (N_170,In_304,In_732);
and U171 (N_171,In_586,In_0);
or U172 (N_172,In_739,In_590);
nand U173 (N_173,In_44,In_190);
or U174 (N_174,In_108,In_319);
and U175 (N_175,In_576,In_218);
and U176 (N_176,In_589,In_199);
nor U177 (N_177,In_400,In_635);
xor U178 (N_178,In_417,In_164);
or U179 (N_179,In_611,In_602);
and U180 (N_180,In_346,In_401);
and U181 (N_181,In_504,In_43);
and U182 (N_182,In_502,In_250);
nor U183 (N_183,In_391,In_445);
nor U184 (N_184,In_608,In_275);
nand U185 (N_185,In_615,In_601);
nand U186 (N_186,In_252,In_553);
or U187 (N_187,In_710,In_556);
nand U188 (N_188,In_481,In_105);
or U189 (N_189,In_83,In_545);
and U190 (N_190,In_140,In_207);
and U191 (N_191,In_623,In_38);
and U192 (N_192,In_570,In_532);
nor U193 (N_193,In_159,In_451);
and U194 (N_194,In_453,In_142);
nand U195 (N_195,In_174,In_256);
and U196 (N_196,In_11,In_724);
or U197 (N_197,In_212,In_323);
and U198 (N_198,In_380,In_4);
and U199 (N_199,In_469,In_582);
nor U200 (N_200,In_648,In_448);
nand U201 (N_201,In_368,In_607);
or U202 (N_202,In_34,In_500);
and U203 (N_203,In_152,In_406);
and U204 (N_204,In_183,In_709);
nor U205 (N_205,In_330,In_78);
and U206 (N_206,In_133,In_56);
or U207 (N_207,In_639,In_77);
or U208 (N_208,In_633,In_22);
and U209 (N_209,In_729,In_155);
and U210 (N_210,In_173,In_492);
nor U211 (N_211,In_211,In_124);
nand U212 (N_212,In_345,In_157);
nor U213 (N_213,In_534,In_329);
nand U214 (N_214,In_75,In_126);
xor U215 (N_215,In_638,In_511);
or U216 (N_216,In_676,In_90);
nor U217 (N_217,In_66,In_728);
xor U218 (N_218,In_232,In_310);
nor U219 (N_219,In_274,In_204);
nand U220 (N_220,In_245,In_27);
nand U221 (N_221,In_327,In_110);
and U222 (N_222,In_51,In_437);
and U223 (N_223,In_219,In_342);
and U224 (N_224,In_16,In_253);
nand U225 (N_225,In_748,In_614);
xor U226 (N_226,In_718,In_427);
xor U227 (N_227,In_678,In_531);
or U228 (N_228,In_452,In_210);
nand U229 (N_229,In_278,In_148);
or U230 (N_230,In_68,In_277);
and U231 (N_231,In_643,In_572);
nor U232 (N_232,In_696,In_358);
nor U233 (N_233,In_514,In_39);
nor U234 (N_234,In_261,In_533);
and U235 (N_235,In_354,In_222);
nor U236 (N_236,In_178,In_574);
or U237 (N_237,In_361,In_376);
or U238 (N_238,In_695,In_381);
and U239 (N_239,In_55,In_165);
nand U240 (N_240,In_181,In_487);
or U241 (N_241,In_661,In_54);
nand U242 (N_242,In_182,In_460);
nor U243 (N_243,In_548,In_450);
or U244 (N_244,In_475,In_518);
nor U245 (N_245,In_302,In_353);
xor U246 (N_246,In_461,In_470);
or U247 (N_247,In_203,In_356);
nand U248 (N_248,In_578,In_396);
nor U249 (N_249,In_271,In_79);
or U250 (N_250,In_700,In_725);
or U251 (N_251,In_166,In_318);
and U252 (N_252,In_660,In_303);
xor U253 (N_253,In_493,In_495);
nand U254 (N_254,In_641,In_626);
nor U255 (N_255,In_620,In_373);
or U256 (N_256,In_653,In_441);
nand U257 (N_257,In_96,In_738);
and U258 (N_258,In_671,In_673);
or U259 (N_259,In_106,In_82);
nor U260 (N_260,In_624,In_667);
or U261 (N_261,In_414,In_720);
or U262 (N_262,In_326,In_294);
or U263 (N_263,In_187,In_241);
and U264 (N_264,In_479,In_554);
or U265 (N_265,In_161,In_175);
xor U266 (N_266,In_372,In_114);
nand U267 (N_267,In_76,In_268);
nand U268 (N_268,In_269,In_550);
and U269 (N_269,In_462,In_287);
nor U270 (N_270,In_276,In_692);
nand U271 (N_271,In_699,In_488);
nand U272 (N_272,In_711,In_188);
nor U273 (N_273,In_215,In_730);
or U274 (N_274,In_722,In_138);
and U275 (N_275,In_433,In_143);
and U276 (N_276,In_388,In_706);
nor U277 (N_277,In_399,In_478);
nand U278 (N_278,In_279,In_619);
nor U279 (N_279,In_131,In_480);
nor U280 (N_280,In_367,In_244);
nor U281 (N_281,In_420,In_1);
or U282 (N_282,In_389,In_220);
and U283 (N_283,In_293,In_507);
nor U284 (N_284,In_698,In_93);
nand U285 (N_285,In_111,In_627);
and U286 (N_286,In_415,In_80);
nand U287 (N_287,In_650,In_742);
nand U288 (N_288,In_335,In_60);
nor U289 (N_289,In_428,In_425);
and U290 (N_290,In_697,In_701);
nor U291 (N_291,In_424,In_6);
nor U292 (N_292,In_324,In_707);
nand U293 (N_293,In_569,In_622);
or U294 (N_294,In_712,In_36);
xnor U295 (N_295,In_513,In_679);
or U296 (N_296,In_365,In_446);
nor U297 (N_297,In_186,In_313);
nand U298 (N_298,In_584,In_547);
nand U299 (N_299,In_18,In_216);
or U300 (N_300,In_196,In_339);
and U301 (N_301,In_130,In_411);
nand U302 (N_302,In_649,In_375);
and U303 (N_303,In_35,In_240);
nor U304 (N_304,In_33,In_731);
and U305 (N_305,In_727,In_224);
nand U306 (N_306,In_374,In_634);
and U307 (N_307,In_744,In_340);
nor U308 (N_308,In_647,In_366);
and U309 (N_309,In_543,In_147);
nand U310 (N_310,In_436,In_139);
and U311 (N_311,In_630,In_629);
and U312 (N_312,In_656,In_681);
nand U313 (N_313,In_315,In_515);
nor U314 (N_314,In_393,In_37);
or U315 (N_315,In_557,In_246);
or U316 (N_316,In_541,In_309);
or U317 (N_317,In_134,In_386);
nand U318 (N_318,In_458,In_328);
or U319 (N_319,In_285,In_206);
nor U320 (N_320,In_682,In_316);
and U321 (N_321,In_409,In_628);
and U322 (N_322,In_46,In_291);
or U323 (N_323,In_497,In_50);
or U324 (N_324,In_577,In_498);
or U325 (N_325,In_378,In_672);
nor U326 (N_326,In_398,In_336);
and U327 (N_327,In_664,In_525);
nand U328 (N_328,In_423,In_349);
nor U329 (N_329,In_52,In_259);
and U330 (N_330,In_251,In_362);
nor U331 (N_331,In_435,In_62);
nand U332 (N_332,In_674,In_193);
and U333 (N_333,In_646,In_13);
nor U334 (N_334,In_658,In_559);
or U335 (N_335,In_357,In_443);
nand U336 (N_336,In_238,In_49);
nor U337 (N_337,In_438,In_297);
or U338 (N_338,In_494,In_63);
and U339 (N_339,In_234,In_308);
nor U340 (N_340,In_734,In_359);
or U341 (N_341,In_474,In_145);
and U342 (N_342,In_526,In_686);
xnor U343 (N_343,In_527,In_510);
and U344 (N_344,In_444,In_101);
or U345 (N_345,In_392,In_283);
nand U346 (N_346,In_73,In_351);
and U347 (N_347,In_747,In_213);
or U348 (N_348,In_567,In_12);
nor U349 (N_349,In_128,In_523);
or U350 (N_350,In_25,In_67);
or U351 (N_351,In_100,In_517);
or U352 (N_352,In_264,In_226);
nor U353 (N_353,In_516,In_288);
nor U354 (N_354,In_348,In_144);
nor U355 (N_355,In_137,In_197);
nand U356 (N_356,In_717,In_223);
or U357 (N_357,In_198,In_270);
nor U358 (N_358,In_72,In_192);
nand U359 (N_359,In_289,In_84);
or U360 (N_360,In_160,In_42);
or U361 (N_361,In_163,In_455);
nor U362 (N_362,In_385,In_248);
nor U363 (N_363,In_596,In_273);
and U364 (N_364,In_733,In_632);
or U365 (N_365,In_384,In_102);
nor U366 (N_366,In_171,In_344);
or U367 (N_367,In_88,In_57);
nor U368 (N_368,In_74,In_231);
nor U369 (N_369,In_704,In_242);
or U370 (N_370,In_47,In_59);
or U371 (N_371,In_563,In_741);
nand U372 (N_372,In_558,In_127);
nor U373 (N_373,In_305,In_434);
and U374 (N_374,In_670,In_609);
and U375 (N_375,In_50,In_328);
nand U376 (N_376,In_275,In_232);
nand U377 (N_377,In_290,In_175);
nor U378 (N_378,In_549,In_375);
and U379 (N_379,In_160,In_181);
nor U380 (N_380,In_76,In_672);
nand U381 (N_381,In_1,In_232);
and U382 (N_382,In_619,In_311);
nand U383 (N_383,In_372,In_471);
and U384 (N_384,In_72,In_126);
or U385 (N_385,In_642,In_526);
or U386 (N_386,In_705,In_518);
nand U387 (N_387,In_566,In_12);
nor U388 (N_388,In_396,In_276);
nor U389 (N_389,In_674,In_490);
and U390 (N_390,In_257,In_141);
nand U391 (N_391,In_362,In_353);
nor U392 (N_392,In_483,In_599);
xnor U393 (N_393,In_468,In_474);
and U394 (N_394,In_279,In_231);
nand U395 (N_395,In_340,In_178);
and U396 (N_396,In_594,In_312);
or U397 (N_397,In_113,In_660);
xnor U398 (N_398,In_616,In_306);
nor U399 (N_399,In_701,In_117);
and U400 (N_400,In_747,In_37);
nand U401 (N_401,In_25,In_81);
nor U402 (N_402,In_588,In_413);
or U403 (N_403,In_278,In_8);
nor U404 (N_404,In_313,In_136);
nand U405 (N_405,In_443,In_458);
and U406 (N_406,In_251,In_116);
nor U407 (N_407,In_337,In_727);
nor U408 (N_408,In_292,In_471);
or U409 (N_409,In_704,In_146);
or U410 (N_410,In_75,In_212);
nand U411 (N_411,In_471,In_138);
nor U412 (N_412,In_387,In_327);
or U413 (N_413,In_444,In_395);
or U414 (N_414,In_700,In_13);
or U415 (N_415,In_739,In_589);
nand U416 (N_416,In_703,In_473);
or U417 (N_417,In_434,In_243);
nor U418 (N_418,In_572,In_2);
nand U419 (N_419,In_529,In_101);
and U420 (N_420,In_36,In_506);
nor U421 (N_421,In_371,In_166);
nor U422 (N_422,In_634,In_459);
or U423 (N_423,In_635,In_363);
xnor U424 (N_424,In_321,In_272);
or U425 (N_425,In_216,In_634);
and U426 (N_426,In_339,In_733);
nor U427 (N_427,In_13,In_300);
or U428 (N_428,In_638,In_211);
nand U429 (N_429,In_543,In_69);
xor U430 (N_430,In_40,In_629);
or U431 (N_431,In_589,In_424);
nor U432 (N_432,In_603,In_704);
and U433 (N_433,In_700,In_727);
nand U434 (N_434,In_282,In_188);
or U435 (N_435,In_134,In_515);
and U436 (N_436,In_628,In_426);
nor U437 (N_437,In_741,In_105);
nand U438 (N_438,In_523,In_300);
nand U439 (N_439,In_508,In_690);
nand U440 (N_440,In_468,In_590);
nand U441 (N_441,In_581,In_423);
or U442 (N_442,In_400,In_696);
and U443 (N_443,In_90,In_195);
and U444 (N_444,In_21,In_296);
nor U445 (N_445,In_154,In_78);
or U446 (N_446,In_606,In_549);
and U447 (N_447,In_0,In_641);
nor U448 (N_448,In_711,In_97);
nor U449 (N_449,In_328,In_200);
or U450 (N_450,In_520,In_171);
nor U451 (N_451,In_83,In_275);
and U452 (N_452,In_318,In_91);
nor U453 (N_453,In_551,In_600);
xnor U454 (N_454,In_727,In_115);
nand U455 (N_455,In_40,In_595);
and U456 (N_456,In_655,In_450);
nand U457 (N_457,In_697,In_66);
nor U458 (N_458,In_95,In_627);
nand U459 (N_459,In_251,In_606);
and U460 (N_460,In_419,In_21);
or U461 (N_461,In_509,In_722);
nor U462 (N_462,In_25,In_673);
nor U463 (N_463,In_94,In_117);
and U464 (N_464,In_383,In_344);
nor U465 (N_465,In_630,In_659);
nor U466 (N_466,In_640,In_526);
and U467 (N_467,In_107,In_703);
nor U468 (N_468,In_256,In_23);
and U469 (N_469,In_221,In_147);
nor U470 (N_470,In_653,In_562);
nand U471 (N_471,In_218,In_589);
and U472 (N_472,In_146,In_404);
nor U473 (N_473,In_725,In_17);
nor U474 (N_474,In_193,In_700);
nor U475 (N_475,In_260,In_274);
and U476 (N_476,In_290,In_149);
nand U477 (N_477,In_424,In_123);
nand U478 (N_478,In_364,In_174);
or U479 (N_479,In_721,In_150);
nor U480 (N_480,In_509,In_203);
or U481 (N_481,In_331,In_742);
or U482 (N_482,In_423,In_214);
and U483 (N_483,In_680,In_64);
or U484 (N_484,In_220,In_377);
nand U485 (N_485,In_533,In_602);
xnor U486 (N_486,In_523,In_209);
or U487 (N_487,In_378,In_744);
or U488 (N_488,In_110,In_25);
nand U489 (N_489,In_608,In_345);
nand U490 (N_490,In_670,In_56);
nand U491 (N_491,In_709,In_716);
nor U492 (N_492,In_86,In_33);
nor U493 (N_493,In_673,In_565);
nor U494 (N_494,In_365,In_336);
or U495 (N_495,In_674,In_132);
or U496 (N_496,In_322,In_491);
nor U497 (N_497,In_439,In_641);
or U498 (N_498,In_358,In_97);
nor U499 (N_499,In_335,In_59);
nor U500 (N_500,N_345,N_357);
or U501 (N_501,N_81,N_48);
or U502 (N_502,N_175,N_335);
and U503 (N_503,N_182,N_117);
and U504 (N_504,N_370,N_312);
and U505 (N_505,N_79,N_39);
or U506 (N_506,N_161,N_342);
nand U507 (N_507,N_405,N_185);
or U508 (N_508,N_91,N_465);
or U509 (N_509,N_383,N_230);
nand U510 (N_510,N_356,N_494);
nor U511 (N_511,N_226,N_74);
and U512 (N_512,N_415,N_401);
and U513 (N_513,N_206,N_111);
and U514 (N_514,N_18,N_470);
nand U515 (N_515,N_426,N_15);
nor U516 (N_516,N_463,N_489);
or U517 (N_517,N_200,N_316);
and U518 (N_518,N_390,N_322);
or U519 (N_519,N_68,N_73);
or U520 (N_520,N_381,N_134);
and U521 (N_521,N_58,N_139);
nor U522 (N_522,N_155,N_268);
or U523 (N_523,N_170,N_121);
nand U524 (N_524,N_8,N_475);
and U525 (N_525,N_309,N_5);
and U526 (N_526,N_481,N_329);
or U527 (N_527,N_246,N_374);
nand U528 (N_528,N_499,N_62);
nand U529 (N_529,N_317,N_44);
nor U530 (N_530,N_37,N_343);
and U531 (N_531,N_416,N_326);
nand U532 (N_532,N_430,N_113);
nand U533 (N_533,N_156,N_496);
or U534 (N_534,N_314,N_266);
nor U535 (N_535,N_320,N_477);
or U536 (N_536,N_131,N_339);
xor U537 (N_537,N_341,N_212);
nor U538 (N_538,N_20,N_307);
nor U539 (N_539,N_225,N_201);
nand U540 (N_540,N_86,N_162);
or U541 (N_541,N_262,N_141);
and U542 (N_542,N_105,N_11);
or U543 (N_543,N_304,N_493);
or U544 (N_544,N_178,N_420);
and U545 (N_545,N_99,N_358);
nand U546 (N_546,N_248,N_97);
nand U547 (N_547,N_172,N_176);
or U548 (N_548,N_61,N_197);
and U549 (N_549,N_330,N_63);
xnor U550 (N_550,N_461,N_64);
or U551 (N_551,N_350,N_360);
and U552 (N_552,N_462,N_362);
nand U553 (N_553,N_336,N_16);
nor U554 (N_554,N_310,N_245);
nor U555 (N_555,N_421,N_261);
or U556 (N_556,N_455,N_491);
nor U557 (N_557,N_154,N_398);
and U558 (N_558,N_215,N_332);
and U559 (N_559,N_236,N_292);
and U560 (N_560,N_387,N_267);
nor U561 (N_561,N_471,N_300);
nand U562 (N_562,N_424,N_19);
nor U563 (N_563,N_67,N_497);
nand U564 (N_564,N_393,N_209);
or U565 (N_565,N_204,N_411);
nand U566 (N_566,N_114,N_190);
nor U567 (N_567,N_194,N_177);
nand U568 (N_568,N_394,N_433);
nand U569 (N_569,N_80,N_273);
nor U570 (N_570,N_253,N_364);
and U571 (N_571,N_66,N_340);
and U572 (N_572,N_102,N_214);
nor U573 (N_573,N_371,N_137);
nor U574 (N_574,N_227,N_346);
nand U575 (N_575,N_363,N_223);
or U576 (N_576,N_419,N_382);
nor U577 (N_577,N_440,N_129);
nand U578 (N_578,N_112,N_31);
nor U579 (N_579,N_338,N_408);
or U580 (N_580,N_232,N_286);
xor U581 (N_581,N_365,N_359);
and U582 (N_582,N_115,N_439);
and U583 (N_583,N_250,N_391);
or U584 (N_584,N_375,N_34);
and U585 (N_585,N_294,N_355);
nand U586 (N_586,N_485,N_168);
and U587 (N_587,N_120,N_95);
and U588 (N_588,N_325,N_380);
or U589 (N_589,N_327,N_219);
nand U590 (N_590,N_229,N_376);
and U591 (N_591,N_98,N_136);
nor U592 (N_592,N_422,N_234);
and U593 (N_593,N_207,N_75);
nor U594 (N_594,N_474,N_196);
and U595 (N_595,N_347,N_349);
and U596 (N_596,N_189,N_438);
nor U597 (N_597,N_71,N_466);
nand U598 (N_598,N_259,N_368);
or U599 (N_599,N_457,N_23);
nand U600 (N_600,N_313,N_93);
nand U601 (N_601,N_452,N_293);
or U602 (N_602,N_96,N_441);
nand U603 (N_603,N_388,N_445);
or U604 (N_604,N_284,N_84);
and U605 (N_605,N_231,N_145);
and U606 (N_606,N_498,N_128);
and U607 (N_607,N_399,N_319);
nand U608 (N_608,N_249,N_255);
nand U609 (N_609,N_331,N_290);
or U610 (N_610,N_472,N_144);
and U611 (N_611,N_397,N_334);
and U612 (N_612,N_151,N_51);
and U613 (N_613,N_198,N_6);
and U614 (N_614,N_33,N_119);
and U615 (N_615,N_403,N_38);
or U616 (N_616,N_417,N_54);
nor U617 (N_617,N_379,N_274);
or U618 (N_618,N_252,N_389);
nor U619 (N_619,N_72,N_431);
or U620 (N_620,N_203,N_402);
and U621 (N_621,N_278,N_427);
and U622 (N_622,N_239,N_409);
nor U623 (N_623,N_40,N_451);
nor U624 (N_624,N_160,N_352);
or U625 (N_625,N_14,N_437);
nand U626 (N_626,N_469,N_432);
or U627 (N_627,N_412,N_218);
or U628 (N_628,N_473,N_264);
nor U629 (N_629,N_413,N_49);
and U630 (N_630,N_276,N_163);
nor U631 (N_631,N_351,N_159);
nor U632 (N_632,N_88,N_354);
nand U633 (N_633,N_164,N_378);
nand U634 (N_634,N_140,N_407);
or U635 (N_635,N_46,N_385);
nor U636 (N_636,N_187,N_444);
nand U637 (N_637,N_251,N_130);
nand U638 (N_638,N_297,N_254);
and U639 (N_639,N_180,N_302);
nand U640 (N_640,N_125,N_205);
nor U641 (N_641,N_256,N_487);
and U642 (N_642,N_386,N_90);
or U643 (N_643,N_202,N_109);
nand U644 (N_644,N_257,N_57);
xor U645 (N_645,N_436,N_495);
or U646 (N_646,N_484,N_324);
or U647 (N_647,N_0,N_282);
or U648 (N_648,N_56,N_344);
and U649 (N_649,N_305,N_60);
or U650 (N_650,N_42,N_106);
nor U651 (N_651,N_443,N_428);
nor U652 (N_652,N_240,N_157);
nor U653 (N_653,N_4,N_29);
or U654 (N_654,N_216,N_132);
or U655 (N_655,N_184,N_9);
nand U656 (N_656,N_315,N_400);
and U657 (N_657,N_287,N_279);
or U658 (N_658,N_83,N_247);
nand U659 (N_659,N_321,N_27);
nand U660 (N_660,N_281,N_147);
nor U661 (N_661,N_480,N_25);
and U662 (N_662,N_92,N_126);
xor U663 (N_663,N_392,N_183);
or U664 (N_664,N_384,N_211);
nor U665 (N_665,N_260,N_486);
nor U666 (N_666,N_78,N_45);
or U667 (N_667,N_10,N_468);
xor U668 (N_668,N_296,N_456);
nor U669 (N_669,N_221,N_453);
nor U670 (N_670,N_446,N_283);
or U671 (N_671,N_337,N_224);
and U672 (N_672,N_241,N_146);
nand U673 (N_673,N_244,N_169);
nand U674 (N_674,N_22,N_373);
xor U675 (N_675,N_77,N_318);
nor U676 (N_676,N_299,N_53);
and U677 (N_677,N_82,N_7);
nor U678 (N_678,N_423,N_333);
or U679 (N_679,N_2,N_116);
nand U680 (N_680,N_165,N_142);
nor U681 (N_681,N_32,N_150);
or U682 (N_682,N_482,N_306);
or U683 (N_683,N_133,N_174);
nor U684 (N_684,N_149,N_65);
nor U685 (N_685,N_17,N_108);
and U686 (N_686,N_328,N_191);
nor U687 (N_687,N_166,N_429);
or U688 (N_688,N_186,N_454);
xor U689 (N_689,N_195,N_30);
xor U690 (N_690,N_24,N_442);
and U691 (N_691,N_28,N_217);
nor U692 (N_692,N_410,N_26);
nor U693 (N_693,N_107,N_89);
and U694 (N_694,N_447,N_483);
or U695 (N_695,N_87,N_353);
or U696 (N_696,N_396,N_348);
nor U697 (N_697,N_476,N_70);
and U698 (N_698,N_270,N_488);
or U699 (N_699,N_171,N_41);
nor U700 (N_700,N_404,N_13);
nand U701 (N_701,N_377,N_269);
and U702 (N_702,N_47,N_289);
or U703 (N_703,N_414,N_76);
nand U704 (N_704,N_308,N_479);
or U705 (N_705,N_213,N_210);
or U706 (N_706,N_21,N_94);
and U707 (N_707,N_311,N_1);
or U708 (N_708,N_242,N_3);
or U709 (N_709,N_50,N_59);
and U710 (N_710,N_179,N_208);
nand U711 (N_711,N_43,N_425);
or U712 (N_712,N_272,N_104);
or U713 (N_713,N_118,N_369);
nand U714 (N_714,N_366,N_173);
and U715 (N_715,N_492,N_271);
nand U716 (N_716,N_291,N_124);
nand U717 (N_717,N_55,N_181);
nor U718 (N_718,N_323,N_235);
or U719 (N_719,N_69,N_52);
and U720 (N_720,N_285,N_193);
and U721 (N_721,N_367,N_103);
nor U722 (N_722,N_418,N_135);
nor U723 (N_723,N_192,N_143);
nor U724 (N_724,N_237,N_228);
or U725 (N_725,N_122,N_406);
nor U726 (N_726,N_490,N_148);
nor U727 (N_727,N_467,N_288);
nand U728 (N_728,N_85,N_361);
nand U729 (N_729,N_298,N_464);
or U730 (N_730,N_280,N_458);
nor U731 (N_731,N_12,N_158);
or U732 (N_732,N_295,N_199);
nand U733 (N_733,N_372,N_123);
xor U734 (N_734,N_101,N_110);
nor U735 (N_735,N_238,N_434);
and U736 (N_736,N_265,N_127);
or U737 (N_737,N_233,N_167);
and U738 (N_738,N_275,N_263);
nor U739 (N_739,N_220,N_277);
or U740 (N_740,N_395,N_243);
or U741 (N_741,N_435,N_152);
xor U742 (N_742,N_36,N_188);
and U743 (N_743,N_258,N_450);
nand U744 (N_744,N_153,N_460);
or U745 (N_745,N_303,N_301);
nor U746 (N_746,N_459,N_448);
and U747 (N_747,N_478,N_138);
nand U748 (N_748,N_100,N_222);
or U749 (N_749,N_35,N_449);
and U750 (N_750,N_456,N_333);
and U751 (N_751,N_485,N_396);
nor U752 (N_752,N_129,N_234);
nor U753 (N_753,N_459,N_265);
and U754 (N_754,N_118,N_370);
nor U755 (N_755,N_317,N_366);
nand U756 (N_756,N_367,N_43);
or U757 (N_757,N_487,N_60);
nand U758 (N_758,N_286,N_483);
nor U759 (N_759,N_130,N_426);
or U760 (N_760,N_231,N_224);
nand U761 (N_761,N_258,N_134);
or U762 (N_762,N_396,N_115);
nand U763 (N_763,N_229,N_297);
and U764 (N_764,N_177,N_184);
nand U765 (N_765,N_201,N_125);
nand U766 (N_766,N_472,N_477);
and U767 (N_767,N_425,N_32);
nand U768 (N_768,N_408,N_319);
and U769 (N_769,N_486,N_495);
and U770 (N_770,N_23,N_113);
nor U771 (N_771,N_376,N_142);
or U772 (N_772,N_41,N_318);
or U773 (N_773,N_164,N_168);
and U774 (N_774,N_40,N_212);
or U775 (N_775,N_147,N_188);
and U776 (N_776,N_321,N_258);
or U777 (N_777,N_51,N_487);
and U778 (N_778,N_215,N_417);
or U779 (N_779,N_9,N_24);
nor U780 (N_780,N_278,N_249);
nand U781 (N_781,N_81,N_446);
and U782 (N_782,N_483,N_322);
nand U783 (N_783,N_498,N_67);
nor U784 (N_784,N_276,N_36);
and U785 (N_785,N_422,N_368);
and U786 (N_786,N_144,N_136);
and U787 (N_787,N_453,N_371);
or U788 (N_788,N_411,N_452);
nand U789 (N_789,N_304,N_52);
and U790 (N_790,N_312,N_233);
or U791 (N_791,N_258,N_487);
or U792 (N_792,N_419,N_479);
nor U793 (N_793,N_351,N_117);
or U794 (N_794,N_248,N_474);
nand U795 (N_795,N_319,N_209);
and U796 (N_796,N_479,N_406);
nand U797 (N_797,N_405,N_26);
and U798 (N_798,N_437,N_482);
nor U799 (N_799,N_474,N_62);
or U800 (N_800,N_67,N_213);
and U801 (N_801,N_273,N_65);
or U802 (N_802,N_143,N_480);
and U803 (N_803,N_103,N_362);
or U804 (N_804,N_405,N_206);
xnor U805 (N_805,N_475,N_225);
or U806 (N_806,N_61,N_446);
or U807 (N_807,N_15,N_26);
or U808 (N_808,N_289,N_491);
or U809 (N_809,N_101,N_166);
nor U810 (N_810,N_149,N_451);
and U811 (N_811,N_79,N_311);
or U812 (N_812,N_242,N_63);
and U813 (N_813,N_244,N_243);
or U814 (N_814,N_458,N_137);
xnor U815 (N_815,N_496,N_84);
nand U816 (N_816,N_493,N_462);
and U817 (N_817,N_245,N_128);
and U818 (N_818,N_347,N_35);
nand U819 (N_819,N_134,N_268);
nor U820 (N_820,N_390,N_161);
or U821 (N_821,N_358,N_9);
or U822 (N_822,N_11,N_164);
nand U823 (N_823,N_116,N_57);
or U824 (N_824,N_480,N_443);
nand U825 (N_825,N_178,N_197);
and U826 (N_826,N_137,N_126);
or U827 (N_827,N_173,N_226);
and U828 (N_828,N_223,N_153);
or U829 (N_829,N_5,N_12);
or U830 (N_830,N_198,N_82);
and U831 (N_831,N_282,N_267);
or U832 (N_832,N_141,N_165);
nand U833 (N_833,N_411,N_226);
nor U834 (N_834,N_136,N_56);
and U835 (N_835,N_20,N_21);
or U836 (N_836,N_208,N_176);
nand U837 (N_837,N_55,N_291);
and U838 (N_838,N_496,N_448);
or U839 (N_839,N_465,N_100);
nor U840 (N_840,N_158,N_121);
nand U841 (N_841,N_284,N_235);
nand U842 (N_842,N_415,N_327);
nor U843 (N_843,N_407,N_229);
nand U844 (N_844,N_52,N_274);
nand U845 (N_845,N_245,N_150);
nor U846 (N_846,N_309,N_338);
and U847 (N_847,N_259,N_254);
and U848 (N_848,N_28,N_289);
and U849 (N_849,N_57,N_403);
and U850 (N_850,N_421,N_35);
or U851 (N_851,N_28,N_450);
or U852 (N_852,N_477,N_154);
nor U853 (N_853,N_33,N_41);
and U854 (N_854,N_142,N_295);
nand U855 (N_855,N_283,N_390);
or U856 (N_856,N_124,N_461);
nand U857 (N_857,N_180,N_286);
nand U858 (N_858,N_175,N_329);
nand U859 (N_859,N_244,N_332);
nand U860 (N_860,N_242,N_64);
and U861 (N_861,N_376,N_498);
nor U862 (N_862,N_109,N_54);
nor U863 (N_863,N_106,N_348);
nor U864 (N_864,N_484,N_175);
and U865 (N_865,N_108,N_36);
or U866 (N_866,N_114,N_63);
nor U867 (N_867,N_440,N_488);
nor U868 (N_868,N_170,N_223);
nor U869 (N_869,N_369,N_416);
nand U870 (N_870,N_322,N_427);
xnor U871 (N_871,N_313,N_309);
nand U872 (N_872,N_367,N_170);
nand U873 (N_873,N_398,N_298);
nor U874 (N_874,N_91,N_271);
or U875 (N_875,N_41,N_302);
and U876 (N_876,N_64,N_224);
nor U877 (N_877,N_298,N_471);
xor U878 (N_878,N_481,N_173);
nor U879 (N_879,N_79,N_462);
or U880 (N_880,N_80,N_55);
xor U881 (N_881,N_257,N_308);
and U882 (N_882,N_483,N_85);
nand U883 (N_883,N_128,N_82);
nor U884 (N_884,N_484,N_43);
or U885 (N_885,N_200,N_420);
and U886 (N_886,N_285,N_459);
nor U887 (N_887,N_360,N_321);
nor U888 (N_888,N_69,N_262);
and U889 (N_889,N_355,N_210);
nand U890 (N_890,N_113,N_320);
nand U891 (N_891,N_358,N_199);
nand U892 (N_892,N_458,N_110);
xnor U893 (N_893,N_354,N_446);
and U894 (N_894,N_130,N_430);
nand U895 (N_895,N_153,N_463);
nand U896 (N_896,N_1,N_106);
and U897 (N_897,N_269,N_241);
or U898 (N_898,N_388,N_273);
or U899 (N_899,N_255,N_108);
nand U900 (N_900,N_382,N_323);
nand U901 (N_901,N_79,N_25);
nor U902 (N_902,N_118,N_357);
nand U903 (N_903,N_170,N_231);
and U904 (N_904,N_201,N_161);
and U905 (N_905,N_247,N_88);
nand U906 (N_906,N_183,N_115);
or U907 (N_907,N_268,N_404);
or U908 (N_908,N_168,N_315);
nor U909 (N_909,N_317,N_304);
and U910 (N_910,N_132,N_305);
xor U911 (N_911,N_361,N_206);
nor U912 (N_912,N_26,N_194);
nor U913 (N_913,N_489,N_477);
nor U914 (N_914,N_84,N_382);
or U915 (N_915,N_338,N_173);
nor U916 (N_916,N_336,N_268);
nor U917 (N_917,N_244,N_349);
or U918 (N_918,N_325,N_443);
or U919 (N_919,N_122,N_151);
nor U920 (N_920,N_233,N_393);
nor U921 (N_921,N_162,N_52);
or U922 (N_922,N_225,N_419);
or U923 (N_923,N_319,N_178);
or U924 (N_924,N_197,N_249);
nand U925 (N_925,N_264,N_412);
nor U926 (N_926,N_234,N_8);
and U927 (N_927,N_239,N_465);
nand U928 (N_928,N_404,N_402);
or U929 (N_929,N_83,N_148);
nor U930 (N_930,N_442,N_206);
nor U931 (N_931,N_55,N_21);
nand U932 (N_932,N_143,N_319);
or U933 (N_933,N_53,N_495);
and U934 (N_934,N_109,N_303);
nor U935 (N_935,N_314,N_381);
xor U936 (N_936,N_154,N_196);
nor U937 (N_937,N_267,N_113);
or U938 (N_938,N_454,N_74);
nor U939 (N_939,N_137,N_300);
or U940 (N_940,N_474,N_264);
or U941 (N_941,N_305,N_300);
nor U942 (N_942,N_191,N_93);
nand U943 (N_943,N_175,N_131);
nor U944 (N_944,N_219,N_347);
or U945 (N_945,N_264,N_395);
or U946 (N_946,N_21,N_345);
nand U947 (N_947,N_3,N_397);
or U948 (N_948,N_420,N_37);
and U949 (N_949,N_296,N_313);
nor U950 (N_950,N_237,N_257);
nand U951 (N_951,N_139,N_175);
nand U952 (N_952,N_276,N_232);
nor U953 (N_953,N_463,N_328);
nand U954 (N_954,N_335,N_460);
nor U955 (N_955,N_221,N_474);
nand U956 (N_956,N_250,N_189);
or U957 (N_957,N_434,N_272);
nor U958 (N_958,N_347,N_332);
nor U959 (N_959,N_482,N_214);
nor U960 (N_960,N_242,N_162);
nand U961 (N_961,N_239,N_347);
or U962 (N_962,N_270,N_29);
nand U963 (N_963,N_373,N_262);
nor U964 (N_964,N_472,N_129);
xor U965 (N_965,N_417,N_463);
nand U966 (N_966,N_173,N_126);
and U967 (N_967,N_227,N_71);
nor U968 (N_968,N_331,N_199);
nand U969 (N_969,N_204,N_447);
nand U970 (N_970,N_224,N_170);
and U971 (N_971,N_418,N_133);
nand U972 (N_972,N_69,N_74);
nor U973 (N_973,N_291,N_495);
xnor U974 (N_974,N_226,N_265);
nand U975 (N_975,N_70,N_181);
nor U976 (N_976,N_155,N_75);
and U977 (N_977,N_348,N_298);
nand U978 (N_978,N_356,N_239);
nor U979 (N_979,N_325,N_496);
and U980 (N_980,N_225,N_170);
nor U981 (N_981,N_466,N_22);
or U982 (N_982,N_256,N_435);
nor U983 (N_983,N_407,N_32);
and U984 (N_984,N_189,N_352);
nor U985 (N_985,N_36,N_205);
nor U986 (N_986,N_245,N_322);
xor U987 (N_987,N_210,N_29);
nand U988 (N_988,N_497,N_72);
nor U989 (N_989,N_92,N_21);
nor U990 (N_990,N_89,N_243);
or U991 (N_991,N_243,N_458);
nand U992 (N_992,N_425,N_378);
nand U993 (N_993,N_379,N_325);
and U994 (N_994,N_216,N_195);
nand U995 (N_995,N_44,N_403);
nand U996 (N_996,N_99,N_141);
nand U997 (N_997,N_423,N_109);
nor U998 (N_998,N_53,N_124);
and U999 (N_999,N_188,N_53);
nand U1000 (N_1000,N_516,N_790);
or U1001 (N_1001,N_542,N_699);
nand U1002 (N_1002,N_566,N_873);
xor U1003 (N_1003,N_593,N_978);
xor U1004 (N_1004,N_786,N_579);
and U1005 (N_1005,N_738,N_961);
and U1006 (N_1006,N_560,N_835);
nor U1007 (N_1007,N_854,N_622);
and U1008 (N_1008,N_728,N_616);
and U1009 (N_1009,N_583,N_595);
and U1010 (N_1010,N_807,N_809);
and U1011 (N_1011,N_685,N_824);
nand U1012 (N_1012,N_505,N_554);
nor U1013 (N_1013,N_735,N_999);
nand U1014 (N_1014,N_906,N_832);
or U1015 (N_1015,N_858,N_651);
and U1016 (N_1016,N_507,N_848);
and U1017 (N_1017,N_925,N_708);
nand U1018 (N_1018,N_633,N_791);
nor U1019 (N_1019,N_747,N_796);
nor U1020 (N_1020,N_888,N_879);
nor U1021 (N_1021,N_751,N_753);
and U1022 (N_1022,N_506,N_909);
or U1023 (N_1023,N_760,N_894);
nor U1024 (N_1024,N_823,N_567);
and U1025 (N_1025,N_581,N_998);
nand U1026 (N_1026,N_818,N_795);
nor U1027 (N_1027,N_676,N_953);
nor U1028 (N_1028,N_997,N_712);
or U1029 (N_1029,N_926,N_526);
nor U1030 (N_1030,N_577,N_821);
nor U1031 (N_1031,N_756,N_922);
or U1032 (N_1032,N_548,N_833);
nor U1033 (N_1033,N_899,N_632);
and U1034 (N_1034,N_981,N_945);
or U1035 (N_1035,N_549,N_752);
nor U1036 (N_1036,N_519,N_544);
or U1037 (N_1037,N_724,N_940);
and U1038 (N_1038,N_564,N_580);
and U1039 (N_1039,N_794,N_606);
nor U1040 (N_1040,N_618,N_895);
nor U1041 (N_1041,N_864,N_501);
nor U1042 (N_1042,N_775,N_810);
or U1043 (N_1043,N_929,N_538);
nand U1044 (N_1044,N_647,N_778);
or U1045 (N_1045,N_770,N_827);
and U1046 (N_1046,N_545,N_524);
nor U1047 (N_1047,N_837,N_784);
nor U1048 (N_1048,N_812,N_903);
and U1049 (N_1049,N_508,N_912);
nand U1050 (N_1050,N_802,N_806);
and U1051 (N_1051,N_570,N_660);
xor U1052 (N_1052,N_740,N_653);
nor U1053 (N_1053,N_748,N_502);
nor U1054 (N_1054,N_512,N_757);
xor U1055 (N_1055,N_594,N_587);
and U1056 (N_1056,N_711,N_522);
and U1057 (N_1057,N_558,N_734);
or U1058 (N_1058,N_630,N_971);
nand U1059 (N_1059,N_596,N_852);
and U1060 (N_1060,N_591,N_772);
nor U1061 (N_1061,N_813,N_541);
or U1062 (N_1062,N_575,N_697);
nor U1063 (N_1063,N_834,N_706);
nand U1064 (N_1064,N_586,N_801);
and U1065 (N_1065,N_950,N_931);
nand U1066 (N_1066,N_627,N_975);
or U1067 (N_1067,N_898,N_987);
and U1068 (N_1068,N_571,N_553);
and U1069 (N_1069,N_543,N_829);
nand U1070 (N_1070,N_880,N_698);
or U1071 (N_1071,N_882,N_709);
nor U1072 (N_1072,N_639,N_762);
or U1073 (N_1073,N_655,N_992);
and U1074 (N_1074,N_608,N_914);
or U1075 (N_1075,N_764,N_675);
nand U1076 (N_1076,N_635,N_642);
xor U1077 (N_1077,N_759,N_517);
or U1078 (N_1078,N_584,N_533);
nand U1079 (N_1079,N_640,N_754);
or U1080 (N_1080,N_849,N_933);
xor U1081 (N_1081,N_695,N_868);
xnor U1082 (N_1082,N_948,N_907);
and U1083 (N_1083,N_787,N_648);
nand U1084 (N_1084,N_979,N_645);
or U1085 (N_1085,N_856,N_831);
and U1086 (N_1086,N_705,N_908);
nand U1087 (N_1087,N_977,N_958);
nand U1088 (N_1088,N_928,N_550);
nand U1089 (N_1089,N_750,N_563);
and U1090 (N_1090,N_511,N_990);
nand U1091 (N_1091,N_681,N_730);
nor U1092 (N_1092,N_718,N_669);
nand U1093 (N_1093,N_703,N_621);
xor U1094 (N_1094,N_902,N_582);
nor U1095 (N_1095,N_599,N_878);
nand U1096 (N_1096,N_561,N_930);
or U1097 (N_1097,N_985,N_889);
and U1098 (N_1098,N_644,N_780);
nand U1099 (N_1099,N_598,N_969);
and U1100 (N_1100,N_634,N_991);
or U1101 (N_1101,N_601,N_717);
nand U1102 (N_1102,N_604,N_671);
and U1103 (N_1103,N_804,N_819);
or U1104 (N_1104,N_901,N_939);
or U1105 (N_1105,N_897,N_528);
or U1106 (N_1106,N_811,N_638);
and U1107 (N_1107,N_741,N_693);
nand U1108 (N_1108,N_947,N_797);
or U1109 (N_1109,N_746,N_624);
or U1110 (N_1110,N_523,N_876);
nor U1111 (N_1111,N_520,N_988);
or U1112 (N_1112,N_518,N_782);
or U1113 (N_1113,N_667,N_905);
or U1114 (N_1114,N_531,N_689);
nor U1115 (N_1115,N_994,N_619);
nand U1116 (N_1116,N_605,N_715);
nor U1117 (N_1117,N_785,N_843);
nand U1118 (N_1118,N_860,N_836);
nor U1119 (N_1119,N_968,N_946);
or U1120 (N_1120,N_921,N_817);
nor U1121 (N_1121,N_870,N_557);
or U1122 (N_1122,N_918,N_589);
nor U1123 (N_1123,N_983,N_504);
nor U1124 (N_1124,N_943,N_960);
nor U1125 (N_1125,N_828,N_736);
nor U1126 (N_1126,N_666,N_949);
nor U1127 (N_1127,N_710,N_919);
nand U1128 (N_1128,N_585,N_840);
nand U1129 (N_1129,N_765,N_920);
nand U1130 (N_1130,N_957,N_989);
or U1131 (N_1131,N_611,N_937);
nor U1132 (N_1132,N_536,N_963);
nand U1133 (N_1133,N_745,N_716);
nor U1134 (N_1134,N_749,N_590);
and U1135 (N_1135,N_934,N_702);
and U1136 (N_1136,N_808,N_515);
or U1137 (N_1137,N_965,N_521);
nor U1138 (N_1138,N_737,N_527);
nand U1139 (N_1139,N_938,N_800);
xor U1140 (N_1140,N_964,N_609);
and U1141 (N_1141,N_652,N_942);
and U1142 (N_1142,N_628,N_683);
nand U1143 (N_1143,N_986,N_534);
nand U1144 (N_1144,N_714,N_851);
or U1145 (N_1145,N_955,N_962);
nand U1146 (N_1146,N_614,N_803);
and U1147 (N_1147,N_867,N_654);
nand U1148 (N_1148,N_911,N_838);
nand U1149 (N_1149,N_610,N_631);
or U1150 (N_1150,N_993,N_670);
or U1151 (N_1151,N_767,N_916);
nor U1152 (N_1152,N_913,N_874);
and U1153 (N_1153,N_673,N_662);
and U1154 (N_1154,N_719,N_691);
nand U1155 (N_1155,N_727,N_869);
or U1156 (N_1156,N_646,N_766);
and U1157 (N_1157,N_830,N_841);
and U1158 (N_1158,N_853,N_742);
nand U1159 (N_1159,N_664,N_863);
and U1160 (N_1160,N_617,N_825);
nor U1161 (N_1161,N_798,N_602);
nor U1162 (N_1162,N_626,N_720);
nor U1163 (N_1163,N_744,N_547);
and U1164 (N_1164,N_540,N_615);
nand U1165 (N_1165,N_551,N_674);
nand U1166 (N_1166,N_915,N_974);
and U1167 (N_1167,N_893,N_886);
or U1168 (N_1168,N_684,N_677);
and U1169 (N_1169,N_578,N_793);
and U1170 (N_1170,N_924,N_773);
nor U1171 (N_1171,N_967,N_984);
and U1172 (N_1172,N_569,N_612);
or U1173 (N_1173,N_771,N_559);
nand U1174 (N_1174,N_855,N_530);
nor U1175 (N_1175,N_845,N_661);
and U1176 (N_1176,N_679,N_696);
nor U1177 (N_1177,N_509,N_537);
nand U1178 (N_1178,N_789,N_733);
nor U1179 (N_1179,N_872,N_625);
nand U1180 (N_1180,N_663,N_763);
nor U1181 (N_1181,N_603,N_844);
nand U1182 (N_1182,N_959,N_755);
nand U1183 (N_1183,N_781,N_866);
nand U1184 (N_1184,N_820,N_643);
or U1185 (N_1185,N_743,N_917);
nand U1186 (N_1186,N_779,N_758);
nand U1187 (N_1187,N_936,N_672);
or U1188 (N_1188,N_503,N_732);
xnor U1189 (N_1189,N_692,N_850);
nor U1190 (N_1190,N_980,N_857);
and U1191 (N_1191,N_970,N_731);
and U1192 (N_1192,N_588,N_686);
nor U1193 (N_1193,N_546,N_885);
nor U1194 (N_1194,N_532,N_552);
or U1195 (N_1195,N_871,N_568);
or U1196 (N_1196,N_613,N_814);
nand U1197 (N_1197,N_707,N_768);
nor U1198 (N_1198,N_805,N_956);
nand U1199 (N_1199,N_713,N_556);
nand U1200 (N_1200,N_881,N_637);
and U1201 (N_1201,N_792,N_839);
xor U1202 (N_1202,N_600,N_761);
and U1203 (N_1203,N_973,N_597);
nor U1204 (N_1204,N_951,N_539);
nor U1205 (N_1205,N_700,N_525);
or U1206 (N_1206,N_900,N_826);
nand U1207 (N_1207,N_500,N_641);
or U1208 (N_1208,N_783,N_776);
and U1209 (N_1209,N_650,N_892);
nand U1210 (N_1210,N_694,N_572);
and U1211 (N_1211,N_799,N_890);
and U1212 (N_1212,N_620,N_510);
or U1213 (N_1213,N_529,N_573);
nand U1214 (N_1214,N_680,N_865);
and U1215 (N_1215,N_636,N_535);
or U1216 (N_1216,N_976,N_690);
or U1217 (N_1217,N_995,N_847);
nor U1218 (N_1218,N_875,N_927);
nor U1219 (N_1219,N_877,N_678);
xnor U1220 (N_1220,N_722,N_859);
nor U1221 (N_1221,N_658,N_944);
or U1222 (N_1222,N_952,N_896);
or U1223 (N_1223,N_665,N_701);
and U1224 (N_1224,N_576,N_996);
or U1225 (N_1225,N_688,N_954);
nor U1226 (N_1226,N_788,N_982);
and U1227 (N_1227,N_846,N_729);
nand U1228 (N_1228,N_562,N_629);
nor U1229 (N_1229,N_887,N_607);
nand U1230 (N_1230,N_514,N_966);
nand U1231 (N_1231,N_972,N_862);
nor U1232 (N_1232,N_769,N_592);
or U1233 (N_1233,N_910,N_656);
nor U1234 (N_1234,N_941,N_842);
nand U1235 (N_1235,N_721,N_777);
or U1236 (N_1236,N_816,N_623);
or U1237 (N_1237,N_565,N_935);
or U1238 (N_1238,N_657,N_659);
nand U1239 (N_1239,N_513,N_861);
nor U1240 (N_1240,N_822,N_682);
nand U1241 (N_1241,N_891,N_932);
nor U1242 (N_1242,N_668,N_704);
and U1243 (N_1243,N_574,N_883);
or U1244 (N_1244,N_774,N_739);
nand U1245 (N_1245,N_555,N_725);
nor U1246 (N_1246,N_904,N_687);
nor U1247 (N_1247,N_884,N_723);
nand U1248 (N_1248,N_923,N_726);
or U1249 (N_1249,N_815,N_649);
and U1250 (N_1250,N_773,N_736);
and U1251 (N_1251,N_591,N_507);
nor U1252 (N_1252,N_793,N_670);
nand U1253 (N_1253,N_817,N_972);
or U1254 (N_1254,N_803,N_870);
and U1255 (N_1255,N_611,N_892);
or U1256 (N_1256,N_778,N_981);
and U1257 (N_1257,N_846,N_937);
nor U1258 (N_1258,N_848,N_815);
and U1259 (N_1259,N_945,N_697);
and U1260 (N_1260,N_862,N_646);
nor U1261 (N_1261,N_758,N_674);
nand U1262 (N_1262,N_591,N_796);
nand U1263 (N_1263,N_536,N_556);
and U1264 (N_1264,N_807,N_526);
or U1265 (N_1265,N_578,N_914);
nor U1266 (N_1266,N_577,N_571);
nand U1267 (N_1267,N_952,N_931);
nand U1268 (N_1268,N_588,N_814);
or U1269 (N_1269,N_601,N_549);
nand U1270 (N_1270,N_848,N_504);
or U1271 (N_1271,N_534,N_673);
or U1272 (N_1272,N_839,N_940);
or U1273 (N_1273,N_753,N_987);
nor U1274 (N_1274,N_569,N_845);
and U1275 (N_1275,N_548,N_665);
or U1276 (N_1276,N_949,N_869);
or U1277 (N_1277,N_760,N_679);
nor U1278 (N_1278,N_851,N_647);
nor U1279 (N_1279,N_808,N_928);
or U1280 (N_1280,N_856,N_652);
and U1281 (N_1281,N_573,N_680);
nor U1282 (N_1282,N_752,N_664);
or U1283 (N_1283,N_983,N_550);
or U1284 (N_1284,N_929,N_712);
or U1285 (N_1285,N_994,N_841);
or U1286 (N_1286,N_702,N_977);
nand U1287 (N_1287,N_617,N_699);
nand U1288 (N_1288,N_972,N_938);
nor U1289 (N_1289,N_946,N_617);
nor U1290 (N_1290,N_664,N_735);
and U1291 (N_1291,N_643,N_695);
and U1292 (N_1292,N_553,N_750);
and U1293 (N_1293,N_763,N_915);
nor U1294 (N_1294,N_536,N_765);
and U1295 (N_1295,N_748,N_909);
or U1296 (N_1296,N_899,N_532);
and U1297 (N_1297,N_575,N_535);
and U1298 (N_1298,N_515,N_821);
nand U1299 (N_1299,N_690,N_568);
or U1300 (N_1300,N_825,N_958);
nand U1301 (N_1301,N_731,N_721);
nor U1302 (N_1302,N_939,N_755);
nor U1303 (N_1303,N_500,N_618);
nor U1304 (N_1304,N_976,N_735);
nand U1305 (N_1305,N_635,N_923);
nand U1306 (N_1306,N_880,N_986);
nand U1307 (N_1307,N_750,N_673);
nor U1308 (N_1308,N_859,N_511);
nor U1309 (N_1309,N_790,N_967);
or U1310 (N_1310,N_547,N_623);
nor U1311 (N_1311,N_941,N_947);
or U1312 (N_1312,N_717,N_969);
and U1313 (N_1313,N_808,N_553);
and U1314 (N_1314,N_548,N_800);
or U1315 (N_1315,N_701,N_903);
or U1316 (N_1316,N_728,N_963);
nor U1317 (N_1317,N_545,N_953);
and U1318 (N_1318,N_789,N_614);
xor U1319 (N_1319,N_975,N_853);
nand U1320 (N_1320,N_612,N_900);
and U1321 (N_1321,N_923,N_926);
nand U1322 (N_1322,N_604,N_736);
and U1323 (N_1323,N_704,N_836);
nor U1324 (N_1324,N_629,N_779);
or U1325 (N_1325,N_701,N_503);
nand U1326 (N_1326,N_998,N_789);
nor U1327 (N_1327,N_930,N_927);
and U1328 (N_1328,N_883,N_691);
or U1329 (N_1329,N_574,N_808);
nor U1330 (N_1330,N_630,N_791);
nand U1331 (N_1331,N_912,N_853);
and U1332 (N_1332,N_996,N_652);
nor U1333 (N_1333,N_876,N_886);
and U1334 (N_1334,N_924,N_663);
nand U1335 (N_1335,N_772,N_628);
nand U1336 (N_1336,N_863,N_588);
or U1337 (N_1337,N_829,N_934);
and U1338 (N_1338,N_923,N_549);
nor U1339 (N_1339,N_810,N_537);
and U1340 (N_1340,N_825,N_853);
or U1341 (N_1341,N_808,N_655);
or U1342 (N_1342,N_752,N_537);
and U1343 (N_1343,N_929,N_609);
and U1344 (N_1344,N_692,N_639);
or U1345 (N_1345,N_810,N_559);
and U1346 (N_1346,N_569,N_995);
or U1347 (N_1347,N_742,N_512);
or U1348 (N_1348,N_926,N_933);
nand U1349 (N_1349,N_554,N_619);
nor U1350 (N_1350,N_889,N_877);
nand U1351 (N_1351,N_796,N_955);
and U1352 (N_1352,N_583,N_657);
or U1353 (N_1353,N_853,N_935);
and U1354 (N_1354,N_797,N_739);
or U1355 (N_1355,N_722,N_857);
nand U1356 (N_1356,N_870,N_521);
nor U1357 (N_1357,N_889,N_942);
and U1358 (N_1358,N_834,N_552);
nand U1359 (N_1359,N_782,N_845);
nor U1360 (N_1360,N_965,N_906);
or U1361 (N_1361,N_632,N_625);
nor U1362 (N_1362,N_802,N_888);
nand U1363 (N_1363,N_871,N_888);
and U1364 (N_1364,N_800,N_523);
nor U1365 (N_1365,N_758,N_619);
nand U1366 (N_1366,N_670,N_687);
nor U1367 (N_1367,N_644,N_674);
and U1368 (N_1368,N_672,N_943);
or U1369 (N_1369,N_882,N_809);
nand U1370 (N_1370,N_537,N_908);
and U1371 (N_1371,N_999,N_873);
nand U1372 (N_1372,N_584,N_620);
or U1373 (N_1373,N_945,N_656);
nand U1374 (N_1374,N_616,N_685);
nand U1375 (N_1375,N_687,N_698);
nand U1376 (N_1376,N_664,N_622);
nand U1377 (N_1377,N_524,N_584);
nand U1378 (N_1378,N_716,N_763);
nor U1379 (N_1379,N_992,N_602);
xor U1380 (N_1380,N_549,N_989);
nand U1381 (N_1381,N_831,N_764);
or U1382 (N_1382,N_835,N_676);
or U1383 (N_1383,N_833,N_884);
xnor U1384 (N_1384,N_768,N_610);
or U1385 (N_1385,N_931,N_534);
nor U1386 (N_1386,N_768,N_613);
nor U1387 (N_1387,N_569,N_883);
or U1388 (N_1388,N_746,N_538);
or U1389 (N_1389,N_612,N_507);
xnor U1390 (N_1390,N_688,N_671);
and U1391 (N_1391,N_961,N_836);
nor U1392 (N_1392,N_673,N_584);
nand U1393 (N_1393,N_592,N_674);
nor U1394 (N_1394,N_803,N_598);
nand U1395 (N_1395,N_516,N_867);
nor U1396 (N_1396,N_904,N_650);
nand U1397 (N_1397,N_645,N_974);
or U1398 (N_1398,N_779,N_682);
nand U1399 (N_1399,N_540,N_569);
or U1400 (N_1400,N_585,N_813);
nor U1401 (N_1401,N_567,N_789);
and U1402 (N_1402,N_511,N_967);
and U1403 (N_1403,N_739,N_652);
nand U1404 (N_1404,N_508,N_536);
nor U1405 (N_1405,N_903,N_972);
and U1406 (N_1406,N_784,N_833);
nor U1407 (N_1407,N_871,N_528);
or U1408 (N_1408,N_960,N_910);
nand U1409 (N_1409,N_885,N_649);
or U1410 (N_1410,N_713,N_776);
or U1411 (N_1411,N_581,N_805);
or U1412 (N_1412,N_840,N_960);
nand U1413 (N_1413,N_780,N_571);
xnor U1414 (N_1414,N_508,N_659);
or U1415 (N_1415,N_547,N_682);
nand U1416 (N_1416,N_751,N_736);
nor U1417 (N_1417,N_511,N_587);
or U1418 (N_1418,N_842,N_900);
nor U1419 (N_1419,N_581,N_735);
nor U1420 (N_1420,N_580,N_880);
or U1421 (N_1421,N_762,N_618);
and U1422 (N_1422,N_832,N_525);
nand U1423 (N_1423,N_590,N_879);
nor U1424 (N_1424,N_647,N_729);
nand U1425 (N_1425,N_989,N_987);
or U1426 (N_1426,N_854,N_573);
or U1427 (N_1427,N_948,N_758);
and U1428 (N_1428,N_641,N_600);
nor U1429 (N_1429,N_687,N_566);
and U1430 (N_1430,N_546,N_768);
and U1431 (N_1431,N_609,N_557);
nor U1432 (N_1432,N_935,N_923);
or U1433 (N_1433,N_580,N_514);
nand U1434 (N_1434,N_556,N_814);
nand U1435 (N_1435,N_864,N_506);
nor U1436 (N_1436,N_585,N_695);
xor U1437 (N_1437,N_818,N_799);
nand U1438 (N_1438,N_925,N_960);
nand U1439 (N_1439,N_991,N_727);
or U1440 (N_1440,N_610,N_785);
nand U1441 (N_1441,N_520,N_637);
nor U1442 (N_1442,N_554,N_909);
nand U1443 (N_1443,N_825,N_664);
and U1444 (N_1444,N_523,N_594);
nand U1445 (N_1445,N_668,N_641);
and U1446 (N_1446,N_565,N_869);
and U1447 (N_1447,N_862,N_939);
nor U1448 (N_1448,N_557,N_709);
nand U1449 (N_1449,N_961,N_913);
and U1450 (N_1450,N_814,N_647);
and U1451 (N_1451,N_567,N_626);
or U1452 (N_1452,N_719,N_853);
and U1453 (N_1453,N_532,N_584);
and U1454 (N_1454,N_836,N_738);
or U1455 (N_1455,N_986,N_780);
or U1456 (N_1456,N_768,N_937);
or U1457 (N_1457,N_832,N_971);
nor U1458 (N_1458,N_639,N_812);
nor U1459 (N_1459,N_718,N_902);
and U1460 (N_1460,N_607,N_667);
and U1461 (N_1461,N_530,N_542);
or U1462 (N_1462,N_701,N_694);
nand U1463 (N_1463,N_859,N_770);
or U1464 (N_1464,N_841,N_658);
nor U1465 (N_1465,N_816,N_999);
or U1466 (N_1466,N_544,N_665);
and U1467 (N_1467,N_770,N_924);
nand U1468 (N_1468,N_646,N_622);
or U1469 (N_1469,N_682,N_515);
nand U1470 (N_1470,N_652,N_617);
nand U1471 (N_1471,N_627,N_948);
and U1472 (N_1472,N_698,N_826);
and U1473 (N_1473,N_878,N_875);
and U1474 (N_1474,N_935,N_550);
nand U1475 (N_1475,N_997,N_988);
nand U1476 (N_1476,N_966,N_911);
and U1477 (N_1477,N_567,N_950);
nor U1478 (N_1478,N_688,N_958);
or U1479 (N_1479,N_940,N_530);
nor U1480 (N_1480,N_968,N_697);
xnor U1481 (N_1481,N_672,N_647);
or U1482 (N_1482,N_589,N_558);
nand U1483 (N_1483,N_917,N_642);
nor U1484 (N_1484,N_780,N_704);
and U1485 (N_1485,N_543,N_990);
xnor U1486 (N_1486,N_733,N_870);
nand U1487 (N_1487,N_815,N_546);
nand U1488 (N_1488,N_622,N_539);
nor U1489 (N_1489,N_713,N_523);
nor U1490 (N_1490,N_658,N_961);
nor U1491 (N_1491,N_530,N_680);
nor U1492 (N_1492,N_517,N_925);
nor U1493 (N_1493,N_601,N_858);
nand U1494 (N_1494,N_605,N_952);
nor U1495 (N_1495,N_509,N_785);
nand U1496 (N_1496,N_921,N_500);
or U1497 (N_1497,N_703,N_699);
nand U1498 (N_1498,N_624,N_560);
nor U1499 (N_1499,N_658,N_822);
and U1500 (N_1500,N_1253,N_1362);
and U1501 (N_1501,N_1066,N_1459);
nand U1502 (N_1502,N_1435,N_1315);
and U1503 (N_1503,N_1180,N_1059);
and U1504 (N_1504,N_1004,N_1283);
nand U1505 (N_1505,N_1421,N_1072);
or U1506 (N_1506,N_1038,N_1102);
and U1507 (N_1507,N_1431,N_1344);
or U1508 (N_1508,N_1101,N_1034);
nand U1509 (N_1509,N_1092,N_1081);
nand U1510 (N_1510,N_1190,N_1017);
or U1511 (N_1511,N_1437,N_1363);
or U1512 (N_1512,N_1274,N_1140);
or U1513 (N_1513,N_1396,N_1058);
or U1514 (N_1514,N_1098,N_1493);
nor U1515 (N_1515,N_1440,N_1353);
nor U1516 (N_1516,N_1231,N_1133);
nand U1517 (N_1517,N_1282,N_1047);
or U1518 (N_1518,N_1216,N_1355);
nand U1519 (N_1519,N_1107,N_1357);
nand U1520 (N_1520,N_1148,N_1365);
nor U1521 (N_1521,N_1436,N_1086);
nand U1522 (N_1522,N_1249,N_1083);
and U1523 (N_1523,N_1377,N_1015);
nand U1524 (N_1524,N_1022,N_1161);
or U1525 (N_1525,N_1224,N_1318);
nand U1526 (N_1526,N_1191,N_1070);
or U1527 (N_1527,N_1491,N_1167);
and U1528 (N_1528,N_1176,N_1263);
nor U1529 (N_1529,N_1169,N_1288);
and U1530 (N_1530,N_1356,N_1040);
nand U1531 (N_1531,N_1379,N_1195);
nor U1532 (N_1532,N_1064,N_1241);
nand U1533 (N_1533,N_1234,N_1123);
and U1534 (N_1534,N_1255,N_1220);
and U1535 (N_1535,N_1346,N_1339);
nor U1536 (N_1536,N_1001,N_1205);
xor U1537 (N_1537,N_1330,N_1380);
nand U1538 (N_1538,N_1397,N_1406);
and U1539 (N_1539,N_1145,N_1067);
or U1540 (N_1540,N_1323,N_1475);
nand U1541 (N_1541,N_1187,N_1046);
nand U1542 (N_1542,N_1413,N_1077);
nor U1543 (N_1543,N_1172,N_1321);
nor U1544 (N_1544,N_1108,N_1432);
or U1545 (N_1545,N_1351,N_1299);
nor U1546 (N_1546,N_1076,N_1014);
or U1547 (N_1547,N_1261,N_1225);
and U1548 (N_1548,N_1018,N_1376);
or U1549 (N_1549,N_1302,N_1236);
and U1550 (N_1550,N_1358,N_1273);
and U1551 (N_1551,N_1174,N_1245);
nand U1552 (N_1552,N_1115,N_1359);
nand U1553 (N_1553,N_1338,N_1259);
nand U1554 (N_1554,N_1229,N_1240);
and U1555 (N_1555,N_1414,N_1345);
nor U1556 (N_1556,N_1449,N_1266);
nor U1557 (N_1557,N_1441,N_1457);
and U1558 (N_1558,N_1294,N_1036);
or U1559 (N_1559,N_1419,N_1178);
nor U1560 (N_1560,N_1157,N_1489);
nor U1561 (N_1561,N_1279,N_1160);
xor U1562 (N_1562,N_1235,N_1027);
and U1563 (N_1563,N_1037,N_1394);
nor U1564 (N_1564,N_1324,N_1139);
nor U1565 (N_1565,N_1199,N_1204);
and U1566 (N_1566,N_1478,N_1292);
and U1567 (N_1567,N_1389,N_1211);
and U1568 (N_1568,N_1320,N_1269);
and U1569 (N_1569,N_1202,N_1331);
or U1570 (N_1570,N_1285,N_1177);
nand U1571 (N_1571,N_1367,N_1369);
nor U1572 (N_1572,N_1024,N_1061);
nor U1573 (N_1573,N_1210,N_1011);
and U1574 (N_1574,N_1163,N_1354);
nor U1575 (N_1575,N_1254,N_1463);
or U1576 (N_1576,N_1122,N_1470);
nor U1577 (N_1577,N_1049,N_1073);
or U1578 (N_1578,N_1458,N_1455);
or U1579 (N_1579,N_1296,N_1252);
or U1580 (N_1580,N_1492,N_1343);
nand U1581 (N_1581,N_1050,N_1010);
or U1582 (N_1582,N_1117,N_1062);
nand U1583 (N_1583,N_1151,N_1247);
and U1584 (N_1584,N_1298,N_1183);
and U1585 (N_1585,N_1422,N_1428);
nand U1586 (N_1586,N_1398,N_1103);
and U1587 (N_1587,N_1232,N_1251);
and U1588 (N_1588,N_1329,N_1392);
nand U1589 (N_1589,N_1287,N_1087);
xor U1590 (N_1590,N_1222,N_1270);
or U1591 (N_1591,N_1276,N_1239);
nand U1592 (N_1592,N_1156,N_1485);
nand U1593 (N_1593,N_1385,N_1041);
nand U1594 (N_1594,N_1184,N_1390);
or U1595 (N_1595,N_1196,N_1469);
nor U1596 (N_1596,N_1483,N_1007);
or U1597 (N_1597,N_1486,N_1141);
and U1598 (N_1598,N_1289,N_1075);
and U1599 (N_1599,N_1314,N_1134);
or U1600 (N_1600,N_1207,N_1124);
nand U1601 (N_1601,N_1429,N_1096);
nor U1602 (N_1602,N_1368,N_1243);
and U1603 (N_1603,N_1130,N_1260);
or U1604 (N_1604,N_1498,N_1456);
nor U1605 (N_1605,N_1472,N_1409);
and U1606 (N_1606,N_1424,N_1056);
and U1607 (N_1607,N_1030,N_1480);
or U1608 (N_1608,N_1106,N_1352);
and U1609 (N_1609,N_1142,N_1048);
or U1610 (N_1610,N_1381,N_1332);
nor U1611 (N_1611,N_1194,N_1111);
nand U1612 (N_1612,N_1479,N_1057);
nand U1613 (N_1613,N_1452,N_1152);
nand U1614 (N_1614,N_1149,N_1182);
and U1615 (N_1615,N_1290,N_1135);
nand U1616 (N_1616,N_1496,N_1063);
and U1617 (N_1617,N_1219,N_1035);
and U1618 (N_1618,N_1109,N_1074);
or U1619 (N_1619,N_1246,N_1039);
nor U1620 (N_1620,N_1188,N_1293);
nand U1621 (N_1621,N_1166,N_1402);
nor U1622 (N_1622,N_1340,N_1291);
and U1623 (N_1623,N_1104,N_1116);
or U1624 (N_1624,N_1304,N_1080);
nor U1625 (N_1625,N_1425,N_1461);
nand U1626 (N_1626,N_1214,N_1230);
and U1627 (N_1627,N_1335,N_1131);
and U1628 (N_1628,N_1325,N_1129);
or U1629 (N_1629,N_1091,N_1113);
nand U1630 (N_1630,N_1069,N_1181);
nor U1631 (N_1631,N_1043,N_1029);
nand U1632 (N_1632,N_1295,N_1447);
nor U1633 (N_1633,N_1258,N_1016);
nand U1634 (N_1634,N_1060,N_1423);
nand U1635 (N_1635,N_1065,N_1426);
or U1636 (N_1636,N_1114,N_1418);
nand U1637 (N_1637,N_1495,N_1451);
nor U1638 (N_1638,N_1159,N_1158);
nand U1639 (N_1639,N_1078,N_1100);
nor U1640 (N_1640,N_1238,N_1226);
nor U1641 (N_1641,N_1006,N_1407);
nand U1642 (N_1642,N_1089,N_1453);
nand U1643 (N_1643,N_1446,N_1484);
nor U1644 (N_1644,N_1053,N_1378);
or U1645 (N_1645,N_1023,N_1126);
nand U1646 (N_1646,N_1179,N_1348);
nor U1647 (N_1647,N_1420,N_1143);
nor U1648 (N_1648,N_1373,N_1054);
and U1649 (N_1649,N_1085,N_1490);
and U1650 (N_1650,N_1044,N_1110);
and U1651 (N_1651,N_1002,N_1383);
nor U1652 (N_1652,N_1164,N_1013);
and U1653 (N_1653,N_1311,N_1248);
nor U1654 (N_1654,N_1444,N_1403);
and U1655 (N_1655,N_1328,N_1300);
nand U1656 (N_1656,N_1105,N_1228);
nand U1657 (N_1657,N_1212,N_1319);
xnor U1658 (N_1658,N_1003,N_1162);
and U1659 (N_1659,N_1218,N_1209);
nand U1660 (N_1660,N_1312,N_1488);
or U1661 (N_1661,N_1374,N_1473);
or U1662 (N_1662,N_1284,N_1317);
or U1663 (N_1663,N_1068,N_1099);
or U1664 (N_1664,N_1280,N_1112);
nand U1665 (N_1665,N_1297,N_1384);
and U1666 (N_1666,N_1136,N_1494);
and U1667 (N_1667,N_1333,N_1272);
nor U1668 (N_1668,N_1071,N_1201);
nor U1669 (N_1669,N_1118,N_1482);
nor U1670 (N_1670,N_1026,N_1005);
and U1671 (N_1671,N_1301,N_1336);
nand U1672 (N_1672,N_1095,N_1477);
nand U1673 (N_1673,N_1009,N_1079);
nor U1674 (N_1674,N_1430,N_1233);
nand U1675 (N_1675,N_1203,N_1371);
xor U1676 (N_1676,N_1208,N_1360);
nand U1677 (N_1677,N_1032,N_1286);
nand U1678 (N_1678,N_1146,N_1445);
or U1679 (N_1679,N_1128,N_1084);
nand U1680 (N_1680,N_1250,N_1237);
nor U1681 (N_1681,N_1185,N_1415);
nand U1682 (N_1682,N_1197,N_1144);
nand U1683 (N_1683,N_1408,N_1055);
and U1684 (N_1684,N_1132,N_1393);
xnor U1685 (N_1685,N_1326,N_1448);
nand U1686 (N_1686,N_1417,N_1227);
nand U1687 (N_1687,N_1313,N_1434);
nor U1688 (N_1688,N_1316,N_1382);
nand U1689 (N_1689,N_1364,N_1334);
and U1690 (N_1690,N_1342,N_1307);
nor U1691 (N_1691,N_1277,N_1168);
nand U1692 (N_1692,N_1337,N_1278);
or U1693 (N_1693,N_1309,N_1082);
and U1694 (N_1694,N_1265,N_1256);
or U1695 (N_1695,N_1045,N_1465);
and U1696 (N_1696,N_1460,N_1186);
nand U1697 (N_1697,N_1012,N_1471);
nand U1698 (N_1698,N_1405,N_1244);
and U1699 (N_1699,N_1042,N_1200);
nand U1700 (N_1700,N_1341,N_1173);
nand U1701 (N_1701,N_1264,N_1093);
nor U1702 (N_1702,N_1147,N_1150);
nor U1703 (N_1703,N_1021,N_1361);
or U1704 (N_1704,N_1387,N_1349);
nor U1705 (N_1705,N_1175,N_1388);
or U1706 (N_1706,N_1443,N_1499);
nor U1707 (N_1707,N_1275,N_1481);
and U1708 (N_1708,N_1033,N_1242);
nor U1709 (N_1709,N_1120,N_1155);
nor U1710 (N_1710,N_1223,N_1327);
or U1711 (N_1711,N_1416,N_1051);
or U1712 (N_1712,N_1020,N_1262);
or U1713 (N_1713,N_1271,N_1281);
or U1714 (N_1714,N_1464,N_1137);
nand U1715 (N_1715,N_1121,N_1410);
and U1716 (N_1716,N_1192,N_1439);
and U1717 (N_1717,N_1399,N_1391);
and U1718 (N_1718,N_1090,N_1450);
and U1719 (N_1719,N_1025,N_1400);
nand U1720 (N_1720,N_1303,N_1462);
and U1721 (N_1721,N_1088,N_1171);
nand U1722 (N_1722,N_1442,N_1487);
or U1723 (N_1723,N_1305,N_1000);
nor U1724 (N_1724,N_1372,N_1154);
and U1725 (N_1725,N_1433,N_1031);
nor U1726 (N_1726,N_1386,N_1094);
and U1727 (N_1727,N_1468,N_1138);
nor U1728 (N_1728,N_1125,N_1427);
nand U1729 (N_1729,N_1350,N_1217);
nand U1730 (N_1730,N_1119,N_1153);
or U1731 (N_1731,N_1474,N_1497);
nand U1732 (N_1732,N_1221,N_1308);
or U1733 (N_1733,N_1476,N_1193);
xor U1734 (N_1734,N_1310,N_1467);
nor U1735 (N_1735,N_1127,N_1411);
or U1736 (N_1736,N_1206,N_1306);
nand U1737 (N_1737,N_1213,N_1401);
and U1738 (N_1738,N_1466,N_1008);
nand U1739 (N_1739,N_1412,N_1028);
and U1740 (N_1740,N_1165,N_1097);
and U1741 (N_1741,N_1215,N_1268);
or U1742 (N_1742,N_1375,N_1395);
nor U1743 (N_1743,N_1170,N_1438);
nor U1744 (N_1744,N_1347,N_1366);
and U1745 (N_1745,N_1189,N_1267);
nand U1746 (N_1746,N_1370,N_1322);
or U1747 (N_1747,N_1257,N_1404);
nor U1748 (N_1748,N_1019,N_1198);
nand U1749 (N_1749,N_1052,N_1454);
xnor U1750 (N_1750,N_1236,N_1140);
or U1751 (N_1751,N_1078,N_1482);
or U1752 (N_1752,N_1014,N_1194);
nor U1753 (N_1753,N_1453,N_1108);
nand U1754 (N_1754,N_1065,N_1132);
xor U1755 (N_1755,N_1139,N_1060);
and U1756 (N_1756,N_1455,N_1245);
and U1757 (N_1757,N_1177,N_1083);
nor U1758 (N_1758,N_1291,N_1350);
nand U1759 (N_1759,N_1243,N_1092);
and U1760 (N_1760,N_1191,N_1083);
and U1761 (N_1761,N_1348,N_1082);
nand U1762 (N_1762,N_1322,N_1299);
or U1763 (N_1763,N_1363,N_1340);
nor U1764 (N_1764,N_1426,N_1240);
or U1765 (N_1765,N_1400,N_1375);
or U1766 (N_1766,N_1432,N_1133);
nor U1767 (N_1767,N_1029,N_1484);
and U1768 (N_1768,N_1171,N_1143);
and U1769 (N_1769,N_1188,N_1447);
nand U1770 (N_1770,N_1071,N_1206);
nor U1771 (N_1771,N_1266,N_1048);
and U1772 (N_1772,N_1331,N_1098);
nor U1773 (N_1773,N_1045,N_1097);
nand U1774 (N_1774,N_1454,N_1217);
nor U1775 (N_1775,N_1370,N_1446);
nand U1776 (N_1776,N_1179,N_1175);
or U1777 (N_1777,N_1337,N_1064);
or U1778 (N_1778,N_1280,N_1148);
nand U1779 (N_1779,N_1060,N_1354);
or U1780 (N_1780,N_1410,N_1108);
nor U1781 (N_1781,N_1272,N_1031);
nand U1782 (N_1782,N_1403,N_1182);
or U1783 (N_1783,N_1493,N_1312);
nor U1784 (N_1784,N_1249,N_1391);
nand U1785 (N_1785,N_1178,N_1438);
nand U1786 (N_1786,N_1307,N_1242);
and U1787 (N_1787,N_1021,N_1145);
and U1788 (N_1788,N_1045,N_1290);
or U1789 (N_1789,N_1349,N_1246);
nor U1790 (N_1790,N_1124,N_1175);
or U1791 (N_1791,N_1267,N_1399);
nor U1792 (N_1792,N_1064,N_1324);
and U1793 (N_1793,N_1098,N_1473);
and U1794 (N_1794,N_1285,N_1245);
and U1795 (N_1795,N_1303,N_1367);
or U1796 (N_1796,N_1098,N_1348);
nand U1797 (N_1797,N_1034,N_1468);
or U1798 (N_1798,N_1416,N_1453);
nand U1799 (N_1799,N_1031,N_1367);
nor U1800 (N_1800,N_1361,N_1303);
and U1801 (N_1801,N_1219,N_1335);
or U1802 (N_1802,N_1207,N_1484);
nor U1803 (N_1803,N_1227,N_1480);
and U1804 (N_1804,N_1188,N_1491);
or U1805 (N_1805,N_1384,N_1457);
nor U1806 (N_1806,N_1167,N_1237);
nand U1807 (N_1807,N_1433,N_1003);
nor U1808 (N_1808,N_1014,N_1324);
nor U1809 (N_1809,N_1458,N_1262);
xnor U1810 (N_1810,N_1366,N_1303);
nor U1811 (N_1811,N_1447,N_1261);
or U1812 (N_1812,N_1380,N_1334);
and U1813 (N_1813,N_1084,N_1039);
and U1814 (N_1814,N_1401,N_1209);
or U1815 (N_1815,N_1340,N_1370);
and U1816 (N_1816,N_1486,N_1142);
and U1817 (N_1817,N_1158,N_1112);
and U1818 (N_1818,N_1358,N_1313);
and U1819 (N_1819,N_1320,N_1240);
and U1820 (N_1820,N_1387,N_1143);
and U1821 (N_1821,N_1438,N_1045);
or U1822 (N_1822,N_1464,N_1297);
and U1823 (N_1823,N_1021,N_1207);
nand U1824 (N_1824,N_1389,N_1314);
nand U1825 (N_1825,N_1118,N_1396);
nor U1826 (N_1826,N_1153,N_1453);
or U1827 (N_1827,N_1453,N_1244);
and U1828 (N_1828,N_1112,N_1486);
or U1829 (N_1829,N_1125,N_1017);
nand U1830 (N_1830,N_1105,N_1185);
and U1831 (N_1831,N_1085,N_1173);
or U1832 (N_1832,N_1219,N_1044);
nor U1833 (N_1833,N_1392,N_1466);
nor U1834 (N_1834,N_1490,N_1113);
or U1835 (N_1835,N_1155,N_1092);
nor U1836 (N_1836,N_1257,N_1168);
nor U1837 (N_1837,N_1392,N_1164);
nand U1838 (N_1838,N_1116,N_1192);
nor U1839 (N_1839,N_1221,N_1481);
nor U1840 (N_1840,N_1202,N_1006);
and U1841 (N_1841,N_1158,N_1102);
and U1842 (N_1842,N_1410,N_1197);
nand U1843 (N_1843,N_1271,N_1361);
nor U1844 (N_1844,N_1441,N_1402);
and U1845 (N_1845,N_1296,N_1131);
nand U1846 (N_1846,N_1291,N_1439);
or U1847 (N_1847,N_1442,N_1437);
and U1848 (N_1848,N_1083,N_1085);
nand U1849 (N_1849,N_1017,N_1066);
and U1850 (N_1850,N_1045,N_1159);
nand U1851 (N_1851,N_1043,N_1349);
and U1852 (N_1852,N_1359,N_1464);
nand U1853 (N_1853,N_1296,N_1140);
or U1854 (N_1854,N_1110,N_1076);
and U1855 (N_1855,N_1217,N_1415);
and U1856 (N_1856,N_1178,N_1405);
or U1857 (N_1857,N_1076,N_1248);
and U1858 (N_1858,N_1459,N_1262);
and U1859 (N_1859,N_1276,N_1229);
xnor U1860 (N_1860,N_1373,N_1343);
and U1861 (N_1861,N_1266,N_1401);
nor U1862 (N_1862,N_1146,N_1336);
and U1863 (N_1863,N_1374,N_1106);
or U1864 (N_1864,N_1078,N_1028);
nor U1865 (N_1865,N_1368,N_1229);
nor U1866 (N_1866,N_1308,N_1471);
and U1867 (N_1867,N_1012,N_1195);
or U1868 (N_1868,N_1094,N_1423);
or U1869 (N_1869,N_1279,N_1353);
and U1870 (N_1870,N_1235,N_1487);
nand U1871 (N_1871,N_1277,N_1142);
nand U1872 (N_1872,N_1347,N_1094);
nor U1873 (N_1873,N_1321,N_1144);
and U1874 (N_1874,N_1062,N_1359);
and U1875 (N_1875,N_1248,N_1056);
and U1876 (N_1876,N_1348,N_1171);
nor U1877 (N_1877,N_1302,N_1498);
and U1878 (N_1878,N_1073,N_1029);
nand U1879 (N_1879,N_1054,N_1159);
xnor U1880 (N_1880,N_1392,N_1341);
and U1881 (N_1881,N_1231,N_1125);
nand U1882 (N_1882,N_1404,N_1033);
and U1883 (N_1883,N_1449,N_1373);
nor U1884 (N_1884,N_1247,N_1060);
nor U1885 (N_1885,N_1392,N_1126);
and U1886 (N_1886,N_1472,N_1156);
nand U1887 (N_1887,N_1071,N_1093);
or U1888 (N_1888,N_1409,N_1369);
or U1889 (N_1889,N_1225,N_1327);
xnor U1890 (N_1890,N_1476,N_1460);
nor U1891 (N_1891,N_1248,N_1493);
or U1892 (N_1892,N_1396,N_1126);
nor U1893 (N_1893,N_1157,N_1356);
or U1894 (N_1894,N_1242,N_1425);
nor U1895 (N_1895,N_1484,N_1472);
nand U1896 (N_1896,N_1126,N_1465);
or U1897 (N_1897,N_1211,N_1420);
and U1898 (N_1898,N_1406,N_1447);
nor U1899 (N_1899,N_1327,N_1202);
and U1900 (N_1900,N_1053,N_1027);
nor U1901 (N_1901,N_1254,N_1477);
or U1902 (N_1902,N_1290,N_1214);
and U1903 (N_1903,N_1309,N_1126);
and U1904 (N_1904,N_1444,N_1339);
nand U1905 (N_1905,N_1346,N_1125);
nor U1906 (N_1906,N_1154,N_1017);
nand U1907 (N_1907,N_1197,N_1183);
and U1908 (N_1908,N_1360,N_1354);
and U1909 (N_1909,N_1401,N_1102);
or U1910 (N_1910,N_1418,N_1066);
and U1911 (N_1911,N_1222,N_1464);
nand U1912 (N_1912,N_1419,N_1043);
or U1913 (N_1913,N_1107,N_1414);
or U1914 (N_1914,N_1306,N_1110);
nand U1915 (N_1915,N_1189,N_1415);
nand U1916 (N_1916,N_1420,N_1170);
nor U1917 (N_1917,N_1407,N_1356);
or U1918 (N_1918,N_1205,N_1455);
nand U1919 (N_1919,N_1339,N_1116);
and U1920 (N_1920,N_1194,N_1211);
or U1921 (N_1921,N_1063,N_1284);
nor U1922 (N_1922,N_1198,N_1392);
and U1923 (N_1923,N_1429,N_1409);
nand U1924 (N_1924,N_1477,N_1201);
nor U1925 (N_1925,N_1376,N_1332);
or U1926 (N_1926,N_1401,N_1409);
nand U1927 (N_1927,N_1322,N_1241);
or U1928 (N_1928,N_1300,N_1033);
nand U1929 (N_1929,N_1092,N_1427);
or U1930 (N_1930,N_1479,N_1491);
or U1931 (N_1931,N_1371,N_1001);
nor U1932 (N_1932,N_1140,N_1174);
nor U1933 (N_1933,N_1352,N_1062);
and U1934 (N_1934,N_1011,N_1027);
and U1935 (N_1935,N_1282,N_1248);
or U1936 (N_1936,N_1473,N_1198);
nand U1937 (N_1937,N_1345,N_1074);
or U1938 (N_1938,N_1396,N_1013);
or U1939 (N_1939,N_1392,N_1124);
or U1940 (N_1940,N_1428,N_1450);
nor U1941 (N_1941,N_1330,N_1414);
nand U1942 (N_1942,N_1156,N_1153);
and U1943 (N_1943,N_1468,N_1304);
and U1944 (N_1944,N_1102,N_1383);
nand U1945 (N_1945,N_1486,N_1342);
and U1946 (N_1946,N_1395,N_1425);
or U1947 (N_1947,N_1387,N_1101);
nand U1948 (N_1948,N_1488,N_1094);
and U1949 (N_1949,N_1214,N_1049);
and U1950 (N_1950,N_1448,N_1064);
or U1951 (N_1951,N_1112,N_1318);
nand U1952 (N_1952,N_1277,N_1324);
nor U1953 (N_1953,N_1341,N_1037);
or U1954 (N_1954,N_1040,N_1180);
or U1955 (N_1955,N_1152,N_1048);
and U1956 (N_1956,N_1255,N_1487);
nand U1957 (N_1957,N_1340,N_1136);
or U1958 (N_1958,N_1018,N_1167);
nor U1959 (N_1959,N_1262,N_1193);
or U1960 (N_1960,N_1433,N_1203);
nand U1961 (N_1961,N_1111,N_1281);
and U1962 (N_1962,N_1494,N_1304);
nand U1963 (N_1963,N_1040,N_1086);
nand U1964 (N_1964,N_1420,N_1044);
nor U1965 (N_1965,N_1400,N_1179);
nand U1966 (N_1966,N_1361,N_1042);
and U1967 (N_1967,N_1174,N_1112);
nand U1968 (N_1968,N_1458,N_1034);
and U1969 (N_1969,N_1422,N_1009);
nor U1970 (N_1970,N_1071,N_1176);
and U1971 (N_1971,N_1331,N_1000);
or U1972 (N_1972,N_1340,N_1267);
or U1973 (N_1973,N_1329,N_1196);
and U1974 (N_1974,N_1379,N_1322);
nor U1975 (N_1975,N_1347,N_1102);
nor U1976 (N_1976,N_1286,N_1473);
nor U1977 (N_1977,N_1061,N_1135);
or U1978 (N_1978,N_1163,N_1425);
nand U1979 (N_1979,N_1120,N_1241);
or U1980 (N_1980,N_1334,N_1001);
and U1981 (N_1981,N_1263,N_1451);
nand U1982 (N_1982,N_1309,N_1294);
nor U1983 (N_1983,N_1451,N_1257);
or U1984 (N_1984,N_1236,N_1155);
or U1985 (N_1985,N_1239,N_1372);
nor U1986 (N_1986,N_1397,N_1151);
xor U1987 (N_1987,N_1214,N_1336);
and U1988 (N_1988,N_1382,N_1104);
or U1989 (N_1989,N_1262,N_1145);
nor U1990 (N_1990,N_1025,N_1116);
or U1991 (N_1991,N_1435,N_1078);
or U1992 (N_1992,N_1417,N_1202);
nand U1993 (N_1993,N_1479,N_1030);
nor U1994 (N_1994,N_1238,N_1119);
or U1995 (N_1995,N_1485,N_1495);
and U1996 (N_1996,N_1290,N_1090);
nand U1997 (N_1997,N_1398,N_1138);
or U1998 (N_1998,N_1121,N_1270);
and U1999 (N_1999,N_1411,N_1177);
nor U2000 (N_2000,N_1512,N_1839);
or U2001 (N_2001,N_1594,N_1816);
nand U2002 (N_2002,N_1564,N_1722);
xor U2003 (N_2003,N_1639,N_1720);
nand U2004 (N_2004,N_1567,N_1606);
and U2005 (N_2005,N_1505,N_1935);
nor U2006 (N_2006,N_1902,N_1581);
or U2007 (N_2007,N_1922,N_1968);
and U2008 (N_2008,N_1970,N_1727);
nor U2009 (N_2009,N_1507,N_1643);
and U2010 (N_2010,N_1633,N_1588);
and U2011 (N_2011,N_1669,N_1928);
or U2012 (N_2012,N_1673,N_1754);
nand U2013 (N_2013,N_1743,N_1768);
xor U2014 (N_2014,N_1526,N_1607);
nand U2015 (N_2015,N_1939,N_1724);
nand U2016 (N_2016,N_1772,N_1738);
nand U2017 (N_2017,N_1561,N_1974);
nor U2018 (N_2018,N_1586,N_1732);
nor U2019 (N_2019,N_1851,N_1551);
or U2020 (N_2020,N_1725,N_1981);
or U2021 (N_2021,N_1773,N_1859);
or U2022 (N_2022,N_1558,N_1863);
and U2023 (N_2023,N_1809,N_1999);
or U2024 (N_2024,N_1637,N_1745);
nor U2025 (N_2025,N_1797,N_1591);
nor U2026 (N_2026,N_1644,N_1589);
nor U2027 (N_2027,N_1697,N_1681);
nor U2028 (N_2028,N_1667,N_1847);
and U2029 (N_2029,N_1876,N_1543);
or U2030 (N_2030,N_1934,N_1880);
nor U2031 (N_2031,N_1580,N_1717);
nor U2032 (N_2032,N_1957,N_1789);
and U2033 (N_2033,N_1593,N_1840);
and U2034 (N_2034,N_1822,N_1729);
nor U2035 (N_2035,N_1846,N_1504);
nand U2036 (N_2036,N_1595,N_1545);
nor U2037 (N_2037,N_1529,N_1574);
nand U2038 (N_2038,N_1665,N_1664);
and U2039 (N_2039,N_1565,N_1975);
nor U2040 (N_2040,N_1523,N_1536);
nor U2041 (N_2041,N_1503,N_1528);
nand U2042 (N_2042,N_1663,N_1763);
nand U2043 (N_2043,N_1857,N_1790);
or U2044 (N_2044,N_1983,N_1780);
nor U2045 (N_2045,N_1573,N_1955);
and U2046 (N_2046,N_1915,N_1609);
and U2047 (N_2047,N_1943,N_1844);
nor U2048 (N_2048,N_1855,N_1774);
nor U2049 (N_2049,N_1766,N_1510);
nor U2050 (N_2050,N_1937,N_1661);
or U2051 (N_2051,N_1638,N_1684);
and U2052 (N_2052,N_1971,N_1810);
and U2053 (N_2053,N_1592,N_1893);
nor U2054 (N_2054,N_1900,N_1597);
and U2055 (N_2055,N_1887,N_1831);
nand U2056 (N_2056,N_1694,N_1730);
nand U2057 (N_2057,N_1531,N_1520);
nand U2058 (N_2058,N_1631,N_1883);
or U2059 (N_2059,N_1628,N_1791);
or U2060 (N_2060,N_1742,N_1995);
nor U2061 (N_2061,N_1660,N_1699);
nor U2062 (N_2062,N_1898,N_1821);
or U2063 (N_2063,N_1712,N_1583);
xor U2064 (N_2064,N_1575,N_1805);
and U2065 (N_2065,N_1614,N_1794);
xor U2066 (N_2066,N_1817,N_1998);
nand U2067 (N_2067,N_1706,N_1576);
or U2068 (N_2068,N_1765,N_1687);
and U2069 (N_2069,N_1711,N_1962);
or U2070 (N_2070,N_1688,N_1918);
or U2071 (N_2071,N_1612,N_1658);
nand U2072 (N_2072,N_1927,N_1501);
nor U2073 (N_2073,N_1866,N_1517);
xnor U2074 (N_2074,N_1987,N_1522);
nand U2075 (N_2075,N_1864,N_1568);
nor U2076 (N_2076,N_1653,N_1779);
nand U2077 (N_2077,N_1823,N_1889);
and U2078 (N_2078,N_1993,N_1740);
and U2079 (N_2079,N_1914,N_1562);
and U2080 (N_2080,N_1716,N_1587);
and U2081 (N_2081,N_1502,N_1841);
nand U2082 (N_2082,N_1544,N_1509);
or U2083 (N_2083,N_1613,N_1682);
nor U2084 (N_2084,N_1845,N_1701);
nand U2085 (N_2085,N_1756,N_1877);
nor U2086 (N_2086,N_1784,N_1842);
and U2087 (N_2087,N_1795,N_1590);
or U2088 (N_2088,N_1611,N_1560);
or U2089 (N_2089,N_1683,N_1903);
or U2090 (N_2090,N_1830,N_1640);
or U2091 (N_2091,N_1750,N_1650);
and U2092 (N_2092,N_1635,N_1541);
and U2093 (N_2093,N_1532,N_1733);
and U2094 (N_2094,N_1698,N_1966);
or U2095 (N_2095,N_1819,N_1619);
nand U2096 (N_2096,N_1746,N_1759);
and U2097 (N_2097,N_1879,N_1555);
or U2098 (N_2098,N_1648,N_1938);
nand U2099 (N_2099,N_1559,N_1972);
nand U2100 (N_2100,N_1894,N_1837);
and U2101 (N_2101,N_1760,N_1812);
nand U2102 (N_2102,N_1806,N_1911);
nor U2103 (N_2103,N_1901,N_1912);
or U2104 (N_2104,N_1882,N_1600);
nand U2105 (N_2105,N_1994,N_1870);
or U2106 (N_2106,N_1788,N_1518);
and U2107 (N_2107,N_1632,N_1655);
and U2108 (N_2108,N_1961,N_1693);
or U2109 (N_2109,N_1832,N_1799);
and U2110 (N_2110,N_1885,N_1524);
or U2111 (N_2111,N_1838,N_1801);
or U2112 (N_2112,N_1519,N_1967);
and U2113 (N_2113,N_1622,N_1548);
nor U2114 (N_2114,N_1959,N_1888);
nand U2115 (N_2115,N_1954,N_1530);
and U2116 (N_2116,N_1807,N_1770);
nor U2117 (N_2117,N_1570,N_1629);
or U2118 (N_2118,N_1925,N_1867);
nand U2119 (N_2119,N_1811,N_1506);
and U2120 (N_2120,N_1679,N_1602);
nor U2121 (N_2121,N_1978,N_1781);
nand U2122 (N_2122,N_1702,N_1621);
nand U2123 (N_2123,N_1956,N_1843);
nor U2124 (N_2124,N_1721,N_1668);
nand U2125 (N_2125,N_1671,N_1976);
and U2126 (N_2126,N_1786,N_1991);
and U2127 (N_2127,N_1834,N_1654);
nor U2128 (N_2128,N_1726,N_1933);
and U2129 (N_2129,N_1945,N_1718);
and U2130 (N_2130,N_1824,N_1744);
nor U2131 (N_2131,N_1748,N_1657);
or U2132 (N_2132,N_1984,N_1990);
nand U2133 (N_2133,N_1949,N_1584);
xor U2134 (N_2134,N_1804,N_1873);
nand U2135 (N_2135,N_1703,N_1680);
nor U2136 (N_2136,N_1800,N_1926);
xor U2137 (N_2137,N_1989,N_1828);
nand U2138 (N_2138,N_1767,N_1758);
or U2139 (N_2139,N_1753,N_1931);
nor U2140 (N_2140,N_1540,N_1757);
and U2141 (N_2141,N_1696,N_1546);
nor U2142 (N_2142,N_1849,N_1869);
nor U2143 (N_2143,N_1850,N_1645);
xor U2144 (N_2144,N_1686,N_1808);
nand U2145 (N_2145,N_1554,N_1656);
and U2146 (N_2146,N_1930,N_1992);
nor U2147 (N_2147,N_1785,N_1936);
or U2148 (N_2148,N_1813,N_1618);
nand U2149 (N_2149,N_1778,N_1920);
nor U2150 (N_2150,N_1921,N_1865);
nor U2151 (N_2151,N_1685,N_1615);
and U2152 (N_2152,N_1690,N_1986);
nand U2153 (N_2153,N_1747,N_1513);
or U2154 (N_2154,N_1895,N_1878);
or U2155 (N_2155,N_1752,N_1695);
nor U2156 (N_2156,N_1700,N_1672);
nor U2157 (N_2157,N_1897,N_1634);
and U2158 (N_2158,N_1985,N_1941);
and U2159 (N_2159,N_1818,N_1979);
nand U2160 (N_2160,N_1674,N_1798);
and U2161 (N_2161,N_1708,N_1527);
nand U2162 (N_2162,N_1907,N_1627);
nand U2163 (N_2163,N_1616,N_1874);
or U2164 (N_2164,N_1860,N_1557);
and U2165 (N_2165,N_1793,N_1741);
nand U2166 (N_2166,N_1596,N_1617);
and U2167 (N_2167,N_1950,N_1511);
or U2168 (N_2168,N_1709,N_1514);
or U2169 (N_2169,N_1910,N_1636);
and U2170 (N_2170,N_1723,N_1649);
or U2171 (N_2171,N_1525,N_1924);
or U2172 (N_2172,N_1641,N_1886);
xnor U2173 (N_2173,N_1556,N_1892);
nand U2174 (N_2174,N_1792,N_1676);
nand U2175 (N_2175,N_1932,N_1533);
and U2176 (N_2176,N_1980,N_1566);
or U2177 (N_2177,N_1929,N_1691);
nor U2178 (N_2178,N_1647,N_1852);
xnor U2179 (N_2179,N_1692,N_1953);
and U2180 (N_2180,N_1735,N_1642);
and U2181 (N_2181,N_1833,N_1751);
or U2182 (N_2182,N_1861,N_1965);
and U2183 (N_2183,N_1731,N_1547);
nand U2184 (N_2184,N_1969,N_1604);
and U2185 (N_2185,N_1964,N_1977);
nand U2186 (N_2186,N_1913,N_1764);
or U2187 (N_2187,N_1670,N_1951);
and U2188 (N_2188,N_1769,N_1906);
and U2189 (N_2189,N_1871,N_1739);
nor U2190 (N_2190,N_1820,N_1973);
nand U2191 (N_2191,N_1827,N_1947);
and U2192 (N_2192,N_1905,N_1908);
or U2193 (N_2193,N_1626,N_1705);
or U2194 (N_2194,N_1610,N_1625);
or U2195 (N_2195,N_1899,N_1630);
or U2196 (N_2196,N_1677,N_1923);
nor U2197 (N_2197,N_1534,N_1940);
or U2198 (N_2198,N_1598,N_1500);
nor U2199 (N_2199,N_1982,N_1952);
or U2200 (N_2200,N_1776,N_1862);
nor U2201 (N_2201,N_1919,N_1891);
and U2202 (N_2202,N_1603,N_1582);
or U2203 (N_2203,N_1854,N_1624);
or U2204 (N_2204,N_1605,N_1563);
or U2205 (N_2205,N_1715,N_1917);
nor U2206 (N_2206,N_1572,N_1749);
and U2207 (N_2207,N_1571,N_1577);
or U2208 (N_2208,N_1796,N_1771);
nand U2209 (N_2209,N_1535,N_1651);
and U2210 (N_2210,N_1539,N_1623);
and U2211 (N_2211,N_1516,N_1652);
nor U2212 (N_2212,N_1707,N_1853);
and U2213 (N_2213,N_1578,N_1552);
or U2214 (N_2214,N_1620,N_1868);
and U2215 (N_2215,N_1777,N_1714);
nand U2216 (N_2216,N_1856,N_1585);
nand U2217 (N_2217,N_1881,N_1996);
and U2218 (N_2218,N_1608,N_1666);
nand U2219 (N_2219,N_1909,N_1550);
nand U2220 (N_2220,N_1787,N_1761);
and U2221 (N_2221,N_1848,N_1825);
or U2222 (N_2222,N_1736,N_1814);
nor U2223 (N_2223,N_1782,N_1803);
nor U2224 (N_2224,N_1508,N_1538);
or U2225 (N_2225,N_1835,N_1569);
or U2226 (N_2226,N_1997,N_1713);
nand U2227 (N_2227,N_1659,N_1601);
and U2228 (N_2228,N_1963,N_1988);
nor U2229 (N_2229,N_1916,N_1890);
nand U2230 (N_2230,N_1944,N_1775);
nor U2231 (N_2231,N_1675,N_1826);
nor U2232 (N_2232,N_1958,N_1802);
and U2233 (N_2233,N_1884,N_1896);
and U2234 (N_2234,N_1678,N_1755);
nand U2235 (N_2235,N_1858,N_1942);
nor U2236 (N_2236,N_1960,N_1704);
nor U2237 (N_2237,N_1662,N_1904);
nand U2238 (N_2238,N_1728,N_1829);
xor U2239 (N_2239,N_1689,N_1599);
or U2240 (N_2240,N_1875,N_1734);
or U2241 (N_2241,N_1737,N_1710);
or U2242 (N_2242,N_1783,N_1553);
nand U2243 (N_2243,N_1836,N_1542);
or U2244 (N_2244,N_1948,N_1549);
and U2245 (N_2245,N_1872,N_1521);
nor U2246 (N_2246,N_1579,N_1537);
nor U2247 (N_2247,N_1719,N_1946);
or U2248 (N_2248,N_1515,N_1646);
nor U2249 (N_2249,N_1815,N_1762);
nor U2250 (N_2250,N_1983,N_1655);
nand U2251 (N_2251,N_1957,N_1683);
nor U2252 (N_2252,N_1733,N_1700);
nand U2253 (N_2253,N_1841,N_1915);
and U2254 (N_2254,N_1892,N_1874);
nor U2255 (N_2255,N_1883,N_1728);
nor U2256 (N_2256,N_1720,N_1739);
and U2257 (N_2257,N_1576,N_1852);
nor U2258 (N_2258,N_1761,N_1610);
or U2259 (N_2259,N_1803,N_1707);
nand U2260 (N_2260,N_1786,N_1745);
nand U2261 (N_2261,N_1586,N_1814);
nor U2262 (N_2262,N_1765,N_1935);
nor U2263 (N_2263,N_1618,N_1536);
nand U2264 (N_2264,N_1838,N_1712);
nand U2265 (N_2265,N_1995,N_1730);
nor U2266 (N_2266,N_1940,N_1727);
nand U2267 (N_2267,N_1906,N_1940);
and U2268 (N_2268,N_1643,N_1872);
nand U2269 (N_2269,N_1880,N_1507);
nor U2270 (N_2270,N_1906,N_1702);
and U2271 (N_2271,N_1758,N_1761);
or U2272 (N_2272,N_1679,N_1768);
nor U2273 (N_2273,N_1986,N_1718);
or U2274 (N_2274,N_1575,N_1881);
nor U2275 (N_2275,N_1733,N_1737);
nand U2276 (N_2276,N_1693,N_1986);
nand U2277 (N_2277,N_1632,N_1898);
and U2278 (N_2278,N_1527,N_1736);
or U2279 (N_2279,N_1889,N_1847);
or U2280 (N_2280,N_1627,N_1710);
and U2281 (N_2281,N_1691,N_1651);
xor U2282 (N_2282,N_1848,N_1618);
and U2283 (N_2283,N_1806,N_1795);
nand U2284 (N_2284,N_1958,N_1701);
nand U2285 (N_2285,N_1583,N_1783);
nand U2286 (N_2286,N_1598,N_1775);
nor U2287 (N_2287,N_1877,N_1656);
xor U2288 (N_2288,N_1577,N_1617);
nor U2289 (N_2289,N_1804,N_1696);
nor U2290 (N_2290,N_1532,N_1775);
nand U2291 (N_2291,N_1764,N_1943);
and U2292 (N_2292,N_1685,N_1795);
nand U2293 (N_2293,N_1676,N_1661);
xnor U2294 (N_2294,N_1872,N_1715);
and U2295 (N_2295,N_1684,N_1921);
nand U2296 (N_2296,N_1935,N_1925);
nor U2297 (N_2297,N_1954,N_1705);
and U2298 (N_2298,N_1562,N_1792);
nor U2299 (N_2299,N_1836,N_1895);
or U2300 (N_2300,N_1587,N_1884);
and U2301 (N_2301,N_1717,N_1524);
and U2302 (N_2302,N_1600,N_1750);
or U2303 (N_2303,N_1953,N_1913);
nor U2304 (N_2304,N_1752,N_1549);
nand U2305 (N_2305,N_1549,N_1849);
and U2306 (N_2306,N_1926,N_1883);
and U2307 (N_2307,N_1778,N_1548);
and U2308 (N_2308,N_1590,N_1698);
or U2309 (N_2309,N_1677,N_1540);
or U2310 (N_2310,N_1947,N_1793);
xor U2311 (N_2311,N_1584,N_1664);
nand U2312 (N_2312,N_1806,N_1819);
nand U2313 (N_2313,N_1818,N_1724);
nor U2314 (N_2314,N_1687,N_1951);
nand U2315 (N_2315,N_1785,N_1662);
nand U2316 (N_2316,N_1630,N_1644);
nand U2317 (N_2317,N_1618,N_1627);
and U2318 (N_2318,N_1656,N_1905);
nand U2319 (N_2319,N_1724,N_1672);
and U2320 (N_2320,N_1753,N_1704);
nand U2321 (N_2321,N_1643,N_1654);
or U2322 (N_2322,N_1985,N_1660);
and U2323 (N_2323,N_1880,N_1886);
and U2324 (N_2324,N_1700,N_1603);
xnor U2325 (N_2325,N_1566,N_1631);
nand U2326 (N_2326,N_1830,N_1821);
nor U2327 (N_2327,N_1706,N_1907);
nor U2328 (N_2328,N_1632,N_1763);
and U2329 (N_2329,N_1720,N_1548);
nor U2330 (N_2330,N_1643,N_1624);
or U2331 (N_2331,N_1664,N_1835);
nand U2332 (N_2332,N_1640,N_1800);
and U2333 (N_2333,N_1620,N_1946);
and U2334 (N_2334,N_1837,N_1937);
nor U2335 (N_2335,N_1567,N_1518);
or U2336 (N_2336,N_1730,N_1864);
or U2337 (N_2337,N_1776,N_1886);
nand U2338 (N_2338,N_1937,N_1891);
nand U2339 (N_2339,N_1547,N_1773);
or U2340 (N_2340,N_1824,N_1879);
or U2341 (N_2341,N_1732,N_1711);
or U2342 (N_2342,N_1758,N_1879);
or U2343 (N_2343,N_1766,N_1753);
and U2344 (N_2344,N_1906,N_1984);
nand U2345 (N_2345,N_1810,N_1782);
or U2346 (N_2346,N_1608,N_1639);
nor U2347 (N_2347,N_1692,N_1836);
and U2348 (N_2348,N_1521,N_1501);
nor U2349 (N_2349,N_1617,N_1741);
or U2350 (N_2350,N_1725,N_1645);
and U2351 (N_2351,N_1590,N_1587);
nor U2352 (N_2352,N_1772,N_1983);
nor U2353 (N_2353,N_1975,N_1768);
or U2354 (N_2354,N_1801,N_1822);
nand U2355 (N_2355,N_1527,N_1668);
or U2356 (N_2356,N_1906,N_1561);
or U2357 (N_2357,N_1853,N_1616);
nor U2358 (N_2358,N_1557,N_1875);
nor U2359 (N_2359,N_1647,N_1687);
nor U2360 (N_2360,N_1800,N_1880);
nor U2361 (N_2361,N_1800,N_1716);
and U2362 (N_2362,N_1812,N_1621);
nor U2363 (N_2363,N_1971,N_1986);
and U2364 (N_2364,N_1642,N_1821);
nor U2365 (N_2365,N_1512,N_1553);
nor U2366 (N_2366,N_1503,N_1602);
nor U2367 (N_2367,N_1735,N_1699);
nand U2368 (N_2368,N_1529,N_1505);
nand U2369 (N_2369,N_1713,N_1979);
nand U2370 (N_2370,N_1755,N_1575);
nor U2371 (N_2371,N_1677,N_1587);
nand U2372 (N_2372,N_1567,N_1521);
nand U2373 (N_2373,N_1629,N_1791);
nor U2374 (N_2374,N_1519,N_1919);
nand U2375 (N_2375,N_1940,N_1692);
and U2376 (N_2376,N_1639,N_1854);
nand U2377 (N_2377,N_1538,N_1844);
nand U2378 (N_2378,N_1821,N_1937);
or U2379 (N_2379,N_1749,N_1552);
xnor U2380 (N_2380,N_1821,N_1991);
nor U2381 (N_2381,N_1688,N_1920);
nor U2382 (N_2382,N_1561,N_1898);
nand U2383 (N_2383,N_1530,N_1882);
nand U2384 (N_2384,N_1982,N_1831);
nand U2385 (N_2385,N_1839,N_1798);
xnor U2386 (N_2386,N_1798,N_1662);
nand U2387 (N_2387,N_1612,N_1642);
nand U2388 (N_2388,N_1738,N_1614);
and U2389 (N_2389,N_1859,N_1869);
nor U2390 (N_2390,N_1841,N_1812);
and U2391 (N_2391,N_1604,N_1914);
nand U2392 (N_2392,N_1590,N_1533);
and U2393 (N_2393,N_1744,N_1628);
nor U2394 (N_2394,N_1513,N_1893);
nand U2395 (N_2395,N_1622,N_1874);
or U2396 (N_2396,N_1824,N_1562);
and U2397 (N_2397,N_1593,N_1516);
nand U2398 (N_2398,N_1964,N_1755);
nor U2399 (N_2399,N_1941,N_1561);
nand U2400 (N_2400,N_1567,N_1734);
xor U2401 (N_2401,N_1702,N_1914);
nor U2402 (N_2402,N_1585,N_1948);
and U2403 (N_2403,N_1952,N_1938);
nand U2404 (N_2404,N_1899,N_1938);
nor U2405 (N_2405,N_1589,N_1637);
nor U2406 (N_2406,N_1776,N_1796);
or U2407 (N_2407,N_1734,N_1848);
nand U2408 (N_2408,N_1750,N_1748);
nand U2409 (N_2409,N_1617,N_1725);
nor U2410 (N_2410,N_1612,N_1617);
and U2411 (N_2411,N_1552,N_1956);
or U2412 (N_2412,N_1831,N_1929);
or U2413 (N_2413,N_1723,N_1654);
or U2414 (N_2414,N_1660,N_1729);
xor U2415 (N_2415,N_1939,N_1673);
nand U2416 (N_2416,N_1953,N_1645);
and U2417 (N_2417,N_1868,N_1701);
or U2418 (N_2418,N_1844,N_1942);
or U2419 (N_2419,N_1832,N_1660);
and U2420 (N_2420,N_1773,N_1724);
xnor U2421 (N_2421,N_1685,N_1701);
nand U2422 (N_2422,N_1827,N_1956);
nand U2423 (N_2423,N_1935,N_1833);
or U2424 (N_2424,N_1810,N_1727);
nor U2425 (N_2425,N_1783,N_1786);
nand U2426 (N_2426,N_1760,N_1608);
nor U2427 (N_2427,N_1511,N_1666);
nor U2428 (N_2428,N_1541,N_1995);
and U2429 (N_2429,N_1641,N_1592);
and U2430 (N_2430,N_1905,N_1628);
nand U2431 (N_2431,N_1764,N_1902);
nand U2432 (N_2432,N_1889,N_1585);
nor U2433 (N_2433,N_1763,N_1810);
xor U2434 (N_2434,N_1741,N_1923);
nand U2435 (N_2435,N_1855,N_1544);
or U2436 (N_2436,N_1652,N_1849);
nand U2437 (N_2437,N_1699,N_1532);
nor U2438 (N_2438,N_1554,N_1993);
or U2439 (N_2439,N_1750,N_1861);
nor U2440 (N_2440,N_1564,N_1862);
nand U2441 (N_2441,N_1504,N_1891);
or U2442 (N_2442,N_1816,N_1972);
or U2443 (N_2443,N_1728,N_1665);
or U2444 (N_2444,N_1591,N_1586);
and U2445 (N_2445,N_1973,N_1869);
nor U2446 (N_2446,N_1685,N_1689);
or U2447 (N_2447,N_1746,N_1548);
nand U2448 (N_2448,N_1976,N_1842);
or U2449 (N_2449,N_1604,N_1575);
or U2450 (N_2450,N_1639,N_1829);
nand U2451 (N_2451,N_1506,N_1921);
nor U2452 (N_2452,N_1897,N_1984);
and U2453 (N_2453,N_1626,N_1507);
and U2454 (N_2454,N_1780,N_1945);
and U2455 (N_2455,N_1539,N_1964);
nand U2456 (N_2456,N_1697,N_1816);
nand U2457 (N_2457,N_1992,N_1656);
and U2458 (N_2458,N_1826,N_1942);
nor U2459 (N_2459,N_1513,N_1619);
nand U2460 (N_2460,N_1610,N_1732);
nand U2461 (N_2461,N_1632,N_1729);
nand U2462 (N_2462,N_1637,N_1843);
and U2463 (N_2463,N_1509,N_1566);
nand U2464 (N_2464,N_1601,N_1766);
nor U2465 (N_2465,N_1847,N_1785);
and U2466 (N_2466,N_1538,N_1716);
nor U2467 (N_2467,N_1545,N_1601);
or U2468 (N_2468,N_1811,N_1943);
or U2469 (N_2469,N_1588,N_1954);
nor U2470 (N_2470,N_1640,N_1863);
or U2471 (N_2471,N_1579,N_1526);
and U2472 (N_2472,N_1614,N_1596);
and U2473 (N_2473,N_1610,N_1970);
or U2474 (N_2474,N_1897,N_1853);
or U2475 (N_2475,N_1815,N_1516);
nand U2476 (N_2476,N_1543,N_1680);
nor U2477 (N_2477,N_1639,N_1935);
and U2478 (N_2478,N_1521,N_1717);
and U2479 (N_2479,N_1605,N_1894);
and U2480 (N_2480,N_1985,N_1836);
nand U2481 (N_2481,N_1582,N_1964);
nand U2482 (N_2482,N_1903,N_1817);
nor U2483 (N_2483,N_1730,N_1909);
or U2484 (N_2484,N_1846,N_1834);
and U2485 (N_2485,N_1531,N_1882);
nand U2486 (N_2486,N_1918,N_1519);
nand U2487 (N_2487,N_1851,N_1976);
and U2488 (N_2488,N_1764,N_1818);
or U2489 (N_2489,N_1901,N_1542);
and U2490 (N_2490,N_1702,N_1507);
nor U2491 (N_2491,N_1981,N_1533);
and U2492 (N_2492,N_1807,N_1900);
nor U2493 (N_2493,N_1974,N_1888);
nand U2494 (N_2494,N_1611,N_1988);
nor U2495 (N_2495,N_1719,N_1817);
nor U2496 (N_2496,N_1896,N_1789);
nor U2497 (N_2497,N_1522,N_1902);
nor U2498 (N_2498,N_1882,N_1870);
nand U2499 (N_2499,N_1814,N_1558);
or U2500 (N_2500,N_2023,N_2002);
nor U2501 (N_2501,N_2054,N_2171);
and U2502 (N_2502,N_2466,N_2018);
nor U2503 (N_2503,N_2307,N_2057);
or U2504 (N_2504,N_2425,N_2136);
xor U2505 (N_2505,N_2281,N_2473);
and U2506 (N_2506,N_2340,N_2488);
nand U2507 (N_2507,N_2456,N_2304);
nand U2508 (N_2508,N_2076,N_2247);
nand U2509 (N_2509,N_2491,N_2090);
nor U2510 (N_2510,N_2036,N_2276);
nor U2511 (N_2511,N_2167,N_2396);
and U2512 (N_2512,N_2052,N_2319);
and U2513 (N_2513,N_2311,N_2221);
nand U2514 (N_2514,N_2370,N_2371);
nand U2515 (N_2515,N_2358,N_2365);
or U2516 (N_2516,N_2441,N_2055);
nor U2517 (N_2517,N_2048,N_2306);
or U2518 (N_2518,N_2046,N_2197);
or U2519 (N_2519,N_2061,N_2015);
nor U2520 (N_2520,N_2176,N_2087);
and U2521 (N_2521,N_2336,N_2434);
xor U2522 (N_2522,N_2085,N_2162);
nand U2523 (N_2523,N_2458,N_2435);
xnor U2524 (N_2524,N_2022,N_2160);
and U2525 (N_2525,N_2344,N_2361);
nand U2526 (N_2526,N_2495,N_2449);
xnor U2527 (N_2527,N_2134,N_2129);
nand U2528 (N_2528,N_2128,N_2075);
nor U2529 (N_2529,N_2418,N_2012);
and U2530 (N_2530,N_2343,N_2337);
and U2531 (N_2531,N_2393,N_2173);
nand U2532 (N_2532,N_2328,N_2367);
nor U2533 (N_2533,N_2230,N_2077);
nand U2534 (N_2534,N_2264,N_2493);
nor U2535 (N_2535,N_2137,N_2364);
and U2536 (N_2536,N_2375,N_2424);
and U2537 (N_2537,N_2121,N_2079);
and U2538 (N_2538,N_2163,N_2170);
or U2539 (N_2539,N_2106,N_2356);
nor U2540 (N_2540,N_2081,N_2334);
nor U2541 (N_2541,N_2420,N_2395);
nand U2542 (N_2542,N_2279,N_2406);
and U2543 (N_2543,N_2013,N_2189);
or U2544 (N_2544,N_2125,N_2383);
and U2545 (N_2545,N_2470,N_2194);
and U2546 (N_2546,N_2417,N_2192);
nor U2547 (N_2547,N_2070,N_2198);
or U2548 (N_2548,N_2296,N_2133);
nand U2549 (N_2549,N_2154,N_2225);
xnor U2550 (N_2550,N_2404,N_2043);
nand U2551 (N_2551,N_2402,N_2056);
nand U2552 (N_2552,N_2032,N_2244);
nor U2553 (N_2553,N_2258,N_2038);
nand U2554 (N_2554,N_2316,N_2411);
nand U2555 (N_2555,N_2138,N_2444);
nand U2556 (N_2556,N_2332,N_2115);
xnor U2557 (N_2557,N_2146,N_2159);
or U2558 (N_2558,N_2041,N_2156);
and U2559 (N_2559,N_2166,N_2219);
or U2560 (N_2560,N_2331,N_2263);
nand U2561 (N_2561,N_2271,N_2432);
nand U2562 (N_2562,N_2130,N_2031);
nand U2563 (N_2563,N_2141,N_2489);
and U2564 (N_2564,N_2408,N_2414);
or U2565 (N_2565,N_2284,N_2468);
or U2566 (N_2566,N_2014,N_2461);
or U2567 (N_2567,N_2283,N_2436);
nor U2568 (N_2568,N_2157,N_2241);
or U2569 (N_2569,N_2481,N_2063);
xor U2570 (N_2570,N_2437,N_2253);
nor U2571 (N_2571,N_2161,N_2153);
xor U2572 (N_2572,N_2428,N_2246);
nand U2573 (N_2573,N_2182,N_2286);
and U2574 (N_2574,N_2155,N_2397);
nand U2575 (N_2575,N_2386,N_2262);
or U2576 (N_2576,N_2302,N_2080);
and U2577 (N_2577,N_2289,N_2037);
nand U2578 (N_2578,N_2103,N_2205);
nor U2579 (N_2579,N_2313,N_2412);
and U2580 (N_2580,N_2423,N_2147);
nand U2581 (N_2581,N_2497,N_2272);
nor U2582 (N_2582,N_2025,N_2116);
or U2583 (N_2583,N_2407,N_2045);
and U2584 (N_2584,N_2342,N_2238);
or U2585 (N_2585,N_2381,N_2255);
or U2586 (N_2586,N_2024,N_2445);
nor U2587 (N_2587,N_2195,N_2148);
nand U2588 (N_2588,N_2360,N_2236);
nand U2589 (N_2589,N_2318,N_2300);
or U2590 (N_2590,N_2474,N_2480);
and U2591 (N_2591,N_2193,N_2299);
and U2592 (N_2592,N_2034,N_2039);
or U2593 (N_2593,N_2355,N_2377);
or U2594 (N_2594,N_2265,N_2359);
nand U2595 (N_2595,N_2073,N_2463);
nor U2596 (N_2596,N_2347,N_2357);
nand U2597 (N_2597,N_2252,N_2292);
and U2598 (N_2598,N_2184,N_2226);
nand U2599 (N_2599,N_2174,N_2450);
nand U2600 (N_2600,N_2006,N_2059);
or U2601 (N_2601,N_2113,N_2310);
and U2602 (N_2602,N_2314,N_2249);
nand U2603 (N_2603,N_2227,N_2308);
or U2604 (N_2604,N_2351,N_2442);
or U2605 (N_2605,N_2260,N_2487);
or U2606 (N_2606,N_2232,N_2295);
and U2607 (N_2607,N_2330,N_2499);
nor U2608 (N_2608,N_2060,N_2496);
nor U2609 (N_2609,N_2020,N_2168);
nand U2610 (N_2610,N_2224,N_2105);
and U2611 (N_2611,N_2362,N_2096);
nand U2612 (N_2612,N_2145,N_2030);
nor U2613 (N_2613,N_2326,N_2151);
and U2614 (N_2614,N_2352,N_2144);
nand U2615 (N_2615,N_2140,N_2349);
nand U2616 (N_2616,N_2421,N_2233);
nor U2617 (N_2617,N_2483,N_2119);
and U2618 (N_2618,N_2380,N_2471);
or U2619 (N_2619,N_2186,N_2250);
nor U2620 (N_2620,N_2329,N_2216);
and U2621 (N_2621,N_2178,N_2467);
or U2622 (N_2622,N_2009,N_2438);
or U2623 (N_2623,N_2212,N_2150);
nor U2624 (N_2624,N_2222,N_2053);
or U2625 (N_2625,N_2234,N_2183);
and U2626 (N_2626,N_2312,N_2203);
or U2627 (N_2627,N_2350,N_2447);
nand U2628 (N_2628,N_2282,N_2069);
xor U2629 (N_2629,N_2218,N_2280);
and U2630 (N_2630,N_2152,N_2430);
or U2631 (N_2631,N_2089,N_2068);
xnor U2632 (N_2632,N_2259,N_2305);
and U2633 (N_2633,N_2142,N_2426);
and U2634 (N_2634,N_2338,N_2172);
and U2635 (N_2635,N_2187,N_2256);
or U2636 (N_2636,N_2223,N_2028);
nand U2637 (N_2637,N_2066,N_2108);
nor U2638 (N_2638,N_2107,N_2100);
nor U2639 (N_2639,N_2165,N_2391);
nor U2640 (N_2640,N_2476,N_2181);
nor U2641 (N_2641,N_2354,N_2242);
or U2642 (N_2642,N_2398,N_2209);
or U2643 (N_2643,N_2095,N_2261);
or U2644 (N_2644,N_2118,N_2084);
nand U2645 (N_2645,N_2062,N_2453);
nand U2646 (N_2646,N_2422,N_2050);
and U2647 (N_2647,N_2029,N_2498);
and U2648 (N_2648,N_2078,N_2429);
and U2649 (N_2649,N_2245,N_2058);
nor U2650 (N_2650,N_2376,N_2124);
or U2651 (N_2651,N_2215,N_2196);
nor U2652 (N_2652,N_2472,N_2237);
nand U2653 (N_2653,N_2044,N_2410);
or U2654 (N_2654,N_2452,N_2290);
and U2655 (N_2655,N_2475,N_2094);
or U2656 (N_2656,N_2372,N_2093);
and U2657 (N_2657,N_2072,N_2287);
or U2658 (N_2658,N_2460,N_2026);
or U2659 (N_2659,N_2179,N_2341);
nor U2660 (N_2660,N_2104,N_2071);
or U2661 (N_2661,N_2158,N_2353);
or U2662 (N_2662,N_2346,N_2019);
and U2663 (N_2663,N_2220,N_2405);
or U2664 (N_2664,N_2114,N_2240);
nor U2665 (N_2665,N_2419,N_2027);
or U2666 (N_2666,N_2016,N_2401);
nand U2667 (N_2667,N_2007,N_2088);
nor U2668 (N_2668,N_2132,N_2228);
nor U2669 (N_2669,N_2469,N_2321);
and U2670 (N_2670,N_2462,N_2214);
and U2671 (N_2671,N_2248,N_2064);
nor U2672 (N_2672,N_2294,N_2035);
nand U2673 (N_2673,N_2243,N_2102);
nand U2674 (N_2674,N_2266,N_2455);
nand U2675 (N_2675,N_2177,N_2049);
or U2676 (N_2676,N_2413,N_2122);
nand U2677 (N_2677,N_2051,N_2099);
nand U2678 (N_2678,N_2086,N_2010);
nand U2679 (N_2679,N_2040,N_2001);
nand U2680 (N_2680,N_2217,N_2004);
and U2681 (N_2681,N_2185,N_2126);
nor U2682 (N_2682,N_2082,N_2439);
nand U2683 (N_2683,N_2399,N_2288);
or U2684 (N_2684,N_2309,N_2169);
xnor U2685 (N_2685,N_2301,N_2005);
or U2686 (N_2686,N_2324,N_2111);
nand U2687 (N_2687,N_2098,N_2327);
nor U2688 (N_2688,N_2494,N_2257);
nor U2689 (N_2689,N_2490,N_2083);
nand U2690 (N_2690,N_2229,N_2433);
xor U2691 (N_2691,N_2394,N_2385);
nand U2692 (N_2692,N_2091,N_2369);
nor U2693 (N_2693,N_2454,N_2191);
or U2694 (N_2694,N_2431,N_2188);
nand U2695 (N_2695,N_2415,N_2202);
and U2696 (N_2696,N_2373,N_2325);
or U2697 (N_2697,N_2251,N_2204);
nand U2698 (N_2698,N_2149,N_2267);
nor U2699 (N_2699,N_2273,N_2291);
or U2700 (N_2700,N_2190,N_2478);
and U2701 (N_2701,N_2275,N_2368);
and U2702 (N_2702,N_2384,N_2274);
nand U2703 (N_2703,N_2123,N_2403);
and U2704 (N_2704,N_2366,N_2000);
nor U2705 (N_2705,N_2235,N_2277);
or U2706 (N_2706,N_2127,N_2363);
nand U2707 (N_2707,N_2033,N_2293);
nor U2708 (N_2708,N_2207,N_2201);
nand U2709 (N_2709,N_2427,N_2479);
or U2710 (N_2710,N_2269,N_2484);
nor U2711 (N_2711,N_2139,N_2416);
and U2712 (N_2712,N_2348,N_2389);
nor U2713 (N_2713,N_2482,N_2448);
and U2714 (N_2714,N_2392,N_2199);
and U2715 (N_2715,N_2200,N_2388);
and U2716 (N_2716,N_2109,N_2297);
nor U2717 (N_2717,N_2042,N_2323);
nand U2718 (N_2718,N_2017,N_2335);
and U2719 (N_2719,N_2477,N_2345);
and U2720 (N_2720,N_2239,N_2213);
nand U2721 (N_2721,N_2131,N_2390);
nor U2722 (N_2722,N_2011,N_2210);
or U2723 (N_2723,N_2315,N_2021);
or U2724 (N_2724,N_2065,N_2175);
nand U2725 (N_2725,N_2101,N_2112);
xor U2726 (N_2726,N_2231,N_2092);
nor U2727 (N_2727,N_2374,N_2008);
and U2728 (N_2728,N_2409,N_2097);
nand U2729 (N_2729,N_2485,N_2464);
nor U2730 (N_2730,N_2067,N_2180);
xor U2731 (N_2731,N_2285,N_2378);
xor U2732 (N_2732,N_2074,N_2440);
or U2733 (N_2733,N_2492,N_2443);
or U2734 (N_2734,N_2457,N_2339);
nand U2735 (N_2735,N_2322,N_2382);
and U2736 (N_2736,N_2143,N_2047);
and U2737 (N_2737,N_2110,N_2320);
nor U2738 (N_2738,N_2003,N_2387);
and U2739 (N_2739,N_2211,N_2268);
xor U2740 (N_2740,N_2333,N_2270);
and U2741 (N_2741,N_2117,N_2486);
nand U2742 (N_2742,N_2120,N_2303);
nor U2743 (N_2743,N_2446,N_2379);
nor U2744 (N_2744,N_2465,N_2206);
or U2745 (N_2745,N_2278,N_2298);
nand U2746 (N_2746,N_2459,N_2400);
nor U2747 (N_2747,N_2451,N_2208);
and U2748 (N_2748,N_2164,N_2317);
and U2749 (N_2749,N_2135,N_2254);
nand U2750 (N_2750,N_2444,N_2362);
nor U2751 (N_2751,N_2166,N_2435);
xnor U2752 (N_2752,N_2157,N_2018);
nand U2753 (N_2753,N_2393,N_2114);
nor U2754 (N_2754,N_2014,N_2005);
nand U2755 (N_2755,N_2072,N_2006);
or U2756 (N_2756,N_2428,N_2251);
and U2757 (N_2757,N_2271,N_2308);
or U2758 (N_2758,N_2221,N_2398);
and U2759 (N_2759,N_2387,N_2201);
nor U2760 (N_2760,N_2004,N_2243);
nor U2761 (N_2761,N_2000,N_2139);
and U2762 (N_2762,N_2267,N_2176);
nand U2763 (N_2763,N_2344,N_2429);
nor U2764 (N_2764,N_2329,N_2138);
nand U2765 (N_2765,N_2317,N_2159);
and U2766 (N_2766,N_2431,N_2197);
nor U2767 (N_2767,N_2248,N_2093);
and U2768 (N_2768,N_2334,N_2389);
and U2769 (N_2769,N_2045,N_2079);
nand U2770 (N_2770,N_2151,N_2351);
and U2771 (N_2771,N_2061,N_2009);
nand U2772 (N_2772,N_2139,N_2173);
nor U2773 (N_2773,N_2283,N_2416);
nor U2774 (N_2774,N_2249,N_2041);
nand U2775 (N_2775,N_2110,N_2064);
nand U2776 (N_2776,N_2284,N_2300);
nand U2777 (N_2777,N_2236,N_2195);
or U2778 (N_2778,N_2435,N_2381);
or U2779 (N_2779,N_2390,N_2479);
or U2780 (N_2780,N_2184,N_2064);
or U2781 (N_2781,N_2001,N_2321);
nand U2782 (N_2782,N_2348,N_2306);
nor U2783 (N_2783,N_2242,N_2265);
nand U2784 (N_2784,N_2164,N_2019);
nor U2785 (N_2785,N_2312,N_2093);
nand U2786 (N_2786,N_2345,N_2229);
and U2787 (N_2787,N_2406,N_2150);
or U2788 (N_2788,N_2406,N_2231);
and U2789 (N_2789,N_2030,N_2397);
xnor U2790 (N_2790,N_2396,N_2140);
nor U2791 (N_2791,N_2403,N_2143);
or U2792 (N_2792,N_2325,N_2422);
or U2793 (N_2793,N_2217,N_2337);
nand U2794 (N_2794,N_2435,N_2453);
or U2795 (N_2795,N_2127,N_2189);
or U2796 (N_2796,N_2482,N_2091);
nand U2797 (N_2797,N_2031,N_2201);
nand U2798 (N_2798,N_2336,N_2454);
or U2799 (N_2799,N_2477,N_2030);
nor U2800 (N_2800,N_2482,N_2073);
or U2801 (N_2801,N_2139,N_2330);
nand U2802 (N_2802,N_2022,N_2366);
and U2803 (N_2803,N_2422,N_2271);
or U2804 (N_2804,N_2101,N_2177);
and U2805 (N_2805,N_2136,N_2069);
and U2806 (N_2806,N_2359,N_2280);
and U2807 (N_2807,N_2063,N_2006);
and U2808 (N_2808,N_2022,N_2024);
and U2809 (N_2809,N_2374,N_2361);
nor U2810 (N_2810,N_2446,N_2020);
and U2811 (N_2811,N_2472,N_2477);
nand U2812 (N_2812,N_2008,N_2160);
nor U2813 (N_2813,N_2297,N_2379);
xnor U2814 (N_2814,N_2130,N_2180);
and U2815 (N_2815,N_2118,N_2211);
or U2816 (N_2816,N_2134,N_2193);
nor U2817 (N_2817,N_2123,N_2432);
and U2818 (N_2818,N_2175,N_2387);
nand U2819 (N_2819,N_2317,N_2133);
nand U2820 (N_2820,N_2175,N_2485);
nand U2821 (N_2821,N_2370,N_2250);
or U2822 (N_2822,N_2014,N_2024);
nand U2823 (N_2823,N_2007,N_2479);
nand U2824 (N_2824,N_2239,N_2339);
nand U2825 (N_2825,N_2212,N_2273);
and U2826 (N_2826,N_2298,N_2489);
and U2827 (N_2827,N_2320,N_2307);
or U2828 (N_2828,N_2257,N_2363);
and U2829 (N_2829,N_2329,N_2479);
nand U2830 (N_2830,N_2319,N_2433);
or U2831 (N_2831,N_2345,N_2132);
nor U2832 (N_2832,N_2457,N_2295);
xnor U2833 (N_2833,N_2477,N_2065);
and U2834 (N_2834,N_2473,N_2292);
xor U2835 (N_2835,N_2139,N_2424);
nor U2836 (N_2836,N_2441,N_2045);
nor U2837 (N_2837,N_2467,N_2036);
or U2838 (N_2838,N_2366,N_2498);
and U2839 (N_2839,N_2220,N_2120);
and U2840 (N_2840,N_2222,N_2485);
nand U2841 (N_2841,N_2163,N_2091);
nor U2842 (N_2842,N_2150,N_2347);
and U2843 (N_2843,N_2398,N_2043);
and U2844 (N_2844,N_2389,N_2056);
nor U2845 (N_2845,N_2425,N_2491);
or U2846 (N_2846,N_2396,N_2181);
and U2847 (N_2847,N_2325,N_2300);
and U2848 (N_2848,N_2011,N_2024);
nand U2849 (N_2849,N_2399,N_2191);
and U2850 (N_2850,N_2034,N_2229);
nor U2851 (N_2851,N_2325,N_2071);
and U2852 (N_2852,N_2356,N_2295);
or U2853 (N_2853,N_2085,N_2053);
and U2854 (N_2854,N_2101,N_2263);
and U2855 (N_2855,N_2098,N_2207);
and U2856 (N_2856,N_2485,N_2390);
and U2857 (N_2857,N_2415,N_2305);
and U2858 (N_2858,N_2378,N_2099);
or U2859 (N_2859,N_2018,N_2418);
nand U2860 (N_2860,N_2161,N_2408);
or U2861 (N_2861,N_2099,N_2435);
nor U2862 (N_2862,N_2158,N_2430);
nor U2863 (N_2863,N_2287,N_2387);
nor U2864 (N_2864,N_2466,N_2072);
or U2865 (N_2865,N_2031,N_2255);
nand U2866 (N_2866,N_2010,N_2257);
or U2867 (N_2867,N_2474,N_2270);
or U2868 (N_2868,N_2488,N_2246);
nor U2869 (N_2869,N_2287,N_2495);
and U2870 (N_2870,N_2179,N_2027);
or U2871 (N_2871,N_2201,N_2048);
or U2872 (N_2872,N_2203,N_2010);
or U2873 (N_2873,N_2419,N_2126);
and U2874 (N_2874,N_2353,N_2458);
and U2875 (N_2875,N_2228,N_2020);
or U2876 (N_2876,N_2392,N_2461);
nor U2877 (N_2877,N_2082,N_2202);
nor U2878 (N_2878,N_2086,N_2416);
and U2879 (N_2879,N_2035,N_2101);
nand U2880 (N_2880,N_2386,N_2164);
nor U2881 (N_2881,N_2461,N_2151);
nor U2882 (N_2882,N_2011,N_2163);
and U2883 (N_2883,N_2405,N_2173);
nand U2884 (N_2884,N_2226,N_2020);
nand U2885 (N_2885,N_2081,N_2309);
nor U2886 (N_2886,N_2386,N_2136);
nand U2887 (N_2887,N_2084,N_2193);
or U2888 (N_2888,N_2118,N_2083);
nor U2889 (N_2889,N_2324,N_2039);
nand U2890 (N_2890,N_2382,N_2059);
or U2891 (N_2891,N_2048,N_2461);
nor U2892 (N_2892,N_2257,N_2373);
nand U2893 (N_2893,N_2321,N_2453);
nor U2894 (N_2894,N_2399,N_2229);
or U2895 (N_2895,N_2398,N_2141);
nor U2896 (N_2896,N_2060,N_2126);
or U2897 (N_2897,N_2049,N_2277);
nand U2898 (N_2898,N_2336,N_2460);
nand U2899 (N_2899,N_2167,N_2344);
or U2900 (N_2900,N_2035,N_2481);
or U2901 (N_2901,N_2163,N_2265);
nor U2902 (N_2902,N_2389,N_2333);
and U2903 (N_2903,N_2145,N_2201);
nand U2904 (N_2904,N_2277,N_2191);
and U2905 (N_2905,N_2167,N_2018);
nor U2906 (N_2906,N_2111,N_2340);
nand U2907 (N_2907,N_2313,N_2042);
nor U2908 (N_2908,N_2244,N_2333);
and U2909 (N_2909,N_2420,N_2364);
and U2910 (N_2910,N_2290,N_2078);
or U2911 (N_2911,N_2416,N_2494);
or U2912 (N_2912,N_2279,N_2014);
nand U2913 (N_2913,N_2009,N_2310);
nand U2914 (N_2914,N_2405,N_2112);
and U2915 (N_2915,N_2132,N_2087);
nand U2916 (N_2916,N_2147,N_2191);
nand U2917 (N_2917,N_2326,N_2042);
nand U2918 (N_2918,N_2186,N_2231);
nor U2919 (N_2919,N_2285,N_2166);
nand U2920 (N_2920,N_2359,N_2226);
and U2921 (N_2921,N_2048,N_2284);
nand U2922 (N_2922,N_2064,N_2361);
or U2923 (N_2923,N_2112,N_2225);
nand U2924 (N_2924,N_2207,N_2334);
and U2925 (N_2925,N_2175,N_2459);
nand U2926 (N_2926,N_2073,N_2379);
or U2927 (N_2927,N_2022,N_2129);
nor U2928 (N_2928,N_2206,N_2331);
xnor U2929 (N_2929,N_2174,N_2307);
or U2930 (N_2930,N_2244,N_2133);
or U2931 (N_2931,N_2398,N_2264);
and U2932 (N_2932,N_2272,N_2016);
or U2933 (N_2933,N_2475,N_2343);
nor U2934 (N_2934,N_2050,N_2360);
and U2935 (N_2935,N_2284,N_2397);
nor U2936 (N_2936,N_2187,N_2200);
nor U2937 (N_2937,N_2313,N_2233);
nor U2938 (N_2938,N_2151,N_2268);
nand U2939 (N_2939,N_2091,N_2323);
and U2940 (N_2940,N_2471,N_2498);
nor U2941 (N_2941,N_2278,N_2096);
nand U2942 (N_2942,N_2443,N_2030);
nand U2943 (N_2943,N_2353,N_2394);
and U2944 (N_2944,N_2153,N_2193);
and U2945 (N_2945,N_2028,N_2442);
and U2946 (N_2946,N_2238,N_2340);
or U2947 (N_2947,N_2461,N_2296);
nor U2948 (N_2948,N_2361,N_2050);
or U2949 (N_2949,N_2130,N_2363);
and U2950 (N_2950,N_2154,N_2456);
nand U2951 (N_2951,N_2051,N_2138);
or U2952 (N_2952,N_2123,N_2355);
nand U2953 (N_2953,N_2350,N_2142);
nor U2954 (N_2954,N_2075,N_2185);
and U2955 (N_2955,N_2364,N_2139);
and U2956 (N_2956,N_2347,N_2479);
nand U2957 (N_2957,N_2199,N_2229);
or U2958 (N_2958,N_2463,N_2284);
xor U2959 (N_2959,N_2353,N_2110);
or U2960 (N_2960,N_2197,N_2120);
nand U2961 (N_2961,N_2145,N_2004);
nor U2962 (N_2962,N_2197,N_2086);
or U2963 (N_2963,N_2395,N_2109);
and U2964 (N_2964,N_2157,N_2316);
or U2965 (N_2965,N_2123,N_2044);
xor U2966 (N_2966,N_2023,N_2418);
and U2967 (N_2967,N_2149,N_2067);
and U2968 (N_2968,N_2403,N_2368);
nand U2969 (N_2969,N_2223,N_2234);
nor U2970 (N_2970,N_2195,N_2006);
and U2971 (N_2971,N_2210,N_2102);
nor U2972 (N_2972,N_2088,N_2107);
and U2973 (N_2973,N_2287,N_2003);
nor U2974 (N_2974,N_2412,N_2291);
xnor U2975 (N_2975,N_2350,N_2388);
nand U2976 (N_2976,N_2350,N_2277);
nor U2977 (N_2977,N_2018,N_2098);
or U2978 (N_2978,N_2008,N_2091);
or U2979 (N_2979,N_2138,N_2344);
and U2980 (N_2980,N_2246,N_2170);
nand U2981 (N_2981,N_2476,N_2463);
or U2982 (N_2982,N_2277,N_2373);
nand U2983 (N_2983,N_2160,N_2455);
or U2984 (N_2984,N_2148,N_2028);
nor U2985 (N_2985,N_2486,N_2197);
nor U2986 (N_2986,N_2288,N_2093);
nor U2987 (N_2987,N_2449,N_2178);
nor U2988 (N_2988,N_2418,N_2101);
nand U2989 (N_2989,N_2222,N_2444);
and U2990 (N_2990,N_2444,N_2066);
nor U2991 (N_2991,N_2356,N_2183);
or U2992 (N_2992,N_2274,N_2188);
nand U2993 (N_2993,N_2017,N_2173);
or U2994 (N_2994,N_2371,N_2122);
xnor U2995 (N_2995,N_2026,N_2272);
or U2996 (N_2996,N_2146,N_2367);
nor U2997 (N_2997,N_2280,N_2437);
nor U2998 (N_2998,N_2277,N_2399);
and U2999 (N_2999,N_2022,N_2282);
and U3000 (N_3000,N_2732,N_2789);
or U3001 (N_3001,N_2999,N_2517);
nor U3002 (N_3002,N_2840,N_2562);
nand U3003 (N_3003,N_2855,N_2996);
xnor U3004 (N_3004,N_2969,N_2706);
nand U3005 (N_3005,N_2971,N_2619);
xor U3006 (N_3006,N_2584,N_2565);
and U3007 (N_3007,N_2776,N_2921);
or U3008 (N_3008,N_2734,N_2575);
nor U3009 (N_3009,N_2653,N_2862);
nand U3010 (N_3010,N_2908,N_2987);
or U3011 (N_3011,N_2590,N_2952);
nand U3012 (N_3012,N_2784,N_2697);
nor U3013 (N_3013,N_2695,N_2633);
and U3014 (N_3014,N_2675,N_2568);
and U3015 (N_3015,N_2544,N_2611);
and U3016 (N_3016,N_2526,N_2765);
nor U3017 (N_3017,N_2851,N_2906);
or U3018 (N_3018,N_2678,N_2842);
and U3019 (N_3019,N_2669,N_2612);
or U3020 (N_3020,N_2539,N_2885);
or U3021 (N_3021,N_2818,N_2747);
xnor U3022 (N_3022,N_2871,N_2586);
or U3023 (N_3023,N_2618,N_2631);
or U3024 (N_3024,N_2945,N_2880);
nand U3025 (N_3025,N_2771,N_2636);
nor U3026 (N_3026,N_2960,N_2897);
nor U3027 (N_3027,N_2929,N_2783);
nand U3028 (N_3028,N_2807,N_2529);
nor U3029 (N_3029,N_2957,N_2810);
or U3030 (N_3030,N_2884,N_2781);
nand U3031 (N_3031,N_2728,N_2931);
nand U3032 (N_3032,N_2941,N_2558);
or U3033 (N_3033,N_2742,N_2853);
nand U3034 (N_3034,N_2890,N_2924);
nor U3035 (N_3035,N_2620,N_2835);
nand U3036 (N_3036,N_2646,N_2573);
nand U3037 (N_3037,N_2591,N_2830);
nor U3038 (N_3038,N_2609,N_2731);
and U3039 (N_3039,N_2702,N_2549);
nor U3040 (N_3040,N_2792,N_2854);
nor U3041 (N_3041,N_2605,N_2927);
xnor U3042 (N_3042,N_2989,N_2814);
or U3043 (N_3043,N_2600,N_2603);
and U3044 (N_3044,N_2938,N_2962);
nand U3045 (N_3045,N_2506,N_2904);
nor U3046 (N_3046,N_2643,N_2704);
nand U3047 (N_3047,N_2505,N_2541);
and U3048 (N_3048,N_2915,N_2629);
nand U3049 (N_3049,N_2576,N_2944);
and U3050 (N_3050,N_2723,N_2658);
and U3051 (N_3051,N_2614,N_2670);
nand U3052 (N_3052,N_2657,N_2640);
or U3053 (N_3053,N_2972,N_2604);
and U3054 (N_3054,N_2910,N_2946);
nor U3055 (N_3055,N_2759,N_2683);
or U3056 (N_3056,N_2812,N_2777);
and U3057 (N_3057,N_2933,N_2616);
or U3058 (N_3058,N_2594,N_2801);
and U3059 (N_3059,N_2543,N_2887);
xor U3060 (N_3060,N_2736,N_2602);
and U3061 (N_3061,N_2902,N_2766);
nand U3062 (N_3062,N_2649,N_2797);
or U3063 (N_3063,N_2552,N_2896);
and U3064 (N_3064,N_2770,N_2644);
nor U3065 (N_3065,N_2507,N_2727);
nand U3066 (N_3066,N_2825,N_2528);
or U3067 (N_3067,N_2716,N_2659);
nor U3068 (N_3068,N_2664,N_2809);
and U3069 (N_3069,N_2918,N_2863);
and U3070 (N_3070,N_2722,N_2523);
and U3071 (N_3071,N_2782,N_2580);
nor U3072 (N_3072,N_2719,N_2870);
nand U3073 (N_3073,N_2866,N_2864);
nor U3074 (N_3074,N_2905,N_2981);
nand U3075 (N_3075,N_2607,N_2881);
and U3076 (N_3076,N_2656,N_2973);
nor U3077 (N_3077,N_2715,N_2739);
xnor U3078 (N_3078,N_2508,N_2845);
nand U3079 (N_3079,N_2796,N_2527);
and U3080 (N_3080,N_2833,N_2743);
nand U3081 (N_3081,N_2628,N_2708);
nand U3082 (N_3082,N_2516,N_2651);
and U3083 (N_3083,N_2705,N_2819);
or U3084 (N_3084,N_2647,N_2699);
nand U3085 (N_3085,N_2613,N_2567);
and U3086 (N_3086,N_2548,N_2998);
and U3087 (N_3087,N_2861,N_2690);
nand U3088 (N_3088,N_2824,N_2554);
xor U3089 (N_3089,N_2556,N_2821);
nand U3090 (N_3090,N_2597,N_2872);
nor U3091 (N_3091,N_2806,N_2542);
nand U3092 (N_3092,N_2698,N_2674);
or U3093 (N_3093,N_2795,N_2688);
and U3094 (N_3094,N_2808,N_2503);
and U3095 (N_3095,N_2986,N_2898);
nor U3096 (N_3096,N_2521,N_2615);
nand U3097 (N_3097,N_2519,N_2522);
or U3098 (N_3098,N_2763,N_2961);
and U3099 (N_3099,N_2679,N_2794);
and U3100 (N_3100,N_2532,N_2930);
nand U3101 (N_3101,N_2687,N_2671);
xnor U3102 (N_3102,N_2970,N_2601);
nand U3103 (N_3103,N_2546,N_2710);
nor U3104 (N_3104,N_2847,N_2919);
and U3105 (N_3105,N_2867,N_2610);
or U3106 (N_3106,N_2949,N_2965);
or U3107 (N_3107,N_2738,N_2790);
or U3108 (N_3108,N_2672,N_2512);
and U3109 (N_3109,N_2788,N_2889);
or U3110 (N_3110,N_2950,N_2983);
nand U3111 (N_3111,N_2684,N_2958);
nand U3112 (N_3112,N_2626,N_2785);
and U3113 (N_3113,N_2622,N_2943);
nand U3114 (N_3114,N_2860,N_2693);
or U3115 (N_3115,N_2883,N_2963);
or U3116 (N_3116,N_2744,N_2892);
or U3117 (N_3117,N_2700,N_2645);
and U3118 (N_3118,N_2572,N_2838);
nand U3119 (N_3119,N_2828,N_2773);
nand U3120 (N_3120,N_2804,N_2694);
or U3121 (N_3121,N_2968,N_2648);
or U3122 (N_3122,N_2879,N_2535);
nand U3123 (N_3123,N_2514,N_2676);
and U3124 (N_3124,N_2893,N_2939);
and U3125 (N_3125,N_2767,N_2638);
or U3126 (N_3126,N_2786,N_2511);
nand U3127 (N_3127,N_2831,N_2899);
and U3128 (N_3128,N_2707,N_2578);
and U3129 (N_3129,N_2811,N_2935);
or U3130 (N_3130,N_2518,N_2746);
xnor U3131 (N_3131,N_2787,N_2752);
nand U3132 (N_3132,N_2625,N_2577);
xnor U3133 (N_3133,N_2967,N_2520);
nand U3134 (N_3134,N_2691,N_2726);
nor U3135 (N_3135,N_2730,N_2689);
xor U3136 (N_3136,N_2954,N_2560);
nor U3137 (N_3137,N_2900,N_2940);
nor U3138 (N_3138,N_2769,N_2641);
and U3139 (N_3139,N_2713,N_2799);
and U3140 (N_3140,N_2780,N_2701);
nand U3141 (N_3141,N_2741,N_2564);
nor U3142 (N_3142,N_2663,N_2757);
nor U3143 (N_3143,N_2778,N_2886);
and U3144 (N_3144,N_2942,N_2875);
nand U3145 (N_3145,N_2920,N_2551);
nand U3146 (N_3146,N_2761,N_2579);
or U3147 (N_3147,N_2895,N_2585);
or U3148 (N_3148,N_2914,N_2668);
nor U3149 (N_3149,N_2545,N_2632);
or U3150 (N_3150,N_2832,N_2922);
or U3151 (N_3151,N_2913,N_2623);
nor U3152 (N_3152,N_2907,N_2829);
and U3153 (N_3153,N_2923,N_2925);
and U3154 (N_3154,N_2729,N_2903);
nor U3155 (N_3155,N_2714,N_2955);
nor U3156 (N_3156,N_2877,N_2849);
or U3157 (N_3157,N_2846,N_2502);
xor U3158 (N_3158,N_2768,N_2841);
and U3159 (N_3159,N_2878,N_2570);
and U3160 (N_3160,N_2839,N_2985);
and U3161 (N_3161,N_2912,N_2677);
or U3162 (N_3162,N_2630,N_2608);
or U3163 (N_3163,N_2587,N_2873);
nand U3164 (N_3164,N_2917,N_2827);
and U3165 (N_3165,N_2803,N_2740);
or U3166 (N_3166,N_2979,N_2990);
and U3167 (N_3167,N_2550,N_2737);
or U3168 (N_3168,N_2667,N_2977);
and U3169 (N_3169,N_2869,N_2956);
and U3170 (N_3170,N_2772,N_2525);
nand U3171 (N_3171,N_2515,N_2660);
nor U3172 (N_3172,N_2639,N_2583);
nor U3173 (N_3173,N_2953,N_2848);
nor U3174 (N_3174,N_2711,N_2569);
or U3175 (N_3175,N_2837,N_2509);
nand U3176 (N_3176,N_2621,N_2748);
or U3177 (N_3177,N_2888,N_2988);
nand U3178 (N_3178,N_2858,N_2533);
nor U3179 (N_3179,N_2595,N_2717);
nor U3180 (N_3180,N_2593,N_2992);
nand U3181 (N_3181,N_2882,N_2978);
and U3182 (N_3182,N_2844,N_2948);
xnor U3183 (N_3183,N_2537,N_2876);
nor U3184 (N_3184,N_2592,N_2530);
or U3185 (N_3185,N_2563,N_2820);
nor U3186 (N_3186,N_2774,N_2926);
nand U3187 (N_3187,N_2642,N_2709);
nor U3188 (N_3188,N_2966,N_2800);
xnor U3189 (N_3189,N_2982,N_2559);
or U3190 (N_3190,N_2534,N_2685);
and U3191 (N_3191,N_2574,N_2637);
and U3192 (N_3192,N_2934,N_2762);
nand U3193 (N_3193,N_2724,N_2813);
or U3194 (N_3194,N_2566,N_2793);
nand U3195 (N_3195,N_2791,N_2928);
nand U3196 (N_3196,N_2857,N_2721);
and U3197 (N_3197,N_2843,N_2513);
nand U3198 (N_3198,N_2817,N_2775);
and U3199 (N_3199,N_2735,N_2712);
nand U3200 (N_3200,N_2661,N_2859);
nor U3201 (N_3201,N_2991,N_2951);
nor U3202 (N_3202,N_2894,N_2681);
nand U3203 (N_3203,N_2536,N_2802);
and U3204 (N_3204,N_2555,N_2606);
xor U3205 (N_3205,N_2703,N_2760);
nor U3206 (N_3206,N_2909,N_2680);
or U3207 (N_3207,N_2836,N_2547);
nand U3208 (N_3208,N_2974,N_2673);
nor U3209 (N_3209,N_2764,N_2538);
nand U3210 (N_3210,N_2852,N_2561);
and U3211 (N_3211,N_2500,N_2682);
or U3212 (N_3212,N_2834,N_2959);
nor U3213 (N_3213,N_2865,N_2891);
or U3214 (N_3214,N_2686,N_2718);
and U3215 (N_3215,N_2634,N_2756);
nand U3216 (N_3216,N_2696,N_2936);
nand U3217 (N_3217,N_2510,N_2755);
nand U3218 (N_3218,N_2850,N_2815);
nor U3219 (N_3219,N_2758,N_2725);
nand U3220 (N_3220,N_2650,N_2582);
and U3221 (N_3221,N_2662,N_2588);
or U3222 (N_3222,N_2652,N_2822);
nand U3223 (N_3223,N_2692,N_2531);
and U3224 (N_3224,N_2964,N_2816);
nor U3225 (N_3225,N_2504,N_2598);
or U3226 (N_3226,N_2733,N_2823);
nand U3227 (N_3227,N_2596,N_2984);
and U3228 (N_3228,N_2911,N_2557);
or U3229 (N_3229,N_2754,N_2524);
nand U3230 (N_3230,N_2995,N_2581);
or U3231 (N_3231,N_2751,N_2798);
nor U3232 (N_3232,N_2937,N_2932);
or U3233 (N_3233,N_2994,N_2666);
nand U3234 (N_3234,N_2753,N_2589);
nand U3235 (N_3235,N_2617,N_2901);
and U3236 (N_3236,N_2997,N_2868);
nor U3237 (N_3237,N_2856,N_2665);
and U3238 (N_3238,N_2805,N_2976);
nor U3239 (N_3239,N_2540,N_2826);
nor U3240 (N_3240,N_2501,N_2980);
and U3241 (N_3241,N_2750,N_2599);
nand U3242 (N_3242,N_2779,N_2720);
nand U3243 (N_3243,N_2947,N_2627);
or U3244 (N_3244,N_2916,N_2749);
and U3245 (N_3245,N_2624,N_2635);
nand U3246 (N_3246,N_2571,N_2655);
and U3247 (N_3247,N_2975,N_2874);
and U3248 (N_3248,N_2993,N_2553);
nor U3249 (N_3249,N_2745,N_2654);
nand U3250 (N_3250,N_2619,N_2823);
nand U3251 (N_3251,N_2982,N_2991);
nor U3252 (N_3252,N_2897,N_2808);
nand U3253 (N_3253,N_2885,N_2518);
nand U3254 (N_3254,N_2650,N_2898);
nand U3255 (N_3255,N_2565,N_2905);
nand U3256 (N_3256,N_2958,N_2615);
nand U3257 (N_3257,N_2897,N_2890);
nor U3258 (N_3258,N_2990,N_2552);
and U3259 (N_3259,N_2780,N_2942);
xnor U3260 (N_3260,N_2737,N_2593);
or U3261 (N_3261,N_2607,N_2619);
nor U3262 (N_3262,N_2593,N_2793);
or U3263 (N_3263,N_2509,N_2761);
nand U3264 (N_3264,N_2521,N_2735);
or U3265 (N_3265,N_2640,N_2501);
or U3266 (N_3266,N_2964,N_2927);
nor U3267 (N_3267,N_2980,N_2534);
and U3268 (N_3268,N_2743,N_2737);
xor U3269 (N_3269,N_2952,N_2638);
nand U3270 (N_3270,N_2755,N_2564);
nand U3271 (N_3271,N_2876,N_2588);
nand U3272 (N_3272,N_2694,N_2880);
nand U3273 (N_3273,N_2701,N_2974);
and U3274 (N_3274,N_2985,N_2733);
nor U3275 (N_3275,N_2986,N_2957);
nor U3276 (N_3276,N_2937,N_2529);
nor U3277 (N_3277,N_2567,N_2547);
or U3278 (N_3278,N_2523,N_2985);
and U3279 (N_3279,N_2898,N_2737);
or U3280 (N_3280,N_2955,N_2590);
nand U3281 (N_3281,N_2765,N_2706);
or U3282 (N_3282,N_2523,N_2850);
nor U3283 (N_3283,N_2669,N_2503);
nor U3284 (N_3284,N_2848,N_2882);
or U3285 (N_3285,N_2819,N_2659);
or U3286 (N_3286,N_2711,N_2696);
and U3287 (N_3287,N_2742,N_2845);
nand U3288 (N_3288,N_2890,N_2783);
nor U3289 (N_3289,N_2928,N_2786);
nor U3290 (N_3290,N_2585,N_2776);
nand U3291 (N_3291,N_2579,N_2588);
or U3292 (N_3292,N_2946,N_2914);
nor U3293 (N_3293,N_2698,N_2787);
or U3294 (N_3294,N_2700,N_2707);
nand U3295 (N_3295,N_2672,N_2959);
or U3296 (N_3296,N_2835,N_2682);
or U3297 (N_3297,N_2921,N_2586);
nand U3298 (N_3298,N_2957,N_2788);
and U3299 (N_3299,N_2538,N_2650);
nor U3300 (N_3300,N_2856,N_2615);
and U3301 (N_3301,N_2798,N_2599);
or U3302 (N_3302,N_2561,N_2777);
and U3303 (N_3303,N_2782,N_2746);
nor U3304 (N_3304,N_2565,N_2576);
and U3305 (N_3305,N_2550,N_2622);
nor U3306 (N_3306,N_2791,N_2885);
or U3307 (N_3307,N_2918,N_2650);
or U3308 (N_3308,N_2780,N_2847);
nor U3309 (N_3309,N_2789,N_2750);
and U3310 (N_3310,N_2697,N_2791);
or U3311 (N_3311,N_2607,N_2721);
nor U3312 (N_3312,N_2850,N_2714);
or U3313 (N_3313,N_2705,N_2895);
or U3314 (N_3314,N_2566,N_2613);
nor U3315 (N_3315,N_2616,N_2738);
nand U3316 (N_3316,N_2961,N_2860);
nor U3317 (N_3317,N_2767,N_2979);
and U3318 (N_3318,N_2814,N_2698);
nor U3319 (N_3319,N_2662,N_2623);
or U3320 (N_3320,N_2722,N_2774);
nor U3321 (N_3321,N_2770,N_2607);
nor U3322 (N_3322,N_2614,N_2831);
nand U3323 (N_3323,N_2798,N_2870);
or U3324 (N_3324,N_2950,N_2649);
nor U3325 (N_3325,N_2559,N_2890);
and U3326 (N_3326,N_2559,N_2977);
or U3327 (N_3327,N_2826,N_2642);
xor U3328 (N_3328,N_2719,N_2688);
nor U3329 (N_3329,N_2735,N_2899);
nor U3330 (N_3330,N_2694,N_2647);
nor U3331 (N_3331,N_2852,N_2722);
and U3332 (N_3332,N_2833,N_2685);
nor U3333 (N_3333,N_2945,N_2690);
and U3334 (N_3334,N_2747,N_2521);
and U3335 (N_3335,N_2662,N_2580);
and U3336 (N_3336,N_2728,N_2505);
nand U3337 (N_3337,N_2752,N_2538);
nor U3338 (N_3338,N_2774,N_2959);
and U3339 (N_3339,N_2823,N_2955);
and U3340 (N_3340,N_2739,N_2534);
nand U3341 (N_3341,N_2996,N_2731);
nor U3342 (N_3342,N_2536,N_2789);
nor U3343 (N_3343,N_2539,N_2942);
and U3344 (N_3344,N_2747,N_2745);
nor U3345 (N_3345,N_2781,N_2740);
and U3346 (N_3346,N_2531,N_2844);
or U3347 (N_3347,N_2630,N_2740);
nor U3348 (N_3348,N_2509,N_2543);
and U3349 (N_3349,N_2691,N_2676);
nor U3350 (N_3350,N_2778,N_2619);
nand U3351 (N_3351,N_2951,N_2937);
or U3352 (N_3352,N_2987,N_2712);
or U3353 (N_3353,N_2979,N_2894);
nor U3354 (N_3354,N_2896,N_2766);
xnor U3355 (N_3355,N_2541,N_2819);
and U3356 (N_3356,N_2731,N_2747);
nor U3357 (N_3357,N_2855,N_2607);
nand U3358 (N_3358,N_2921,N_2762);
or U3359 (N_3359,N_2908,N_2611);
nand U3360 (N_3360,N_2765,N_2582);
or U3361 (N_3361,N_2771,N_2954);
or U3362 (N_3362,N_2661,N_2541);
nand U3363 (N_3363,N_2816,N_2777);
nor U3364 (N_3364,N_2789,N_2870);
nor U3365 (N_3365,N_2851,N_2585);
nand U3366 (N_3366,N_2594,N_2658);
or U3367 (N_3367,N_2680,N_2688);
nand U3368 (N_3368,N_2546,N_2851);
nand U3369 (N_3369,N_2756,N_2977);
or U3370 (N_3370,N_2847,N_2835);
and U3371 (N_3371,N_2978,N_2617);
nand U3372 (N_3372,N_2771,N_2735);
or U3373 (N_3373,N_2539,N_2774);
and U3374 (N_3374,N_2535,N_2952);
nor U3375 (N_3375,N_2528,N_2558);
nor U3376 (N_3376,N_2985,N_2730);
and U3377 (N_3377,N_2521,N_2763);
or U3378 (N_3378,N_2676,N_2824);
nand U3379 (N_3379,N_2689,N_2642);
or U3380 (N_3380,N_2666,N_2553);
nor U3381 (N_3381,N_2615,N_2845);
and U3382 (N_3382,N_2711,N_2926);
or U3383 (N_3383,N_2919,N_2833);
nor U3384 (N_3384,N_2620,N_2630);
and U3385 (N_3385,N_2753,N_2911);
or U3386 (N_3386,N_2884,N_2710);
nor U3387 (N_3387,N_2686,N_2853);
xor U3388 (N_3388,N_2856,N_2502);
or U3389 (N_3389,N_2933,N_2736);
and U3390 (N_3390,N_2806,N_2931);
and U3391 (N_3391,N_2974,N_2716);
nor U3392 (N_3392,N_2614,N_2777);
or U3393 (N_3393,N_2943,N_2984);
nand U3394 (N_3394,N_2700,N_2607);
nor U3395 (N_3395,N_2702,N_2821);
and U3396 (N_3396,N_2804,N_2842);
nand U3397 (N_3397,N_2596,N_2674);
and U3398 (N_3398,N_2753,N_2676);
nand U3399 (N_3399,N_2833,N_2925);
and U3400 (N_3400,N_2605,N_2764);
nand U3401 (N_3401,N_2909,N_2858);
nand U3402 (N_3402,N_2896,N_2720);
nor U3403 (N_3403,N_2775,N_2680);
nand U3404 (N_3404,N_2639,N_2693);
and U3405 (N_3405,N_2791,N_2507);
or U3406 (N_3406,N_2879,N_2725);
or U3407 (N_3407,N_2771,N_2935);
and U3408 (N_3408,N_2789,N_2801);
nand U3409 (N_3409,N_2750,N_2972);
or U3410 (N_3410,N_2643,N_2604);
and U3411 (N_3411,N_2772,N_2944);
nor U3412 (N_3412,N_2582,N_2842);
or U3413 (N_3413,N_2909,N_2609);
and U3414 (N_3414,N_2694,N_2763);
and U3415 (N_3415,N_2854,N_2639);
nand U3416 (N_3416,N_2637,N_2772);
nand U3417 (N_3417,N_2728,N_2972);
nor U3418 (N_3418,N_2680,N_2641);
xnor U3419 (N_3419,N_2976,N_2913);
and U3420 (N_3420,N_2606,N_2619);
nand U3421 (N_3421,N_2756,N_2972);
or U3422 (N_3422,N_2678,N_2865);
nor U3423 (N_3423,N_2784,N_2891);
nand U3424 (N_3424,N_2637,N_2805);
and U3425 (N_3425,N_2810,N_2854);
and U3426 (N_3426,N_2535,N_2523);
or U3427 (N_3427,N_2639,N_2757);
nor U3428 (N_3428,N_2913,N_2636);
and U3429 (N_3429,N_2831,N_2890);
nand U3430 (N_3430,N_2545,N_2744);
or U3431 (N_3431,N_2551,N_2931);
or U3432 (N_3432,N_2617,N_2837);
nor U3433 (N_3433,N_2515,N_2632);
nor U3434 (N_3434,N_2971,N_2639);
nand U3435 (N_3435,N_2926,N_2702);
nand U3436 (N_3436,N_2842,N_2676);
nand U3437 (N_3437,N_2975,N_2959);
and U3438 (N_3438,N_2701,N_2805);
or U3439 (N_3439,N_2677,N_2540);
and U3440 (N_3440,N_2651,N_2588);
nand U3441 (N_3441,N_2694,N_2833);
nor U3442 (N_3442,N_2559,N_2967);
and U3443 (N_3443,N_2801,N_2764);
nor U3444 (N_3444,N_2634,N_2658);
nand U3445 (N_3445,N_2565,N_2935);
or U3446 (N_3446,N_2631,N_2520);
or U3447 (N_3447,N_2745,N_2934);
or U3448 (N_3448,N_2719,N_2935);
and U3449 (N_3449,N_2803,N_2822);
nor U3450 (N_3450,N_2886,N_2690);
or U3451 (N_3451,N_2698,N_2762);
nand U3452 (N_3452,N_2742,N_2680);
and U3453 (N_3453,N_2577,N_2883);
or U3454 (N_3454,N_2742,N_2624);
nor U3455 (N_3455,N_2912,N_2527);
and U3456 (N_3456,N_2910,N_2935);
nor U3457 (N_3457,N_2572,N_2912);
or U3458 (N_3458,N_2710,N_2591);
and U3459 (N_3459,N_2844,N_2797);
nand U3460 (N_3460,N_2811,N_2784);
or U3461 (N_3461,N_2763,N_2689);
nor U3462 (N_3462,N_2979,N_2754);
and U3463 (N_3463,N_2678,N_2539);
or U3464 (N_3464,N_2885,N_2838);
xnor U3465 (N_3465,N_2681,N_2880);
nand U3466 (N_3466,N_2560,N_2784);
xor U3467 (N_3467,N_2799,N_2608);
nand U3468 (N_3468,N_2651,N_2523);
and U3469 (N_3469,N_2946,N_2547);
or U3470 (N_3470,N_2524,N_2523);
and U3471 (N_3471,N_2579,N_2529);
nand U3472 (N_3472,N_2964,N_2750);
nand U3473 (N_3473,N_2587,N_2743);
nand U3474 (N_3474,N_2557,N_2540);
nand U3475 (N_3475,N_2882,N_2582);
nor U3476 (N_3476,N_2915,N_2841);
nor U3477 (N_3477,N_2731,N_2755);
nor U3478 (N_3478,N_2591,N_2657);
or U3479 (N_3479,N_2866,N_2945);
nand U3480 (N_3480,N_2964,N_2701);
nand U3481 (N_3481,N_2700,N_2926);
or U3482 (N_3482,N_2528,N_2712);
or U3483 (N_3483,N_2874,N_2888);
or U3484 (N_3484,N_2657,N_2967);
and U3485 (N_3485,N_2809,N_2751);
nand U3486 (N_3486,N_2742,N_2695);
or U3487 (N_3487,N_2679,N_2641);
nor U3488 (N_3488,N_2583,N_2935);
and U3489 (N_3489,N_2633,N_2735);
nor U3490 (N_3490,N_2852,N_2617);
and U3491 (N_3491,N_2779,N_2610);
nor U3492 (N_3492,N_2987,N_2704);
nand U3493 (N_3493,N_2864,N_2659);
nor U3494 (N_3494,N_2827,N_2779);
and U3495 (N_3495,N_2682,N_2856);
and U3496 (N_3496,N_2945,N_2693);
nand U3497 (N_3497,N_2666,N_2984);
and U3498 (N_3498,N_2554,N_2976);
or U3499 (N_3499,N_2694,N_2735);
or U3500 (N_3500,N_3260,N_3417);
and U3501 (N_3501,N_3169,N_3450);
nand U3502 (N_3502,N_3423,N_3144);
or U3503 (N_3503,N_3394,N_3140);
or U3504 (N_3504,N_3411,N_3383);
nand U3505 (N_3505,N_3181,N_3385);
or U3506 (N_3506,N_3465,N_3063);
nand U3507 (N_3507,N_3053,N_3022);
nor U3508 (N_3508,N_3012,N_3173);
nor U3509 (N_3509,N_3490,N_3284);
nand U3510 (N_3510,N_3250,N_3248);
and U3511 (N_3511,N_3076,N_3015);
nor U3512 (N_3512,N_3066,N_3337);
and U3513 (N_3513,N_3048,N_3007);
and U3514 (N_3514,N_3440,N_3480);
nand U3515 (N_3515,N_3200,N_3094);
or U3516 (N_3516,N_3213,N_3400);
xor U3517 (N_3517,N_3230,N_3239);
nand U3518 (N_3518,N_3122,N_3183);
nor U3519 (N_3519,N_3280,N_3439);
xor U3520 (N_3520,N_3001,N_3038);
and U3521 (N_3521,N_3121,N_3023);
nand U3522 (N_3522,N_3311,N_3244);
nand U3523 (N_3523,N_3072,N_3095);
nor U3524 (N_3524,N_3231,N_3389);
or U3525 (N_3525,N_3410,N_3170);
or U3526 (N_3526,N_3387,N_3356);
nand U3527 (N_3527,N_3426,N_3415);
or U3528 (N_3528,N_3224,N_3442);
nor U3529 (N_3529,N_3055,N_3069);
or U3530 (N_3530,N_3264,N_3358);
and U3531 (N_3531,N_3204,N_3029);
or U3532 (N_3532,N_3236,N_3077);
nand U3533 (N_3533,N_3452,N_3273);
nor U3534 (N_3534,N_3042,N_3335);
and U3535 (N_3535,N_3475,N_3134);
or U3536 (N_3536,N_3303,N_3176);
nand U3537 (N_3537,N_3379,N_3263);
or U3538 (N_3538,N_3314,N_3476);
nand U3539 (N_3539,N_3296,N_3292);
nor U3540 (N_3540,N_3243,N_3018);
nor U3541 (N_3541,N_3371,N_3110);
nand U3542 (N_3542,N_3154,N_3276);
or U3543 (N_3543,N_3354,N_3348);
xnor U3544 (N_3544,N_3179,N_3395);
or U3545 (N_3545,N_3216,N_3499);
xnor U3546 (N_3546,N_3207,N_3002);
nor U3547 (N_3547,N_3044,N_3454);
and U3548 (N_3548,N_3482,N_3028);
and U3549 (N_3549,N_3218,N_3267);
nor U3550 (N_3550,N_3255,N_3211);
xor U3551 (N_3551,N_3148,N_3494);
nor U3552 (N_3552,N_3266,N_3268);
nor U3553 (N_3553,N_3471,N_3115);
or U3554 (N_3554,N_3363,N_3135);
nor U3555 (N_3555,N_3413,N_3486);
and U3556 (N_3556,N_3232,N_3295);
and U3557 (N_3557,N_3103,N_3456);
nand U3558 (N_3558,N_3437,N_3330);
nor U3559 (N_3559,N_3381,N_3393);
nand U3560 (N_3560,N_3131,N_3418);
and U3561 (N_3561,N_3234,N_3424);
nor U3562 (N_3562,N_3191,N_3489);
nor U3563 (N_3563,N_3453,N_3013);
nor U3564 (N_3564,N_3441,N_3136);
nand U3565 (N_3565,N_3065,N_3321);
nand U3566 (N_3566,N_3229,N_3287);
and U3567 (N_3567,N_3014,N_3118);
or U3568 (N_3568,N_3138,N_3034);
and U3569 (N_3569,N_3327,N_3345);
or U3570 (N_3570,N_3195,N_3035);
or U3571 (N_3571,N_3214,N_3443);
nor U3572 (N_3572,N_3074,N_3225);
or U3573 (N_3573,N_3297,N_3388);
and U3574 (N_3574,N_3332,N_3343);
or U3575 (N_3575,N_3054,N_3305);
nand U3576 (N_3576,N_3275,N_3087);
nand U3577 (N_3577,N_3483,N_3472);
and U3578 (N_3578,N_3198,N_3317);
nand U3579 (N_3579,N_3081,N_3460);
nor U3580 (N_3580,N_3091,N_3033);
or U3581 (N_3581,N_3376,N_3261);
xor U3582 (N_3582,N_3329,N_3270);
and U3583 (N_3583,N_3272,N_3090);
nor U3584 (N_3584,N_3206,N_3127);
nand U3585 (N_3585,N_3399,N_3036);
or U3586 (N_3586,N_3432,N_3257);
nor U3587 (N_3587,N_3215,N_3402);
nand U3588 (N_3588,N_3162,N_3451);
and U3589 (N_3589,N_3386,N_3006);
nor U3590 (N_3590,N_3166,N_3313);
nand U3591 (N_3591,N_3347,N_3228);
nor U3592 (N_3592,N_3188,N_3219);
and U3593 (N_3593,N_3120,N_3189);
or U3594 (N_3594,N_3227,N_3333);
xnor U3595 (N_3595,N_3368,N_3458);
or U3596 (N_3596,N_3378,N_3068);
nand U3597 (N_3597,N_3496,N_3338);
nor U3598 (N_3598,N_3274,N_3146);
or U3599 (N_3599,N_3320,N_3186);
or U3600 (N_3600,N_3051,N_3283);
nand U3601 (N_3601,N_3220,N_3449);
or U3602 (N_3602,N_3010,N_3059);
nand U3603 (N_3603,N_3308,N_3431);
or U3604 (N_3604,N_3180,N_3205);
and U3605 (N_3605,N_3123,N_3380);
nor U3606 (N_3606,N_3089,N_3253);
and U3607 (N_3607,N_3047,N_3056);
or U3608 (N_3608,N_3491,N_3160);
or U3609 (N_3609,N_3102,N_3252);
and U3610 (N_3610,N_3011,N_3428);
and U3611 (N_3611,N_3375,N_3184);
or U3612 (N_3612,N_3340,N_3299);
nand U3613 (N_3613,N_3174,N_3377);
and U3614 (N_3614,N_3039,N_3132);
nand U3615 (N_3615,N_3269,N_3407);
and U3616 (N_3616,N_3082,N_3294);
or U3617 (N_3617,N_3382,N_3466);
nand U3618 (N_3618,N_3290,N_3182);
nand U3619 (N_3619,N_3446,N_3457);
nand U3620 (N_3620,N_3390,N_3488);
nor U3621 (N_3621,N_3073,N_3238);
or U3622 (N_3622,N_3414,N_3366);
or U3623 (N_3623,N_3030,N_3492);
nor U3624 (N_3624,N_3125,N_3331);
and U3625 (N_3625,N_3481,N_3425);
nand U3626 (N_3626,N_3282,N_3126);
nor U3627 (N_3627,N_3097,N_3326);
or U3628 (N_3628,N_3445,N_3062);
nand U3629 (N_3629,N_3279,N_3406);
xnor U3630 (N_3630,N_3470,N_3298);
or U3631 (N_3631,N_3421,N_3222);
nor U3632 (N_3632,N_3459,N_3412);
nand U3633 (N_3633,N_3083,N_3108);
nand U3634 (N_3634,N_3350,N_3075);
and U3635 (N_3635,N_3467,N_3278);
and U3636 (N_3636,N_3060,N_3000);
nand U3637 (N_3637,N_3133,N_3474);
nand U3638 (N_3638,N_3145,N_3004);
nor U3639 (N_3639,N_3455,N_3142);
or U3640 (N_3640,N_3397,N_3361);
nand U3641 (N_3641,N_3288,N_3009);
nand U3642 (N_3642,N_3405,N_3237);
and U3643 (N_3643,N_3319,N_3016);
and U3644 (N_3644,N_3346,N_3433);
xnor U3645 (N_3645,N_3316,N_3367);
and U3646 (N_3646,N_3365,N_3178);
or U3647 (N_3647,N_3357,N_3438);
xor U3648 (N_3648,N_3372,N_3084);
nand U3649 (N_3649,N_3334,N_3289);
nor U3650 (N_3650,N_3223,N_3344);
and U3651 (N_3651,N_3301,N_3221);
nor U3652 (N_3652,N_3444,N_3351);
xnor U3653 (N_3653,N_3151,N_3141);
nor U3654 (N_3654,N_3109,N_3139);
and U3655 (N_3655,N_3107,N_3265);
nand U3656 (N_3656,N_3271,N_3309);
or U3657 (N_3657,N_3155,N_3208);
and U3658 (N_3658,N_3281,N_3398);
or U3659 (N_3659,N_3190,N_3040);
xnor U3660 (N_3660,N_3307,N_3461);
nor U3661 (N_3661,N_3067,N_3021);
and U3662 (N_3662,N_3106,N_3088);
and U3663 (N_3663,N_3360,N_3177);
nor U3664 (N_3664,N_3027,N_3403);
and U3665 (N_3665,N_3262,N_3247);
nand U3666 (N_3666,N_3008,N_3468);
nor U3667 (N_3667,N_3165,N_3434);
xor U3668 (N_3668,N_3187,N_3032);
nand U3669 (N_3669,N_3369,N_3005);
or U3670 (N_3670,N_3064,N_3105);
and U3671 (N_3671,N_3037,N_3167);
and U3672 (N_3672,N_3342,N_3241);
nor U3673 (N_3673,N_3302,N_3242);
nor U3674 (N_3674,N_3098,N_3341);
and U3675 (N_3675,N_3485,N_3355);
nor U3676 (N_3676,N_3349,N_3384);
xor U3677 (N_3677,N_3196,N_3058);
nor U3678 (N_3678,N_3312,N_3277);
or U3679 (N_3679,N_3240,N_3202);
or U3680 (N_3680,N_3130,N_3199);
or U3681 (N_3681,N_3479,N_3464);
nand U3682 (N_3682,N_3112,N_3153);
or U3683 (N_3683,N_3128,N_3306);
or U3684 (N_3684,N_3099,N_3364);
and U3685 (N_3685,N_3093,N_3448);
nand U3686 (N_3686,N_3259,N_3129);
or U3687 (N_3687,N_3353,N_3324);
nand U3688 (N_3688,N_3404,N_3019);
and U3689 (N_3689,N_3429,N_3246);
and U3690 (N_3690,N_3416,N_3463);
and U3691 (N_3691,N_3249,N_3256);
or U3692 (N_3692,N_3025,N_3373);
nand U3693 (N_3693,N_3408,N_3370);
or U3694 (N_3694,N_3100,N_3079);
nand U3695 (N_3695,N_3003,N_3043);
or U3696 (N_3696,N_3147,N_3210);
nor U3697 (N_3697,N_3172,N_3116);
nor U3698 (N_3698,N_3310,N_3286);
and U3699 (N_3699,N_3285,N_3447);
nor U3700 (N_3700,N_3396,N_3362);
and U3701 (N_3701,N_3427,N_3104);
nand U3702 (N_3702,N_3150,N_3031);
and U3703 (N_3703,N_3462,N_3080);
or U3704 (N_3704,N_3113,N_3436);
or U3705 (N_3705,N_3124,N_3085);
nand U3706 (N_3706,N_3304,N_3478);
and U3707 (N_3707,N_3185,N_3157);
nor U3708 (N_3708,N_3175,N_3137);
nand U3709 (N_3709,N_3114,N_3339);
nand U3710 (N_3710,N_3020,N_3487);
nor U3711 (N_3711,N_3493,N_3469);
nor U3712 (N_3712,N_3092,N_3057);
xor U3713 (N_3713,N_3096,N_3171);
and U3714 (N_3714,N_3070,N_3061);
and U3715 (N_3715,N_3049,N_3209);
nand U3716 (N_3716,N_3024,N_3315);
and U3717 (N_3717,N_3193,N_3473);
nand U3718 (N_3718,N_3291,N_3158);
or U3719 (N_3719,N_3235,N_3119);
nor U3720 (N_3720,N_3194,N_3226);
nor U3721 (N_3721,N_3325,N_3420);
and U3722 (N_3722,N_3159,N_3071);
and U3723 (N_3723,N_3201,N_3101);
nor U3724 (N_3724,N_3156,N_3328);
nor U3725 (N_3725,N_3323,N_3117);
or U3726 (N_3726,N_3197,N_3391);
and U3727 (N_3727,N_3017,N_3258);
and U3728 (N_3728,N_3168,N_3161);
and U3729 (N_3729,N_3245,N_3322);
nor U3730 (N_3730,N_3293,N_3435);
nand U3731 (N_3731,N_3318,N_3352);
nor U3732 (N_3732,N_3422,N_3374);
or U3733 (N_3733,N_3233,N_3484);
and U3734 (N_3734,N_3041,N_3149);
nand U3735 (N_3735,N_3359,N_3143);
xor U3736 (N_3736,N_3217,N_3050);
nor U3737 (N_3737,N_3212,N_3300);
nor U3738 (N_3738,N_3045,N_3409);
xnor U3739 (N_3739,N_3392,N_3497);
nor U3740 (N_3740,N_3336,N_3046);
or U3741 (N_3741,N_3477,N_3495);
nor U3742 (N_3742,N_3419,N_3192);
nor U3743 (N_3743,N_3111,N_3430);
and U3744 (N_3744,N_3052,N_3203);
nor U3745 (N_3745,N_3251,N_3401);
nor U3746 (N_3746,N_3086,N_3026);
nand U3747 (N_3747,N_3152,N_3163);
and U3748 (N_3748,N_3498,N_3164);
and U3749 (N_3749,N_3078,N_3254);
nor U3750 (N_3750,N_3033,N_3253);
nor U3751 (N_3751,N_3335,N_3344);
or U3752 (N_3752,N_3047,N_3416);
nor U3753 (N_3753,N_3299,N_3398);
and U3754 (N_3754,N_3382,N_3069);
and U3755 (N_3755,N_3100,N_3432);
nand U3756 (N_3756,N_3491,N_3066);
nand U3757 (N_3757,N_3192,N_3251);
and U3758 (N_3758,N_3473,N_3499);
nor U3759 (N_3759,N_3489,N_3399);
nand U3760 (N_3760,N_3228,N_3492);
or U3761 (N_3761,N_3225,N_3446);
nor U3762 (N_3762,N_3467,N_3242);
nand U3763 (N_3763,N_3431,N_3015);
nand U3764 (N_3764,N_3127,N_3235);
nor U3765 (N_3765,N_3273,N_3071);
nand U3766 (N_3766,N_3408,N_3410);
nand U3767 (N_3767,N_3153,N_3150);
nand U3768 (N_3768,N_3001,N_3168);
or U3769 (N_3769,N_3078,N_3082);
or U3770 (N_3770,N_3423,N_3461);
nor U3771 (N_3771,N_3295,N_3328);
nor U3772 (N_3772,N_3479,N_3174);
nor U3773 (N_3773,N_3270,N_3493);
nand U3774 (N_3774,N_3198,N_3473);
or U3775 (N_3775,N_3214,N_3361);
or U3776 (N_3776,N_3117,N_3456);
and U3777 (N_3777,N_3269,N_3014);
nor U3778 (N_3778,N_3193,N_3135);
nor U3779 (N_3779,N_3099,N_3464);
and U3780 (N_3780,N_3263,N_3465);
nand U3781 (N_3781,N_3077,N_3189);
nand U3782 (N_3782,N_3078,N_3471);
and U3783 (N_3783,N_3376,N_3416);
nand U3784 (N_3784,N_3043,N_3397);
nor U3785 (N_3785,N_3034,N_3388);
and U3786 (N_3786,N_3212,N_3221);
nor U3787 (N_3787,N_3063,N_3276);
or U3788 (N_3788,N_3479,N_3444);
or U3789 (N_3789,N_3458,N_3275);
or U3790 (N_3790,N_3309,N_3264);
and U3791 (N_3791,N_3117,N_3311);
nand U3792 (N_3792,N_3267,N_3113);
nand U3793 (N_3793,N_3343,N_3101);
nor U3794 (N_3794,N_3009,N_3469);
nand U3795 (N_3795,N_3488,N_3340);
and U3796 (N_3796,N_3283,N_3255);
nor U3797 (N_3797,N_3039,N_3394);
and U3798 (N_3798,N_3436,N_3498);
or U3799 (N_3799,N_3276,N_3459);
nor U3800 (N_3800,N_3125,N_3487);
nand U3801 (N_3801,N_3478,N_3198);
and U3802 (N_3802,N_3299,N_3203);
or U3803 (N_3803,N_3445,N_3125);
and U3804 (N_3804,N_3178,N_3414);
nand U3805 (N_3805,N_3468,N_3062);
or U3806 (N_3806,N_3459,N_3333);
nand U3807 (N_3807,N_3406,N_3493);
nand U3808 (N_3808,N_3286,N_3285);
and U3809 (N_3809,N_3323,N_3447);
nand U3810 (N_3810,N_3122,N_3416);
and U3811 (N_3811,N_3019,N_3136);
nand U3812 (N_3812,N_3226,N_3409);
or U3813 (N_3813,N_3411,N_3106);
nand U3814 (N_3814,N_3302,N_3121);
nor U3815 (N_3815,N_3339,N_3295);
and U3816 (N_3816,N_3008,N_3417);
nand U3817 (N_3817,N_3399,N_3245);
nand U3818 (N_3818,N_3199,N_3177);
and U3819 (N_3819,N_3453,N_3470);
and U3820 (N_3820,N_3032,N_3099);
or U3821 (N_3821,N_3032,N_3393);
xor U3822 (N_3822,N_3190,N_3478);
or U3823 (N_3823,N_3404,N_3162);
or U3824 (N_3824,N_3318,N_3180);
nor U3825 (N_3825,N_3416,N_3444);
and U3826 (N_3826,N_3293,N_3129);
or U3827 (N_3827,N_3397,N_3150);
and U3828 (N_3828,N_3079,N_3039);
nor U3829 (N_3829,N_3469,N_3301);
or U3830 (N_3830,N_3326,N_3436);
nand U3831 (N_3831,N_3176,N_3137);
and U3832 (N_3832,N_3413,N_3339);
nand U3833 (N_3833,N_3427,N_3341);
nand U3834 (N_3834,N_3371,N_3069);
nand U3835 (N_3835,N_3063,N_3105);
nor U3836 (N_3836,N_3151,N_3244);
nor U3837 (N_3837,N_3132,N_3468);
nor U3838 (N_3838,N_3493,N_3183);
nor U3839 (N_3839,N_3379,N_3443);
nor U3840 (N_3840,N_3416,N_3477);
and U3841 (N_3841,N_3396,N_3203);
nor U3842 (N_3842,N_3270,N_3196);
or U3843 (N_3843,N_3171,N_3271);
nand U3844 (N_3844,N_3019,N_3393);
and U3845 (N_3845,N_3112,N_3240);
nand U3846 (N_3846,N_3270,N_3220);
nand U3847 (N_3847,N_3175,N_3307);
and U3848 (N_3848,N_3018,N_3006);
nand U3849 (N_3849,N_3052,N_3475);
nand U3850 (N_3850,N_3478,N_3431);
and U3851 (N_3851,N_3424,N_3143);
and U3852 (N_3852,N_3301,N_3349);
and U3853 (N_3853,N_3305,N_3380);
or U3854 (N_3854,N_3162,N_3322);
and U3855 (N_3855,N_3171,N_3005);
nand U3856 (N_3856,N_3073,N_3050);
or U3857 (N_3857,N_3363,N_3231);
or U3858 (N_3858,N_3235,N_3360);
or U3859 (N_3859,N_3015,N_3405);
or U3860 (N_3860,N_3031,N_3073);
and U3861 (N_3861,N_3161,N_3116);
or U3862 (N_3862,N_3279,N_3060);
and U3863 (N_3863,N_3070,N_3138);
nor U3864 (N_3864,N_3345,N_3388);
and U3865 (N_3865,N_3471,N_3335);
and U3866 (N_3866,N_3324,N_3200);
nor U3867 (N_3867,N_3372,N_3154);
or U3868 (N_3868,N_3104,N_3399);
nor U3869 (N_3869,N_3161,N_3211);
and U3870 (N_3870,N_3191,N_3465);
nor U3871 (N_3871,N_3362,N_3424);
nand U3872 (N_3872,N_3253,N_3430);
nand U3873 (N_3873,N_3498,N_3221);
or U3874 (N_3874,N_3097,N_3416);
or U3875 (N_3875,N_3212,N_3100);
nand U3876 (N_3876,N_3107,N_3344);
nor U3877 (N_3877,N_3138,N_3093);
or U3878 (N_3878,N_3157,N_3054);
and U3879 (N_3879,N_3027,N_3397);
or U3880 (N_3880,N_3429,N_3008);
nand U3881 (N_3881,N_3495,N_3370);
nor U3882 (N_3882,N_3033,N_3007);
nand U3883 (N_3883,N_3186,N_3250);
nor U3884 (N_3884,N_3402,N_3459);
nand U3885 (N_3885,N_3156,N_3361);
nor U3886 (N_3886,N_3050,N_3392);
or U3887 (N_3887,N_3325,N_3005);
nor U3888 (N_3888,N_3102,N_3165);
and U3889 (N_3889,N_3458,N_3118);
xor U3890 (N_3890,N_3373,N_3077);
or U3891 (N_3891,N_3073,N_3115);
nand U3892 (N_3892,N_3425,N_3477);
nand U3893 (N_3893,N_3148,N_3365);
and U3894 (N_3894,N_3040,N_3067);
nand U3895 (N_3895,N_3097,N_3062);
or U3896 (N_3896,N_3228,N_3270);
nand U3897 (N_3897,N_3114,N_3006);
nand U3898 (N_3898,N_3228,N_3313);
xnor U3899 (N_3899,N_3082,N_3243);
or U3900 (N_3900,N_3062,N_3106);
or U3901 (N_3901,N_3311,N_3114);
or U3902 (N_3902,N_3050,N_3440);
nand U3903 (N_3903,N_3173,N_3279);
nor U3904 (N_3904,N_3259,N_3176);
nand U3905 (N_3905,N_3103,N_3489);
and U3906 (N_3906,N_3303,N_3247);
nand U3907 (N_3907,N_3137,N_3282);
nand U3908 (N_3908,N_3016,N_3403);
nand U3909 (N_3909,N_3071,N_3414);
and U3910 (N_3910,N_3323,N_3494);
and U3911 (N_3911,N_3321,N_3290);
and U3912 (N_3912,N_3421,N_3311);
and U3913 (N_3913,N_3091,N_3467);
nor U3914 (N_3914,N_3300,N_3179);
and U3915 (N_3915,N_3015,N_3394);
or U3916 (N_3916,N_3035,N_3022);
and U3917 (N_3917,N_3326,N_3049);
nor U3918 (N_3918,N_3181,N_3375);
or U3919 (N_3919,N_3167,N_3041);
or U3920 (N_3920,N_3291,N_3317);
nand U3921 (N_3921,N_3374,N_3045);
or U3922 (N_3922,N_3307,N_3073);
nor U3923 (N_3923,N_3010,N_3055);
nand U3924 (N_3924,N_3226,N_3292);
or U3925 (N_3925,N_3054,N_3165);
and U3926 (N_3926,N_3305,N_3484);
or U3927 (N_3927,N_3254,N_3398);
or U3928 (N_3928,N_3470,N_3025);
and U3929 (N_3929,N_3154,N_3164);
nand U3930 (N_3930,N_3190,N_3417);
or U3931 (N_3931,N_3383,N_3448);
nor U3932 (N_3932,N_3089,N_3392);
nor U3933 (N_3933,N_3260,N_3416);
xor U3934 (N_3934,N_3383,N_3254);
and U3935 (N_3935,N_3036,N_3233);
nor U3936 (N_3936,N_3056,N_3439);
nor U3937 (N_3937,N_3307,N_3198);
or U3938 (N_3938,N_3118,N_3287);
or U3939 (N_3939,N_3264,N_3069);
nor U3940 (N_3940,N_3067,N_3228);
or U3941 (N_3941,N_3287,N_3452);
or U3942 (N_3942,N_3026,N_3210);
and U3943 (N_3943,N_3402,N_3292);
or U3944 (N_3944,N_3371,N_3467);
nand U3945 (N_3945,N_3201,N_3348);
xnor U3946 (N_3946,N_3441,N_3225);
or U3947 (N_3947,N_3311,N_3068);
nor U3948 (N_3948,N_3393,N_3391);
nor U3949 (N_3949,N_3347,N_3353);
and U3950 (N_3950,N_3282,N_3142);
nand U3951 (N_3951,N_3394,N_3049);
nor U3952 (N_3952,N_3218,N_3170);
nor U3953 (N_3953,N_3104,N_3430);
nand U3954 (N_3954,N_3052,N_3303);
and U3955 (N_3955,N_3220,N_3341);
nor U3956 (N_3956,N_3075,N_3184);
nor U3957 (N_3957,N_3294,N_3415);
nand U3958 (N_3958,N_3206,N_3113);
nand U3959 (N_3959,N_3291,N_3280);
nand U3960 (N_3960,N_3456,N_3160);
and U3961 (N_3961,N_3298,N_3106);
nor U3962 (N_3962,N_3454,N_3243);
or U3963 (N_3963,N_3089,N_3091);
nand U3964 (N_3964,N_3312,N_3060);
nand U3965 (N_3965,N_3028,N_3481);
nor U3966 (N_3966,N_3392,N_3036);
nor U3967 (N_3967,N_3150,N_3243);
nor U3968 (N_3968,N_3102,N_3440);
and U3969 (N_3969,N_3288,N_3266);
or U3970 (N_3970,N_3164,N_3427);
and U3971 (N_3971,N_3190,N_3471);
or U3972 (N_3972,N_3284,N_3240);
and U3973 (N_3973,N_3147,N_3415);
nor U3974 (N_3974,N_3328,N_3249);
and U3975 (N_3975,N_3446,N_3409);
or U3976 (N_3976,N_3081,N_3126);
nor U3977 (N_3977,N_3267,N_3252);
nand U3978 (N_3978,N_3344,N_3360);
or U3979 (N_3979,N_3001,N_3421);
nor U3980 (N_3980,N_3307,N_3471);
nor U3981 (N_3981,N_3144,N_3136);
nand U3982 (N_3982,N_3091,N_3103);
nand U3983 (N_3983,N_3233,N_3144);
and U3984 (N_3984,N_3147,N_3219);
nor U3985 (N_3985,N_3343,N_3346);
and U3986 (N_3986,N_3135,N_3128);
xor U3987 (N_3987,N_3400,N_3477);
xnor U3988 (N_3988,N_3331,N_3092);
and U3989 (N_3989,N_3464,N_3367);
or U3990 (N_3990,N_3466,N_3388);
and U3991 (N_3991,N_3046,N_3437);
xnor U3992 (N_3992,N_3137,N_3395);
nand U3993 (N_3993,N_3212,N_3408);
nand U3994 (N_3994,N_3138,N_3030);
and U3995 (N_3995,N_3066,N_3247);
or U3996 (N_3996,N_3236,N_3464);
or U3997 (N_3997,N_3310,N_3483);
nand U3998 (N_3998,N_3111,N_3419);
nand U3999 (N_3999,N_3151,N_3296);
nand U4000 (N_4000,N_3639,N_3794);
or U4001 (N_4001,N_3961,N_3737);
nand U4002 (N_4002,N_3753,N_3568);
and U4003 (N_4003,N_3971,N_3975);
or U4004 (N_4004,N_3716,N_3887);
or U4005 (N_4005,N_3651,N_3670);
and U4006 (N_4006,N_3710,N_3813);
nor U4007 (N_4007,N_3880,N_3997);
and U4008 (N_4008,N_3626,N_3560);
nand U4009 (N_4009,N_3635,N_3634);
and U4010 (N_4010,N_3974,N_3614);
or U4011 (N_4011,N_3889,N_3522);
nand U4012 (N_4012,N_3657,N_3902);
or U4013 (N_4013,N_3760,N_3698);
and U4014 (N_4014,N_3680,N_3621);
or U4015 (N_4015,N_3615,N_3801);
or U4016 (N_4016,N_3798,N_3994);
nor U4017 (N_4017,N_3714,N_3517);
nor U4018 (N_4018,N_3838,N_3816);
or U4019 (N_4019,N_3868,N_3793);
or U4020 (N_4020,N_3799,N_3664);
and U4021 (N_4021,N_3862,N_3843);
or U4022 (N_4022,N_3756,N_3542);
nand U4023 (N_4023,N_3589,N_3539);
and U4024 (N_4024,N_3774,N_3941);
nand U4025 (N_4025,N_3612,N_3649);
nand U4026 (N_4026,N_3518,N_3511);
nor U4027 (N_4027,N_3688,N_3565);
or U4028 (N_4028,N_3908,N_3643);
and U4029 (N_4029,N_3556,N_3527);
nor U4030 (N_4030,N_3863,N_3625);
and U4031 (N_4031,N_3602,N_3805);
nand U4032 (N_4032,N_3755,N_3828);
nand U4033 (N_4033,N_3747,N_3502);
or U4034 (N_4034,N_3700,N_3787);
and U4035 (N_4035,N_3748,N_3576);
or U4036 (N_4036,N_3582,N_3967);
nor U4037 (N_4037,N_3687,N_3622);
or U4038 (N_4038,N_3662,N_3544);
nand U4039 (N_4039,N_3830,N_3965);
or U4040 (N_4040,N_3978,N_3734);
nor U4041 (N_4041,N_3531,N_3865);
nor U4042 (N_4042,N_3987,N_3730);
nand U4043 (N_4043,N_3583,N_3786);
nor U4044 (N_4044,N_3746,N_3937);
and U4045 (N_4045,N_3877,N_3699);
nor U4046 (N_4046,N_3628,N_3872);
and U4047 (N_4047,N_3864,N_3999);
or U4048 (N_4048,N_3882,N_3919);
nand U4049 (N_4049,N_3766,N_3564);
and U4050 (N_4050,N_3982,N_3593);
nand U4051 (N_4051,N_3510,N_3546);
nand U4052 (N_4052,N_3859,N_3802);
nor U4053 (N_4053,N_3520,N_3618);
nor U4054 (N_4054,N_3806,N_3550);
and U4055 (N_4055,N_3599,N_3848);
and U4056 (N_4056,N_3610,N_3731);
and U4057 (N_4057,N_3638,N_3811);
or U4058 (N_4058,N_3726,N_3577);
nand U4059 (N_4059,N_3860,N_3948);
nand U4060 (N_4060,N_3934,N_3895);
or U4061 (N_4061,N_3765,N_3815);
and U4062 (N_4062,N_3888,N_3630);
or U4063 (N_4063,N_3823,N_3529);
and U4064 (N_4064,N_3856,N_3917);
and U4065 (N_4065,N_3789,N_3600);
nor U4066 (N_4066,N_3744,N_3822);
and U4067 (N_4067,N_3950,N_3585);
xor U4068 (N_4068,N_3866,N_3892);
nand U4069 (N_4069,N_3833,N_3525);
nand U4070 (N_4070,N_3549,N_3619);
nand U4071 (N_4071,N_3508,N_3944);
nor U4072 (N_4072,N_3795,N_3690);
and U4073 (N_4073,N_3901,N_3749);
or U4074 (N_4074,N_3504,N_3711);
nand U4075 (N_4075,N_3613,N_3562);
and U4076 (N_4076,N_3963,N_3706);
nand U4077 (N_4077,N_3738,N_3952);
and U4078 (N_4078,N_3691,N_3792);
nor U4079 (N_4079,N_3905,N_3874);
and U4080 (N_4080,N_3921,N_3608);
nor U4081 (N_4081,N_3935,N_3705);
nand U4082 (N_4082,N_3678,N_3962);
and U4083 (N_4083,N_3909,N_3587);
or U4084 (N_4084,N_3574,N_3954);
or U4085 (N_4085,N_3557,N_3910);
nor U4086 (N_4086,N_3671,N_3646);
nor U4087 (N_4087,N_3841,N_3637);
or U4088 (N_4088,N_3767,N_3885);
nand U4089 (N_4089,N_3972,N_3993);
or U4090 (N_4090,N_3837,N_3809);
nor U4091 (N_4091,N_3543,N_3829);
nor U4092 (N_4092,N_3826,N_3985);
nor U4093 (N_4093,N_3672,N_3778);
nand U4094 (N_4094,N_3553,N_3769);
nor U4095 (N_4095,N_3790,N_3729);
or U4096 (N_4096,N_3929,N_3605);
nor U4097 (N_4097,N_3505,N_3976);
nor U4098 (N_4098,N_3697,N_3572);
xnor U4099 (N_4099,N_3911,N_3580);
or U4100 (N_4100,N_3675,N_3509);
and U4101 (N_4101,N_3873,N_3567);
nand U4102 (N_4102,N_3658,N_3846);
or U4103 (N_4103,N_3578,N_3953);
and U4104 (N_4104,N_3853,N_3930);
and U4105 (N_4105,N_3652,N_3835);
nand U4106 (N_4106,N_3918,N_3717);
nand U4107 (N_4107,N_3904,N_3640);
nor U4108 (N_4108,N_3852,N_3762);
and U4109 (N_4109,N_3513,N_3581);
or U4110 (N_4110,N_3596,N_3530);
or U4111 (N_4111,N_3536,N_3552);
and U4112 (N_4112,N_3712,N_3588);
nand U4113 (N_4113,N_3839,N_3736);
nor U4114 (N_4114,N_3590,N_3685);
nand U4115 (N_4115,N_3973,N_3526);
nand U4116 (N_4116,N_3740,N_3931);
nand U4117 (N_4117,N_3551,N_3654);
nor U4118 (N_4118,N_3607,N_3884);
nor U4119 (N_4119,N_3849,N_3724);
and U4120 (N_4120,N_3927,N_3850);
nand U4121 (N_4121,N_3673,N_3983);
or U4122 (N_4122,N_3840,N_3779);
and U4123 (N_4123,N_3629,N_3913);
nand U4124 (N_4124,N_3641,N_3503);
nand U4125 (N_4125,N_3660,N_3689);
nand U4126 (N_4126,N_3532,N_3869);
nor U4127 (N_4127,N_3570,N_3514);
and U4128 (N_4128,N_3598,N_3571);
nand U4129 (N_4129,N_3939,N_3970);
or U4130 (N_4130,N_3507,N_3896);
or U4131 (N_4131,N_3986,N_3777);
or U4132 (N_4132,N_3964,N_3594);
nand U4133 (N_4133,N_3878,N_3897);
and U4134 (N_4134,N_3783,N_3844);
nand U4135 (N_4135,N_3788,N_3524);
or U4136 (N_4136,N_3745,N_3611);
and U4137 (N_4137,N_3782,N_3752);
or U4138 (N_4138,N_3655,N_3928);
xnor U4139 (N_4139,N_3692,N_3940);
and U4140 (N_4140,N_3701,N_3956);
or U4141 (N_4141,N_3616,N_3569);
xor U4142 (N_4142,N_3523,N_3758);
nor U4143 (N_4143,N_3707,N_3728);
nor U4144 (N_4144,N_3647,N_3883);
nor U4145 (N_4145,N_3780,N_3926);
and U4146 (N_4146,N_3923,N_3721);
or U4147 (N_4147,N_3946,N_3770);
or U4148 (N_4148,N_3968,N_3945);
and U4149 (N_4149,N_3659,N_3665);
nand U4150 (N_4150,N_3591,N_3784);
or U4151 (N_4151,N_3879,N_3703);
or U4152 (N_4152,N_3669,N_3667);
or U4153 (N_4153,N_3501,N_3521);
and U4154 (N_4154,N_3741,N_3771);
nand U4155 (N_4155,N_3966,N_3609);
and U4156 (N_4156,N_3847,N_3535);
or U4157 (N_4157,N_3915,N_3814);
and U4158 (N_4158,N_3891,N_3506);
and U4159 (N_4159,N_3559,N_3555);
or U4160 (N_4160,N_3713,N_3995);
or U4161 (N_4161,N_3980,N_3633);
nor U4162 (N_4162,N_3955,N_3554);
nand U4163 (N_4163,N_3754,N_3558);
and U4164 (N_4164,N_3836,N_3733);
and U4165 (N_4165,N_3781,N_3695);
and U4166 (N_4166,N_3515,N_3674);
nor U4167 (N_4167,N_3653,N_3694);
nor U4168 (N_4168,N_3606,N_3871);
and U4169 (N_4169,N_3797,N_3682);
and U4170 (N_4170,N_3750,N_3907);
nor U4171 (N_4171,N_3947,N_3881);
or U4172 (N_4172,N_3988,N_3597);
nand U4173 (N_4173,N_3776,N_3761);
or U4174 (N_4174,N_3916,N_3854);
and U4175 (N_4175,N_3894,N_3870);
nor U4176 (N_4176,N_3704,N_3832);
nor U4177 (N_4177,N_3725,N_3584);
and U4178 (N_4178,N_3764,N_3732);
nand U4179 (N_4179,N_3791,N_3723);
or U4180 (N_4180,N_3533,N_3912);
nor U4181 (N_4181,N_3735,N_3996);
nor U4182 (N_4182,N_3825,N_3709);
nand U4183 (N_4183,N_3932,N_3545);
nor U4184 (N_4184,N_3785,N_3632);
and U4185 (N_4185,N_3943,N_3537);
nand U4186 (N_4186,N_3715,N_3893);
and U4187 (N_4187,N_3684,N_3739);
nand U4188 (N_4188,N_3959,N_3817);
nand U4189 (N_4189,N_3623,N_3627);
nand U4190 (N_4190,N_3696,N_3708);
and U4191 (N_4191,N_3851,N_3679);
nand U4192 (N_4192,N_3548,N_3775);
or U4193 (N_4193,N_3656,N_3743);
nor U4194 (N_4194,N_3821,N_3681);
nand U4195 (N_4195,N_3924,N_3936);
nand U4196 (N_4196,N_3516,N_3796);
nand U4197 (N_4197,N_3922,N_3845);
nand U4198 (N_4198,N_3620,N_3960);
and U4199 (N_4199,N_3636,N_3800);
nor U4200 (N_4200,N_3981,N_3899);
nand U4201 (N_4201,N_3876,N_3759);
or U4202 (N_4202,N_3858,N_3538);
and U4203 (N_4203,N_3722,N_3834);
nor U4204 (N_4204,N_3903,N_3803);
and U4205 (N_4205,N_3818,N_3683);
and U4206 (N_4206,N_3603,N_3650);
nand U4207 (N_4207,N_3592,N_3686);
xor U4208 (N_4208,N_3842,N_3566);
or U4209 (N_4209,N_3855,N_3804);
nor U4210 (N_4210,N_3949,N_3595);
or U4211 (N_4211,N_3512,N_3768);
nor U4212 (N_4212,N_3977,N_3773);
and U4213 (N_4213,N_3648,N_3617);
and U4214 (N_4214,N_3819,N_3751);
nand U4215 (N_4215,N_3933,N_3742);
nand U4216 (N_4216,N_3989,N_3604);
nor U4217 (N_4217,N_3958,N_3875);
nand U4218 (N_4218,N_3575,N_3601);
and U4219 (N_4219,N_3719,N_3624);
and U4220 (N_4220,N_3957,N_3676);
and U4221 (N_4221,N_3718,N_3519);
nand U4222 (N_4222,N_3942,N_3693);
nor U4223 (N_4223,N_3702,N_3857);
nand U4224 (N_4224,N_3720,N_3808);
nand U4225 (N_4225,N_3661,N_3563);
or U4226 (N_4226,N_3668,N_3772);
and U4227 (N_4227,N_3900,N_3807);
nand U4228 (N_4228,N_3642,N_3991);
nor U4229 (N_4229,N_3528,N_3663);
or U4230 (N_4230,N_3914,N_3886);
and U4231 (N_4231,N_3969,N_3992);
and U4232 (N_4232,N_3631,N_3979);
nor U4233 (N_4233,N_3861,N_3920);
nor U4234 (N_4234,N_3561,N_3763);
nor U4235 (N_4235,N_3500,N_3810);
and U4236 (N_4236,N_3890,N_3824);
nor U4237 (N_4237,N_3831,N_3540);
or U4238 (N_4238,N_3541,N_3898);
and U4239 (N_4239,N_3645,N_3573);
and U4240 (N_4240,N_3820,N_3984);
nor U4241 (N_4241,N_3666,N_3867);
or U4242 (N_4242,N_3951,N_3925);
and U4243 (N_4243,N_3998,N_3644);
nor U4244 (N_4244,N_3727,N_3586);
nand U4245 (N_4245,N_3579,N_3534);
or U4246 (N_4246,N_3812,N_3990);
and U4247 (N_4247,N_3938,N_3757);
and U4248 (N_4248,N_3677,N_3906);
nor U4249 (N_4249,N_3827,N_3547);
nand U4250 (N_4250,N_3532,N_3600);
and U4251 (N_4251,N_3905,N_3833);
nor U4252 (N_4252,N_3943,N_3946);
nor U4253 (N_4253,N_3611,N_3858);
and U4254 (N_4254,N_3828,N_3781);
nor U4255 (N_4255,N_3597,N_3637);
and U4256 (N_4256,N_3825,N_3788);
xor U4257 (N_4257,N_3914,N_3533);
or U4258 (N_4258,N_3925,N_3959);
nand U4259 (N_4259,N_3740,N_3610);
or U4260 (N_4260,N_3719,N_3707);
and U4261 (N_4261,N_3849,N_3623);
and U4262 (N_4262,N_3975,N_3888);
nor U4263 (N_4263,N_3891,N_3855);
nor U4264 (N_4264,N_3988,N_3711);
nor U4265 (N_4265,N_3963,N_3894);
nand U4266 (N_4266,N_3683,N_3515);
nand U4267 (N_4267,N_3576,N_3921);
nor U4268 (N_4268,N_3870,N_3620);
nor U4269 (N_4269,N_3894,N_3944);
and U4270 (N_4270,N_3876,N_3732);
nor U4271 (N_4271,N_3765,N_3926);
nand U4272 (N_4272,N_3853,N_3983);
xnor U4273 (N_4273,N_3599,N_3696);
or U4274 (N_4274,N_3629,N_3561);
and U4275 (N_4275,N_3586,N_3684);
nor U4276 (N_4276,N_3671,N_3752);
and U4277 (N_4277,N_3787,N_3526);
nand U4278 (N_4278,N_3502,N_3916);
nor U4279 (N_4279,N_3597,N_3564);
xor U4280 (N_4280,N_3946,N_3590);
or U4281 (N_4281,N_3535,N_3654);
or U4282 (N_4282,N_3605,N_3639);
and U4283 (N_4283,N_3757,N_3593);
nor U4284 (N_4284,N_3974,N_3541);
or U4285 (N_4285,N_3630,N_3699);
nand U4286 (N_4286,N_3771,N_3911);
nand U4287 (N_4287,N_3630,N_3534);
and U4288 (N_4288,N_3596,N_3976);
or U4289 (N_4289,N_3624,N_3934);
nor U4290 (N_4290,N_3506,N_3774);
and U4291 (N_4291,N_3641,N_3925);
and U4292 (N_4292,N_3873,N_3940);
and U4293 (N_4293,N_3513,N_3545);
nand U4294 (N_4294,N_3776,N_3527);
and U4295 (N_4295,N_3717,N_3783);
nor U4296 (N_4296,N_3628,N_3572);
nor U4297 (N_4297,N_3635,N_3927);
and U4298 (N_4298,N_3779,N_3926);
and U4299 (N_4299,N_3831,N_3926);
or U4300 (N_4300,N_3777,N_3868);
nand U4301 (N_4301,N_3743,N_3630);
nand U4302 (N_4302,N_3851,N_3810);
and U4303 (N_4303,N_3797,N_3811);
and U4304 (N_4304,N_3654,N_3925);
and U4305 (N_4305,N_3821,N_3750);
or U4306 (N_4306,N_3582,N_3763);
or U4307 (N_4307,N_3876,N_3677);
and U4308 (N_4308,N_3790,N_3710);
or U4309 (N_4309,N_3690,N_3626);
xor U4310 (N_4310,N_3622,N_3594);
nor U4311 (N_4311,N_3937,N_3955);
or U4312 (N_4312,N_3691,N_3722);
or U4313 (N_4313,N_3669,N_3599);
nor U4314 (N_4314,N_3946,N_3618);
nor U4315 (N_4315,N_3681,N_3987);
nor U4316 (N_4316,N_3847,N_3684);
nor U4317 (N_4317,N_3536,N_3777);
and U4318 (N_4318,N_3740,N_3601);
or U4319 (N_4319,N_3726,N_3751);
nor U4320 (N_4320,N_3908,N_3597);
or U4321 (N_4321,N_3575,N_3885);
or U4322 (N_4322,N_3637,N_3886);
nand U4323 (N_4323,N_3793,N_3630);
nand U4324 (N_4324,N_3989,N_3760);
and U4325 (N_4325,N_3808,N_3695);
nand U4326 (N_4326,N_3611,N_3722);
and U4327 (N_4327,N_3524,N_3844);
nor U4328 (N_4328,N_3818,N_3815);
and U4329 (N_4329,N_3658,N_3898);
nand U4330 (N_4330,N_3853,N_3794);
and U4331 (N_4331,N_3905,N_3782);
nor U4332 (N_4332,N_3669,N_3754);
or U4333 (N_4333,N_3542,N_3910);
or U4334 (N_4334,N_3558,N_3965);
nand U4335 (N_4335,N_3673,N_3751);
and U4336 (N_4336,N_3605,N_3624);
nor U4337 (N_4337,N_3803,N_3738);
nand U4338 (N_4338,N_3511,N_3877);
and U4339 (N_4339,N_3508,N_3891);
or U4340 (N_4340,N_3639,N_3764);
and U4341 (N_4341,N_3589,N_3927);
or U4342 (N_4342,N_3517,N_3586);
and U4343 (N_4343,N_3812,N_3943);
or U4344 (N_4344,N_3773,N_3520);
and U4345 (N_4345,N_3944,N_3904);
nor U4346 (N_4346,N_3702,N_3696);
or U4347 (N_4347,N_3773,N_3523);
nor U4348 (N_4348,N_3514,N_3926);
and U4349 (N_4349,N_3966,N_3910);
or U4350 (N_4350,N_3580,N_3776);
nand U4351 (N_4351,N_3711,N_3779);
nor U4352 (N_4352,N_3837,N_3732);
nand U4353 (N_4353,N_3534,N_3748);
xnor U4354 (N_4354,N_3783,N_3504);
nor U4355 (N_4355,N_3955,N_3863);
or U4356 (N_4356,N_3725,N_3693);
nand U4357 (N_4357,N_3747,N_3847);
nand U4358 (N_4358,N_3725,N_3556);
and U4359 (N_4359,N_3769,N_3754);
nor U4360 (N_4360,N_3696,N_3712);
and U4361 (N_4361,N_3619,N_3748);
and U4362 (N_4362,N_3953,N_3643);
and U4363 (N_4363,N_3574,N_3926);
nand U4364 (N_4364,N_3833,N_3603);
nor U4365 (N_4365,N_3931,N_3600);
nand U4366 (N_4366,N_3681,N_3615);
or U4367 (N_4367,N_3877,N_3732);
and U4368 (N_4368,N_3939,N_3868);
and U4369 (N_4369,N_3655,N_3884);
nor U4370 (N_4370,N_3503,N_3733);
nor U4371 (N_4371,N_3752,N_3824);
nand U4372 (N_4372,N_3663,N_3802);
or U4373 (N_4373,N_3762,N_3790);
and U4374 (N_4374,N_3909,N_3872);
nor U4375 (N_4375,N_3747,N_3842);
or U4376 (N_4376,N_3845,N_3964);
or U4377 (N_4377,N_3508,N_3585);
nor U4378 (N_4378,N_3672,N_3738);
nor U4379 (N_4379,N_3920,N_3955);
nand U4380 (N_4380,N_3712,N_3769);
nand U4381 (N_4381,N_3997,N_3573);
nor U4382 (N_4382,N_3804,N_3900);
and U4383 (N_4383,N_3857,N_3875);
nand U4384 (N_4384,N_3506,N_3942);
or U4385 (N_4385,N_3520,N_3575);
nor U4386 (N_4386,N_3549,N_3828);
xnor U4387 (N_4387,N_3706,N_3815);
or U4388 (N_4388,N_3798,N_3972);
or U4389 (N_4389,N_3566,N_3647);
nand U4390 (N_4390,N_3948,N_3532);
nand U4391 (N_4391,N_3582,N_3781);
nand U4392 (N_4392,N_3554,N_3909);
nor U4393 (N_4393,N_3566,N_3790);
and U4394 (N_4394,N_3589,N_3884);
nand U4395 (N_4395,N_3542,N_3918);
and U4396 (N_4396,N_3779,N_3933);
nor U4397 (N_4397,N_3968,N_3781);
and U4398 (N_4398,N_3680,N_3507);
and U4399 (N_4399,N_3790,N_3878);
nor U4400 (N_4400,N_3813,N_3747);
nor U4401 (N_4401,N_3839,N_3890);
or U4402 (N_4402,N_3733,N_3740);
or U4403 (N_4403,N_3503,N_3517);
or U4404 (N_4404,N_3623,N_3980);
nand U4405 (N_4405,N_3865,N_3501);
xor U4406 (N_4406,N_3747,N_3749);
or U4407 (N_4407,N_3556,N_3557);
and U4408 (N_4408,N_3945,N_3655);
nand U4409 (N_4409,N_3781,N_3833);
or U4410 (N_4410,N_3850,N_3735);
and U4411 (N_4411,N_3986,N_3869);
nand U4412 (N_4412,N_3526,N_3809);
xor U4413 (N_4413,N_3980,N_3774);
and U4414 (N_4414,N_3942,N_3523);
nand U4415 (N_4415,N_3861,N_3839);
nor U4416 (N_4416,N_3850,N_3546);
or U4417 (N_4417,N_3575,N_3992);
nand U4418 (N_4418,N_3679,N_3994);
nand U4419 (N_4419,N_3606,N_3740);
nor U4420 (N_4420,N_3579,N_3866);
nand U4421 (N_4421,N_3583,N_3907);
or U4422 (N_4422,N_3688,N_3761);
and U4423 (N_4423,N_3893,N_3760);
nand U4424 (N_4424,N_3643,N_3533);
nand U4425 (N_4425,N_3630,N_3665);
and U4426 (N_4426,N_3830,N_3560);
and U4427 (N_4427,N_3545,N_3993);
nor U4428 (N_4428,N_3618,N_3851);
or U4429 (N_4429,N_3915,N_3810);
and U4430 (N_4430,N_3681,N_3995);
or U4431 (N_4431,N_3799,N_3919);
nand U4432 (N_4432,N_3581,N_3625);
nor U4433 (N_4433,N_3984,N_3894);
nor U4434 (N_4434,N_3887,N_3777);
and U4435 (N_4435,N_3827,N_3582);
nand U4436 (N_4436,N_3955,N_3867);
nand U4437 (N_4437,N_3774,N_3809);
and U4438 (N_4438,N_3924,N_3519);
xor U4439 (N_4439,N_3882,N_3950);
or U4440 (N_4440,N_3820,N_3885);
nand U4441 (N_4441,N_3670,N_3744);
or U4442 (N_4442,N_3774,N_3683);
or U4443 (N_4443,N_3952,N_3596);
or U4444 (N_4444,N_3907,N_3855);
and U4445 (N_4445,N_3602,N_3609);
nand U4446 (N_4446,N_3885,N_3928);
and U4447 (N_4447,N_3925,N_3882);
and U4448 (N_4448,N_3560,N_3656);
and U4449 (N_4449,N_3914,N_3503);
xor U4450 (N_4450,N_3515,N_3656);
nand U4451 (N_4451,N_3772,N_3555);
or U4452 (N_4452,N_3712,N_3985);
nand U4453 (N_4453,N_3718,N_3560);
and U4454 (N_4454,N_3755,N_3762);
and U4455 (N_4455,N_3563,N_3529);
nor U4456 (N_4456,N_3827,N_3974);
nand U4457 (N_4457,N_3927,N_3883);
and U4458 (N_4458,N_3717,N_3702);
and U4459 (N_4459,N_3597,N_3933);
and U4460 (N_4460,N_3571,N_3612);
nand U4461 (N_4461,N_3832,N_3801);
and U4462 (N_4462,N_3960,N_3701);
nor U4463 (N_4463,N_3921,N_3657);
nor U4464 (N_4464,N_3547,N_3989);
nand U4465 (N_4465,N_3733,N_3537);
nor U4466 (N_4466,N_3569,N_3905);
nor U4467 (N_4467,N_3722,N_3805);
nand U4468 (N_4468,N_3563,N_3536);
nand U4469 (N_4469,N_3930,N_3993);
and U4470 (N_4470,N_3556,N_3943);
or U4471 (N_4471,N_3741,N_3514);
nor U4472 (N_4472,N_3806,N_3534);
and U4473 (N_4473,N_3761,N_3720);
and U4474 (N_4474,N_3799,N_3683);
or U4475 (N_4475,N_3791,N_3974);
nand U4476 (N_4476,N_3686,N_3643);
or U4477 (N_4477,N_3697,N_3622);
or U4478 (N_4478,N_3658,N_3962);
nand U4479 (N_4479,N_3527,N_3578);
and U4480 (N_4480,N_3605,N_3838);
or U4481 (N_4481,N_3728,N_3987);
or U4482 (N_4482,N_3513,N_3757);
nor U4483 (N_4483,N_3830,N_3752);
and U4484 (N_4484,N_3899,N_3782);
nand U4485 (N_4485,N_3925,N_3915);
or U4486 (N_4486,N_3773,N_3519);
or U4487 (N_4487,N_3649,N_3901);
nand U4488 (N_4488,N_3551,N_3965);
or U4489 (N_4489,N_3585,N_3609);
and U4490 (N_4490,N_3780,N_3775);
nor U4491 (N_4491,N_3529,N_3678);
nand U4492 (N_4492,N_3725,N_3858);
or U4493 (N_4493,N_3537,N_3634);
and U4494 (N_4494,N_3982,N_3608);
nor U4495 (N_4495,N_3962,N_3996);
nand U4496 (N_4496,N_3863,N_3533);
and U4497 (N_4497,N_3849,N_3634);
and U4498 (N_4498,N_3642,N_3938);
or U4499 (N_4499,N_3831,N_3966);
nand U4500 (N_4500,N_4258,N_4375);
nand U4501 (N_4501,N_4453,N_4473);
xor U4502 (N_4502,N_4043,N_4178);
nor U4503 (N_4503,N_4196,N_4168);
and U4504 (N_4504,N_4463,N_4040);
or U4505 (N_4505,N_4144,N_4143);
or U4506 (N_4506,N_4136,N_4413);
and U4507 (N_4507,N_4187,N_4309);
and U4508 (N_4508,N_4365,N_4278);
nor U4509 (N_4509,N_4363,N_4414);
nor U4510 (N_4510,N_4210,N_4435);
nand U4511 (N_4511,N_4337,N_4117);
and U4512 (N_4512,N_4298,N_4087);
nor U4513 (N_4513,N_4247,N_4222);
nand U4514 (N_4514,N_4150,N_4038);
and U4515 (N_4515,N_4124,N_4377);
xnor U4516 (N_4516,N_4497,N_4049);
or U4517 (N_4517,N_4367,N_4475);
nor U4518 (N_4518,N_4307,N_4319);
and U4519 (N_4519,N_4304,N_4105);
nand U4520 (N_4520,N_4209,N_4442);
nand U4521 (N_4521,N_4181,N_4244);
and U4522 (N_4522,N_4107,N_4020);
nor U4523 (N_4523,N_4190,N_4028);
nand U4524 (N_4524,N_4132,N_4163);
nand U4525 (N_4525,N_4385,N_4321);
or U4526 (N_4526,N_4418,N_4013);
or U4527 (N_4527,N_4230,N_4391);
and U4528 (N_4528,N_4311,N_4289);
nand U4529 (N_4529,N_4341,N_4395);
nor U4530 (N_4530,N_4201,N_4416);
nand U4531 (N_4531,N_4283,N_4408);
or U4532 (N_4532,N_4001,N_4432);
and U4533 (N_4533,N_4084,N_4380);
and U4534 (N_4534,N_4184,N_4382);
or U4535 (N_4535,N_4110,N_4215);
or U4536 (N_4536,N_4131,N_4271);
nor U4537 (N_4537,N_4447,N_4485);
nand U4538 (N_4538,N_4401,N_4138);
and U4539 (N_4539,N_4329,N_4156);
and U4540 (N_4540,N_4441,N_4290);
nand U4541 (N_4541,N_4188,N_4157);
and U4542 (N_4542,N_4465,N_4220);
or U4543 (N_4543,N_4387,N_4456);
nor U4544 (N_4544,N_4285,N_4360);
or U4545 (N_4545,N_4388,N_4114);
nor U4546 (N_4546,N_4088,N_4098);
nor U4547 (N_4547,N_4279,N_4440);
nor U4548 (N_4548,N_4356,N_4005);
nor U4549 (N_4549,N_4364,N_4228);
nand U4550 (N_4550,N_4019,N_4306);
and U4551 (N_4551,N_4482,N_4390);
and U4552 (N_4552,N_4488,N_4434);
nor U4553 (N_4553,N_4324,N_4151);
nand U4554 (N_4554,N_4268,N_4249);
and U4555 (N_4555,N_4185,N_4255);
nor U4556 (N_4556,N_4443,N_4075);
nor U4557 (N_4557,N_4393,N_4097);
nor U4558 (N_4558,N_4152,N_4396);
nor U4559 (N_4559,N_4345,N_4242);
or U4560 (N_4560,N_4464,N_4133);
nor U4561 (N_4561,N_4373,N_4113);
nand U4562 (N_4562,N_4016,N_4027);
and U4563 (N_4563,N_4240,N_4112);
or U4564 (N_4564,N_4137,N_4366);
and U4565 (N_4565,N_4014,N_4331);
and U4566 (N_4566,N_4404,N_4468);
and U4567 (N_4567,N_4351,N_4427);
xor U4568 (N_4568,N_4284,N_4323);
nor U4569 (N_4569,N_4409,N_4370);
nor U4570 (N_4570,N_4122,N_4039);
nor U4571 (N_4571,N_4164,N_4257);
nor U4572 (N_4572,N_4402,N_4426);
nand U4573 (N_4573,N_4352,N_4275);
nand U4574 (N_4574,N_4357,N_4287);
or U4575 (N_4575,N_4080,N_4081);
or U4576 (N_4576,N_4448,N_4481);
or U4577 (N_4577,N_4291,N_4498);
and U4578 (N_4578,N_4006,N_4221);
nor U4579 (N_4579,N_4116,N_4262);
and U4580 (N_4580,N_4276,N_4436);
and U4581 (N_4581,N_4135,N_4322);
nand U4582 (N_4582,N_4047,N_4389);
and U4583 (N_4583,N_4051,N_4336);
nor U4584 (N_4584,N_4310,N_4328);
or U4585 (N_4585,N_4035,N_4159);
and U4586 (N_4586,N_4302,N_4126);
xnor U4587 (N_4587,N_4096,N_4374);
nor U4588 (N_4588,N_4073,N_4089);
nand U4589 (N_4589,N_4252,N_4248);
and U4590 (N_4590,N_4338,N_4076);
nor U4591 (N_4591,N_4277,N_4095);
or U4592 (N_4592,N_4128,N_4292);
nor U4593 (N_4593,N_4381,N_4063);
and U4594 (N_4594,N_4079,N_4218);
nor U4595 (N_4595,N_4224,N_4476);
xor U4596 (N_4596,N_4213,N_4272);
and U4597 (N_4597,N_4194,N_4176);
nor U4598 (N_4598,N_4359,N_4216);
nand U4599 (N_4599,N_4241,N_4118);
or U4600 (N_4600,N_4246,N_4266);
nand U4601 (N_4601,N_4055,N_4398);
nand U4602 (N_4602,N_4265,N_4412);
nand U4603 (N_4603,N_4177,N_4334);
and U4604 (N_4604,N_4149,N_4183);
nand U4605 (N_4605,N_4108,N_4003);
nor U4606 (N_4606,N_4036,N_4446);
nand U4607 (N_4607,N_4263,N_4361);
or U4608 (N_4608,N_4399,N_4032);
and U4609 (N_4609,N_4332,N_4077);
or U4610 (N_4610,N_4392,N_4227);
nand U4611 (N_4611,N_4010,N_4444);
nor U4612 (N_4612,N_4160,N_4474);
and U4613 (N_4613,N_4494,N_4109);
nand U4614 (N_4614,N_4161,N_4471);
and U4615 (N_4615,N_4425,N_4411);
nor U4616 (N_4616,N_4140,N_4064);
xor U4617 (N_4617,N_4312,N_4034);
or U4618 (N_4618,N_4031,N_4417);
or U4619 (N_4619,N_4335,N_4451);
nor U4620 (N_4620,N_4033,N_4026);
nand U4621 (N_4621,N_4061,N_4008);
nor U4622 (N_4622,N_4171,N_4460);
nor U4623 (N_4623,N_4368,N_4078);
and U4624 (N_4624,N_4214,N_4457);
nor U4625 (N_4625,N_4025,N_4251);
nand U4626 (N_4626,N_4407,N_4330);
and U4627 (N_4627,N_4123,N_4069);
and U4628 (N_4628,N_4383,N_4226);
nor U4629 (N_4629,N_4455,N_4207);
or U4630 (N_4630,N_4466,N_4231);
and U4631 (N_4631,N_4467,N_4121);
or U4632 (N_4632,N_4023,N_4091);
nor U4633 (N_4633,N_4045,N_4486);
nand U4634 (N_4634,N_4483,N_4420);
nand U4635 (N_4635,N_4256,N_4301);
and U4636 (N_4636,N_4155,N_4119);
and U4637 (N_4637,N_4294,N_4090);
nor U4638 (N_4638,N_4379,N_4115);
xor U4639 (N_4639,N_4030,N_4139);
nand U4640 (N_4640,N_4303,N_4470);
and U4641 (N_4641,N_4437,N_4146);
nand U4642 (N_4642,N_4093,N_4172);
or U4643 (N_4643,N_4259,N_4315);
nor U4644 (N_4644,N_4410,N_4102);
or U4645 (N_4645,N_4250,N_4120);
or U4646 (N_4646,N_4261,N_4491);
nand U4647 (N_4647,N_4449,N_4358);
nor U4648 (N_4648,N_4354,N_4326);
nor U4649 (N_4649,N_4142,N_4169);
and U4650 (N_4650,N_4127,N_4000);
nor U4651 (N_4651,N_4254,N_4293);
xnor U4652 (N_4652,N_4267,N_4104);
nor U4653 (N_4653,N_4349,N_4197);
or U4654 (N_4654,N_4342,N_4433);
and U4655 (N_4655,N_4074,N_4092);
or U4656 (N_4656,N_4371,N_4340);
nand U4657 (N_4657,N_4052,N_4492);
nor U4658 (N_4658,N_4200,N_4439);
nand U4659 (N_4659,N_4067,N_4384);
nor U4660 (N_4660,N_4192,N_4376);
or U4661 (N_4661,N_4461,N_4495);
nand U4662 (N_4662,N_4145,N_4101);
nor U4663 (N_4663,N_4348,N_4297);
nor U4664 (N_4664,N_4445,N_4308);
nor U4665 (N_4665,N_4239,N_4273);
and U4666 (N_4666,N_4191,N_4166);
or U4667 (N_4667,N_4170,N_4062);
and U4668 (N_4668,N_4086,N_4499);
nand U4669 (N_4669,N_4496,N_4158);
and U4670 (N_4670,N_4421,N_4288);
or U4671 (N_4671,N_4422,N_4217);
nand U4672 (N_4672,N_4477,N_4462);
nor U4673 (N_4673,N_4232,N_4175);
or U4674 (N_4674,N_4179,N_4129);
or U4675 (N_4675,N_4204,N_4180);
or U4676 (N_4676,N_4094,N_4346);
nor U4677 (N_4677,N_4487,N_4205);
or U4678 (N_4678,N_4264,N_4369);
or U4679 (N_4679,N_4225,N_4056);
nand U4680 (N_4680,N_4295,N_4148);
nor U4681 (N_4681,N_4208,N_4431);
nor U4682 (N_4682,N_4193,N_4206);
nor U4683 (N_4683,N_4423,N_4037);
nand U4684 (N_4684,N_4068,N_4182);
xnor U4685 (N_4685,N_4245,N_4058);
and U4686 (N_4686,N_4362,N_4054);
and U4687 (N_4687,N_4313,N_4378);
or U4688 (N_4688,N_4424,N_4484);
nor U4689 (N_4689,N_4198,N_4282);
nand U4690 (N_4690,N_4203,N_4022);
nand U4691 (N_4691,N_4071,N_4333);
or U4692 (N_4692,N_4042,N_4141);
nand U4693 (N_4693,N_4317,N_4320);
or U4694 (N_4694,N_4325,N_4235);
or U4695 (N_4695,N_4286,N_4134);
nor U4696 (N_4696,N_4048,N_4314);
xor U4697 (N_4697,N_4017,N_4186);
or U4698 (N_4698,N_4029,N_4478);
or U4699 (N_4699,N_4355,N_4270);
nand U4700 (N_4700,N_4438,N_4386);
or U4701 (N_4701,N_4004,N_4070);
nor U4702 (N_4702,N_4253,N_4237);
and U4703 (N_4703,N_4002,N_4162);
or U4704 (N_4704,N_4012,N_4147);
nor U4705 (N_4705,N_4007,N_4274);
and U4706 (N_4706,N_4327,N_4125);
or U4707 (N_4707,N_4299,N_4099);
and U4708 (N_4708,N_4472,N_4238);
nor U4709 (N_4709,N_4415,N_4165);
and U4710 (N_4710,N_4479,N_4085);
or U4711 (N_4711,N_4212,N_4189);
nand U4712 (N_4712,N_4173,N_4344);
nand U4713 (N_4713,N_4452,N_4400);
and U4714 (N_4714,N_4174,N_4397);
nand U4715 (N_4715,N_4103,N_4280);
and U4716 (N_4716,N_4153,N_4300);
and U4717 (N_4717,N_4044,N_4018);
nand U4718 (N_4718,N_4202,N_4234);
nand U4719 (N_4719,N_4243,N_4458);
or U4720 (N_4720,N_4490,N_4480);
nor U4721 (N_4721,N_4233,N_4223);
nor U4722 (N_4722,N_4195,N_4429);
and U4723 (N_4723,N_4372,N_4339);
nor U4724 (N_4724,N_4130,N_4350);
xor U4725 (N_4725,N_4024,N_4343);
or U4726 (N_4726,N_4229,N_4111);
and U4727 (N_4727,N_4100,N_4347);
nor U4728 (N_4728,N_4083,N_4260);
and U4729 (N_4729,N_4053,N_4459);
nor U4730 (N_4730,N_4199,N_4060);
nand U4731 (N_4731,N_4236,N_4305);
and U4732 (N_4732,N_4082,N_4021);
or U4733 (N_4733,N_4430,N_4489);
nand U4734 (N_4734,N_4219,N_4065);
nand U4735 (N_4735,N_4419,N_4450);
or U4736 (N_4736,N_4059,N_4394);
and U4737 (N_4737,N_4072,N_4106);
or U4738 (N_4738,N_4318,N_4269);
nor U4739 (N_4739,N_4211,N_4154);
and U4740 (N_4740,N_4009,N_4316);
or U4741 (N_4741,N_4167,N_4406);
or U4742 (N_4742,N_4281,N_4046);
or U4743 (N_4743,N_4066,N_4011);
or U4744 (N_4744,N_4493,N_4057);
or U4745 (N_4745,N_4403,N_4454);
xnor U4746 (N_4746,N_4405,N_4428);
nand U4747 (N_4747,N_4041,N_4015);
nand U4748 (N_4748,N_4296,N_4050);
nand U4749 (N_4749,N_4353,N_4469);
or U4750 (N_4750,N_4005,N_4339);
and U4751 (N_4751,N_4017,N_4387);
nand U4752 (N_4752,N_4050,N_4461);
and U4753 (N_4753,N_4102,N_4387);
nand U4754 (N_4754,N_4316,N_4036);
nand U4755 (N_4755,N_4031,N_4101);
nand U4756 (N_4756,N_4340,N_4355);
and U4757 (N_4757,N_4454,N_4463);
or U4758 (N_4758,N_4365,N_4465);
nand U4759 (N_4759,N_4099,N_4389);
or U4760 (N_4760,N_4279,N_4031);
and U4761 (N_4761,N_4487,N_4499);
nor U4762 (N_4762,N_4303,N_4062);
or U4763 (N_4763,N_4337,N_4300);
nand U4764 (N_4764,N_4237,N_4375);
and U4765 (N_4765,N_4262,N_4467);
or U4766 (N_4766,N_4083,N_4098);
nand U4767 (N_4767,N_4204,N_4194);
nor U4768 (N_4768,N_4101,N_4128);
nand U4769 (N_4769,N_4184,N_4192);
xnor U4770 (N_4770,N_4219,N_4309);
or U4771 (N_4771,N_4240,N_4152);
nand U4772 (N_4772,N_4390,N_4205);
nor U4773 (N_4773,N_4496,N_4082);
or U4774 (N_4774,N_4232,N_4479);
nor U4775 (N_4775,N_4386,N_4271);
and U4776 (N_4776,N_4069,N_4011);
or U4777 (N_4777,N_4218,N_4207);
or U4778 (N_4778,N_4392,N_4409);
or U4779 (N_4779,N_4195,N_4458);
nor U4780 (N_4780,N_4269,N_4308);
nor U4781 (N_4781,N_4170,N_4226);
or U4782 (N_4782,N_4370,N_4013);
and U4783 (N_4783,N_4168,N_4198);
nor U4784 (N_4784,N_4188,N_4344);
nand U4785 (N_4785,N_4472,N_4174);
nand U4786 (N_4786,N_4473,N_4131);
nand U4787 (N_4787,N_4316,N_4369);
or U4788 (N_4788,N_4475,N_4462);
and U4789 (N_4789,N_4310,N_4186);
nand U4790 (N_4790,N_4286,N_4446);
and U4791 (N_4791,N_4470,N_4279);
or U4792 (N_4792,N_4068,N_4263);
nand U4793 (N_4793,N_4137,N_4193);
xor U4794 (N_4794,N_4038,N_4050);
or U4795 (N_4795,N_4215,N_4217);
nor U4796 (N_4796,N_4118,N_4406);
nand U4797 (N_4797,N_4216,N_4245);
nor U4798 (N_4798,N_4174,N_4030);
or U4799 (N_4799,N_4198,N_4351);
nor U4800 (N_4800,N_4227,N_4139);
nor U4801 (N_4801,N_4118,N_4396);
or U4802 (N_4802,N_4350,N_4200);
nor U4803 (N_4803,N_4182,N_4040);
or U4804 (N_4804,N_4444,N_4232);
nand U4805 (N_4805,N_4427,N_4282);
nor U4806 (N_4806,N_4184,N_4222);
or U4807 (N_4807,N_4412,N_4072);
nor U4808 (N_4808,N_4023,N_4008);
and U4809 (N_4809,N_4268,N_4023);
nor U4810 (N_4810,N_4301,N_4460);
nand U4811 (N_4811,N_4123,N_4356);
or U4812 (N_4812,N_4085,N_4100);
nand U4813 (N_4813,N_4431,N_4025);
nor U4814 (N_4814,N_4408,N_4282);
or U4815 (N_4815,N_4248,N_4249);
nor U4816 (N_4816,N_4102,N_4055);
nor U4817 (N_4817,N_4374,N_4033);
or U4818 (N_4818,N_4164,N_4029);
and U4819 (N_4819,N_4305,N_4111);
nand U4820 (N_4820,N_4171,N_4008);
or U4821 (N_4821,N_4037,N_4151);
or U4822 (N_4822,N_4234,N_4451);
xnor U4823 (N_4823,N_4087,N_4209);
nand U4824 (N_4824,N_4279,N_4292);
nand U4825 (N_4825,N_4244,N_4379);
or U4826 (N_4826,N_4403,N_4339);
and U4827 (N_4827,N_4162,N_4210);
and U4828 (N_4828,N_4389,N_4424);
nand U4829 (N_4829,N_4051,N_4115);
and U4830 (N_4830,N_4244,N_4306);
nor U4831 (N_4831,N_4216,N_4136);
and U4832 (N_4832,N_4330,N_4108);
nor U4833 (N_4833,N_4309,N_4266);
and U4834 (N_4834,N_4264,N_4465);
or U4835 (N_4835,N_4250,N_4033);
nand U4836 (N_4836,N_4451,N_4291);
nand U4837 (N_4837,N_4436,N_4409);
or U4838 (N_4838,N_4345,N_4187);
and U4839 (N_4839,N_4176,N_4335);
and U4840 (N_4840,N_4345,N_4264);
and U4841 (N_4841,N_4441,N_4142);
and U4842 (N_4842,N_4182,N_4026);
nand U4843 (N_4843,N_4262,N_4328);
nor U4844 (N_4844,N_4027,N_4316);
nor U4845 (N_4845,N_4464,N_4448);
nor U4846 (N_4846,N_4428,N_4033);
or U4847 (N_4847,N_4004,N_4486);
nor U4848 (N_4848,N_4363,N_4117);
and U4849 (N_4849,N_4190,N_4016);
nand U4850 (N_4850,N_4162,N_4462);
xnor U4851 (N_4851,N_4144,N_4130);
nand U4852 (N_4852,N_4040,N_4460);
nand U4853 (N_4853,N_4432,N_4474);
nand U4854 (N_4854,N_4104,N_4131);
or U4855 (N_4855,N_4188,N_4151);
or U4856 (N_4856,N_4131,N_4486);
nand U4857 (N_4857,N_4180,N_4365);
or U4858 (N_4858,N_4212,N_4306);
or U4859 (N_4859,N_4042,N_4138);
or U4860 (N_4860,N_4113,N_4182);
nor U4861 (N_4861,N_4084,N_4335);
nor U4862 (N_4862,N_4128,N_4035);
or U4863 (N_4863,N_4348,N_4175);
nor U4864 (N_4864,N_4370,N_4251);
and U4865 (N_4865,N_4240,N_4364);
nand U4866 (N_4866,N_4074,N_4240);
nand U4867 (N_4867,N_4152,N_4022);
nor U4868 (N_4868,N_4278,N_4404);
nor U4869 (N_4869,N_4049,N_4044);
nor U4870 (N_4870,N_4408,N_4032);
nor U4871 (N_4871,N_4016,N_4436);
nor U4872 (N_4872,N_4371,N_4108);
nor U4873 (N_4873,N_4028,N_4298);
nor U4874 (N_4874,N_4237,N_4401);
or U4875 (N_4875,N_4472,N_4321);
or U4876 (N_4876,N_4097,N_4281);
xor U4877 (N_4877,N_4102,N_4358);
and U4878 (N_4878,N_4410,N_4161);
and U4879 (N_4879,N_4020,N_4159);
nand U4880 (N_4880,N_4255,N_4013);
nor U4881 (N_4881,N_4154,N_4265);
and U4882 (N_4882,N_4251,N_4459);
or U4883 (N_4883,N_4338,N_4497);
nor U4884 (N_4884,N_4289,N_4425);
nor U4885 (N_4885,N_4099,N_4364);
and U4886 (N_4886,N_4088,N_4179);
and U4887 (N_4887,N_4168,N_4308);
nand U4888 (N_4888,N_4402,N_4274);
nor U4889 (N_4889,N_4193,N_4142);
or U4890 (N_4890,N_4117,N_4247);
and U4891 (N_4891,N_4072,N_4275);
nand U4892 (N_4892,N_4291,N_4151);
and U4893 (N_4893,N_4262,N_4234);
nor U4894 (N_4894,N_4476,N_4294);
and U4895 (N_4895,N_4159,N_4443);
nor U4896 (N_4896,N_4334,N_4371);
nor U4897 (N_4897,N_4484,N_4077);
and U4898 (N_4898,N_4499,N_4062);
and U4899 (N_4899,N_4252,N_4120);
nor U4900 (N_4900,N_4101,N_4329);
or U4901 (N_4901,N_4071,N_4191);
and U4902 (N_4902,N_4196,N_4058);
nand U4903 (N_4903,N_4377,N_4136);
or U4904 (N_4904,N_4230,N_4324);
and U4905 (N_4905,N_4088,N_4437);
or U4906 (N_4906,N_4023,N_4481);
and U4907 (N_4907,N_4093,N_4359);
nand U4908 (N_4908,N_4016,N_4166);
nor U4909 (N_4909,N_4142,N_4306);
nor U4910 (N_4910,N_4310,N_4082);
or U4911 (N_4911,N_4214,N_4429);
and U4912 (N_4912,N_4423,N_4190);
or U4913 (N_4913,N_4174,N_4093);
nand U4914 (N_4914,N_4496,N_4367);
nor U4915 (N_4915,N_4157,N_4124);
nor U4916 (N_4916,N_4254,N_4098);
nand U4917 (N_4917,N_4315,N_4177);
and U4918 (N_4918,N_4465,N_4328);
nand U4919 (N_4919,N_4008,N_4179);
or U4920 (N_4920,N_4179,N_4440);
and U4921 (N_4921,N_4087,N_4027);
and U4922 (N_4922,N_4363,N_4435);
or U4923 (N_4923,N_4005,N_4103);
nand U4924 (N_4924,N_4109,N_4346);
and U4925 (N_4925,N_4210,N_4412);
or U4926 (N_4926,N_4076,N_4319);
and U4927 (N_4927,N_4361,N_4498);
nand U4928 (N_4928,N_4388,N_4309);
nor U4929 (N_4929,N_4091,N_4465);
nand U4930 (N_4930,N_4420,N_4111);
and U4931 (N_4931,N_4167,N_4380);
or U4932 (N_4932,N_4337,N_4057);
nand U4933 (N_4933,N_4305,N_4366);
nand U4934 (N_4934,N_4270,N_4056);
nand U4935 (N_4935,N_4288,N_4196);
or U4936 (N_4936,N_4298,N_4180);
and U4937 (N_4937,N_4164,N_4225);
nor U4938 (N_4938,N_4455,N_4316);
nor U4939 (N_4939,N_4302,N_4369);
nand U4940 (N_4940,N_4342,N_4237);
and U4941 (N_4941,N_4094,N_4442);
nor U4942 (N_4942,N_4107,N_4248);
nor U4943 (N_4943,N_4120,N_4096);
and U4944 (N_4944,N_4282,N_4304);
or U4945 (N_4945,N_4385,N_4071);
or U4946 (N_4946,N_4080,N_4470);
nor U4947 (N_4947,N_4383,N_4339);
nor U4948 (N_4948,N_4301,N_4188);
and U4949 (N_4949,N_4419,N_4479);
or U4950 (N_4950,N_4200,N_4354);
and U4951 (N_4951,N_4116,N_4040);
nor U4952 (N_4952,N_4496,N_4469);
nand U4953 (N_4953,N_4479,N_4362);
nor U4954 (N_4954,N_4073,N_4488);
or U4955 (N_4955,N_4488,N_4147);
nor U4956 (N_4956,N_4017,N_4272);
or U4957 (N_4957,N_4413,N_4004);
nand U4958 (N_4958,N_4479,N_4358);
nand U4959 (N_4959,N_4297,N_4209);
xor U4960 (N_4960,N_4427,N_4073);
nand U4961 (N_4961,N_4245,N_4073);
or U4962 (N_4962,N_4021,N_4198);
or U4963 (N_4963,N_4190,N_4059);
nor U4964 (N_4964,N_4099,N_4234);
and U4965 (N_4965,N_4258,N_4057);
or U4966 (N_4966,N_4000,N_4262);
xnor U4967 (N_4967,N_4363,N_4394);
and U4968 (N_4968,N_4303,N_4444);
nand U4969 (N_4969,N_4448,N_4115);
and U4970 (N_4970,N_4271,N_4029);
nor U4971 (N_4971,N_4448,N_4384);
nor U4972 (N_4972,N_4383,N_4452);
nor U4973 (N_4973,N_4009,N_4104);
nand U4974 (N_4974,N_4189,N_4426);
nor U4975 (N_4975,N_4482,N_4315);
and U4976 (N_4976,N_4222,N_4414);
nand U4977 (N_4977,N_4431,N_4373);
and U4978 (N_4978,N_4098,N_4164);
and U4979 (N_4979,N_4213,N_4081);
nor U4980 (N_4980,N_4395,N_4210);
or U4981 (N_4981,N_4091,N_4365);
nor U4982 (N_4982,N_4189,N_4434);
or U4983 (N_4983,N_4390,N_4044);
nand U4984 (N_4984,N_4074,N_4115);
nor U4985 (N_4985,N_4129,N_4153);
and U4986 (N_4986,N_4120,N_4354);
nor U4987 (N_4987,N_4115,N_4313);
xnor U4988 (N_4988,N_4198,N_4414);
or U4989 (N_4989,N_4089,N_4415);
or U4990 (N_4990,N_4164,N_4186);
or U4991 (N_4991,N_4253,N_4492);
or U4992 (N_4992,N_4428,N_4476);
nor U4993 (N_4993,N_4051,N_4128);
nor U4994 (N_4994,N_4077,N_4253);
nand U4995 (N_4995,N_4370,N_4452);
and U4996 (N_4996,N_4427,N_4061);
nor U4997 (N_4997,N_4328,N_4098);
nand U4998 (N_4998,N_4258,N_4324);
xor U4999 (N_4999,N_4310,N_4396);
nand UO_0 (O_0,N_4695,N_4711);
and UO_1 (O_1,N_4837,N_4925);
nor UO_2 (O_2,N_4567,N_4657);
and UO_3 (O_3,N_4787,N_4861);
nand UO_4 (O_4,N_4819,N_4656);
or UO_5 (O_5,N_4870,N_4991);
and UO_6 (O_6,N_4669,N_4697);
nand UO_7 (O_7,N_4826,N_4782);
nand UO_8 (O_8,N_4962,N_4548);
and UO_9 (O_9,N_4974,N_4586);
nand UO_10 (O_10,N_4642,N_4676);
or UO_11 (O_11,N_4988,N_4628);
or UO_12 (O_12,N_4707,N_4747);
and UO_13 (O_13,N_4599,N_4802);
and UO_14 (O_14,N_4886,N_4850);
nand UO_15 (O_15,N_4934,N_4938);
nor UO_16 (O_16,N_4994,N_4705);
and UO_17 (O_17,N_4767,N_4763);
or UO_18 (O_18,N_4738,N_4739);
nand UO_19 (O_19,N_4954,N_4791);
and UO_20 (O_20,N_4950,N_4955);
nor UO_21 (O_21,N_4724,N_4872);
nor UO_22 (O_22,N_4587,N_4947);
and UO_23 (O_23,N_4948,N_4523);
or UO_24 (O_24,N_4919,N_4671);
and UO_25 (O_25,N_4893,N_4990);
and UO_26 (O_26,N_4881,N_4598);
nor UO_27 (O_27,N_4627,N_4744);
and UO_28 (O_28,N_4976,N_4588);
nor UO_29 (O_29,N_4923,N_4924);
nand UO_30 (O_30,N_4666,N_4559);
nand UO_31 (O_31,N_4971,N_4832);
nand UO_32 (O_32,N_4603,N_4970);
nor UO_33 (O_33,N_4932,N_4633);
or UO_34 (O_34,N_4665,N_4883);
and UO_35 (O_35,N_4765,N_4838);
nor UO_36 (O_36,N_4735,N_4847);
or UO_37 (O_37,N_4898,N_4564);
and UO_38 (O_38,N_4681,N_4888);
nor UO_39 (O_39,N_4961,N_4756);
nor UO_40 (O_40,N_4785,N_4877);
nand UO_41 (O_41,N_4736,N_4640);
nand UO_42 (O_42,N_4800,N_4538);
nand UO_43 (O_43,N_4933,N_4967);
and UO_44 (O_44,N_4814,N_4986);
or UO_45 (O_45,N_4605,N_4606);
nor UO_46 (O_46,N_4788,N_4664);
or UO_47 (O_47,N_4981,N_4778);
nor UO_48 (O_48,N_4698,N_4508);
xor UO_49 (O_49,N_4966,N_4550);
nor UO_50 (O_50,N_4648,N_4719);
nor UO_51 (O_51,N_4912,N_4515);
and UO_52 (O_52,N_4764,N_4636);
and UO_53 (O_53,N_4983,N_4793);
nor UO_54 (O_54,N_4649,N_4944);
or UO_55 (O_55,N_4833,N_4821);
nor UO_56 (O_56,N_4634,N_4687);
xor UO_57 (O_57,N_4600,N_4609);
nor UO_58 (O_58,N_4722,N_4834);
nand UO_59 (O_59,N_4901,N_4549);
and UO_60 (O_60,N_4561,N_4558);
nor UO_61 (O_61,N_4854,N_4593);
or UO_62 (O_62,N_4980,N_4964);
xor UO_63 (O_63,N_4867,N_4957);
xor UO_64 (O_64,N_4562,N_4859);
or UO_65 (O_65,N_4841,N_4998);
nand UO_66 (O_66,N_4750,N_4995);
nor UO_67 (O_67,N_4701,N_4873);
nor UO_68 (O_68,N_4942,N_4706);
or UO_69 (O_69,N_4977,N_4720);
and UO_70 (O_70,N_4613,N_4978);
and UO_71 (O_71,N_4848,N_4668);
or UO_72 (O_72,N_4553,N_4928);
nand UO_73 (O_73,N_4647,N_4969);
and UO_74 (O_74,N_4540,N_4709);
nand UO_75 (O_75,N_4547,N_4997);
nand UO_76 (O_76,N_4616,N_4560);
and UO_77 (O_77,N_4646,N_4611);
or UO_78 (O_78,N_4895,N_4573);
nor UO_79 (O_79,N_4694,N_4989);
and UO_80 (O_80,N_4725,N_4885);
or UO_81 (O_81,N_4541,N_4945);
nand UO_82 (O_82,N_4604,N_4535);
or UO_83 (O_83,N_4731,N_4805);
nor UO_84 (O_84,N_4830,N_4690);
or UO_85 (O_85,N_4512,N_4552);
nor UO_86 (O_86,N_4825,N_4817);
or UO_87 (O_87,N_4855,N_4811);
or UO_88 (O_88,N_4503,N_4776);
or UO_89 (O_89,N_4596,N_4777);
nand UO_90 (O_90,N_4622,N_4670);
nor UO_91 (O_91,N_4715,N_4931);
and UO_92 (O_92,N_4520,N_4984);
nand UO_93 (O_93,N_4810,N_4632);
and UO_94 (O_94,N_4638,N_4816);
nand UO_95 (O_95,N_4526,N_4953);
and UO_96 (O_96,N_4685,N_4792);
nand UO_97 (O_97,N_4799,N_4884);
and UO_98 (O_98,N_4740,N_4667);
and UO_99 (O_99,N_4992,N_4982);
nor UO_100 (O_100,N_4557,N_4581);
nand UO_101 (O_101,N_4631,N_4514);
nand UO_102 (O_102,N_4653,N_4568);
nand UO_103 (O_103,N_4660,N_4614);
and UO_104 (O_104,N_4835,N_4892);
or UO_105 (O_105,N_4516,N_4539);
and UO_106 (O_106,N_4863,N_4659);
and UO_107 (O_107,N_4839,N_4882);
or UO_108 (O_108,N_4975,N_4713);
nand UO_109 (O_109,N_4796,N_4852);
and UO_110 (O_110,N_4965,N_4688);
nand UO_111 (O_111,N_4758,N_4663);
or UO_112 (O_112,N_4645,N_4607);
and UO_113 (O_113,N_4987,N_4973);
nand UO_114 (O_114,N_4595,N_4643);
xnor UO_115 (O_115,N_4730,N_4570);
nand UO_116 (O_116,N_4718,N_4755);
nand UO_117 (O_117,N_4789,N_4522);
and UO_118 (O_118,N_4536,N_4673);
and UO_119 (O_119,N_4909,N_4921);
nor UO_120 (O_120,N_4617,N_4531);
nand UO_121 (O_121,N_4906,N_4807);
or UO_122 (O_122,N_4639,N_4780);
nor UO_123 (O_123,N_4786,N_4517);
nor UO_124 (O_124,N_4565,N_4704);
and UO_125 (O_125,N_4678,N_4521);
nand UO_126 (O_126,N_4630,N_4662);
xor UO_127 (O_127,N_4554,N_4712);
and UO_128 (O_128,N_4504,N_4551);
or UO_129 (O_129,N_4626,N_4537);
nand UO_130 (O_130,N_4745,N_4917);
nor UO_131 (O_131,N_4529,N_4920);
and UO_132 (O_132,N_4576,N_4904);
nand UO_133 (O_133,N_4675,N_4737);
nor UO_134 (O_134,N_4686,N_4635);
nand UO_135 (O_135,N_4556,N_4612);
or UO_136 (O_136,N_4829,N_4996);
nand UO_137 (O_137,N_4899,N_4571);
nand UO_138 (O_138,N_4768,N_4672);
and UO_139 (O_139,N_4913,N_4615);
and UO_140 (O_140,N_4922,N_4851);
nand UO_141 (O_141,N_4702,N_4849);
and UO_142 (O_142,N_4519,N_4623);
nor UO_143 (O_143,N_4812,N_4692);
nor UO_144 (O_144,N_4710,N_4887);
and UO_145 (O_145,N_4908,N_4751);
and UO_146 (O_146,N_4869,N_4907);
nor UO_147 (O_147,N_4813,N_4960);
and UO_148 (O_148,N_4771,N_4809);
nand UO_149 (O_149,N_4524,N_4930);
and UO_150 (O_150,N_4746,N_4579);
xor UO_151 (O_151,N_4620,N_4696);
nor UO_152 (O_152,N_4741,N_4716);
or UO_153 (O_153,N_4896,N_4608);
nand UO_154 (O_154,N_4584,N_4822);
or UO_155 (O_155,N_4530,N_4952);
or UO_156 (O_156,N_4815,N_4858);
nand UO_157 (O_157,N_4618,N_4940);
or UO_158 (O_158,N_4625,N_4889);
nand UO_159 (O_159,N_4781,N_4582);
nor UO_160 (O_160,N_4784,N_4985);
nor UO_161 (O_161,N_4958,N_4594);
and UO_162 (O_162,N_4684,N_4823);
nand UO_163 (O_163,N_4926,N_4871);
nand UO_164 (O_164,N_4546,N_4937);
nand UO_165 (O_165,N_4875,N_4773);
nor UO_166 (O_166,N_4533,N_4742);
nor UO_167 (O_167,N_4689,N_4699);
or UO_168 (O_168,N_4801,N_4808);
nor UO_169 (O_169,N_4574,N_4602);
nand UO_170 (O_170,N_4790,N_4677);
nand UO_171 (O_171,N_4629,N_4703);
or UO_172 (O_172,N_4693,N_4769);
nor UO_173 (O_173,N_4654,N_4916);
nor UO_174 (O_174,N_4717,N_4874);
nand UO_175 (O_175,N_4783,N_4624);
nand UO_176 (O_176,N_4798,N_4759);
or UO_177 (O_177,N_4846,N_4655);
and UO_178 (O_178,N_4972,N_4824);
and UO_179 (O_179,N_4866,N_4569);
and UO_180 (O_180,N_4806,N_4856);
nor UO_181 (O_181,N_4864,N_4840);
and UO_182 (O_182,N_4910,N_4532);
or UO_183 (O_183,N_4865,N_4591);
or UO_184 (O_184,N_4658,N_4652);
or UO_185 (O_185,N_4610,N_4661);
nand UO_186 (O_186,N_4506,N_4525);
or UO_187 (O_187,N_4897,N_4827);
nand UO_188 (O_188,N_4754,N_4585);
nor UO_189 (O_189,N_4803,N_4580);
or UO_190 (O_190,N_4733,N_4949);
or UO_191 (O_191,N_4510,N_4583);
nand UO_192 (O_192,N_4843,N_4844);
and UO_193 (O_193,N_4727,N_4749);
nand UO_194 (O_194,N_4507,N_4728);
or UO_195 (O_195,N_4939,N_4641);
and UO_196 (O_196,N_4891,N_4723);
nor UO_197 (O_197,N_4878,N_4774);
or UO_198 (O_198,N_4578,N_4726);
nand UO_199 (O_199,N_4820,N_4589);
or UO_200 (O_200,N_4753,N_4505);
and UO_201 (O_201,N_4757,N_4857);
and UO_202 (O_202,N_4592,N_4518);
and UO_203 (O_203,N_4818,N_4779);
or UO_204 (O_204,N_4650,N_4831);
and UO_205 (O_205,N_4963,N_4601);
nand UO_206 (O_206,N_4880,N_4979);
or UO_207 (O_207,N_4879,N_4894);
nor UO_208 (O_208,N_4918,N_4683);
and UO_209 (O_209,N_4743,N_4761);
nand UO_210 (O_210,N_4619,N_4674);
nor UO_211 (O_211,N_4959,N_4914);
and UO_212 (O_212,N_4842,N_4902);
nand UO_213 (O_213,N_4797,N_4714);
nand UO_214 (O_214,N_4577,N_4734);
and UO_215 (O_215,N_4691,N_4951);
nor UO_216 (O_216,N_4682,N_4563);
or UO_217 (O_217,N_4905,N_4766);
nor UO_218 (O_218,N_4501,N_4566);
or UO_219 (O_219,N_4509,N_4502);
and UO_220 (O_220,N_4943,N_4936);
and UO_221 (O_221,N_4590,N_4500);
and UO_222 (O_222,N_4935,N_4968);
nand UO_223 (O_223,N_4956,N_4545);
nor UO_224 (O_224,N_4544,N_4637);
or UO_225 (O_225,N_4679,N_4804);
and UO_226 (O_226,N_4915,N_4543);
and UO_227 (O_227,N_4721,N_4770);
and UO_228 (O_228,N_4862,N_4795);
or UO_229 (O_229,N_4644,N_4941);
xnor UO_230 (O_230,N_4900,N_4762);
and UO_231 (O_231,N_4794,N_4772);
and UO_232 (O_232,N_4527,N_4993);
nand UO_233 (O_233,N_4700,N_4876);
nand UO_234 (O_234,N_4597,N_4890);
and UO_235 (O_235,N_4621,N_4828);
nand UO_236 (O_236,N_4572,N_4752);
and UO_237 (O_237,N_4732,N_4511);
and UO_238 (O_238,N_4836,N_4845);
nor UO_239 (O_239,N_4999,N_4927);
nor UO_240 (O_240,N_4946,N_4680);
or UO_241 (O_241,N_4651,N_4748);
nand UO_242 (O_242,N_4853,N_4513);
and UO_243 (O_243,N_4555,N_4528);
or UO_244 (O_244,N_4729,N_4860);
and UO_245 (O_245,N_4760,N_4542);
and UO_246 (O_246,N_4929,N_4868);
nand UO_247 (O_247,N_4575,N_4708);
nand UO_248 (O_248,N_4534,N_4775);
and UO_249 (O_249,N_4911,N_4903);
or UO_250 (O_250,N_4582,N_4961);
nand UO_251 (O_251,N_4919,N_4585);
and UO_252 (O_252,N_4853,N_4981);
or UO_253 (O_253,N_4974,N_4840);
xor UO_254 (O_254,N_4563,N_4565);
and UO_255 (O_255,N_4938,N_4960);
and UO_256 (O_256,N_4500,N_4988);
or UO_257 (O_257,N_4828,N_4829);
or UO_258 (O_258,N_4663,N_4850);
nor UO_259 (O_259,N_4813,N_4965);
nor UO_260 (O_260,N_4563,N_4799);
and UO_261 (O_261,N_4513,N_4882);
nor UO_262 (O_262,N_4786,N_4606);
nor UO_263 (O_263,N_4858,N_4924);
nor UO_264 (O_264,N_4801,N_4679);
nor UO_265 (O_265,N_4677,N_4787);
nand UO_266 (O_266,N_4696,N_4660);
xor UO_267 (O_267,N_4883,N_4566);
xor UO_268 (O_268,N_4807,N_4561);
xor UO_269 (O_269,N_4718,N_4711);
nand UO_270 (O_270,N_4834,N_4610);
or UO_271 (O_271,N_4585,N_4855);
and UO_272 (O_272,N_4705,N_4708);
or UO_273 (O_273,N_4947,N_4655);
nor UO_274 (O_274,N_4838,N_4705);
nor UO_275 (O_275,N_4576,N_4920);
and UO_276 (O_276,N_4705,N_4930);
nand UO_277 (O_277,N_4595,N_4824);
nand UO_278 (O_278,N_4961,N_4868);
and UO_279 (O_279,N_4762,N_4631);
or UO_280 (O_280,N_4842,N_4853);
nand UO_281 (O_281,N_4808,N_4605);
xor UO_282 (O_282,N_4898,N_4651);
nor UO_283 (O_283,N_4539,N_4587);
nor UO_284 (O_284,N_4654,N_4586);
nor UO_285 (O_285,N_4735,N_4675);
or UO_286 (O_286,N_4516,N_4741);
and UO_287 (O_287,N_4957,N_4720);
nor UO_288 (O_288,N_4648,N_4680);
nor UO_289 (O_289,N_4625,N_4556);
or UO_290 (O_290,N_4502,N_4635);
or UO_291 (O_291,N_4856,N_4631);
and UO_292 (O_292,N_4667,N_4790);
or UO_293 (O_293,N_4891,N_4848);
or UO_294 (O_294,N_4509,N_4622);
and UO_295 (O_295,N_4719,N_4876);
or UO_296 (O_296,N_4778,N_4886);
xor UO_297 (O_297,N_4730,N_4860);
or UO_298 (O_298,N_4910,N_4584);
nand UO_299 (O_299,N_4992,N_4540);
nand UO_300 (O_300,N_4827,N_4722);
and UO_301 (O_301,N_4627,N_4780);
nand UO_302 (O_302,N_4745,N_4865);
nand UO_303 (O_303,N_4564,N_4827);
or UO_304 (O_304,N_4873,N_4869);
or UO_305 (O_305,N_4745,N_4777);
nor UO_306 (O_306,N_4997,N_4756);
nand UO_307 (O_307,N_4586,N_4650);
nand UO_308 (O_308,N_4624,N_4765);
nor UO_309 (O_309,N_4727,N_4750);
and UO_310 (O_310,N_4830,N_4897);
or UO_311 (O_311,N_4656,N_4883);
nand UO_312 (O_312,N_4538,N_4787);
and UO_313 (O_313,N_4561,N_4727);
nand UO_314 (O_314,N_4979,N_4737);
and UO_315 (O_315,N_4841,N_4666);
or UO_316 (O_316,N_4796,N_4623);
and UO_317 (O_317,N_4711,N_4540);
nand UO_318 (O_318,N_4998,N_4763);
nand UO_319 (O_319,N_4941,N_4764);
xor UO_320 (O_320,N_4749,N_4568);
nand UO_321 (O_321,N_4858,N_4581);
nand UO_322 (O_322,N_4935,N_4816);
or UO_323 (O_323,N_4865,N_4762);
or UO_324 (O_324,N_4548,N_4583);
nand UO_325 (O_325,N_4873,N_4824);
nor UO_326 (O_326,N_4938,N_4529);
nor UO_327 (O_327,N_4873,N_4697);
or UO_328 (O_328,N_4945,N_4719);
nand UO_329 (O_329,N_4726,N_4959);
and UO_330 (O_330,N_4652,N_4830);
nor UO_331 (O_331,N_4994,N_4615);
nand UO_332 (O_332,N_4518,N_4676);
nor UO_333 (O_333,N_4654,N_4695);
nor UO_334 (O_334,N_4983,N_4591);
nor UO_335 (O_335,N_4589,N_4641);
and UO_336 (O_336,N_4964,N_4912);
nor UO_337 (O_337,N_4755,N_4861);
nor UO_338 (O_338,N_4812,N_4600);
and UO_339 (O_339,N_4574,N_4630);
nand UO_340 (O_340,N_4642,N_4962);
nand UO_341 (O_341,N_4701,N_4559);
nand UO_342 (O_342,N_4580,N_4576);
nor UO_343 (O_343,N_4927,N_4977);
nand UO_344 (O_344,N_4756,N_4975);
and UO_345 (O_345,N_4560,N_4719);
nor UO_346 (O_346,N_4669,N_4832);
nand UO_347 (O_347,N_4542,N_4955);
nand UO_348 (O_348,N_4982,N_4776);
and UO_349 (O_349,N_4949,N_4770);
nor UO_350 (O_350,N_4996,N_4934);
and UO_351 (O_351,N_4993,N_4941);
and UO_352 (O_352,N_4856,N_4784);
nand UO_353 (O_353,N_4536,N_4691);
and UO_354 (O_354,N_4599,N_4772);
nor UO_355 (O_355,N_4762,N_4788);
or UO_356 (O_356,N_4801,N_4744);
and UO_357 (O_357,N_4883,N_4827);
and UO_358 (O_358,N_4752,N_4676);
or UO_359 (O_359,N_4992,N_4841);
nand UO_360 (O_360,N_4838,N_4715);
nor UO_361 (O_361,N_4972,N_4637);
or UO_362 (O_362,N_4732,N_4935);
and UO_363 (O_363,N_4767,N_4852);
nand UO_364 (O_364,N_4817,N_4978);
and UO_365 (O_365,N_4970,N_4700);
and UO_366 (O_366,N_4568,N_4832);
nor UO_367 (O_367,N_4843,N_4541);
nand UO_368 (O_368,N_4922,N_4599);
nand UO_369 (O_369,N_4781,N_4615);
nor UO_370 (O_370,N_4922,N_4739);
or UO_371 (O_371,N_4564,N_4674);
nor UO_372 (O_372,N_4842,N_4804);
nor UO_373 (O_373,N_4862,N_4522);
and UO_374 (O_374,N_4920,N_4636);
and UO_375 (O_375,N_4616,N_4986);
nor UO_376 (O_376,N_4523,N_4854);
nor UO_377 (O_377,N_4791,N_4818);
or UO_378 (O_378,N_4747,N_4966);
and UO_379 (O_379,N_4523,N_4982);
or UO_380 (O_380,N_4507,N_4919);
or UO_381 (O_381,N_4842,N_4639);
nor UO_382 (O_382,N_4726,N_4697);
nor UO_383 (O_383,N_4999,N_4797);
nand UO_384 (O_384,N_4503,N_4653);
nand UO_385 (O_385,N_4793,N_4630);
or UO_386 (O_386,N_4643,N_4558);
nor UO_387 (O_387,N_4607,N_4512);
nand UO_388 (O_388,N_4897,N_4772);
nor UO_389 (O_389,N_4928,N_4715);
nand UO_390 (O_390,N_4765,N_4939);
and UO_391 (O_391,N_4983,N_4529);
and UO_392 (O_392,N_4541,N_4719);
nand UO_393 (O_393,N_4892,N_4803);
nor UO_394 (O_394,N_4581,N_4866);
and UO_395 (O_395,N_4988,N_4966);
xor UO_396 (O_396,N_4762,N_4813);
nor UO_397 (O_397,N_4694,N_4689);
nor UO_398 (O_398,N_4647,N_4719);
nand UO_399 (O_399,N_4632,N_4639);
and UO_400 (O_400,N_4546,N_4691);
nor UO_401 (O_401,N_4599,N_4605);
or UO_402 (O_402,N_4674,N_4933);
and UO_403 (O_403,N_4508,N_4739);
or UO_404 (O_404,N_4567,N_4797);
nand UO_405 (O_405,N_4889,N_4529);
nor UO_406 (O_406,N_4993,N_4840);
nand UO_407 (O_407,N_4559,N_4726);
nand UO_408 (O_408,N_4539,N_4970);
nor UO_409 (O_409,N_4680,N_4869);
nor UO_410 (O_410,N_4882,N_4730);
nand UO_411 (O_411,N_4577,N_4939);
or UO_412 (O_412,N_4553,N_4767);
or UO_413 (O_413,N_4740,N_4858);
or UO_414 (O_414,N_4585,N_4848);
or UO_415 (O_415,N_4919,N_4907);
xor UO_416 (O_416,N_4859,N_4844);
nand UO_417 (O_417,N_4761,N_4995);
and UO_418 (O_418,N_4753,N_4586);
and UO_419 (O_419,N_4938,N_4979);
xnor UO_420 (O_420,N_4887,N_4621);
nor UO_421 (O_421,N_4977,N_4988);
nor UO_422 (O_422,N_4889,N_4826);
or UO_423 (O_423,N_4697,N_4734);
nand UO_424 (O_424,N_4753,N_4939);
nor UO_425 (O_425,N_4810,N_4977);
xnor UO_426 (O_426,N_4749,N_4629);
and UO_427 (O_427,N_4969,N_4623);
nand UO_428 (O_428,N_4559,N_4690);
nand UO_429 (O_429,N_4633,N_4524);
nor UO_430 (O_430,N_4665,N_4594);
or UO_431 (O_431,N_4815,N_4725);
and UO_432 (O_432,N_4537,N_4589);
nor UO_433 (O_433,N_4975,N_4838);
nor UO_434 (O_434,N_4637,N_4833);
nand UO_435 (O_435,N_4568,N_4656);
and UO_436 (O_436,N_4972,N_4885);
nor UO_437 (O_437,N_4680,N_4555);
nand UO_438 (O_438,N_4999,N_4693);
nand UO_439 (O_439,N_4600,N_4867);
nor UO_440 (O_440,N_4730,N_4781);
and UO_441 (O_441,N_4889,N_4778);
nand UO_442 (O_442,N_4808,N_4921);
and UO_443 (O_443,N_4526,N_4684);
nand UO_444 (O_444,N_4569,N_4735);
nor UO_445 (O_445,N_4697,N_4645);
nor UO_446 (O_446,N_4597,N_4942);
nor UO_447 (O_447,N_4931,N_4871);
and UO_448 (O_448,N_4943,N_4762);
xnor UO_449 (O_449,N_4661,N_4562);
nand UO_450 (O_450,N_4973,N_4539);
and UO_451 (O_451,N_4734,N_4952);
or UO_452 (O_452,N_4651,N_4868);
nand UO_453 (O_453,N_4646,N_4804);
nand UO_454 (O_454,N_4904,N_4699);
and UO_455 (O_455,N_4630,N_4832);
and UO_456 (O_456,N_4529,N_4615);
nand UO_457 (O_457,N_4737,N_4780);
nor UO_458 (O_458,N_4661,N_4772);
or UO_459 (O_459,N_4822,N_4897);
nand UO_460 (O_460,N_4599,N_4951);
nor UO_461 (O_461,N_4612,N_4999);
and UO_462 (O_462,N_4875,N_4902);
nand UO_463 (O_463,N_4969,N_4602);
and UO_464 (O_464,N_4790,N_4639);
and UO_465 (O_465,N_4770,N_4571);
nand UO_466 (O_466,N_4567,N_4932);
and UO_467 (O_467,N_4517,N_4747);
nor UO_468 (O_468,N_4810,N_4803);
nor UO_469 (O_469,N_4936,N_4947);
nand UO_470 (O_470,N_4658,N_4856);
nor UO_471 (O_471,N_4521,N_4835);
or UO_472 (O_472,N_4978,N_4681);
nor UO_473 (O_473,N_4860,N_4792);
nor UO_474 (O_474,N_4759,N_4855);
or UO_475 (O_475,N_4811,N_4822);
nand UO_476 (O_476,N_4747,N_4932);
nor UO_477 (O_477,N_4830,N_4528);
nor UO_478 (O_478,N_4694,N_4628);
nor UO_479 (O_479,N_4814,N_4766);
and UO_480 (O_480,N_4633,N_4574);
or UO_481 (O_481,N_4567,N_4978);
and UO_482 (O_482,N_4997,N_4765);
nor UO_483 (O_483,N_4718,N_4562);
and UO_484 (O_484,N_4988,N_4722);
nand UO_485 (O_485,N_4547,N_4771);
nor UO_486 (O_486,N_4567,N_4606);
nand UO_487 (O_487,N_4656,N_4764);
nand UO_488 (O_488,N_4636,N_4639);
xor UO_489 (O_489,N_4635,N_4761);
and UO_490 (O_490,N_4722,N_4680);
or UO_491 (O_491,N_4714,N_4709);
xnor UO_492 (O_492,N_4627,N_4929);
or UO_493 (O_493,N_4800,N_4561);
nor UO_494 (O_494,N_4674,N_4854);
and UO_495 (O_495,N_4569,N_4793);
nand UO_496 (O_496,N_4626,N_4896);
nor UO_497 (O_497,N_4959,N_4757);
and UO_498 (O_498,N_4916,N_4658);
or UO_499 (O_499,N_4696,N_4551);
and UO_500 (O_500,N_4882,N_4640);
nor UO_501 (O_501,N_4503,N_4559);
or UO_502 (O_502,N_4853,N_4792);
nand UO_503 (O_503,N_4655,N_4768);
and UO_504 (O_504,N_4558,N_4765);
nand UO_505 (O_505,N_4578,N_4539);
nor UO_506 (O_506,N_4740,N_4737);
nor UO_507 (O_507,N_4859,N_4539);
nand UO_508 (O_508,N_4975,N_4963);
nor UO_509 (O_509,N_4653,N_4954);
nor UO_510 (O_510,N_4537,N_4927);
nand UO_511 (O_511,N_4658,N_4623);
nor UO_512 (O_512,N_4655,N_4987);
and UO_513 (O_513,N_4894,N_4861);
nor UO_514 (O_514,N_4892,N_4773);
nand UO_515 (O_515,N_4768,N_4514);
nor UO_516 (O_516,N_4556,N_4743);
nand UO_517 (O_517,N_4789,N_4881);
nor UO_518 (O_518,N_4662,N_4538);
nand UO_519 (O_519,N_4964,N_4875);
or UO_520 (O_520,N_4583,N_4912);
nand UO_521 (O_521,N_4623,N_4555);
or UO_522 (O_522,N_4503,N_4605);
or UO_523 (O_523,N_4871,N_4653);
or UO_524 (O_524,N_4688,N_4886);
or UO_525 (O_525,N_4578,N_4543);
and UO_526 (O_526,N_4937,N_4689);
nand UO_527 (O_527,N_4667,N_4522);
nand UO_528 (O_528,N_4587,N_4788);
xor UO_529 (O_529,N_4618,N_4860);
nor UO_530 (O_530,N_4946,N_4934);
nor UO_531 (O_531,N_4705,N_4852);
nor UO_532 (O_532,N_4594,N_4886);
or UO_533 (O_533,N_4766,N_4850);
nand UO_534 (O_534,N_4602,N_4533);
or UO_535 (O_535,N_4905,N_4509);
nor UO_536 (O_536,N_4826,N_4747);
or UO_537 (O_537,N_4502,N_4767);
nand UO_538 (O_538,N_4796,N_4567);
and UO_539 (O_539,N_4772,N_4873);
nor UO_540 (O_540,N_4829,N_4677);
or UO_541 (O_541,N_4722,N_4773);
nand UO_542 (O_542,N_4733,N_4516);
or UO_543 (O_543,N_4640,N_4791);
and UO_544 (O_544,N_4789,N_4721);
or UO_545 (O_545,N_4752,N_4640);
nand UO_546 (O_546,N_4858,N_4631);
and UO_547 (O_547,N_4783,N_4635);
or UO_548 (O_548,N_4530,N_4566);
and UO_549 (O_549,N_4693,N_4775);
or UO_550 (O_550,N_4568,N_4933);
nand UO_551 (O_551,N_4769,N_4535);
or UO_552 (O_552,N_4555,N_4777);
and UO_553 (O_553,N_4743,N_4924);
nand UO_554 (O_554,N_4518,N_4673);
nor UO_555 (O_555,N_4964,N_4670);
or UO_556 (O_556,N_4584,N_4978);
or UO_557 (O_557,N_4634,N_4615);
and UO_558 (O_558,N_4552,N_4740);
nor UO_559 (O_559,N_4909,N_4541);
nor UO_560 (O_560,N_4599,N_4654);
nand UO_561 (O_561,N_4929,N_4752);
or UO_562 (O_562,N_4796,N_4898);
nand UO_563 (O_563,N_4972,N_4750);
nor UO_564 (O_564,N_4837,N_4712);
nor UO_565 (O_565,N_4925,N_4733);
or UO_566 (O_566,N_4518,N_4910);
and UO_567 (O_567,N_4958,N_4897);
nand UO_568 (O_568,N_4668,N_4978);
nor UO_569 (O_569,N_4837,N_4685);
nor UO_570 (O_570,N_4982,N_4695);
nand UO_571 (O_571,N_4711,N_4623);
nor UO_572 (O_572,N_4650,N_4537);
nor UO_573 (O_573,N_4732,N_4906);
nand UO_574 (O_574,N_4566,N_4573);
nand UO_575 (O_575,N_4694,N_4912);
and UO_576 (O_576,N_4712,N_4668);
and UO_577 (O_577,N_4554,N_4878);
and UO_578 (O_578,N_4841,N_4872);
nor UO_579 (O_579,N_4626,N_4977);
nor UO_580 (O_580,N_4599,N_4985);
nor UO_581 (O_581,N_4501,N_4912);
or UO_582 (O_582,N_4726,N_4609);
or UO_583 (O_583,N_4965,N_4611);
and UO_584 (O_584,N_4904,N_4735);
nand UO_585 (O_585,N_4675,N_4538);
nand UO_586 (O_586,N_4530,N_4760);
xnor UO_587 (O_587,N_4681,N_4807);
or UO_588 (O_588,N_4698,N_4707);
nor UO_589 (O_589,N_4563,N_4886);
nand UO_590 (O_590,N_4685,N_4714);
nor UO_591 (O_591,N_4824,N_4532);
and UO_592 (O_592,N_4972,N_4514);
or UO_593 (O_593,N_4836,N_4902);
nand UO_594 (O_594,N_4546,N_4536);
or UO_595 (O_595,N_4976,N_4999);
or UO_596 (O_596,N_4773,N_4508);
and UO_597 (O_597,N_4945,N_4675);
nand UO_598 (O_598,N_4992,N_4885);
nor UO_599 (O_599,N_4970,N_4503);
or UO_600 (O_600,N_4839,N_4710);
nand UO_601 (O_601,N_4527,N_4649);
nor UO_602 (O_602,N_4847,N_4643);
or UO_603 (O_603,N_4884,N_4716);
or UO_604 (O_604,N_4544,N_4605);
nand UO_605 (O_605,N_4562,N_4949);
nor UO_606 (O_606,N_4898,N_4730);
nand UO_607 (O_607,N_4904,N_4868);
nand UO_608 (O_608,N_4507,N_4560);
nand UO_609 (O_609,N_4520,N_4751);
or UO_610 (O_610,N_4925,N_4649);
or UO_611 (O_611,N_4979,N_4631);
nor UO_612 (O_612,N_4841,N_4879);
and UO_613 (O_613,N_4897,N_4847);
and UO_614 (O_614,N_4615,N_4644);
and UO_615 (O_615,N_4889,N_4554);
and UO_616 (O_616,N_4697,N_4609);
nor UO_617 (O_617,N_4874,N_4715);
and UO_618 (O_618,N_4859,N_4722);
nor UO_619 (O_619,N_4502,N_4994);
or UO_620 (O_620,N_4813,N_4854);
and UO_621 (O_621,N_4824,N_4759);
nand UO_622 (O_622,N_4553,N_4799);
or UO_623 (O_623,N_4806,N_4575);
nor UO_624 (O_624,N_4672,N_4754);
nand UO_625 (O_625,N_4626,N_4800);
and UO_626 (O_626,N_4992,N_4895);
nor UO_627 (O_627,N_4757,N_4750);
nand UO_628 (O_628,N_4501,N_4706);
nor UO_629 (O_629,N_4779,N_4954);
and UO_630 (O_630,N_4727,N_4947);
nand UO_631 (O_631,N_4669,N_4985);
nor UO_632 (O_632,N_4880,N_4996);
and UO_633 (O_633,N_4807,N_4704);
nand UO_634 (O_634,N_4620,N_4576);
and UO_635 (O_635,N_4889,N_4820);
nand UO_636 (O_636,N_4896,N_4934);
or UO_637 (O_637,N_4804,N_4641);
or UO_638 (O_638,N_4809,N_4946);
or UO_639 (O_639,N_4972,N_4827);
xnor UO_640 (O_640,N_4853,N_4807);
or UO_641 (O_641,N_4632,N_4702);
nand UO_642 (O_642,N_4638,N_4937);
xnor UO_643 (O_643,N_4826,N_4727);
or UO_644 (O_644,N_4833,N_4916);
and UO_645 (O_645,N_4614,N_4864);
and UO_646 (O_646,N_4618,N_4953);
nand UO_647 (O_647,N_4793,N_4703);
nand UO_648 (O_648,N_4582,N_4788);
nor UO_649 (O_649,N_4884,N_4766);
and UO_650 (O_650,N_4828,N_4703);
nor UO_651 (O_651,N_4819,N_4709);
and UO_652 (O_652,N_4804,N_4909);
and UO_653 (O_653,N_4645,N_4503);
nand UO_654 (O_654,N_4975,N_4930);
or UO_655 (O_655,N_4941,N_4802);
or UO_656 (O_656,N_4636,N_4811);
nand UO_657 (O_657,N_4624,N_4691);
or UO_658 (O_658,N_4691,N_4556);
nand UO_659 (O_659,N_4700,N_4771);
nand UO_660 (O_660,N_4996,N_4855);
nor UO_661 (O_661,N_4619,N_4868);
nor UO_662 (O_662,N_4847,N_4956);
or UO_663 (O_663,N_4843,N_4979);
nor UO_664 (O_664,N_4860,N_4731);
and UO_665 (O_665,N_4913,N_4908);
or UO_666 (O_666,N_4815,N_4624);
or UO_667 (O_667,N_4507,N_4513);
nor UO_668 (O_668,N_4923,N_4943);
nor UO_669 (O_669,N_4816,N_4784);
or UO_670 (O_670,N_4791,N_4785);
nand UO_671 (O_671,N_4775,N_4864);
and UO_672 (O_672,N_4584,N_4671);
nor UO_673 (O_673,N_4604,N_4705);
nor UO_674 (O_674,N_4693,N_4666);
or UO_675 (O_675,N_4615,N_4895);
or UO_676 (O_676,N_4612,N_4903);
nor UO_677 (O_677,N_4606,N_4648);
and UO_678 (O_678,N_4671,N_4524);
nand UO_679 (O_679,N_4858,N_4951);
and UO_680 (O_680,N_4700,N_4960);
or UO_681 (O_681,N_4805,N_4920);
or UO_682 (O_682,N_4680,N_4848);
nand UO_683 (O_683,N_4711,N_4924);
nand UO_684 (O_684,N_4516,N_4973);
and UO_685 (O_685,N_4874,N_4997);
nand UO_686 (O_686,N_4904,N_4665);
or UO_687 (O_687,N_4602,N_4525);
nor UO_688 (O_688,N_4995,N_4556);
and UO_689 (O_689,N_4994,N_4799);
and UO_690 (O_690,N_4523,N_4626);
nand UO_691 (O_691,N_4934,N_4625);
or UO_692 (O_692,N_4802,N_4706);
and UO_693 (O_693,N_4707,N_4953);
or UO_694 (O_694,N_4770,N_4745);
nand UO_695 (O_695,N_4877,N_4589);
nand UO_696 (O_696,N_4523,N_4896);
nor UO_697 (O_697,N_4679,N_4559);
nor UO_698 (O_698,N_4914,N_4841);
nand UO_699 (O_699,N_4647,N_4829);
or UO_700 (O_700,N_4889,N_4965);
or UO_701 (O_701,N_4685,N_4859);
nor UO_702 (O_702,N_4938,N_4972);
nor UO_703 (O_703,N_4797,N_4966);
and UO_704 (O_704,N_4974,N_4737);
or UO_705 (O_705,N_4800,N_4607);
nor UO_706 (O_706,N_4979,N_4939);
or UO_707 (O_707,N_4769,N_4654);
and UO_708 (O_708,N_4981,N_4661);
or UO_709 (O_709,N_4909,N_4691);
or UO_710 (O_710,N_4793,N_4735);
xor UO_711 (O_711,N_4504,N_4664);
and UO_712 (O_712,N_4548,N_4626);
nand UO_713 (O_713,N_4535,N_4801);
nor UO_714 (O_714,N_4762,N_4843);
nor UO_715 (O_715,N_4801,N_4938);
nor UO_716 (O_716,N_4514,N_4906);
nand UO_717 (O_717,N_4711,N_4659);
or UO_718 (O_718,N_4854,N_4500);
and UO_719 (O_719,N_4675,N_4713);
and UO_720 (O_720,N_4725,N_4503);
or UO_721 (O_721,N_4586,N_4799);
or UO_722 (O_722,N_4613,N_4686);
nand UO_723 (O_723,N_4837,N_4640);
nand UO_724 (O_724,N_4801,N_4641);
or UO_725 (O_725,N_4946,N_4838);
or UO_726 (O_726,N_4892,N_4864);
nand UO_727 (O_727,N_4500,N_4705);
and UO_728 (O_728,N_4600,N_4783);
and UO_729 (O_729,N_4666,N_4572);
or UO_730 (O_730,N_4946,N_4547);
or UO_731 (O_731,N_4712,N_4748);
or UO_732 (O_732,N_4961,N_4626);
nand UO_733 (O_733,N_4989,N_4541);
and UO_734 (O_734,N_4570,N_4500);
nand UO_735 (O_735,N_4671,N_4548);
and UO_736 (O_736,N_4888,N_4987);
and UO_737 (O_737,N_4993,N_4666);
nand UO_738 (O_738,N_4686,N_4528);
nand UO_739 (O_739,N_4796,N_4577);
nor UO_740 (O_740,N_4710,N_4587);
xnor UO_741 (O_741,N_4932,N_4862);
nor UO_742 (O_742,N_4767,N_4643);
xnor UO_743 (O_743,N_4640,N_4503);
or UO_744 (O_744,N_4801,N_4663);
nand UO_745 (O_745,N_4639,N_4606);
and UO_746 (O_746,N_4516,N_4856);
and UO_747 (O_747,N_4898,N_4866);
nor UO_748 (O_748,N_4578,N_4694);
nand UO_749 (O_749,N_4576,N_4761);
nor UO_750 (O_750,N_4577,N_4895);
nor UO_751 (O_751,N_4512,N_4513);
and UO_752 (O_752,N_4803,N_4670);
and UO_753 (O_753,N_4572,N_4704);
or UO_754 (O_754,N_4668,N_4803);
nor UO_755 (O_755,N_4878,N_4785);
or UO_756 (O_756,N_4923,N_4671);
and UO_757 (O_757,N_4508,N_4613);
nand UO_758 (O_758,N_4627,N_4935);
and UO_759 (O_759,N_4567,N_4585);
and UO_760 (O_760,N_4754,N_4896);
and UO_761 (O_761,N_4648,N_4850);
and UO_762 (O_762,N_4871,N_4701);
xnor UO_763 (O_763,N_4765,N_4754);
nor UO_764 (O_764,N_4718,N_4783);
and UO_765 (O_765,N_4603,N_4610);
or UO_766 (O_766,N_4558,N_4748);
nor UO_767 (O_767,N_4957,N_4608);
nand UO_768 (O_768,N_4594,N_4915);
or UO_769 (O_769,N_4741,N_4894);
nand UO_770 (O_770,N_4687,N_4932);
or UO_771 (O_771,N_4843,N_4857);
nor UO_772 (O_772,N_4679,N_4787);
nor UO_773 (O_773,N_4694,N_4817);
or UO_774 (O_774,N_4955,N_4613);
nand UO_775 (O_775,N_4764,N_4618);
and UO_776 (O_776,N_4639,N_4756);
and UO_777 (O_777,N_4797,N_4731);
nor UO_778 (O_778,N_4982,N_4723);
nand UO_779 (O_779,N_4911,N_4730);
nand UO_780 (O_780,N_4907,N_4624);
and UO_781 (O_781,N_4699,N_4914);
or UO_782 (O_782,N_4986,N_4647);
and UO_783 (O_783,N_4990,N_4641);
and UO_784 (O_784,N_4967,N_4527);
and UO_785 (O_785,N_4900,N_4891);
nand UO_786 (O_786,N_4711,N_4527);
and UO_787 (O_787,N_4902,N_4571);
or UO_788 (O_788,N_4769,N_4812);
nand UO_789 (O_789,N_4722,N_4615);
or UO_790 (O_790,N_4912,N_4995);
nand UO_791 (O_791,N_4612,N_4856);
and UO_792 (O_792,N_4914,N_4884);
xor UO_793 (O_793,N_4529,N_4885);
nand UO_794 (O_794,N_4584,N_4531);
and UO_795 (O_795,N_4535,N_4533);
nor UO_796 (O_796,N_4861,N_4942);
nor UO_797 (O_797,N_4844,N_4862);
nand UO_798 (O_798,N_4730,N_4994);
or UO_799 (O_799,N_4682,N_4502);
or UO_800 (O_800,N_4990,N_4772);
nand UO_801 (O_801,N_4911,N_4974);
and UO_802 (O_802,N_4541,N_4587);
xor UO_803 (O_803,N_4806,N_4839);
nor UO_804 (O_804,N_4671,N_4624);
and UO_805 (O_805,N_4879,N_4885);
nand UO_806 (O_806,N_4970,N_4811);
nor UO_807 (O_807,N_4936,N_4774);
nand UO_808 (O_808,N_4592,N_4795);
or UO_809 (O_809,N_4534,N_4682);
nor UO_810 (O_810,N_4917,N_4828);
nand UO_811 (O_811,N_4589,N_4817);
nand UO_812 (O_812,N_4527,N_4546);
and UO_813 (O_813,N_4523,N_4827);
or UO_814 (O_814,N_4896,N_4839);
nand UO_815 (O_815,N_4864,N_4587);
nor UO_816 (O_816,N_4719,N_4584);
and UO_817 (O_817,N_4646,N_4766);
nand UO_818 (O_818,N_4742,N_4758);
or UO_819 (O_819,N_4919,N_4980);
and UO_820 (O_820,N_4943,N_4803);
or UO_821 (O_821,N_4840,N_4942);
nand UO_822 (O_822,N_4529,N_4537);
or UO_823 (O_823,N_4759,N_4501);
or UO_824 (O_824,N_4575,N_4865);
and UO_825 (O_825,N_4948,N_4783);
nor UO_826 (O_826,N_4531,N_4654);
or UO_827 (O_827,N_4929,N_4592);
or UO_828 (O_828,N_4738,N_4672);
nor UO_829 (O_829,N_4880,N_4707);
nor UO_830 (O_830,N_4723,N_4520);
nand UO_831 (O_831,N_4763,N_4915);
nand UO_832 (O_832,N_4936,N_4941);
and UO_833 (O_833,N_4927,N_4953);
or UO_834 (O_834,N_4534,N_4956);
or UO_835 (O_835,N_4719,N_4531);
and UO_836 (O_836,N_4965,N_4549);
or UO_837 (O_837,N_4717,N_4801);
nand UO_838 (O_838,N_4980,N_4735);
nor UO_839 (O_839,N_4868,N_4957);
nor UO_840 (O_840,N_4920,N_4881);
nor UO_841 (O_841,N_4664,N_4974);
nand UO_842 (O_842,N_4591,N_4970);
and UO_843 (O_843,N_4543,N_4940);
and UO_844 (O_844,N_4580,N_4703);
nor UO_845 (O_845,N_4705,N_4791);
or UO_846 (O_846,N_4791,N_4707);
or UO_847 (O_847,N_4851,N_4853);
nand UO_848 (O_848,N_4903,N_4845);
nand UO_849 (O_849,N_4987,N_4986);
nor UO_850 (O_850,N_4813,N_4667);
nor UO_851 (O_851,N_4515,N_4901);
xor UO_852 (O_852,N_4707,N_4580);
nor UO_853 (O_853,N_4811,N_4530);
and UO_854 (O_854,N_4746,N_4989);
nand UO_855 (O_855,N_4839,N_4632);
or UO_856 (O_856,N_4594,N_4923);
or UO_857 (O_857,N_4899,N_4761);
nand UO_858 (O_858,N_4971,N_4803);
or UO_859 (O_859,N_4892,N_4841);
nor UO_860 (O_860,N_4847,N_4757);
nand UO_861 (O_861,N_4700,N_4553);
and UO_862 (O_862,N_4616,N_4621);
or UO_863 (O_863,N_4510,N_4600);
or UO_864 (O_864,N_4946,N_4585);
xor UO_865 (O_865,N_4867,N_4816);
nor UO_866 (O_866,N_4913,N_4592);
nor UO_867 (O_867,N_4759,N_4544);
or UO_868 (O_868,N_4826,N_4709);
nor UO_869 (O_869,N_4625,N_4776);
and UO_870 (O_870,N_4683,N_4991);
nor UO_871 (O_871,N_4558,N_4636);
and UO_872 (O_872,N_4632,N_4522);
nor UO_873 (O_873,N_4777,N_4847);
and UO_874 (O_874,N_4700,N_4506);
and UO_875 (O_875,N_4937,N_4625);
or UO_876 (O_876,N_4609,N_4629);
nand UO_877 (O_877,N_4846,N_4865);
xnor UO_878 (O_878,N_4665,N_4791);
or UO_879 (O_879,N_4958,N_4571);
or UO_880 (O_880,N_4632,N_4538);
or UO_881 (O_881,N_4944,N_4886);
or UO_882 (O_882,N_4619,N_4550);
nor UO_883 (O_883,N_4920,N_4831);
nand UO_884 (O_884,N_4557,N_4509);
and UO_885 (O_885,N_4737,N_4755);
nand UO_886 (O_886,N_4771,N_4974);
nor UO_887 (O_887,N_4853,N_4542);
or UO_888 (O_888,N_4679,N_4589);
nand UO_889 (O_889,N_4796,N_4654);
and UO_890 (O_890,N_4555,N_4605);
nor UO_891 (O_891,N_4602,N_4975);
nand UO_892 (O_892,N_4590,N_4851);
nand UO_893 (O_893,N_4789,N_4685);
nand UO_894 (O_894,N_4863,N_4829);
nor UO_895 (O_895,N_4958,N_4819);
and UO_896 (O_896,N_4751,N_4533);
or UO_897 (O_897,N_4641,N_4856);
and UO_898 (O_898,N_4964,N_4660);
nor UO_899 (O_899,N_4880,N_4833);
nor UO_900 (O_900,N_4920,N_4808);
nor UO_901 (O_901,N_4733,N_4673);
and UO_902 (O_902,N_4715,N_4542);
nor UO_903 (O_903,N_4735,N_4850);
xor UO_904 (O_904,N_4513,N_4912);
or UO_905 (O_905,N_4584,N_4705);
nor UO_906 (O_906,N_4550,N_4696);
nand UO_907 (O_907,N_4695,N_4914);
and UO_908 (O_908,N_4677,N_4673);
nor UO_909 (O_909,N_4864,N_4774);
or UO_910 (O_910,N_4559,N_4785);
nor UO_911 (O_911,N_4735,N_4859);
or UO_912 (O_912,N_4805,N_4847);
nor UO_913 (O_913,N_4588,N_4755);
and UO_914 (O_914,N_4841,N_4681);
or UO_915 (O_915,N_4646,N_4740);
and UO_916 (O_916,N_4685,N_4936);
and UO_917 (O_917,N_4645,N_4891);
and UO_918 (O_918,N_4890,N_4515);
nand UO_919 (O_919,N_4518,N_4688);
nand UO_920 (O_920,N_4853,N_4564);
or UO_921 (O_921,N_4636,N_4619);
or UO_922 (O_922,N_4737,N_4870);
nor UO_923 (O_923,N_4687,N_4988);
nand UO_924 (O_924,N_4637,N_4985);
and UO_925 (O_925,N_4937,N_4912);
and UO_926 (O_926,N_4852,N_4509);
nand UO_927 (O_927,N_4702,N_4708);
and UO_928 (O_928,N_4526,N_4767);
or UO_929 (O_929,N_4694,N_4796);
nand UO_930 (O_930,N_4858,N_4526);
nor UO_931 (O_931,N_4587,N_4564);
nand UO_932 (O_932,N_4998,N_4507);
or UO_933 (O_933,N_4732,N_4698);
xor UO_934 (O_934,N_4858,N_4929);
nand UO_935 (O_935,N_4570,N_4600);
nor UO_936 (O_936,N_4601,N_4690);
or UO_937 (O_937,N_4869,N_4615);
or UO_938 (O_938,N_4752,N_4610);
nand UO_939 (O_939,N_4736,N_4789);
or UO_940 (O_940,N_4533,N_4571);
nand UO_941 (O_941,N_4784,N_4797);
nand UO_942 (O_942,N_4505,N_4772);
nor UO_943 (O_943,N_4520,N_4640);
and UO_944 (O_944,N_4555,N_4951);
or UO_945 (O_945,N_4767,N_4999);
and UO_946 (O_946,N_4638,N_4783);
and UO_947 (O_947,N_4988,N_4823);
nand UO_948 (O_948,N_4562,N_4557);
nor UO_949 (O_949,N_4534,N_4504);
nor UO_950 (O_950,N_4582,N_4668);
nand UO_951 (O_951,N_4909,N_4900);
nand UO_952 (O_952,N_4794,N_4588);
nor UO_953 (O_953,N_4760,N_4600);
or UO_954 (O_954,N_4506,N_4789);
nand UO_955 (O_955,N_4546,N_4588);
and UO_956 (O_956,N_4711,N_4910);
nor UO_957 (O_957,N_4893,N_4917);
nor UO_958 (O_958,N_4723,N_4803);
and UO_959 (O_959,N_4571,N_4823);
or UO_960 (O_960,N_4693,N_4521);
and UO_961 (O_961,N_4665,N_4854);
nand UO_962 (O_962,N_4897,N_4981);
nand UO_963 (O_963,N_4507,N_4631);
and UO_964 (O_964,N_4967,N_4873);
nor UO_965 (O_965,N_4976,N_4606);
or UO_966 (O_966,N_4657,N_4964);
nor UO_967 (O_967,N_4585,N_4554);
xnor UO_968 (O_968,N_4612,N_4878);
and UO_969 (O_969,N_4793,N_4694);
nor UO_970 (O_970,N_4821,N_4818);
or UO_971 (O_971,N_4517,N_4550);
nor UO_972 (O_972,N_4677,N_4649);
nor UO_973 (O_973,N_4518,N_4571);
nand UO_974 (O_974,N_4556,N_4684);
nand UO_975 (O_975,N_4952,N_4903);
nand UO_976 (O_976,N_4894,N_4892);
or UO_977 (O_977,N_4927,N_4617);
nor UO_978 (O_978,N_4968,N_4846);
and UO_979 (O_979,N_4935,N_4537);
nand UO_980 (O_980,N_4680,N_4902);
or UO_981 (O_981,N_4896,N_4909);
or UO_982 (O_982,N_4784,N_4502);
nand UO_983 (O_983,N_4922,N_4844);
nand UO_984 (O_984,N_4938,N_4929);
or UO_985 (O_985,N_4763,N_4700);
nand UO_986 (O_986,N_4730,N_4877);
and UO_987 (O_987,N_4947,N_4814);
nor UO_988 (O_988,N_4564,N_4943);
or UO_989 (O_989,N_4604,N_4798);
and UO_990 (O_990,N_4604,N_4829);
nand UO_991 (O_991,N_4718,N_4732);
or UO_992 (O_992,N_4623,N_4583);
and UO_993 (O_993,N_4775,N_4582);
nor UO_994 (O_994,N_4529,N_4543);
nor UO_995 (O_995,N_4591,N_4879);
or UO_996 (O_996,N_4846,N_4561);
or UO_997 (O_997,N_4925,N_4667);
or UO_998 (O_998,N_4584,N_4536);
or UO_999 (O_999,N_4513,N_4689);
endmodule