module basic_750_5000_1000_2_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2504,N_2505,N_2506,N_2507,N_2509,N_2510,N_2511,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2523,N_2524,N_2525,N_2526,N_2527,N_2529,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2538,N_2539,N_2540,N_2542,N_2543,N_2544,N_2546,N_2547,N_2548,N_2549,N_2552,N_2553,N_2554,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2600,N_2601,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2626,N_2628,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2648,N_2649,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2662,N_2663,N_2664,N_2665,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2676,N_2677,N_2678,N_2679,N_2681,N_2682,N_2683,N_2685,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2694,N_2695,N_2697,N_2699,N_2700,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2711,N_2712,N_2713,N_2714,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2724,N_2726,N_2727,N_2728,N_2730,N_2732,N_2733,N_2734,N_2735,N_2736,N_2738,N_2739,N_2740,N_2741,N_2743,N_2744,N_2745,N_2749,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2768,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2778,N_2779,N_2780,N_2781,N_2782,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2827,N_2828,N_2829,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2839,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2849,N_2850,N_2851,N_2852,N_2853,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2876,N_2878,N_2879,N_2880,N_2882,N_2885,N_2886,N_2888,N_2889,N_2890,N_2891,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2912,N_2913,N_2914,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2925,N_2927,N_2928,N_2929,N_2930,N_2933,N_2934,N_2935,N_2939,N_2941,N_2943,N_2945,N_2946,N_2947,N_2948,N_2951,N_2952,N_2953,N_2955,N_2956,N_2957,N_2958,N_2959,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2984,N_2987,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2999,N_3000,N_3001,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3021,N_3022,N_3023,N_3024,N_3026,N_3028,N_3029,N_3030,N_3033,N_3034,N_3035,N_3036,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3054,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3075,N_3076,N_3078,N_3079,N_3081,N_3083,N_3085,N_3087,N_3088,N_3090,N_3091,N_3092,N_3093,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3106,N_3108,N_3109,N_3110,N_3111,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3121,N_3122,N_3124,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3155,N_3157,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3168,N_3169,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3190,N_3191,N_3192,N_3193,N_3194,N_3196,N_3197,N_3198,N_3199,N_3200,N_3202,N_3204,N_3205,N_3206,N_3207,N_3208,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3226,N_3227,N_3228,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3311,N_3312,N_3313,N_3315,N_3317,N_3319,N_3320,N_3321,N_3323,N_3325,N_3326,N_3327,N_3328,N_3330,N_3331,N_3333,N_3334,N_3335,N_3336,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3363,N_3364,N_3365,N_3366,N_3367,N_3370,N_3371,N_3372,N_3373,N_3374,N_3376,N_3377,N_3378,N_3379,N_3380,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3392,N_3393,N_3394,N_3395,N_3397,N_3398,N_3399,N_3401,N_3402,N_3403,N_3404,N_3405,N_3408,N_3409,N_3412,N_3413,N_3414,N_3415,N_3416,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3435,N_3436,N_3438,N_3439,N_3440,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3481,N_3482,N_3483,N_3484,N_3485,N_3487,N_3488,N_3489,N_3490,N_3491,N_3493,N_3494,N_3495,N_3496,N_3497,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3506,N_3507,N_3508,N_3513,N_3514,N_3515,N_3516,N_3517,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3527,N_3528,N_3529,N_3531,N_3534,N_3535,N_3537,N_3538,N_3539,N_3540,N_3542,N_3543,N_3544,N_3545,N_3548,N_3549,N_3550,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3564,N_3565,N_3566,N_3567,N_3568,N_3571,N_3572,N_3573,N_3574,N_3575,N_3577,N_3578,N_3579,N_3580,N_3582,N_3583,N_3584,N_3586,N_3587,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3601,N_3602,N_3604,N_3605,N_3606,N_3608,N_3609,N_3610,N_3611,N_3613,N_3614,N_3615,N_3616,N_3620,N_3623,N_3624,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3653,N_3654,N_3655,N_3656,N_3658,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3667,N_3668,N_3672,N_3673,N_3674,N_3676,N_3678,N_3679,N_3681,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3692,N_3693,N_3694,N_3695,N_3697,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3724,N_3725,N_3726,N_3727,N_3729,N_3733,N_3734,N_3736,N_3737,N_3738,N_3739,N_3743,N_3744,N_3745,N_3746,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3757,N_3758,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3773,N_3774,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3783,N_3784,N_3785,N_3786,N_3787,N_3789,N_3791,N_3792,N_3793,N_3794,N_3795,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3809,N_3810,N_3811,N_3813,N_3814,N_3815,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3824,N_3826,N_3828,N_3829,N_3830,N_3831,N_3833,N_3834,N_3835,N_3837,N_3838,N_3839,N_3840,N_3842,N_3844,N_3845,N_3847,N_3848,N_3849,N_3850,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3861,N_3862,N_3864,N_3865,N_3866,N_3867,N_3868,N_3870,N_3871,N_3872,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3883,N_3884,N_3887,N_3888,N_3890,N_3891,N_3892,N_3893,N_3895,N_3896,N_3897,N_3898,N_3899,N_3903,N_3904,N_3905,N_3906,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3920,N_3921,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3943,N_3944,N_3945,N_3946,N_3949,N_3950,N_3951,N_3953,N_3954,N_3955,N_3956,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3991,N_3992,N_3994,N_3995,N_3996,N_3997,N_3998,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4021,N_4022,N_4023,N_4024,N_4025,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4049,N_4050,N_4051,N_4052,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4072,N_4073,N_4075,N_4077,N_4080,N_4082,N_4083,N_4084,N_4085,N_4086,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4096,N_4097,N_4098,N_4101,N_4102,N_4103,N_4105,N_4106,N_4107,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4122,N_4123,N_4124,N_4125,N_4128,N_4129,N_4130,N_4132,N_4133,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4143,N_4144,N_4146,N_4147,N_4148,N_4149,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4164,N_4166,N_4167,N_4168,N_4169,N_4170,N_4173,N_4174,N_4176,N_4178,N_4179,N_4180,N_4181,N_4182,N_4184,N_4185,N_4186,N_4188,N_4190,N_4193,N_4194,N_4196,N_4197,N_4198,N_4199,N_4200,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4213,N_4214,N_4215,N_4218,N_4219,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4228,N_4229,N_4231,N_4232,N_4233,N_4234,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4254,N_4255,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4285,N_4286,N_4287,N_4288,N_4289,N_4291,N_4292,N_4293,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4321,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4335,N_4337,N_4338,N_4340,N_4341,N_4342,N_4345,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4374,N_4375,N_4376,N_4377,N_4379,N_4380,N_4381,N_4382,N_4384,N_4385,N_4386,N_4388,N_4390,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4401,N_4402,N_4403,N_4404,N_4405,N_4408,N_4409,N_4410,N_4411,N_4412,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4421,N_4422,N_4423,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4460,N_4462,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4483,N_4484,N_4485,N_4487,N_4488,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4499,N_4500,N_4502,N_4504,N_4505,N_4507,N_4509,N_4510,N_4511,N_4512,N_4514,N_4515,N_4516,N_4517,N_4518,N_4520,N_4521,N_4522,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4534,N_4535,N_4536,N_4538,N_4539,N_4540,N_4542,N_4543,N_4544,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4569,N_4570,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4583,N_4584,N_4586,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4617,N_4618,N_4619,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4633,N_4634,N_4635,N_4636,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4659,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4717,N_4718,N_4720,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4731,N_4732,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4750,N_4751,N_4753,N_4754,N_4756,N_4757,N_4758,N_4759,N_4760,N_4762,N_4763,N_4766,N_4768,N_4769,N_4770,N_4771,N_4773,N_4774,N_4776,N_4778,N_4779,N_4780,N_4782,N_4784,N_4786,N_4787,N_4788,N_4789,N_4790,N_4792,N_4795,N_4796,N_4797,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4809,N_4810,N_4811,N_4812,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4822,N_4823,N_4824,N_4825,N_4827,N_4828,N_4829,N_4830,N_4832,N_4834,N_4835,N_4838,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4864,N_4865,N_4868,N_4869,N_4870,N_4872,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4881,N_4882,N_4883,N_4886,N_4887,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4908,N_4910,N_4913,N_4914,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4949,N_4952,N_4953,N_4955,N_4956,N_4957,N_4960,N_4961,N_4962,N_4963,N_4964,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4975,N_4976,N_4977,N_4978,N_4982,N_4983,N_4984,N_4986,N_4987,N_4989,N_4990,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997;
or U0 (N_0,In_162,In_676);
nor U1 (N_1,In_576,In_43);
and U2 (N_2,In_595,In_610);
nand U3 (N_3,In_195,In_149);
and U4 (N_4,In_292,In_56);
and U5 (N_5,In_244,In_531);
nor U6 (N_6,In_142,In_358);
nor U7 (N_7,In_689,In_287);
nand U8 (N_8,In_50,In_713);
or U9 (N_9,In_667,In_49);
and U10 (N_10,In_746,In_282);
or U11 (N_11,In_410,In_550);
or U12 (N_12,In_545,In_7);
xnor U13 (N_13,In_202,In_293);
nor U14 (N_14,In_328,In_4);
xnor U15 (N_15,In_586,In_183);
nand U16 (N_16,In_106,In_38);
and U17 (N_17,In_716,In_683);
nand U18 (N_18,In_724,In_647);
and U19 (N_19,In_53,In_267);
nor U20 (N_20,In_290,In_416);
and U21 (N_21,In_268,In_294);
or U22 (N_22,In_697,In_568);
and U23 (N_23,In_632,In_74);
and U24 (N_24,In_216,In_366);
nor U25 (N_25,In_34,In_717);
or U26 (N_26,In_318,In_602);
or U27 (N_27,In_609,In_289);
nor U28 (N_28,In_262,In_670);
and U29 (N_29,In_377,In_515);
nor U30 (N_30,In_574,In_329);
xor U31 (N_31,In_508,In_370);
or U32 (N_32,In_728,In_68);
nor U33 (N_33,In_415,In_431);
and U34 (N_34,In_529,In_107);
and U35 (N_35,In_631,In_427);
or U36 (N_36,In_10,In_198);
and U37 (N_37,In_348,In_164);
or U38 (N_38,In_743,In_354);
nor U39 (N_39,In_503,In_692);
xnor U40 (N_40,In_448,In_662);
nand U41 (N_41,In_365,In_691);
or U42 (N_42,In_470,In_19);
nand U43 (N_43,In_710,In_690);
nand U44 (N_44,In_501,In_133);
xor U45 (N_45,In_606,In_104);
nor U46 (N_46,In_234,In_35);
and U47 (N_47,In_32,In_89);
and U48 (N_48,In_504,In_205);
or U49 (N_49,In_168,In_126);
nor U50 (N_50,In_409,In_578);
nand U51 (N_51,In_740,In_621);
or U52 (N_52,In_270,In_475);
or U53 (N_53,In_140,In_417);
or U54 (N_54,In_558,In_170);
nand U55 (N_55,In_203,In_384);
xor U56 (N_56,In_519,In_197);
nand U57 (N_57,In_63,In_642);
and U58 (N_58,In_257,In_594);
and U59 (N_59,In_639,In_671);
or U60 (N_60,In_590,In_269);
and U61 (N_61,In_483,In_31);
and U62 (N_62,In_587,In_402);
nor U63 (N_63,In_230,In_464);
xor U64 (N_64,In_744,In_544);
nand U65 (N_65,In_397,In_458);
nor U66 (N_66,In_525,In_633);
xor U67 (N_67,In_444,In_300);
xnor U68 (N_68,In_733,In_86);
or U69 (N_69,In_357,In_301);
nor U70 (N_70,In_138,In_556);
and U71 (N_71,In_252,In_232);
nand U72 (N_72,In_605,In_339);
or U73 (N_73,In_509,In_628);
xnor U74 (N_74,In_122,In_565);
nand U75 (N_75,In_109,In_79);
nand U76 (N_76,In_258,In_323);
nand U77 (N_77,In_93,In_616);
nand U78 (N_78,In_66,In_306);
xor U79 (N_79,In_12,In_271);
and U80 (N_80,In_111,In_607);
nor U81 (N_81,In_430,In_152);
and U82 (N_82,In_481,In_71);
and U83 (N_83,In_314,In_277);
xnor U84 (N_84,In_611,In_584);
or U85 (N_85,In_285,In_378);
and U86 (N_86,In_286,In_645);
and U87 (N_87,In_562,In_487);
or U88 (N_88,In_100,In_461);
and U89 (N_89,In_346,In_406);
or U90 (N_90,In_390,In_695);
and U91 (N_91,In_185,In_128);
nand U92 (N_92,In_711,In_121);
and U93 (N_93,In_426,In_403);
nor U94 (N_94,In_251,In_182);
xnor U95 (N_95,In_491,In_579);
nor U96 (N_96,In_72,In_553);
xor U97 (N_97,In_414,In_5);
nand U98 (N_98,In_331,In_714);
and U99 (N_99,In_433,In_736);
and U100 (N_100,In_557,In_489);
nor U101 (N_101,In_404,In_60);
nor U102 (N_102,In_523,In_564);
or U103 (N_103,In_14,In_687);
or U104 (N_104,In_9,In_153);
or U105 (N_105,In_591,In_239);
nor U106 (N_106,In_0,In_210);
nor U107 (N_107,In_208,In_259);
and U108 (N_108,In_572,In_37);
xnor U109 (N_109,In_280,In_64);
or U110 (N_110,In_219,In_337);
xor U111 (N_111,In_209,In_712);
xnor U112 (N_112,In_547,In_310);
or U113 (N_113,In_13,In_455);
xor U114 (N_114,In_349,In_147);
nand U115 (N_115,In_83,In_419);
or U116 (N_116,In_187,In_211);
nand U117 (N_117,In_120,In_673);
and U118 (N_118,In_52,In_469);
and U119 (N_119,In_243,In_46);
or U120 (N_120,In_151,In_54);
and U121 (N_121,In_541,In_125);
and U122 (N_122,In_641,In_206);
xnor U123 (N_123,In_375,In_669);
nand U124 (N_124,In_486,In_70);
xor U125 (N_125,In_478,In_178);
or U126 (N_126,In_413,In_604);
nor U127 (N_127,In_305,In_472);
or U128 (N_128,In_696,In_663);
or U129 (N_129,In_175,In_500);
or U130 (N_130,In_302,In_601);
xnor U131 (N_131,In_352,In_296);
nand U132 (N_132,In_116,In_423);
xor U133 (N_133,In_563,In_615);
nor U134 (N_134,In_40,In_304);
and U135 (N_135,In_23,In_598);
xor U136 (N_136,In_437,In_193);
xor U137 (N_137,In_391,In_599);
and U138 (N_138,In_388,In_272);
xor U139 (N_139,In_261,In_582);
xor U140 (N_140,In_399,In_537);
and U141 (N_141,In_657,In_189);
xor U142 (N_142,In_473,In_221);
or U143 (N_143,In_372,In_614);
or U144 (N_144,In_82,In_634);
xnor U145 (N_145,In_492,In_659);
nand U146 (N_146,In_253,In_629);
xnor U147 (N_147,In_24,In_677);
xnor U148 (N_148,In_429,In_192);
nor U149 (N_149,In_364,In_362);
xnor U150 (N_150,In_368,In_465);
xnor U151 (N_151,In_456,In_434);
xnor U152 (N_152,In_560,In_725);
or U153 (N_153,In_278,In_741);
and U154 (N_154,In_200,In_581);
nand U155 (N_155,In_668,In_11);
or U156 (N_156,In_682,In_117);
nand U157 (N_157,In_99,In_105);
nor U158 (N_158,In_432,In_196);
nand U159 (N_159,In_17,In_171);
nand U160 (N_160,In_87,In_3);
xnor U161 (N_161,In_41,In_227);
and U162 (N_162,In_367,In_451);
nand U163 (N_163,In_180,In_55);
nor U164 (N_164,In_317,In_307);
nand U165 (N_165,In_651,In_490);
nand U166 (N_166,In_254,In_226);
xor U167 (N_167,In_466,In_181);
and U168 (N_168,In_25,In_439);
xnor U169 (N_169,In_308,In_436);
nand U170 (N_170,In_485,In_30);
xor U171 (N_171,In_204,In_660);
and U172 (N_172,In_283,In_446);
xor U173 (N_173,In_161,In_699);
nor U174 (N_174,In_163,In_493);
nand U175 (N_175,In_319,In_569);
nand U176 (N_176,In_47,In_527);
xor U177 (N_177,In_597,In_176);
nor U178 (N_178,In_518,In_148);
and U179 (N_179,In_135,In_21);
nor U180 (N_180,In_245,In_543);
and U181 (N_181,In_412,In_476);
nand U182 (N_182,In_327,In_542);
or U183 (N_183,In_652,In_588);
nor U184 (N_184,In_603,In_680);
xor U185 (N_185,In_459,In_441);
nor U186 (N_186,In_457,In_347);
or U187 (N_187,In_732,In_383);
xor U188 (N_188,In_637,In_702);
and U189 (N_189,In_284,In_114);
or U190 (N_190,In_749,In_727);
nand U191 (N_191,In_173,In_635);
nand U192 (N_192,In_108,In_396);
nor U193 (N_193,In_145,In_242);
nand U194 (N_194,In_540,In_693);
nor U195 (N_195,In_585,In_745);
nor U196 (N_196,In_119,In_511);
nor U197 (N_197,In_29,In_371);
or U198 (N_198,In_684,In_548);
xor U199 (N_199,In_309,In_36);
nand U200 (N_200,In_169,In_342);
nand U201 (N_201,In_613,In_129);
nand U202 (N_202,In_250,In_75);
nor U203 (N_203,In_344,In_103);
or U204 (N_204,In_76,In_561);
or U205 (N_205,In_505,In_194);
or U206 (N_206,In_520,In_57);
nand U207 (N_207,In_172,In_449);
xnor U208 (N_208,In_256,In_167);
nor U209 (N_209,In_554,In_705);
nand U210 (N_210,In_379,In_665);
nand U211 (N_211,In_722,In_132);
nand U212 (N_212,In_648,In_653);
or U213 (N_213,In_322,In_731);
nand U214 (N_214,In_273,In_229);
nor U215 (N_215,In_217,In_228);
nor U216 (N_216,In_235,In_596);
and U217 (N_217,In_526,In_333);
and U218 (N_218,In_361,In_382);
and U219 (N_219,In_452,In_275);
nor U220 (N_220,In_462,In_559);
nand U221 (N_221,In_157,In_199);
nor U222 (N_222,In_207,In_643);
xor U223 (N_223,In_685,In_535);
nor U224 (N_224,In_482,In_2);
or U225 (N_225,In_737,In_566);
and U226 (N_226,In_664,In_626);
xnor U227 (N_227,In_549,In_401);
and U228 (N_228,In_137,In_263);
xnor U229 (N_229,In_742,In_67);
or U230 (N_230,In_69,In_646);
nor U231 (N_231,In_369,In_356);
nor U232 (N_232,In_654,In_341);
nand U233 (N_233,In_471,In_620);
or U234 (N_234,In_240,In_246);
or U235 (N_235,In_389,In_376);
nand U236 (N_236,In_386,In_479);
xor U237 (N_237,In_315,In_655);
xor U238 (N_238,In_360,In_650);
or U239 (N_239,In_191,In_92);
xor U240 (N_240,In_530,In_61);
xnor U241 (N_241,In_218,In_65);
xnor U242 (N_242,In_58,In_484);
xor U243 (N_243,In_570,In_332);
and U244 (N_244,In_698,In_186);
and U245 (N_245,In_514,In_343);
nor U246 (N_246,In_480,In_592);
nand U247 (N_247,In_291,In_735);
or U248 (N_248,In_720,In_624);
and U249 (N_249,In_334,In_644);
and U250 (N_250,In_666,In_498);
and U251 (N_251,In_59,In_640);
and U252 (N_252,In_719,In_276);
nor U253 (N_253,In_238,In_345);
nand U254 (N_254,In_101,In_623);
nand U255 (N_255,In_335,In_324);
or U256 (N_256,In_336,In_700);
nor U257 (N_257,In_715,In_730);
xnor U258 (N_258,In_679,In_27);
or U259 (N_259,In_454,In_395);
xnor U260 (N_260,In_688,In_201);
and U261 (N_261,In_723,In_381);
or U262 (N_262,In_447,In_577);
and U263 (N_263,In_709,In_88);
nand U264 (N_264,In_474,In_48);
xnor U265 (N_265,In_625,In_747);
nor U266 (N_266,In_81,In_215);
xnor U267 (N_267,In_130,In_297);
and U268 (N_268,In_134,In_408);
and U269 (N_269,In_538,In_636);
and U270 (N_270,In_532,In_467);
nand U271 (N_271,In_77,In_442);
or U272 (N_272,In_627,In_154);
xor U273 (N_273,In_214,In_115);
nor U274 (N_274,In_313,In_589);
nand U275 (N_275,In_704,In_96);
and U276 (N_276,In_223,In_139);
and U277 (N_277,In_353,In_143);
or U278 (N_278,In_113,In_718);
nor U279 (N_279,In_600,In_748);
xor U280 (N_280,In_363,In_110);
nor U281 (N_281,In_438,In_39);
nand U282 (N_282,In_721,In_84);
xnor U283 (N_283,In_144,In_411);
or U284 (N_284,In_661,In_340);
nand U285 (N_285,In_184,In_51);
xnor U286 (N_286,In_80,In_734);
nor U287 (N_287,In_141,In_1);
xor U288 (N_288,In_619,In_512);
xnor U289 (N_289,In_160,In_499);
or U290 (N_290,In_460,In_533);
nand U291 (N_291,In_298,In_443);
nor U292 (N_292,In_255,In_179);
or U293 (N_293,In_150,In_708);
nand U294 (N_294,In_274,In_539);
nor U295 (N_295,In_468,In_233);
nor U296 (N_296,In_649,In_146);
or U297 (N_297,In_312,In_303);
or U298 (N_298,In_316,In_502);
or U299 (N_299,In_44,In_617);
nand U300 (N_300,In_488,In_536);
xor U301 (N_301,In_320,In_15);
nand U302 (N_302,In_311,In_445);
and U303 (N_303,In_98,In_612);
or U304 (N_304,In_95,In_422);
xor U305 (N_305,In_321,In_495);
nand U306 (N_306,In_729,In_236);
and U307 (N_307,In_156,In_16);
nor U308 (N_308,In_97,In_656);
xor U309 (N_309,In_392,In_580);
or U310 (N_310,In_131,In_299);
nor U311 (N_311,In_220,In_90);
and U312 (N_312,In_213,In_738);
and U313 (N_313,In_188,In_418);
xnor U314 (N_314,In_249,In_573);
xnor U315 (N_315,In_45,In_94);
xnor U316 (N_316,In_393,In_583);
or U317 (N_317,In_112,In_552);
or U318 (N_318,In_516,In_359);
and U319 (N_319,In_279,In_6);
xor U320 (N_320,In_513,In_477);
nor U321 (N_321,In_62,In_288);
or U322 (N_322,In_506,In_224);
and U323 (N_323,In_517,In_571);
and U324 (N_324,In_212,In_190);
and U325 (N_325,In_701,In_593);
nor U326 (N_326,In_703,In_102);
nand U327 (N_327,In_546,In_380);
and U328 (N_328,In_237,In_450);
nand U329 (N_329,In_534,In_507);
or U330 (N_330,In_707,In_266);
and U331 (N_331,In_28,In_630);
and U332 (N_332,In_225,In_231);
xor U333 (N_333,In_350,In_241);
or U334 (N_334,In_265,In_165);
nand U335 (N_335,In_177,In_524);
nor U336 (N_336,In_78,In_330);
nor U337 (N_337,In_351,In_510);
nand U338 (N_338,In_706,In_326);
nor U339 (N_339,In_166,In_118);
or U340 (N_340,In_678,In_374);
and U341 (N_341,In_295,In_521);
and U342 (N_342,In_528,In_494);
and U343 (N_343,In_400,In_281);
or U344 (N_344,In_394,In_425);
or U345 (N_345,In_123,In_608);
or U346 (N_346,In_497,In_420);
nor U347 (N_347,In_42,In_174);
or U348 (N_348,In_739,In_575);
nor U349 (N_349,In_385,In_622);
or U350 (N_350,In_158,In_373);
or U351 (N_351,In_355,In_638);
nand U352 (N_352,In_18,In_248);
nor U353 (N_353,In_222,In_387);
nor U354 (N_354,In_694,In_555);
or U355 (N_355,In_567,In_428);
nor U356 (N_356,In_338,In_136);
xnor U357 (N_357,In_618,In_681);
nor U358 (N_358,In_405,In_91);
nand U359 (N_359,In_159,In_440);
xor U360 (N_360,In_8,In_22);
and U361 (N_361,In_325,In_421);
nand U362 (N_362,In_424,In_127);
nor U363 (N_363,In_33,In_85);
xor U364 (N_364,In_73,In_726);
nand U365 (N_365,In_260,In_453);
and U366 (N_366,In_551,In_674);
nand U367 (N_367,In_26,In_398);
xor U368 (N_368,In_686,In_463);
and U369 (N_369,In_496,In_124);
xnor U370 (N_370,In_658,In_407);
nor U371 (N_371,In_435,In_247);
nor U372 (N_372,In_264,In_522);
or U373 (N_373,In_20,In_155);
or U374 (N_374,In_675,In_672);
xor U375 (N_375,In_16,In_372);
xnor U376 (N_376,In_417,In_605);
and U377 (N_377,In_499,In_428);
and U378 (N_378,In_472,In_535);
and U379 (N_379,In_488,In_156);
and U380 (N_380,In_398,In_298);
xor U381 (N_381,In_186,In_646);
and U382 (N_382,In_557,In_635);
xor U383 (N_383,In_294,In_276);
nor U384 (N_384,In_68,In_645);
or U385 (N_385,In_581,In_484);
and U386 (N_386,In_136,In_426);
and U387 (N_387,In_689,In_739);
and U388 (N_388,In_581,In_351);
or U389 (N_389,In_575,In_89);
xor U390 (N_390,In_666,In_567);
and U391 (N_391,In_602,In_137);
xor U392 (N_392,In_150,In_428);
or U393 (N_393,In_406,In_456);
or U394 (N_394,In_449,In_237);
or U395 (N_395,In_62,In_500);
or U396 (N_396,In_381,In_279);
nor U397 (N_397,In_514,In_365);
nand U398 (N_398,In_22,In_306);
xnor U399 (N_399,In_401,In_747);
and U400 (N_400,In_144,In_329);
nor U401 (N_401,In_187,In_254);
nand U402 (N_402,In_393,In_494);
and U403 (N_403,In_142,In_511);
xnor U404 (N_404,In_597,In_639);
nand U405 (N_405,In_294,In_329);
nor U406 (N_406,In_262,In_725);
or U407 (N_407,In_593,In_408);
nor U408 (N_408,In_36,In_505);
xnor U409 (N_409,In_457,In_465);
or U410 (N_410,In_620,In_24);
and U411 (N_411,In_672,In_691);
or U412 (N_412,In_448,In_436);
and U413 (N_413,In_708,In_397);
and U414 (N_414,In_613,In_739);
nand U415 (N_415,In_529,In_570);
nand U416 (N_416,In_608,In_232);
nand U417 (N_417,In_679,In_342);
or U418 (N_418,In_674,In_139);
nand U419 (N_419,In_63,In_421);
and U420 (N_420,In_507,In_327);
nor U421 (N_421,In_322,In_617);
xnor U422 (N_422,In_405,In_398);
xnor U423 (N_423,In_95,In_576);
or U424 (N_424,In_334,In_543);
and U425 (N_425,In_261,In_724);
and U426 (N_426,In_454,In_741);
and U427 (N_427,In_162,In_485);
xor U428 (N_428,In_453,In_391);
and U429 (N_429,In_572,In_485);
and U430 (N_430,In_39,In_117);
xnor U431 (N_431,In_333,In_708);
nand U432 (N_432,In_604,In_382);
nor U433 (N_433,In_557,In_246);
xnor U434 (N_434,In_112,In_224);
and U435 (N_435,In_431,In_110);
nor U436 (N_436,In_2,In_69);
xnor U437 (N_437,In_436,In_19);
nor U438 (N_438,In_700,In_541);
xnor U439 (N_439,In_142,In_295);
or U440 (N_440,In_481,In_418);
and U441 (N_441,In_697,In_648);
nor U442 (N_442,In_469,In_515);
and U443 (N_443,In_150,In_204);
xnor U444 (N_444,In_406,In_80);
nor U445 (N_445,In_507,In_659);
and U446 (N_446,In_115,In_376);
nand U447 (N_447,In_421,In_302);
and U448 (N_448,In_394,In_735);
nor U449 (N_449,In_28,In_580);
nand U450 (N_450,In_735,In_594);
and U451 (N_451,In_221,In_399);
nor U452 (N_452,In_170,In_682);
and U453 (N_453,In_597,In_708);
and U454 (N_454,In_87,In_460);
xor U455 (N_455,In_679,In_618);
and U456 (N_456,In_631,In_609);
and U457 (N_457,In_356,In_276);
or U458 (N_458,In_43,In_590);
xor U459 (N_459,In_174,In_581);
nor U460 (N_460,In_252,In_103);
and U461 (N_461,In_127,In_144);
nand U462 (N_462,In_324,In_249);
or U463 (N_463,In_561,In_110);
nand U464 (N_464,In_190,In_157);
xor U465 (N_465,In_287,In_635);
nor U466 (N_466,In_406,In_250);
or U467 (N_467,In_235,In_119);
and U468 (N_468,In_637,In_421);
and U469 (N_469,In_413,In_455);
or U470 (N_470,In_56,In_746);
xnor U471 (N_471,In_247,In_56);
and U472 (N_472,In_358,In_286);
nor U473 (N_473,In_501,In_402);
and U474 (N_474,In_643,In_221);
xnor U475 (N_475,In_272,In_688);
nand U476 (N_476,In_225,In_289);
or U477 (N_477,In_631,In_623);
nand U478 (N_478,In_344,In_144);
and U479 (N_479,In_584,In_524);
nand U480 (N_480,In_410,In_587);
and U481 (N_481,In_437,In_474);
xnor U482 (N_482,In_282,In_636);
and U483 (N_483,In_127,In_147);
nor U484 (N_484,In_411,In_517);
or U485 (N_485,In_460,In_72);
or U486 (N_486,In_420,In_60);
xnor U487 (N_487,In_375,In_631);
or U488 (N_488,In_23,In_719);
nand U489 (N_489,In_276,In_226);
or U490 (N_490,In_494,In_498);
nor U491 (N_491,In_596,In_253);
and U492 (N_492,In_25,In_26);
or U493 (N_493,In_637,In_728);
xor U494 (N_494,In_286,In_529);
or U495 (N_495,In_53,In_162);
or U496 (N_496,In_605,In_570);
xor U497 (N_497,In_275,In_499);
or U498 (N_498,In_634,In_578);
nand U499 (N_499,In_98,In_303);
or U500 (N_500,In_299,In_263);
xnor U501 (N_501,In_335,In_559);
or U502 (N_502,In_291,In_458);
nand U503 (N_503,In_232,In_308);
xor U504 (N_504,In_237,In_602);
xor U505 (N_505,In_158,In_564);
nor U506 (N_506,In_550,In_250);
and U507 (N_507,In_276,In_199);
and U508 (N_508,In_198,In_4);
xor U509 (N_509,In_314,In_551);
nand U510 (N_510,In_88,In_180);
nand U511 (N_511,In_639,In_181);
or U512 (N_512,In_195,In_612);
xor U513 (N_513,In_173,In_648);
nor U514 (N_514,In_299,In_494);
and U515 (N_515,In_399,In_688);
and U516 (N_516,In_606,In_272);
and U517 (N_517,In_657,In_231);
nand U518 (N_518,In_662,In_274);
or U519 (N_519,In_402,In_22);
nor U520 (N_520,In_206,In_707);
nor U521 (N_521,In_258,In_102);
or U522 (N_522,In_335,In_386);
nand U523 (N_523,In_406,In_309);
nor U524 (N_524,In_675,In_702);
or U525 (N_525,In_312,In_209);
or U526 (N_526,In_388,In_594);
nor U527 (N_527,In_511,In_159);
nand U528 (N_528,In_183,In_423);
nor U529 (N_529,In_105,In_507);
nor U530 (N_530,In_166,In_631);
and U531 (N_531,In_390,In_121);
xor U532 (N_532,In_331,In_500);
xnor U533 (N_533,In_704,In_281);
and U534 (N_534,In_496,In_546);
and U535 (N_535,In_516,In_254);
or U536 (N_536,In_325,In_413);
and U537 (N_537,In_214,In_216);
and U538 (N_538,In_96,In_574);
xor U539 (N_539,In_246,In_355);
nor U540 (N_540,In_262,In_519);
xor U541 (N_541,In_547,In_617);
nand U542 (N_542,In_688,In_288);
and U543 (N_543,In_384,In_504);
xnor U544 (N_544,In_380,In_157);
nor U545 (N_545,In_298,In_411);
nand U546 (N_546,In_191,In_315);
or U547 (N_547,In_485,In_699);
nand U548 (N_548,In_565,In_346);
and U549 (N_549,In_154,In_103);
or U550 (N_550,In_439,In_219);
xor U551 (N_551,In_121,In_4);
and U552 (N_552,In_504,In_580);
or U553 (N_553,In_524,In_672);
xor U554 (N_554,In_525,In_287);
xnor U555 (N_555,In_259,In_129);
nand U556 (N_556,In_630,In_369);
xor U557 (N_557,In_259,In_246);
nor U558 (N_558,In_638,In_371);
nor U559 (N_559,In_502,In_311);
nor U560 (N_560,In_571,In_211);
or U561 (N_561,In_203,In_515);
nand U562 (N_562,In_484,In_316);
xnor U563 (N_563,In_606,In_560);
xor U564 (N_564,In_185,In_76);
xor U565 (N_565,In_260,In_17);
nand U566 (N_566,In_725,In_253);
nand U567 (N_567,In_247,In_501);
nor U568 (N_568,In_10,In_508);
xnor U569 (N_569,In_331,In_126);
xnor U570 (N_570,In_155,In_283);
nor U571 (N_571,In_608,In_517);
nand U572 (N_572,In_283,In_670);
xor U573 (N_573,In_654,In_477);
or U574 (N_574,In_71,In_547);
xnor U575 (N_575,In_445,In_631);
and U576 (N_576,In_298,In_50);
nand U577 (N_577,In_463,In_386);
nor U578 (N_578,In_446,In_467);
nand U579 (N_579,In_244,In_552);
and U580 (N_580,In_310,In_622);
nor U581 (N_581,In_89,In_255);
xnor U582 (N_582,In_147,In_570);
and U583 (N_583,In_449,In_705);
or U584 (N_584,In_505,In_740);
or U585 (N_585,In_644,In_279);
and U586 (N_586,In_526,In_719);
nor U587 (N_587,In_673,In_587);
and U588 (N_588,In_504,In_3);
nor U589 (N_589,In_544,In_695);
nor U590 (N_590,In_165,In_412);
or U591 (N_591,In_175,In_698);
or U592 (N_592,In_746,In_348);
and U593 (N_593,In_80,In_31);
xnor U594 (N_594,In_738,In_445);
xor U595 (N_595,In_346,In_398);
or U596 (N_596,In_456,In_258);
or U597 (N_597,In_379,In_609);
or U598 (N_598,In_682,In_555);
or U599 (N_599,In_717,In_14);
or U600 (N_600,In_73,In_149);
xor U601 (N_601,In_303,In_158);
nand U602 (N_602,In_312,In_543);
nor U603 (N_603,In_248,In_127);
and U604 (N_604,In_695,In_208);
or U605 (N_605,In_526,In_624);
nand U606 (N_606,In_48,In_52);
xnor U607 (N_607,In_613,In_395);
nand U608 (N_608,In_468,In_579);
or U609 (N_609,In_136,In_501);
nor U610 (N_610,In_35,In_683);
nand U611 (N_611,In_618,In_644);
xnor U612 (N_612,In_577,In_572);
xor U613 (N_613,In_477,In_661);
or U614 (N_614,In_210,In_185);
or U615 (N_615,In_49,In_265);
nor U616 (N_616,In_439,In_170);
nor U617 (N_617,In_624,In_683);
and U618 (N_618,In_700,In_627);
xor U619 (N_619,In_496,In_223);
nand U620 (N_620,In_292,In_267);
or U621 (N_621,In_109,In_449);
nand U622 (N_622,In_598,In_725);
nand U623 (N_623,In_321,In_510);
or U624 (N_624,In_102,In_130);
nand U625 (N_625,In_475,In_317);
nand U626 (N_626,In_489,In_501);
or U627 (N_627,In_428,In_58);
nand U628 (N_628,In_38,In_37);
and U629 (N_629,In_523,In_496);
nor U630 (N_630,In_346,In_555);
or U631 (N_631,In_687,In_433);
or U632 (N_632,In_232,In_662);
nor U633 (N_633,In_720,In_62);
nand U634 (N_634,In_676,In_230);
and U635 (N_635,In_122,In_130);
and U636 (N_636,In_151,In_389);
and U637 (N_637,In_111,In_683);
nand U638 (N_638,In_739,In_130);
and U639 (N_639,In_533,In_366);
and U640 (N_640,In_622,In_684);
and U641 (N_641,In_256,In_631);
or U642 (N_642,In_370,In_441);
nor U643 (N_643,In_376,In_422);
nor U644 (N_644,In_219,In_155);
xnor U645 (N_645,In_306,In_258);
and U646 (N_646,In_329,In_468);
or U647 (N_647,In_231,In_223);
or U648 (N_648,In_298,In_158);
and U649 (N_649,In_314,In_27);
and U650 (N_650,In_515,In_131);
or U651 (N_651,In_262,In_643);
or U652 (N_652,In_328,In_537);
or U653 (N_653,In_672,In_552);
nand U654 (N_654,In_623,In_425);
nand U655 (N_655,In_526,In_147);
and U656 (N_656,In_234,In_709);
or U657 (N_657,In_449,In_485);
nand U658 (N_658,In_358,In_74);
and U659 (N_659,In_676,In_262);
nor U660 (N_660,In_455,In_660);
nand U661 (N_661,In_714,In_419);
nor U662 (N_662,In_624,In_295);
and U663 (N_663,In_247,In_274);
or U664 (N_664,In_285,In_346);
or U665 (N_665,In_604,In_531);
nand U666 (N_666,In_481,In_41);
nor U667 (N_667,In_583,In_698);
nor U668 (N_668,In_150,In_384);
xor U669 (N_669,In_632,In_662);
xnor U670 (N_670,In_711,In_339);
nor U671 (N_671,In_515,In_619);
xor U672 (N_672,In_737,In_253);
nand U673 (N_673,In_191,In_605);
nand U674 (N_674,In_100,In_482);
nand U675 (N_675,In_163,In_99);
nor U676 (N_676,In_573,In_344);
xnor U677 (N_677,In_524,In_190);
nor U678 (N_678,In_4,In_355);
xnor U679 (N_679,In_446,In_41);
and U680 (N_680,In_129,In_433);
xnor U681 (N_681,In_671,In_425);
xor U682 (N_682,In_452,In_175);
nand U683 (N_683,In_403,In_316);
and U684 (N_684,In_605,In_26);
nand U685 (N_685,In_103,In_720);
and U686 (N_686,In_369,In_178);
nand U687 (N_687,In_448,In_186);
xor U688 (N_688,In_691,In_578);
nand U689 (N_689,In_217,In_27);
nand U690 (N_690,In_447,In_402);
nand U691 (N_691,In_13,In_159);
nand U692 (N_692,In_733,In_278);
xnor U693 (N_693,In_371,In_703);
or U694 (N_694,In_448,In_417);
and U695 (N_695,In_304,In_228);
nand U696 (N_696,In_679,In_114);
xor U697 (N_697,In_539,In_236);
nand U698 (N_698,In_723,In_328);
nand U699 (N_699,In_488,In_153);
xor U700 (N_700,In_59,In_268);
nor U701 (N_701,In_573,In_394);
xor U702 (N_702,In_87,In_667);
nor U703 (N_703,In_526,In_189);
and U704 (N_704,In_157,In_111);
nor U705 (N_705,In_589,In_382);
nand U706 (N_706,In_308,In_116);
and U707 (N_707,In_125,In_287);
and U708 (N_708,In_113,In_726);
and U709 (N_709,In_249,In_200);
nor U710 (N_710,In_186,In_718);
nand U711 (N_711,In_308,In_722);
nor U712 (N_712,In_495,In_736);
nor U713 (N_713,In_709,In_575);
nor U714 (N_714,In_409,In_55);
or U715 (N_715,In_35,In_139);
and U716 (N_716,In_604,In_392);
xnor U717 (N_717,In_651,In_504);
nand U718 (N_718,In_529,In_598);
xnor U719 (N_719,In_428,In_268);
xnor U720 (N_720,In_680,In_6);
xnor U721 (N_721,In_381,In_332);
and U722 (N_722,In_337,In_423);
nand U723 (N_723,In_113,In_571);
xnor U724 (N_724,In_280,In_740);
and U725 (N_725,In_340,In_264);
and U726 (N_726,In_29,In_409);
xor U727 (N_727,In_469,In_429);
and U728 (N_728,In_457,In_274);
or U729 (N_729,In_322,In_140);
or U730 (N_730,In_530,In_738);
nand U731 (N_731,In_669,In_523);
and U732 (N_732,In_318,In_96);
nand U733 (N_733,In_643,In_593);
or U734 (N_734,In_383,In_26);
and U735 (N_735,In_423,In_194);
nor U736 (N_736,In_426,In_375);
nand U737 (N_737,In_681,In_159);
or U738 (N_738,In_664,In_360);
nor U739 (N_739,In_124,In_553);
nand U740 (N_740,In_144,In_33);
xor U741 (N_741,In_175,In_19);
and U742 (N_742,In_521,In_578);
nor U743 (N_743,In_478,In_724);
nand U744 (N_744,In_625,In_143);
nor U745 (N_745,In_130,In_124);
nor U746 (N_746,In_728,In_696);
nor U747 (N_747,In_668,In_17);
and U748 (N_748,In_415,In_263);
and U749 (N_749,In_350,In_628);
and U750 (N_750,In_731,In_719);
xor U751 (N_751,In_168,In_726);
and U752 (N_752,In_432,In_636);
or U753 (N_753,In_640,In_373);
xor U754 (N_754,In_153,In_497);
nor U755 (N_755,In_374,In_238);
and U756 (N_756,In_480,In_400);
and U757 (N_757,In_680,In_195);
nand U758 (N_758,In_314,In_212);
and U759 (N_759,In_60,In_373);
or U760 (N_760,In_236,In_26);
nor U761 (N_761,In_192,In_438);
and U762 (N_762,In_500,In_109);
and U763 (N_763,In_601,In_671);
nand U764 (N_764,In_728,In_400);
and U765 (N_765,In_356,In_172);
and U766 (N_766,In_636,In_116);
nand U767 (N_767,In_574,In_168);
and U768 (N_768,In_158,In_131);
nor U769 (N_769,In_512,In_729);
xor U770 (N_770,In_706,In_196);
xnor U771 (N_771,In_335,In_623);
and U772 (N_772,In_312,In_332);
and U773 (N_773,In_202,In_697);
and U774 (N_774,In_501,In_588);
or U775 (N_775,In_123,In_524);
nand U776 (N_776,In_204,In_520);
and U777 (N_777,In_137,In_505);
and U778 (N_778,In_607,In_72);
xnor U779 (N_779,In_435,In_367);
xnor U780 (N_780,In_78,In_394);
nand U781 (N_781,In_467,In_31);
or U782 (N_782,In_717,In_589);
nand U783 (N_783,In_670,In_577);
and U784 (N_784,In_527,In_274);
nand U785 (N_785,In_121,In_509);
xor U786 (N_786,In_630,In_284);
xor U787 (N_787,In_702,In_304);
nor U788 (N_788,In_385,In_478);
nand U789 (N_789,In_80,In_326);
or U790 (N_790,In_121,In_700);
nand U791 (N_791,In_125,In_123);
xnor U792 (N_792,In_50,In_118);
nand U793 (N_793,In_332,In_349);
nand U794 (N_794,In_10,In_650);
nand U795 (N_795,In_237,In_353);
xnor U796 (N_796,In_531,In_236);
nand U797 (N_797,In_498,In_113);
nand U798 (N_798,In_129,In_711);
or U799 (N_799,In_667,In_104);
and U800 (N_800,In_701,In_434);
nor U801 (N_801,In_273,In_381);
or U802 (N_802,In_603,In_744);
or U803 (N_803,In_631,In_149);
xor U804 (N_804,In_281,In_395);
xor U805 (N_805,In_326,In_228);
xnor U806 (N_806,In_312,In_402);
nor U807 (N_807,In_393,In_447);
or U808 (N_808,In_554,In_352);
or U809 (N_809,In_509,In_117);
nor U810 (N_810,In_148,In_368);
nand U811 (N_811,In_524,In_625);
nor U812 (N_812,In_126,In_215);
and U813 (N_813,In_157,In_154);
nand U814 (N_814,In_651,In_151);
xor U815 (N_815,In_429,In_336);
nor U816 (N_816,In_673,In_588);
xor U817 (N_817,In_519,In_729);
or U818 (N_818,In_52,In_117);
nor U819 (N_819,In_135,In_74);
or U820 (N_820,In_200,In_492);
nand U821 (N_821,In_335,In_164);
and U822 (N_822,In_359,In_177);
xnor U823 (N_823,In_478,In_297);
nand U824 (N_824,In_112,In_355);
nor U825 (N_825,In_564,In_357);
nor U826 (N_826,In_746,In_623);
nor U827 (N_827,In_580,In_675);
and U828 (N_828,In_191,In_665);
nor U829 (N_829,In_550,In_336);
nor U830 (N_830,In_70,In_148);
nand U831 (N_831,In_503,In_457);
and U832 (N_832,In_703,In_536);
nand U833 (N_833,In_269,In_33);
and U834 (N_834,In_220,In_335);
nor U835 (N_835,In_448,In_50);
xnor U836 (N_836,In_180,In_462);
or U837 (N_837,In_209,In_460);
or U838 (N_838,In_415,In_723);
nor U839 (N_839,In_160,In_114);
nor U840 (N_840,In_160,In_563);
xor U841 (N_841,In_297,In_41);
nand U842 (N_842,In_702,In_542);
nor U843 (N_843,In_631,In_248);
or U844 (N_844,In_285,In_151);
and U845 (N_845,In_518,In_631);
nor U846 (N_846,In_393,In_426);
nor U847 (N_847,In_199,In_81);
xor U848 (N_848,In_580,In_194);
and U849 (N_849,In_124,In_172);
nand U850 (N_850,In_251,In_297);
nand U851 (N_851,In_537,In_327);
and U852 (N_852,In_728,In_422);
and U853 (N_853,In_310,In_446);
nor U854 (N_854,In_629,In_326);
or U855 (N_855,In_635,In_477);
nor U856 (N_856,In_315,In_196);
nor U857 (N_857,In_565,In_375);
nand U858 (N_858,In_207,In_483);
and U859 (N_859,In_142,In_563);
or U860 (N_860,In_287,In_105);
nand U861 (N_861,In_180,In_379);
xnor U862 (N_862,In_189,In_240);
nor U863 (N_863,In_534,In_46);
or U864 (N_864,In_441,In_9);
nor U865 (N_865,In_708,In_645);
and U866 (N_866,In_192,In_635);
nand U867 (N_867,In_709,In_535);
and U868 (N_868,In_553,In_318);
or U869 (N_869,In_27,In_62);
nor U870 (N_870,In_483,In_381);
nor U871 (N_871,In_571,In_538);
nand U872 (N_872,In_464,In_23);
and U873 (N_873,In_174,In_334);
nor U874 (N_874,In_715,In_248);
nor U875 (N_875,In_443,In_521);
nor U876 (N_876,In_148,In_722);
nand U877 (N_877,In_350,In_464);
or U878 (N_878,In_646,In_682);
nand U879 (N_879,In_428,In_69);
nand U880 (N_880,In_197,In_421);
nor U881 (N_881,In_418,In_740);
and U882 (N_882,In_332,In_229);
nand U883 (N_883,In_453,In_443);
or U884 (N_884,In_18,In_499);
nor U885 (N_885,In_362,In_172);
and U886 (N_886,In_125,In_1);
xnor U887 (N_887,In_397,In_564);
and U888 (N_888,In_587,In_225);
xor U889 (N_889,In_282,In_576);
nand U890 (N_890,In_18,In_29);
nor U891 (N_891,In_475,In_714);
nor U892 (N_892,In_249,In_389);
and U893 (N_893,In_679,In_15);
nand U894 (N_894,In_84,In_557);
or U895 (N_895,In_325,In_730);
nand U896 (N_896,In_203,In_390);
or U897 (N_897,In_676,In_37);
and U898 (N_898,In_587,In_637);
xor U899 (N_899,In_474,In_528);
nand U900 (N_900,In_290,In_107);
and U901 (N_901,In_438,In_688);
xnor U902 (N_902,In_536,In_133);
nor U903 (N_903,In_344,In_48);
and U904 (N_904,In_135,In_707);
nor U905 (N_905,In_392,In_660);
nor U906 (N_906,In_390,In_553);
nand U907 (N_907,In_362,In_136);
xnor U908 (N_908,In_277,In_496);
and U909 (N_909,In_324,In_635);
and U910 (N_910,In_33,In_37);
xnor U911 (N_911,In_459,In_606);
nand U912 (N_912,In_205,In_301);
nand U913 (N_913,In_460,In_722);
or U914 (N_914,In_657,In_615);
nand U915 (N_915,In_60,In_667);
or U916 (N_916,In_55,In_732);
nor U917 (N_917,In_446,In_231);
and U918 (N_918,In_199,In_568);
nand U919 (N_919,In_102,In_734);
or U920 (N_920,In_413,In_308);
xnor U921 (N_921,In_589,In_442);
nand U922 (N_922,In_654,In_716);
nand U923 (N_923,In_314,In_411);
nand U924 (N_924,In_647,In_328);
xor U925 (N_925,In_402,In_367);
nand U926 (N_926,In_567,In_531);
and U927 (N_927,In_743,In_478);
or U928 (N_928,In_191,In_465);
nor U929 (N_929,In_50,In_246);
nor U930 (N_930,In_638,In_115);
and U931 (N_931,In_343,In_510);
xnor U932 (N_932,In_410,In_533);
nand U933 (N_933,In_106,In_446);
nor U934 (N_934,In_586,In_613);
or U935 (N_935,In_532,In_476);
and U936 (N_936,In_721,In_635);
nand U937 (N_937,In_47,In_601);
nor U938 (N_938,In_749,In_557);
and U939 (N_939,In_247,In_678);
nor U940 (N_940,In_623,In_381);
xor U941 (N_941,In_743,In_156);
xnor U942 (N_942,In_592,In_104);
and U943 (N_943,In_244,In_324);
and U944 (N_944,In_473,In_499);
nand U945 (N_945,In_530,In_184);
and U946 (N_946,In_106,In_411);
or U947 (N_947,In_308,In_200);
xor U948 (N_948,In_527,In_37);
xnor U949 (N_949,In_18,In_749);
or U950 (N_950,In_429,In_658);
xor U951 (N_951,In_671,In_185);
nand U952 (N_952,In_469,In_331);
nor U953 (N_953,In_491,In_224);
and U954 (N_954,In_519,In_605);
or U955 (N_955,In_651,In_515);
and U956 (N_956,In_152,In_445);
and U957 (N_957,In_639,In_33);
and U958 (N_958,In_343,In_658);
and U959 (N_959,In_493,In_370);
and U960 (N_960,In_406,In_430);
xor U961 (N_961,In_267,In_356);
nand U962 (N_962,In_657,In_402);
nand U963 (N_963,In_114,In_557);
xor U964 (N_964,In_159,In_414);
xor U965 (N_965,In_716,In_468);
xnor U966 (N_966,In_179,In_536);
xnor U967 (N_967,In_9,In_50);
nor U968 (N_968,In_624,In_420);
and U969 (N_969,In_661,In_155);
xor U970 (N_970,In_450,In_15);
or U971 (N_971,In_203,In_414);
or U972 (N_972,In_259,In_104);
xor U973 (N_973,In_577,In_94);
and U974 (N_974,In_158,In_527);
nor U975 (N_975,In_605,In_526);
and U976 (N_976,In_607,In_25);
xnor U977 (N_977,In_639,In_519);
and U978 (N_978,In_586,In_232);
nand U979 (N_979,In_543,In_267);
nor U980 (N_980,In_353,In_436);
nor U981 (N_981,In_55,In_667);
xnor U982 (N_982,In_56,In_78);
xor U983 (N_983,In_561,In_529);
and U984 (N_984,In_113,In_439);
nand U985 (N_985,In_77,In_6);
nand U986 (N_986,In_701,In_730);
nor U987 (N_987,In_610,In_397);
xor U988 (N_988,In_30,In_349);
and U989 (N_989,In_379,In_205);
xnor U990 (N_990,In_342,In_283);
or U991 (N_991,In_703,In_265);
and U992 (N_992,In_104,In_83);
and U993 (N_993,In_246,In_441);
and U994 (N_994,In_257,In_563);
xnor U995 (N_995,In_444,In_458);
xnor U996 (N_996,In_115,In_473);
nor U997 (N_997,In_16,In_136);
xor U998 (N_998,In_76,In_459);
or U999 (N_999,In_674,In_511);
and U1000 (N_1000,In_9,In_8);
or U1001 (N_1001,In_11,In_568);
nor U1002 (N_1002,In_296,In_646);
xor U1003 (N_1003,In_388,In_45);
nand U1004 (N_1004,In_492,In_644);
xor U1005 (N_1005,In_58,In_355);
and U1006 (N_1006,In_612,In_739);
xnor U1007 (N_1007,In_24,In_372);
nor U1008 (N_1008,In_684,In_674);
nor U1009 (N_1009,In_59,In_577);
and U1010 (N_1010,In_594,In_88);
or U1011 (N_1011,In_622,In_722);
nor U1012 (N_1012,In_240,In_662);
and U1013 (N_1013,In_441,In_542);
or U1014 (N_1014,In_330,In_340);
xnor U1015 (N_1015,In_525,In_308);
xnor U1016 (N_1016,In_125,In_586);
and U1017 (N_1017,In_669,In_526);
xnor U1018 (N_1018,In_664,In_224);
or U1019 (N_1019,In_602,In_112);
nor U1020 (N_1020,In_204,In_180);
nor U1021 (N_1021,In_129,In_128);
nor U1022 (N_1022,In_343,In_435);
nor U1023 (N_1023,In_663,In_674);
nor U1024 (N_1024,In_110,In_51);
and U1025 (N_1025,In_432,In_81);
xor U1026 (N_1026,In_575,In_43);
nor U1027 (N_1027,In_178,In_528);
xnor U1028 (N_1028,In_238,In_30);
nor U1029 (N_1029,In_140,In_263);
xor U1030 (N_1030,In_276,In_1);
or U1031 (N_1031,In_77,In_546);
nand U1032 (N_1032,In_260,In_154);
xor U1033 (N_1033,In_86,In_60);
xnor U1034 (N_1034,In_320,In_635);
or U1035 (N_1035,In_668,In_240);
nor U1036 (N_1036,In_330,In_285);
or U1037 (N_1037,In_438,In_274);
xnor U1038 (N_1038,In_7,In_687);
or U1039 (N_1039,In_407,In_343);
xor U1040 (N_1040,In_181,In_568);
xnor U1041 (N_1041,In_461,In_718);
nand U1042 (N_1042,In_172,In_34);
nor U1043 (N_1043,In_661,In_275);
or U1044 (N_1044,In_416,In_680);
xnor U1045 (N_1045,In_173,In_10);
and U1046 (N_1046,In_551,In_719);
nand U1047 (N_1047,In_115,In_306);
or U1048 (N_1048,In_161,In_350);
nand U1049 (N_1049,In_711,In_722);
and U1050 (N_1050,In_653,In_13);
and U1051 (N_1051,In_549,In_184);
nor U1052 (N_1052,In_335,In_137);
or U1053 (N_1053,In_154,In_725);
xor U1054 (N_1054,In_514,In_94);
or U1055 (N_1055,In_541,In_340);
xor U1056 (N_1056,In_738,In_576);
nand U1057 (N_1057,In_478,In_270);
nor U1058 (N_1058,In_669,In_154);
xor U1059 (N_1059,In_109,In_32);
and U1060 (N_1060,In_525,In_298);
nor U1061 (N_1061,In_5,In_655);
xnor U1062 (N_1062,In_76,In_384);
nor U1063 (N_1063,In_597,In_703);
or U1064 (N_1064,In_35,In_169);
or U1065 (N_1065,In_241,In_8);
nand U1066 (N_1066,In_289,In_661);
xor U1067 (N_1067,In_24,In_468);
nand U1068 (N_1068,In_139,In_152);
nand U1069 (N_1069,In_39,In_608);
nor U1070 (N_1070,In_707,In_87);
or U1071 (N_1071,In_126,In_720);
nor U1072 (N_1072,In_416,In_696);
nor U1073 (N_1073,In_556,In_728);
nor U1074 (N_1074,In_745,In_511);
and U1075 (N_1075,In_256,In_495);
nand U1076 (N_1076,In_624,In_144);
nand U1077 (N_1077,In_429,In_419);
xnor U1078 (N_1078,In_394,In_736);
or U1079 (N_1079,In_273,In_298);
nor U1080 (N_1080,In_230,In_219);
nor U1081 (N_1081,In_407,In_232);
or U1082 (N_1082,In_177,In_229);
xnor U1083 (N_1083,In_415,In_591);
nand U1084 (N_1084,In_249,In_578);
nor U1085 (N_1085,In_83,In_19);
nor U1086 (N_1086,In_701,In_605);
or U1087 (N_1087,In_78,In_186);
xnor U1088 (N_1088,In_682,In_747);
or U1089 (N_1089,In_326,In_246);
nand U1090 (N_1090,In_467,In_128);
and U1091 (N_1091,In_315,In_677);
or U1092 (N_1092,In_299,In_310);
nor U1093 (N_1093,In_568,In_487);
or U1094 (N_1094,In_749,In_378);
and U1095 (N_1095,In_512,In_471);
nand U1096 (N_1096,In_644,In_265);
nand U1097 (N_1097,In_515,In_261);
xor U1098 (N_1098,In_732,In_179);
xnor U1099 (N_1099,In_576,In_496);
nor U1100 (N_1100,In_150,In_480);
nand U1101 (N_1101,In_599,In_40);
and U1102 (N_1102,In_476,In_367);
nand U1103 (N_1103,In_703,In_606);
nor U1104 (N_1104,In_552,In_149);
nor U1105 (N_1105,In_430,In_688);
xor U1106 (N_1106,In_134,In_672);
or U1107 (N_1107,In_392,In_597);
nand U1108 (N_1108,In_586,In_568);
nor U1109 (N_1109,In_429,In_340);
nor U1110 (N_1110,In_374,In_104);
nor U1111 (N_1111,In_105,In_340);
or U1112 (N_1112,In_404,In_254);
nand U1113 (N_1113,In_687,In_661);
and U1114 (N_1114,In_332,In_333);
or U1115 (N_1115,In_314,In_8);
nor U1116 (N_1116,In_78,In_155);
and U1117 (N_1117,In_9,In_685);
nor U1118 (N_1118,In_710,In_619);
xor U1119 (N_1119,In_546,In_175);
and U1120 (N_1120,In_464,In_337);
or U1121 (N_1121,In_441,In_102);
nor U1122 (N_1122,In_578,In_232);
nand U1123 (N_1123,In_589,In_143);
xnor U1124 (N_1124,In_132,In_520);
nor U1125 (N_1125,In_221,In_127);
nand U1126 (N_1126,In_333,In_564);
and U1127 (N_1127,In_397,In_123);
xnor U1128 (N_1128,In_271,In_398);
nor U1129 (N_1129,In_532,In_259);
nor U1130 (N_1130,In_357,In_181);
nor U1131 (N_1131,In_97,In_431);
xor U1132 (N_1132,In_53,In_250);
xnor U1133 (N_1133,In_594,In_59);
nor U1134 (N_1134,In_157,In_8);
or U1135 (N_1135,In_451,In_245);
nand U1136 (N_1136,In_612,In_525);
or U1137 (N_1137,In_385,In_498);
and U1138 (N_1138,In_696,In_655);
or U1139 (N_1139,In_403,In_309);
nand U1140 (N_1140,In_343,In_191);
nand U1141 (N_1141,In_177,In_155);
xnor U1142 (N_1142,In_34,In_588);
nand U1143 (N_1143,In_168,In_483);
or U1144 (N_1144,In_698,In_191);
nand U1145 (N_1145,In_297,In_218);
or U1146 (N_1146,In_66,In_88);
and U1147 (N_1147,In_408,In_740);
xnor U1148 (N_1148,In_105,In_539);
nand U1149 (N_1149,In_249,In_641);
and U1150 (N_1150,In_699,In_209);
and U1151 (N_1151,In_3,In_297);
xor U1152 (N_1152,In_454,In_707);
xnor U1153 (N_1153,In_40,In_494);
nand U1154 (N_1154,In_612,In_386);
xnor U1155 (N_1155,In_290,In_14);
or U1156 (N_1156,In_184,In_665);
xnor U1157 (N_1157,In_324,In_114);
and U1158 (N_1158,In_97,In_624);
and U1159 (N_1159,In_427,In_467);
or U1160 (N_1160,In_711,In_661);
nand U1161 (N_1161,In_640,In_607);
or U1162 (N_1162,In_539,In_637);
xnor U1163 (N_1163,In_446,In_656);
xor U1164 (N_1164,In_555,In_295);
nand U1165 (N_1165,In_633,In_5);
xnor U1166 (N_1166,In_118,In_548);
nand U1167 (N_1167,In_711,In_688);
and U1168 (N_1168,In_505,In_68);
xor U1169 (N_1169,In_442,In_103);
nor U1170 (N_1170,In_729,In_574);
nor U1171 (N_1171,In_252,In_199);
xor U1172 (N_1172,In_254,In_13);
and U1173 (N_1173,In_201,In_690);
nand U1174 (N_1174,In_483,In_45);
nor U1175 (N_1175,In_21,In_737);
or U1176 (N_1176,In_195,In_742);
xnor U1177 (N_1177,In_127,In_42);
xor U1178 (N_1178,In_595,In_335);
and U1179 (N_1179,In_645,In_588);
and U1180 (N_1180,In_354,In_736);
and U1181 (N_1181,In_349,In_319);
nor U1182 (N_1182,In_652,In_730);
xnor U1183 (N_1183,In_10,In_668);
and U1184 (N_1184,In_230,In_525);
or U1185 (N_1185,In_719,In_412);
nand U1186 (N_1186,In_322,In_505);
nand U1187 (N_1187,In_586,In_209);
xor U1188 (N_1188,In_25,In_710);
nand U1189 (N_1189,In_160,In_605);
nand U1190 (N_1190,In_67,In_661);
or U1191 (N_1191,In_22,In_500);
and U1192 (N_1192,In_418,In_218);
xor U1193 (N_1193,In_487,In_185);
and U1194 (N_1194,In_523,In_332);
xnor U1195 (N_1195,In_579,In_623);
and U1196 (N_1196,In_389,In_81);
and U1197 (N_1197,In_530,In_453);
nand U1198 (N_1198,In_708,In_474);
or U1199 (N_1199,In_284,In_422);
nor U1200 (N_1200,In_144,In_256);
nand U1201 (N_1201,In_98,In_451);
or U1202 (N_1202,In_611,In_180);
nand U1203 (N_1203,In_159,In_342);
or U1204 (N_1204,In_139,In_600);
or U1205 (N_1205,In_398,In_565);
nor U1206 (N_1206,In_372,In_616);
or U1207 (N_1207,In_84,In_135);
and U1208 (N_1208,In_70,In_534);
nand U1209 (N_1209,In_362,In_353);
or U1210 (N_1210,In_198,In_217);
and U1211 (N_1211,In_286,In_517);
and U1212 (N_1212,In_314,In_487);
nor U1213 (N_1213,In_678,In_256);
nand U1214 (N_1214,In_229,In_361);
xor U1215 (N_1215,In_36,In_655);
and U1216 (N_1216,In_291,In_561);
nand U1217 (N_1217,In_455,In_171);
or U1218 (N_1218,In_578,In_161);
and U1219 (N_1219,In_122,In_672);
and U1220 (N_1220,In_518,In_69);
xnor U1221 (N_1221,In_328,In_429);
xnor U1222 (N_1222,In_475,In_5);
and U1223 (N_1223,In_202,In_499);
and U1224 (N_1224,In_677,In_666);
xnor U1225 (N_1225,In_363,In_148);
nor U1226 (N_1226,In_58,In_235);
xnor U1227 (N_1227,In_409,In_393);
nand U1228 (N_1228,In_558,In_22);
nand U1229 (N_1229,In_44,In_523);
nand U1230 (N_1230,In_458,In_55);
and U1231 (N_1231,In_159,In_626);
or U1232 (N_1232,In_704,In_604);
or U1233 (N_1233,In_60,In_225);
and U1234 (N_1234,In_129,In_330);
xnor U1235 (N_1235,In_485,In_170);
and U1236 (N_1236,In_422,In_605);
nand U1237 (N_1237,In_499,In_336);
or U1238 (N_1238,In_256,In_342);
or U1239 (N_1239,In_584,In_731);
nand U1240 (N_1240,In_240,In_171);
and U1241 (N_1241,In_182,In_115);
or U1242 (N_1242,In_648,In_743);
xnor U1243 (N_1243,In_32,In_129);
nand U1244 (N_1244,In_84,In_748);
nand U1245 (N_1245,In_279,In_714);
and U1246 (N_1246,In_737,In_15);
nand U1247 (N_1247,In_402,In_673);
nand U1248 (N_1248,In_739,In_176);
nor U1249 (N_1249,In_212,In_44);
nand U1250 (N_1250,In_129,In_599);
or U1251 (N_1251,In_667,In_571);
or U1252 (N_1252,In_95,In_370);
xnor U1253 (N_1253,In_749,In_259);
or U1254 (N_1254,In_603,In_140);
and U1255 (N_1255,In_743,In_373);
or U1256 (N_1256,In_459,In_590);
xor U1257 (N_1257,In_418,In_745);
xor U1258 (N_1258,In_304,In_127);
and U1259 (N_1259,In_511,In_592);
and U1260 (N_1260,In_210,In_316);
or U1261 (N_1261,In_438,In_494);
xnor U1262 (N_1262,In_592,In_39);
xor U1263 (N_1263,In_486,In_576);
or U1264 (N_1264,In_486,In_327);
nand U1265 (N_1265,In_299,In_485);
nand U1266 (N_1266,In_342,In_210);
or U1267 (N_1267,In_625,In_576);
and U1268 (N_1268,In_179,In_332);
nor U1269 (N_1269,In_542,In_699);
and U1270 (N_1270,In_576,In_54);
xnor U1271 (N_1271,In_46,In_98);
nor U1272 (N_1272,In_455,In_634);
nor U1273 (N_1273,In_689,In_514);
and U1274 (N_1274,In_55,In_741);
nor U1275 (N_1275,In_509,In_694);
nand U1276 (N_1276,In_87,In_383);
nor U1277 (N_1277,In_250,In_661);
nor U1278 (N_1278,In_390,In_489);
xnor U1279 (N_1279,In_326,In_588);
nand U1280 (N_1280,In_292,In_409);
nand U1281 (N_1281,In_349,In_695);
and U1282 (N_1282,In_523,In_487);
nor U1283 (N_1283,In_530,In_12);
xnor U1284 (N_1284,In_2,In_472);
nor U1285 (N_1285,In_746,In_328);
nand U1286 (N_1286,In_742,In_276);
and U1287 (N_1287,In_588,In_640);
or U1288 (N_1288,In_575,In_74);
and U1289 (N_1289,In_286,In_118);
nand U1290 (N_1290,In_503,In_206);
and U1291 (N_1291,In_602,In_721);
nand U1292 (N_1292,In_46,In_246);
or U1293 (N_1293,In_240,In_436);
and U1294 (N_1294,In_368,In_113);
or U1295 (N_1295,In_528,In_725);
nand U1296 (N_1296,In_381,In_680);
xor U1297 (N_1297,In_419,In_597);
or U1298 (N_1298,In_695,In_16);
nor U1299 (N_1299,In_506,In_153);
xor U1300 (N_1300,In_5,In_744);
or U1301 (N_1301,In_65,In_109);
or U1302 (N_1302,In_601,In_220);
nor U1303 (N_1303,In_488,In_596);
nand U1304 (N_1304,In_692,In_648);
nor U1305 (N_1305,In_583,In_98);
and U1306 (N_1306,In_174,In_308);
nand U1307 (N_1307,In_420,In_193);
or U1308 (N_1308,In_211,In_93);
nor U1309 (N_1309,In_471,In_289);
nand U1310 (N_1310,In_284,In_549);
or U1311 (N_1311,In_703,In_611);
xnor U1312 (N_1312,In_553,In_567);
xnor U1313 (N_1313,In_473,In_289);
nor U1314 (N_1314,In_37,In_274);
nand U1315 (N_1315,In_740,In_609);
and U1316 (N_1316,In_618,In_445);
nor U1317 (N_1317,In_107,In_300);
xnor U1318 (N_1318,In_631,In_664);
nor U1319 (N_1319,In_615,In_603);
nand U1320 (N_1320,In_536,In_238);
xnor U1321 (N_1321,In_251,In_436);
and U1322 (N_1322,In_407,In_333);
nand U1323 (N_1323,In_744,In_206);
and U1324 (N_1324,In_672,In_721);
and U1325 (N_1325,In_645,In_444);
xor U1326 (N_1326,In_52,In_421);
and U1327 (N_1327,In_362,In_706);
or U1328 (N_1328,In_671,In_8);
and U1329 (N_1329,In_592,In_308);
and U1330 (N_1330,In_386,In_398);
nor U1331 (N_1331,In_15,In_600);
xor U1332 (N_1332,In_634,In_535);
xor U1333 (N_1333,In_336,In_410);
and U1334 (N_1334,In_631,In_70);
and U1335 (N_1335,In_457,In_740);
or U1336 (N_1336,In_265,In_2);
nand U1337 (N_1337,In_184,In_83);
xnor U1338 (N_1338,In_326,In_695);
or U1339 (N_1339,In_401,In_411);
xnor U1340 (N_1340,In_248,In_662);
nor U1341 (N_1341,In_720,In_676);
xor U1342 (N_1342,In_75,In_108);
nor U1343 (N_1343,In_552,In_108);
and U1344 (N_1344,In_566,In_571);
and U1345 (N_1345,In_301,In_83);
or U1346 (N_1346,In_464,In_557);
nor U1347 (N_1347,In_70,In_709);
nor U1348 (N_1348,In_485,In_197);
nor U1349 (N_1349,In_305,In_202);
nor U1350 (N_1350,In_458,In_507);
and U1351 (N_1351,In_736,In_155);
nand U1352 (N_1352,In_92,In_533);
nor U1353 (N_1353,In_590,In_339);
or U1354 (N_1354,In_584,In_334);
nand U1355 (N_1355,In_662,In_724);
nor U1356 (N_1356,In_306,In_746);
nor U1357 (N_1357,In_537,In_137);
xnor U1358 (N_1358,In_203,In_506);
xor U1359 (N_1359,In_559,In_370);
nor U1360 (N_1360,In_675,In_605);
nand U1361 (N_1361,In_285,In_212);
or U1362 (N_1362,In_469,In_514);
or U1363 (N_1363,In_638,In_362);
nand U1364 (N_1364,In_670,In_340);
xnor U1365 (N_1365,In_442,In_556);
or U1366 (N_1366,In_87,In_240);
xnor U1367 (N_1367,In_627,In_264);
nor U1368 (N_1368,In_289,In_717);
or U1369 (N_1369,In_252,In_399);
nand U1370 (N_1370,In_502,In_472);
xnor U1371 (N_1371,In_685,In_410);
or U1372 (N_1372,In_143,In_179);
and U1373 (N_1373,In_641,In_434);
nor U1374 (N_1374,In_429,In_263);
nand U1375 (N_1375,In_729,In_728);
xnor U1376 (N_1376,In_18,In_88);
or U1377 (N_1377,In_613,In_399);
nand U1378 (N_1378,In_599,In_344);
xnor U1379 (N_1379,In_394,In_90);
nand U1380 (N_1380,In_137,In_318);
nand U1381 (N_1381,In_150,In_288);
xnor U1382 (N_1382,In_416,In_705);
or U1383 (N_1383,In_8,In_14);
xor U1384 (N_1384,In_85,In_40);
nor U1385 (N_1385,In_399,In_393);
or U1386 (N_1386,In_272,In_583);
and U1387 (N_1387,In_628,In_66);
or U1388 (N_1388,In_205,In_509);
nor U1389 (N_1389,In_483,In_311);
and U1390 (N_1390,In_556,In_126);
or U1391 (N_1391,In_91,In_628);
or U1392 (N_1392,In_342,In_284);
nor U1393 (N_1393,In_455,In_422);
xnor U1394 (N_1394,In_145,In_254);
and U1395 (N_1395,In_688,In_181);
nor U1396 (N_1396,In_538,In_232);
nor U1397 (N_1397,In_194,In_527);
and U1398 (N_1398,In_445,In_170);
nor U1399 (N_1399,In_354,In_480);
nand U1400 (N_1400,In_729,In_499);
xor U1401 (N_1401,In_66,In_682);
xnor U1402 (N_1402,In_392,In_304);
nor U1403 (N_1403,In_680,In_553);
nor U1404 (N_1404,In_174,In_711);
or U1405 (N_1405,In_613,In_154);
or U1406 (N_1406,In_587,In_82);
or U1407 (N_1407,In_215,In_443);
xnor U1408 (N_1408,In_709,In_527);
xor U1409 (N_1409,In_464,In_319);
and U1410 (N_1410,In_214,In_647);
nor U1411 (N_1411,In_714,In_389);
or U1412 (N_1412,In_193,In_552);
xnor U1413 (N_1413,In_385,In_503);
nor U1414 (N_1414,In_567,In_82);
nand U1415 (N_1415,In_640,In_416);
nand U1416 (N_1416,In_1,In_414);
nor U1417 (N_1417,In_380,In_478);
nor U1418 (N_1418,In_143,In_552);
and U1419 (N_1419,In_492,In_172);
or U1420 (N_1420,In_313,In_340);
and U1421 (N_1421,In_521,In_482);
nor U1422 (N_1422,In_180,In_597);
nor U1423 (N_1423,In_715,In_646);
xnor U1424 (N_1424,In_85,In_611);
and U1425 (N_1425,In_131,In_657);
or U1426 (N_1426,In_24,In_103);
nand U1427 (N_1427,In_263,In_567);
nand U1428 (N_1428,In_344,In_511);
nand U1429 (N_1429,In_573,In_501);
nor U1430 (N_1430,In_460,In_449);
nand U1431 (N_1431,In_213,In_22);
nor U1432 (N_1432,In_335,In_40);
xnor U1433 (N_1433,In_252,In_269);
xnor U1434 (N_1434,In_408,In_17);
and U1435 (N_1435,In_353,In_175);
and U1436 (N_1436,In_35,In_556);
or U1437 (N_1437,In_191,In_327);
nor U1438 (N_1438,In_412,In_229);
xor U1439 (N_1439,In_692,In_571);
nand U1440 (N_1440,In_373,In_261);
or U1441 (N_1441,In_77,In_395);
xnor U1442 (N_1442,In_335,In_460);
nor U1443 (N_1443,In_705,In_491);
xnor U1444 (N_1444,In_227,In_697);
xor U1445 (N_1445,In_89,In_134);
nand U1446 (N_1446,In_710,In_64);
and U1447 (N_1447,In_423,In_484);
nand U1448 (N_1448,In_189,In_356);
and U1449 (N_1449,In_71,In_709);
xor U1450 (N_1450,In_347,In_142);
nor U1451 (N_1451,In_329,In_206);
or U1452 (N_1452,In_360,In_732);
xnor U1453 (N_1453,In_386,In_629);
xnor U1454 (N_1454,In_128,In_494);
or U1455 (N_1455,In_455,In_207);
xor U1456 (N_1456,In_510,In_276);
nor U1457 (N_1457,In_414,In_408);
nor U1458 (N_1458,In_334,In_563);
nor U1459 (N_1459,In_64,In_656);
or U1460 (N_1460,In_741,In_117);
or U1461 (N_1461,In_73,In_48);
and U1462 (N_1462,In_286,In_259);
or U1463 (N_1463,In_214,In_490);
and U1464 (N_1464,In_135,In_91);
and U1465 (N_1465,In_594,In_304);
nand U1466 (N_1466,In_486,In_60);
and U1467 (N_1467,In_609,In_590);
xor U1468 (N_1468,In_627,In_67);
and U1469 (N_1469,In_317,In_352);
nor U1470 (N_1470,In_243,In_439);
or U1471 (N_1471,In_144,In_106);
nand U1472 (N_1472,In_446,In_704);
xnor U1473 (N_1473,In_3,In_347);
and U1474 (N_1474,In_396,In_56);
or U1475 (N_1475,In_315,In_503);
nor U1476 (N_1476,In_145,In_186);
and U1477 (N_1477,In_479,In_464);
or U1478 (N_1478,In_498,In_723);
nand U1479 (N_1479,In_733,In_736);
and U1480 (N_1480,In_644,In_508);
xor U1481 (N_1481,In_335,In_478);
or U1482 (N_1482,In_124,In_418);
and U1483 (N_1483,In_354,In_286);
xnor U1484 (N_1484,In_677,In_662);
or U1485 (N_1485,In_709,In_255);
and U1486 (N_1486,In_734,In_188);
or U1487 (N_1487,In_191,In_338);
nand U1488 (N_1488,In_421,In_106);
nand U1489 (N_1489,In_474,In_436);
and U1490 (N_1490,In_518,In_684);
xnor U1491 (N_1491,In_220,In_73);
nor U1492 (N_1492,In_186,In_492);
xnor U1493 (N_1493,In_561,In_582);
nand U1494 (N_1494,In_569,In_34);
and U1495 (N_1495,In_365,In_156);
nor U1496 (N_1496,In_7,In_340);
nand U1497 (N_1497,In_106,In_108);
nand U1498 (N_1498,In_85,In_155);
xor U1499 (N_1499,In_616,In_517);
nand U1500 (N_1500,In_398,In_357);
xnor U1501 (N_1501,In_17,In_264);
nand U1502 (N_1502,In_245,In_395);
and U1503 (N_1503,In_174,In_91);
and U1504 (N_1504,In_137,In_735);
nand U1505 (N_1505,In_647,In_87);
nor U1506 (N_1506,In_724,In_403);
and U1507 (N_1507,In_441,In_77);
xnor U1508 (N_1508,In_694,In_253);
nor U1509 (N_1509,In_564,In_162);
nor U1510 (N_1510,In_219,In_513);
or U1511 (N_1511,In_110,In_508);
nand U1512 (N_1512,In_255,In_223);
and U1513 (N_1513,In_536,In_468);
xor U1514 (N_1514,In_626,In_222);
xor U1515 (N_1515,In_436,In_665);
and U1516 (N_1516,In_299,In_201);
nand U1517 (N_1517,In_117,In_628);
and U1518 (N_1518,In_104,In_24);
xnor U1519 (N_1519,In_398,In_3);
and U1520 (N_1520,In_12,In_718);
nor U1521 (N_1521,In_459,In_222);
nor U1522 (N_1522,In_185,In_209);
nor U1523 (N_1523,In_625,In_598);
xnor U1524 (N_1524,In_31,In_29);
or U1525 (N_1525,In_621,In_398);
nor U1526 (N_1526,In_49,In_734);
xor U1527 (N_1527,In_142,In_167);
xnor U1528 (N_1528,In_211,In_646);
nor U1529 (N_1529,In_225,In_220);
xor U1530 (N_1530,In_584,In_442);
and U1531 (N_1531,In_37,In_713);
xnor U1532 (N_1532,In_59,In_443);
nand U1533 (N_1533,In_226,In_127);
nor U1534 (N_1534,In_271,In_298);
xnor U1535 (N_1535,In_408,In_77);
nor U1536 (N_1536,In_238,In_359);
nor U1537 (N_1537,In_182,In_85);
and U1538 (N_1538,In_593,In_317);
nand U1539 (N_1539,In_200,In_342);
and U1540 (N_1540,In_116,In_340);
xnor U1541 (N_1541,In_581,In_686);
xor U1542 (N_1542,In_462,In_359);
and U1543 (N_1543,In_257,In_537);
and U1544 (N_1544,In_523,In_615);
xor U1545 (N_1545,In_590,In_434);
xor U1546 (N_1546,In_666,In_413);
nand U1547 (N_1547,In_333,In_341);
nand U1548 (N_1548,In_451,In_550);
nor U1549 (N_1549,In_237,In_63);
xnor U1550 (N_1550,In_232,In_714);
or U1551 (N_1551,In_733,In_472);
nand U1552 (N_1552,In_690,In_658);
or U1553 (N_1553,In_183,In_204);
or U1554 (N_1554,In_449,In_745);
nand U1555 (N_1555,In_171,In_322);
and U1556 (N_1556,In_59,In_107);
nor U1557 (N_1557,In_569,In_457);
and U1558 (N_1558,In_22,In_211);
nand U1559 (N_1559,In_20,In_487);
and U1560 (N_1560,In_382,In_168);
or U1561 (N_1561,In_592,In_703);
xnor U1562 (N_1562,In_631,In_489);
xnor U1563 (N_1563,In_544,In_310);
or U1564 (N_1564,In_247,In_736);
nor U1565 (N_1565,In_748,In_213);
or U1566 (N_1566,In_336,In_676);
or U1567 (N_1567,In_27,In_21);
xor U1568 (N_1568,In_703,In_488);
and U1569 (N_1569,In_391,In_644);
xnor U1570 (N_1570,In_79,In_168);
or U1571 (N_1571,In_115,In_78);
nor U1572 (N_1572,In_712,In_182);
xor U1573 (N_1573,In_534,In_639);
nor U1574 (N_1574,In_715,In_289);
xor U1575 (N_1575,In_521,In_167);
and U1576 (N_1576,In_353,In_570);
xor U1577 (N_1577,In_686,In_523);
nor U1578 (N_1578,In_119,In_743);
and U1579 (N_1579,In_50,In_500);
and U1580 (N_1580,In_584,In_336);
or U1581 (N_1581,In_450,In_118);
nand U1582 (N_1582,In_15,In_667);
nor U1583 (N_1583,In_348,In_747);
nor U1584 (N_1584,In_717,In_438);
xnor U1585 (N_1585,In_227,In_346);
nor U1586 (N_1586,In_73,In_180);
or U1587 (N_1587,In_391,In_510);
and U1588 (N_1588,In_251,In_326);
or U1589 (N_1589,In_592,In_60);
or U1590 (N_1590,In_262,In_651);
xor U1591 (N_1591,In_191,In_289);
nand U1592 (N_1592,In_546,In_218);
and U1593 (N_1593,In_462,In_455);
and U1594 (N_1594,In_460,In_603);
nor U1595 (N_1595,In_712,In_102);
or U1596 (N_1596,In_122,In_270);
nand U1597 (N_1597,In_460,In_595);
or U1598 (N_1598,In_258,In_443);
nand U1599 (N_1599,In_64,In_409);
nor U1600 (N_1600,In_154,In_642);
xor U1601 (N_1601,In_441,In_657);
nand U1602 (N_1602,In_608,In_498);
nand U1603 (N_1603,In_642,In_507);
or U1604 (N_1604,In_243,In_587);
or U1605 (N_1605,In_525,In_464);
or U1606 (N_1606,In_658,In_6);
nand U1607 (N_1607,In_157,In_18);
or U1608 (N_1608,In_543,In_29);
xor U1609 (N_1609,In_528,In_271);
and U1610 (N_1610,In_667,In_141);
and U1611 (N_1611,In_488,In_641);
nand U1612 (N_1612,In_477,In_677);
or U1613 (N_1613,In_607,In_448);
xor U1614 (N_1614,In_496,In_744);
nor U1615 (N_1615,In_132,In_1);
or U1616 (N_1616,In_316,In_402);
xor U1617 (N_1617,In_71,In_446);
nor U1618 (N_1618,In_563,In_260);
or U1619 (N_1619,In_506,In_368);
or U1620 (N_1620,In_612,In_246);
nand U1621 (N_1621,In_477,In_644);
xnor U1622 (N_1622,In_603,In_240);
nor U1623 (N_1623,In_233,In_318);
nor U1624 (N_1624,In_695,In_500);
and U1625 (N_1625,In_589,In_712);
or U1626 (N_1626,In_658,In_340);
or U1627 (N_1627,In_56,In_156);
and U1628 (N_1628,In_431,In_83);
and U1629 (N_1629,In_354,In_160);
or U1630 (N_1630,In_509,In_26);
and U1631 (N_1631,In_658,In_533);
nor U1632 (N_1632,In_71,In_42);
nand U1633 (N_1633,In_426,In_92);
or U1634 (N_1634,In_442,In_186);
xor U1635 (N_1635,In_411,In_243);
or U1636 (N_1636,In_623,In_588);
or U1637 (N_1637,In_56,In_622);
and U1638 (N_1638,In_601,In_605);
nand U1639 (N_1639,In_627,In_373);
nand U1640 (N_1640,In_208,In_424);
nor U1641 (N_1641,In_361,In_232);
or U1642 (N_1642,In_211,In_537);
nand U1643 (N_1643,In_690,In_115);
nor U1644 (N_1644,In_392,In_544);
and U1645 (N_1645,In_329,In_563);
nor U1646 (N_1646,In_656,In_705);
nand U1647 (N_1647,In_444,In_393);
nor U1648 (N_1648,In_239,In_257);
xnor U1649 (N_1649,In_119,In_242);
and U1650 (N_1650,In_645,In_36);
nor U1651 (N_1651,In_513,In_278);
or U1652 (N_1652,In_104,In_564);
nand U1653 (N_1653,In_455,In_620);
nand U1654 (N_1654,In_262,In_95);
or U1655 (N_1655,In_322,In_541);
or U1656 (N_1656,In_156,In_409);
nor U1657 (N_1657,In_279,In_351);
xnor U1658 (N_1658,In_373,In_259);
or U1659 (N_1659,In_317,In_695);
or U1660 (N_1660,In_354,In_442);
xnor U1661 (N_1661,In_622,In_288);
xnor U1662 (N_1662,In_581,In_466);
xnor U1663 (N_1663,In_128,In_549);
and U1664 (N_1664,In_497,In_558);
nor U1665 (N_1665,In_337,In_199);
nand U1666 (N_1666,In_547,In_515);
or U1667 (N_1667,In_227,In_596);
nor U1668 (N_1668,In_36,In_218);
nand U1669 (N_1669,In_313,In_152);
nor U1670 (N_1670,In_157,In_3);
xor U1671 (N_1671,In_550,In_601);
xor U1672 (N_1672,In_438,In_650);
nor U1673 (N_1673,In_520,In_162);
nor U1674 (N_1674,In_11,In_316);
xor U1675 (N_1675,In_325,In_732);
xnor U1676 (N_1676,In_78,In_30);
or U1677 (N_1677,In_675,In_525);
nor U1678 (N_1678,In_73,In_178);
nor U1679 (N_1679,In_134,In_735);
nand U1680 (N_1680,In_22,In_442);
and U1681 (N_1681,In_488,In_70);
and U1682 (N_1682,In_166,In_19);
and U1683 (N_1683,In_524,In_241);
and U1684 (N_1684,In_513,In_397);
nor U1685 (N_1685,In_28,In_602);
xor U1686 (N_1686,In_284,In_151);
xor U1687 (N_1687,In_547,In_296);
nand U1688 (N_1688,In_196,In_465);
nand U1689 (N_1689,In_43,In_542);
and U1690 (N_1690,In_292,In_469);
or U1691 (N_1691,In_583,In_689);
xor U1692 (N_1692,In_14,In_292);
xnor U1693 (N_1693,In_444,In_590);
nor U1694 (N_1694,In_333,In_365);
xnor U1695 (N_1695,In_348,In_702);
or U1696 (N_1696,In_675,In_116);
or U1697 (N_1697,In_83,In_380);
or U1698 (N_1698,In_546,In_217);
xnor U1699 (N_1699,In_386,In_221);
xor U1700 (N_1700,In_271,In_267);
xor U1701 (N_1701,In_45,In_152);
xnor U1702 (N_1702,In_469,In_710);
xnor U1703 (N_1703,In_129,In_467);
nor U1704 (N_1704,In_35,In_96);
xor U1705 (N_1705,In_155,In_3);
or U1706 (N_1706,In_658,In_411);
or U1707 (N_1707,In_74,In_47);
nand U1708 (N_1708,In_178,In_171);
and U1709 (N_1709,In_674,In_712);
nand U1710 (N_1710,In_483,In_657);
and U1711 (N_1711,In_184,In_714);
nand U1712 (N_1712,In_645,In_594);
nand U1713 (N_1713,In_204,In_132);
nor U1714 (N_1714,In_716,In_652);
xor U1715 (N_1715,In_123,In_159);
nor U1716 (N_1716,In_28,In_40);
nand U1717 (N_1717,In_229,In_737);
xor U1718 (N_1718,In_332,In_662);
nor U1719 (N_1719,In_302,In_534);
xor U1720 (N_1720,In_471,In_468);
or U1721 (N_1721,In_341,In_736);
or U1722 (N_1722,In_516,In_717);
and U1723 (N_1723,In_517,In_88);
or U1724 (N_1724,In_563,In_688);
or U1725 (N_1725,In_542,In_82);
nor U1726 (N_1726,In_453,In_536);
nand U1727 (N_1727,In_69,In_96);
nand U1728 (N_1728,In_178,In_22);
nand U1729 (N_1729,In_195,In_13);
nor U1730 (N_1730,In_431,In_518);
xnor U1731 (N_1731,In_536,In_134);
or U1732 (N_1732,In_347,In_161);
and U1733 (N_1733,In_196,In_353);
xnor U1734 (N_1734,In_680,In_437);
nand U1735 (N_1735,In_430,In_10);
or U1736 (N_1736,In_153,In_373);
and U1737 (N_1737,In_271,In_427);
or U1738 (N_1738,In_63,In_83);
or U1739 (N_1739,In_73,In_11);
and U1740 (N_1740,In_456,In_122);
or U1741 (N_1741,In_336,In_306);
or U1742 (N_1742,In_251,In_644);
nand U1743 (N_1743,In_57,In_303);
xor U1744 (N_1744,In_100,In_473);
or U1745 (N_1745,In_246,In_740);
and U1746 (N_1746,In_601,In_291);
xnor U1747 (N_1747,In_362,In_417);
xnor U1748 (N_1748,In_77,In_527);
and U1749 (N_1749,In_362,In_384);
nand U1750 (N_1750,In_659,In_686);
xnor U1751 (N_1751,In_619,In_615);
nand U1752 (N_1752,In_222,In_438);
and U1753 (N_1753,In_283,In_109);
nand U1754 (N_1754,In_395,In_33);
or U1755 (N_1755,In_720,In_279);
nand U1756 (N_1756,In_414,In_731);
xor U1757 (N_1757,In_681,In_289);
nor U1758 (N_1758,In_8,In_190);
and U1759 (N_1759,In_570,In_380);
or U1760 (N_1760,In_634,In_226);
and U1761 (N_1761,In_454,In_490);
and U1762 (N_1762,In_316,In_724);
and U1763 (N_1763,In_676,In_661);
xor U1764 (N_1764,In_607,In_736);
and U1765 (N_1765,In_98,In_653);
and U1766 (N_1766,In_563,In_436);
nand U1767 (N_1767,In_353,In_317);
nor U1768 (N_1768,In_353,In_35);
xor U1769 (N_1769,In_207,In_701);
nand U1770 (N_1770,In_641,In_179);
or U1771 (N_1771,In_124,In_402);
xnor U1772 (N_1772,In_712,In_297);
nand U1773 (N_1773,In_706,In_38);
xnor U1774 (N_1774,In_279,In_310);
and U1775 (N_1775,In_166,In_384);
and U1776 (N_1776,In_190,In_531);
nand U1777 (N_1777,In_305,In_408);
and U1778 (N_1778,In_228,In_246);
xnor U1779 (N_1779,In_493,In_383);
xor U1780 (N_1780,In_622,In_235);
nand U1781 (N_1781,In_46,In_632);
or U1782 (N_1782,In_34,In_10);
and U1783 (N_1783,In_305,In_500);
or U1784 (N_1784,In_439,In_647);
xnor U1785 (N_1785,In_38,In_162);
nor U1786 (N_1786,In_178,In_305);
nor U1787 (N_1787,In_184,In_52);
xnor U1788 (N_1788,In_468,In_741);
nor U1789 (N_1789,In_348,In_649);
and U1790 (N_1790,In_217,In_278);
nor U1791 (N_1791,In_53,In_684);
nor U1792 (N_1792,In_446,In_435);
xor U1793 (N_1793,In_351,In_246);
or U1794 (N_1794,In_462,In_681);
and U1795 (N_1795,In_581,In_435);
or U1796 (N_1796,In_451,In_248);
or U1797 (N_1797,In_315,In_425);
nor U1798 (N_1798,In_160,In_102);
nor U1799 (N_1799,In_557,In_524);
or U1800 (N_1800,In_341,In_129);
and U1801 (N_1801,In_647,In_157);
and U1802 (N_1802,In_398,In_598);
nand U1803 (N_1803,In_18,In_536);
or U1804 (N_1804,In_659,In_246);
nor U1805 (N_1805,In_353,In_43);
xnor U1806 (N_1806,In_461,In_412);
xor U1807 (N_1807,In_585,In_646);
nor U1808 (N_1808,In_46,In_35);
nand U1809 (N_1809,In_623,In_6);
xor U1810 (N_1810,In_32,In_737);
or U1811 (N_1811,In_416,In_562);
xor U1812 (N_1812,In_56,In_164);
and U1813 (N_1813,In_620,In_77);
and U1814 (N_1814,In_159,In_648);
or U1815 (N_1815,In_516,In_313);
or U1816 (N_1816,In_452,In_388);
or U1817 (N_1817,In_594,In_442);
and U1818 (N_1818,In_408,In_55);
or U1819 (N_1819,In_321,In_379);
and U1820 (N_1820,In_180,In_13);
and U1821 (N_1821,In_314,In_344);
or U1822 (N_1822,In_526,In_124);
or U1823 (N_1823,In_572,In_429);
nor U1824 (N_1824,In_400,In_152);
nor U1825 (N_1825,In_507,In_583);
nor U1826 (N_1826,In_591,In_283);
xor U1827 (N_1827,In_720,In_282);
xor U1828 (N_1828,In_494,In_196);
nand U1829 (N_1829,In_25,In_197);
nand U1830 (N_1830,In_556,In_699);
nand U1831 (N_1831,In_700,In_221);
nor U1832 (N_1832,In_252,In_258);
nand U1833 (N_1833,In_613,In_0);
or U1834 (N_1834,In_621,In_166);
nor U1835 (N_1835,In_153,In_484);
and U1836 (N_1836,In_363,In_186);
nand U1837 (N_1837,In_704,In_195);
xor U1838 (N_1838,In_578,In_205);
nand U1839 (N_1839,In_439,In_464);
and U1840 (N_1840,In_45,In_444);
or U1841 (N_1841,In_415,In_608);
nand U1842 (N_1842,In_716,In_692);
nand U1843 (N_1843,In_58,In_434);
xnor U1844 (N_1844,In_136,In_76);
xnor U1845 (N_1845,In_447,In_413);
xnor U1846 (N_1846,In_484,In_491);
nor U1847 (N_1847,In_64,In_347);
and U1848 (N_1848,In_701,In_660);
and U1849 (N_1849,In_72,In_335);
nor U1850 (N_1850,In_136,In_189);
xor U1851 (N_1851,In_298,In_447);
or U1852 (N_1852,In_39,In_458);
and U1853 (N_1853,In_516,In_155);
or U1854 (N_1854,In_384,In_640);
nand U1855 (N_1855,In_546,In_649);
nor U1856 (N_1856,In_240,In_209);
nor U1857 (N_1857,In_528,In_651);
xnor U1858 (N_1858,In_479,In_164);
and U1859 (N_1859,In_707,In_382);
or U1860 (N_1860,In_732,In_703);
nor U1861 (N_1861,In_264,In_177);
nor U1862 (N_1862,In_735,In_241);
nand U1863 (N_1863,In_12,In_182);
xnor U1864 (N_1864,In_627,In_522);
and U1865 (N_1865,In_6,In_266);
or U1866 (N_1866,In_600,In_21);
or U1867 (N_1867,In_456,In_143);
xnor U1868 (N_1868,In_544,In_327);
nor U1869 (N_1869,In_620,In_331);
and U1870 (N_1870,In_270,In_242);
nor U1871 (N_1871,In_506,In_691);
or U1872 (N_1872,In_84,In_711);
nor U1873 (N_1873,In_726,In_651);
nor U1874 (N_1874,In_672,In_59);
xnor U1875 (N_1875,In_6,In_669);
and U1876 (N_1876,In_233,In_78);
or U1877 (N_1877,In_399,In_259);
or U1878 (N_1878,In_321,In_281);
nand U1879 (N_1879,In_192,In_154);
nor U1880 (N_1880,In_221,In_584);
and U1881 (N_1881,In_401,In_665);
nand U1882 (N_1882,In_473,In_677);
nand U1883 (N_1883,In_236,In_208);
nand U1884 (N_1884,In_381,In_91);
nor U1885 (N_1885,In_345,In_234);
nor U1886 (N_1886,In_76,In_106);
or U1887 (N_1887,In_432,In_233);
and U1888 (N_1888,In_528,In_199);
and U1889 (N_1889,In_314,In_101);
nor U1890 (N_1890,In_65,In_476);
or U1891 (N_1891,In_457,In_35);
and U1892 (N_1892,In_288,In_414);
xor U1893 (N_1893,In_16,In_532);
xnor U1894 (N_1894,In_624,In_451);
and U1895 (N_1895,In_554,In_148);
nand U1896 (N_1896,In_677,In_249);
nor U1897 (N_1897,In_35,In_354);
xnor U1898 (N_1898,In_308,In_212);
or U1899 (N_1899,In_36,In_526);
and U1900 (N_1900,In_156,In_485);
or U1901 (N_1901,In_33,In_535);
xnor U1902 (N_1902,In_730,In_708);
and U1903 (N_1903,In_342,In_676);
nand U1904 (N_1904,In_137,In_165);
xnor U1905 (N_1905,In_161,In_568);
or U1906 (N_1906,In_122,In_32);
nor U1907 (N_1907,In_591,In_563);
nand U1908 (N_1908,In_569,In_733);
and U1909 (N_1909,In_272,In_290);
or U1910 (N_1910,In_119,In_590);
and U1911 (N_1911,In_76,In_93);
nor U1912 (N_1912,In_10,In_626);
nand U1913 (N_1913,In_243,In_16);
nor U1914 (N_1914,In_502,In_303);
nor U1915 (N_1915,In_605,In_513);
xnor U1916 (N_1916,In_191,In_115);
and U1917 (N_1917,In_229,In_388);
nand U1918 (N_1918,In_377,In_96);
or U1919 (N_1919,In_357,In_653);
nand U1920 (N_1920,In_677,In_531);
and U1921 (N_1921,In_622,In_657);
nand U1922 (N_1922,In_4,In_721);
and U1923 (N_1923,In_36,In_1);
nand U1924 (N_1924,In_313,In_289);
nor U1925 (N_1925,In_500,In_506);
or U1926 (N_1926,In_595,In_641);
or U1927 (N_1927,In_239,In_504);
nor U1928 (N_1928,In_34,In_272);
or U1929 (N_1929,In_176,In_124);
xor U1930 (N_1930,In_713,In_366);
and U1931 (N_1931,In_634,In_258);
xor U1932 (N_1932,In_31,In_309);
or U1933 (N_1933,In_466,In_704);
or U1934 (N_1934,In_655,In_446);
and U1935 (N_1935,In_182,In_622);
nand U1936 (N_1936,In_398,In_432);
or U1937 (N_1937,In_270,In_292);
nor U1938 (N_1938,In_482,In_601);
or U1939 (N_1939,In_46,In_740);
and U1940 (N_1940,In_692,In_318);
nor U1941 (N_1941,In_604,In_334);
and U1942 (N_1942,In_615,In_673);
nand U1943 (N_1943,In_375,In_509);
xnor U1944 (N_1944,In_566,In_125);
and U1945 (N_1945,In_231,In_133);
or U1946 (N_1946,In_114,In_708);
nor U1947 (N_1947,In_63,In_113);
xor U1948 (N_1948,In_234,In_313);
xor U1949 (N_1949,In_348,In_128);
and U1950 (N_1950,In_435,In_262);
and U1951 (N_1951,In_644,In_195);
or U1952 (N_1952,In_587,In_101);
and U1953 (N_1953,In_78,In_109);
nor U1954 (N_1954,In_492,In_314);
and U1955 (N_1955,In_42,In_114);
nor U1956 (N_1956,In_694,In_511);
nor U1957 (N_1957,In_657,In_507);
nand U1958 (N_1958,In_209,In_564);
nor U1959 (N_1959,In_447,In_594);
and U1960 (N_1960,In_449,In_61);
xnor U1961 (N_1961,In_84,In_235);
or U1962 (N_1962,In_200,In_128);
or U1963 (N_1963,In_90,In_210);
nor U1964 (N_1964,In_447,In_739);
xnor U1965 (N_1965,In_625,In_685);
nor U1966 (N_1966,In_101,In_651);
xnor U1967 (N_1967,In_677,In_45);
xor U1968 (N_1968,In_598,In_666);
xnor U1969 (N_1969,In_572,In_161);
nand U1970 (N_1970,In_723,In_615);
nor U1971 (N_1971,In_620,In_212);
nor U1972 (N_1972,In_451,In_336);
xor U1973 (N_1973,In_309,In_196);
xor U1974 (N_1974,In_35,In_246);
or U1975 (N_1975,In_35,In_728);
nand U1976 (N_1976,In_85,In_422);
or U1977 (N_1977,In_705,In_282);
nor U1978 (N_1978,In_343,In_640);
nand U1979 (N_1979,In_488,In_299);
nand U1980 (N_1980,In_457,In_166);
and U1981 (N_1981,In_249,In_399);
nand U1982 (N_1982,In_198,In_99);
nand U1983 (N_1983,In_516,In_295);
and U1984 (N_1984,In_515,In_451);
or U1985 (N_1985,In_475,In_471);
nor U1986 (N_1986,In_295,In_5);
xor U1987 (N_1987,In_386,In_37);
or U1988 (N_1988,In_674,In_203);
nor U1989 (N_1989,In_179,In_202);
or U1990 (N_1990,In_542,In_216);
nand U1991 (N_1991,In_166,In_175);
or U1992 (N_1992,In_373,In_247);
nand U1993 (N_1993,In_719,In_136);
nand U1994 (N_1994,In_647,In_285);
nand U1995 (N_1995,In_467,In_525);
nand U1996 (N_1996,In_545,In_563);
and U1997 (N_1997,In_607,In_104);
and U1998 (N_1998,In_145,In_0);
or U1999 (N_1999,In_31,In_130);
nand U2000 (N_2000,In_128,In_219);
nand U2001 (N_2001,In_748,In_129);
nand U2002 (N_2002,In_414,In_728);
and U2003 (N_2003,In_181,In_501);
xor U2004 (N_2004,In_147,In_697);
and U2005 (N_2005,In_336,In_728);
nand U2006 (N_2006,In_257,In_280);
nor U2007 (N_2007,In_544,In_635);
nand U2008 (N_2008,In_176,In_321);
nand U2009 (N_2009,In_661,In_560);
or U2010 (N_2010,In_161,In_133);
or U2011 (N_2011,In_721,In_536);
or U2012 (N_2012,In_429,In_168);
or U2013 (N_2013,In_290,In_239);
nand U2014 (N_2014,In_371,In_282);
and U2015 (N_2015,In_56,In_57);
and U2016 (N_2016,In_314,In_436);
and U2017 (N_2017,In_680,In_13);
and U2018 (N_2018,In_375,In_584);
or U2019 (N_2019,In_543,In_210);
and U2020 (N_2020,In_70,In_446);
xnor U2021 (N_2021,In_464,In_470);
and U2022 (N_2022,In_97,In_84);
nand U2023 (N_2023,In_309,In_363);
and U2024 (N_2024,In_19,In_719);
xor U2025 (N_2025,In_162,In_688);
and U2026 (N_2026,In_421,In_182);
and U2027 (N_2027,In_194,In_639);
xor U2028 (N_2028,In_546,In_148);
nor U2029 (N_2029,In_643,In_248);
and U2030 (N_2030,In_726,In_454);
xnor U2031 (N_2031,In_694,In_156);
nand U2032 (N_2032,In_289,In_435);
or U2033 (N_2033,In_636,In_571);
and U2034 (N_2034,In_728,In_75);
or U2035 (N_2035,In_202,In_446);
and U2036 (N_2036,In_53,In_172);
xnor U2037 (N_2037,In_204,In_227);
nor U2038 (N_2038,In_251,In_211);
nor U2039 (N_2039,In_252,In_627);
nor U2040 (N_2040,In_395,In_147);
xor U2041 (N_2041,In_575,In_305);
nand U2042 (N_2042,In_696,In_381);
nor U2043 (N_2043,In_713,In_480);
and U2044 (N_2044,In_538,In_746);
or U2045 (N_2045,In_665,In_391);
nor U2046 (N_2046,In_525,In_50);
and U2047 (N_2047,In_289,In_583);
or U2048 (N_2048,In_410,In_294);
nor U2049 (N_2049,In_35,In_363);
and U2050 (N_2050,In_703,In_303);
nor U2051 (N_2051,In_55,In_33);
xor U2052 (N_2052,In_529,In_259);
nand U2053 (N_2053,In_116,In_394);
and U2054 (N_2054,In_241,In_292);
or U2055 (N_2055,In_735,In_726);
xor U2056 (N_2056,In_517,In_695);
nand U2057 (N_2057,In_240,In_722);
xor U2058 (N_2058,In_48,In_348);
nor U2059 (N_2059,In_240,In_466);
and U2060 (N_2060,In_176,In_18);
nor U2061 (N_2061,In_189,In_624);
nor U2062 (N_2062,In_716,In_268);
xor U2063 (N_2063,In_352,In_441);
nor U2064 (N_2064,In_605,In_182);
xnor U2065 (N_2065,In_492,In_211);
or U2066 (N_2066,In_571,In_322);
or U2067 (N_2067,In_679,In_160);
xor U2068 (N_2068,In_364,In_324);
or U2069 (N_2069,In_556,In_665);
or U2070 (N_2070,In_289,In_196);
or U2071 (N_2071,In_681,In_96);
nand U2072 (N_2072,In_215,In_393);
and U2073 (N_2073,In_562,In_444);
nor U2074 (N_2074,In_150,In_724);
xor U2075 (N_2075,In_744,In_351);
nand U2076 (N_2076,In_231,In_715);
nor U2077 (N_2077,In_297,In_663);
and U2078 (N_2078,In_101,In_33);
or U2079 (N_2079,In_733,In_250);
and U2080 (N_2080,In_482,In_416);
xor U2081 (N_2081,In_200,In_616);
xor U2082 (N_2082,In_177,In_685);
and U2083 (N_2083,In_551,In_350);
or U2084 (N_2084,In_626,In_178);
and U2085 (N_2085,In_504,In_476);
nand U2086 (N_2086,In_238,In_126);
or U2087 (N_2087,In_442,In_213);
and U2088 (N_2088,In_695,In_384);
nand U2089 (N_2089,In_566,In_485);
nand U2090 (N_2090,In_94,In_222);
xnor U2091 (N_2091,In_70,In_579);
xnor U2092 (N_2092,In_119,In_289);
and U2093 (N_2093,In_639,In_507);
xor U2094 (N_2094,In_721,In_553);
and U2095 (N_2095,In_568,In_373);
xor U2096 (N_2096,In_73,In_462);
nor U2097 (N_2097,In_221,In_64);
nor U2098 (N_2098,In_280,In_679);
or U2099 (N_2099,In_207,In_558);
xor U2100 (N_2100,In_697,In_128);
nand U2101 (N_2101,In_128,In_56);
xor U2102 (N_2102,In_19,In_614);
nor U2103 (N_2103,In_720,In_697);
xnor U2104 (N_2104,In_590,In_535);
xnor U2105 (N_2105,In_588,In_383);
nand U2106 (N_2106,In_99,In_319);
and U2107 (N_2107,In_113,In_180);
or U2108 (N_2108,In_586,In_643);
xnor U2109 (N_2109,In_363,In_334);
and U2110 (N_2110,In_68,In_574);
nand U2111 (N_2111,In_42,In_351);
and U2112 (N_2112,In_14,In_559);
and U2113 (N_2113,In_288,In_283);
and U2114 (N_2114,In_664,In_720);
xnor U2115 (N_2115,In_449,In_116);
nand U2116 (N_2116,In_686,In_416);
nand U2117 (N_2117,In_26,In_639);
and U2118 (N_2118,In_197,In_616);
nand U2119 (N_2119,In_74,In_601);
or U2120 (N_2120,In_85,In_462);
nor U2121 (N_2121,In_430,In_172);
and U2122 (N_2122,In_435,In_538);
nand U2123 (N_2123,In_266,In_730);
nor U2124 (N_2124,In_126,In_49);
nor U2125 (N_2125,In_195,In_115);
or U2126 (N_2126,In_579,In_37);
and U2127 (N_2127,In_605,In_246);
nand U2128 (N_2128,In_517,In_630);
and U2129 (N_2129,In_515,In_747);
nor U2130 (N_2130,In_9,In_687);
xnor U2131 (N_2131,In_521,In_614);
and U2132 (N_2132,In_240,In_81);
xnor U2133 (N_2133,In_165,In_102);
nor U2134 (N_2134,In_360,In_616);
and U2135 (N_2135,In_448,In_409);
nor U2136 (N_2136,In_194,In_312);
or U2137 (N_2137,In_694,In_722);
nand U2138 (N_2138,In_274,In_692);
or U2139 (N_2139,In_119,In_679);
and U2140 (N_2140,In_132,In_87);
nor U2141 (N_2141,In_610,In_468);
nand U2142 (N_2142,In_427,In_42);
nand U2143 (N_2143,In_234,In_308);
and U2144 (N_2144,In_63,In_182);
nand U2145 (N_2145,In_283,In_238);
nor U2146 (N_2146,In_241,In_48);
nor U2147 (N_2147,In_74,In_696);
or U2148 (N_2148,In_544,In_318);
nand U2149 (N_2149,In_584,In_644);
nor U2150 (N_2150,In_640,In_262);
xnor U2151 (N_2151,In_324,In_332);
nor U2152 (N_2152,In_310,In_369);
nor U2153 (N_2153,In_331,In_621);
or U2154 (N_2154,In_575,In_399);
nor U2155 (N_2155,In_674,In_61);
nand U2156 (N_2156,In_520,In_703);
nor U2157 (N_2157,In_729,In_461);
and U2158 (N_2158,In_358,In_196);
and U2159 (N_2159,In_528,In_0);
or U2160 (N_2160,In_161,In_58);
or U2161 (N_2161,In_530,In_625);
nand U2162 (N_2162,In_717,In_660);
nor U2163 (N_2163,In_519,In_371);
and U2164 (N_2164,In_0,In_531);
nand U2165 (N_2165,In_607,In_484);
or U2166 (N_2166,In_745,In_324);
xnor U2167 (N_2167,In_741,In_408);
xor U2168 (N_2168,In_635,In_658);
nor U2169 (N_2169,In_436,In_486);
or U2170 (N_2170,In_326,In_605);
and U2171 (N_2171,In_301,In_534);
and U2172 (N_2172,In_704,In_730);
nor U2173 (N_2173,In_591,In_128);
xnor U2174 (N_2174,In_396,In_592);
nor U2175 (N_2175,In_95,In_703);
and U2176 (N_2176,In_373,In_336);
and U2177 (N_2177,In_30,In_464);
nor U2178 (N_2178,In_421,In_117);
nand U2179 (N_2179,In_583,In_16);
nor U2180 (N_2180,In_587,In_312);
nor U2181 (N_2181,In_663,In_693);
or U2182 (N_2182,In_296,In_188);
nor U2183 (N_2183,In_728,In_98);
nand U2184 (N_2184,In_552,In_498);
nor U2185 (N_2185,In_301,In_593);
nor U2186 (N_2186,In_684,In_77);
and U2187 (N_2187,In_87,In_733);
and U2188 (N_2188,In_101,In_196);
nor U2189 (N_2189,In_592,In_519);
and U2190 (N_2190,In_483,In_66);
nor U2191 (N_2191,In_673,In_660);
nand U2192 (N_2192,In_550,In_388);
and U2193 (N_2193,In_509,In_508);
xnor U2194 (N_2194,In_730,In_349);
nor U2195 (N_2195,In_23,In_351);
nor U2196 (N_2196,In_12,In_28);
nor U2197 (N_2197,In_34,In_69);
nor U2198 (N_2198,In_724,In_700);
nand U2199 (N_2199,In_718,In_520);
and U2200 (N_2200,In_251,In_164);
and U2201 (N_2201,In_55,In_520);
nand U2202 (N_2202,In_479,In_640);
xor U2203 (N_2203,In_396,In_348);
nor U2204 (N_2204,In_514,In_121);
xor U2205 (N_2205,In_537,In_177);
nor U2206 (N_2206,In_631,In_338);
or U2207 (N_2207,In_292,In_379);
xor U2208 (N_2208,In_556,In_648);
nor U2209 (N_2209,In_33,In_440);
nand U2210 (N_2210,In_1,In_113);
nand U2211 (N_2211,In_587,In_387);
xor U2212 (N_2212,In_186,In_459);
nand U2213 (N_2213,In_193,In_112);
and U2214 (N_2214,In_19,In_711);
nor U2215 (N_2215,In_310,In_264);
and U2216 (N_2216,In_439,In_304);
nor U2217 (N_2217,In_734,In_94);
xor U2218 (N_2218,In_91,In_422);
or U2219 (N_2219,In_271,In_482);
xor U2220 (N_2220,In_86,In_378);
xor U2221 (N_2221,In_495,In_719);
and U2222 (N_2222,In_402,In_315);
or U2223 (N_2223,In_502,In_254);
xnor U2224 (N_2224,In_385,In_304);
or U2225 (N_2225,In_579,In_127);
nand U2226 (N_2226,In_130,In_603);
nor U2227 (N_2227,In_352,In_585);
xor U2228 (N_2228,In_367,In_529);
and U2229 (N_2229,In_25,In_160);
and U2230 (N_2230,In_328,In_708);
nor U2231 (N_2231,In_171,In_565);
xor U2232 (N_2232,In_555,In_96);
or U2233 (N_2233,In_283,In_56);
nand U2234 (N_2234,In_256,In_203);
or U2235 (N_2235,In_79,In_499);
nor U2236 (N_2236,In_33,In_486);
xnor U2237 (N_2237,In_169,In_250);
and U2238 (N_2238,In_498,In_512);
nand U2239 (N_2239,In_138,In_499);
nand U2240 (N_2240,In_368,In_505);
xnor U2241 (N_2241,In_367,In_228);
nand U2242 (N_2242,In_262,In_663);
nor U2243 (N_2243,In_511,In_453);
or U2244 (N_2244,In_673,In_727);
and U2245 (N_2245,In_456,In_377);
nand U2246 (N_2246,In_221,In_68);
and U2247 (N_2247,In_521,In_186);
or U2248 (N_2248,In_104,In_620);
and U2249 (N_2249,In_33,In_470);
xnor U2250 (N_2250,In_563,In_423);
nand U2251 (N_2251,In_435,In_432);
or U2252 (N_2252,In_529,In_44);
or U2253 (N_2253,In_265,In_699);
and U2254 (N_2254,In_55,In_279);
and U2255 (N_2255,In_488,In_638);
and U2256 (N_2256,In_8,In_564);
xor U2257 (N_2257,In_93,In_726);
or U2258 (N_2258,In_184,In_537);
nor U2259 (N_2259,In_685,In_622);
or U2260 (N_2260,In_618,In_675);
and U2261 (N_2261,In_722,In_174);
or U2262 (N_2262,In_250,In_428);
and U2263 (N_2263,In_516,In_549);
xor U2264 (N_2264,In_95,In_98);
xor U2265 (N_2265,In_683,In_292);
nand U2266 (N_2266,In_147,In_706);
xnor U2267 (N_2267,In_549,In_112);
or U2268 (N_2268,In_530,In_564);
xnor U2269 (N_2269,In_525,In_727);
and U2270 (N_2270,In_187,In_478);
nand U2271 (N_2271,In_397,In_559);
xnor U2272 (N_2272,In_178,In_283);
and U2273 (N_2273,In_539,In_48);
or U2274 (N_2274,In_59,In_708);
or U2275 (N_2275,In_368,In_402);
or U2276 (N_2276,In_95,In_152);
nor U2277 (N_2277,In_452,In_243);
and U2278 (N_2278,In_548,In_487);
and U2279 (N_2279,In_215,In_429);
and U2280 (N_2280,In_193,In_733);
nand U2281 (N_2281,In_221,In_163);
or U2282 (N_2282,In_562,In_386);
or U2283 (N_2283,In_68,In_138);
nor U2284 (N_2284,In_628,In_165);
xor U2285 (N_2285,In_728,In_619);
or U2286 (N_2286,In_78,In_448);
nor U2287 (N_2287,In_408,In_444);
xnor U2288 (N_2288,In_333,In_294);
nand U2289 (N_2289,In_694,In_207);
and U2290 (N_2290,In_253,In_686);
nand U2291 (N_2291,In_656,In_676);
xor U2292 (N_2292,In_504,In_228);
xnor U2293 (N_2293,In_418,In_8);
and U2294 (N_2294,In_513,In_673);
nor U2295 (N_2295,In_70,In_381);
and U2296 (N_2296,In_438,In_136);
and U2297 (N_2297,In_24,In_308);
nor U2298 (N_2298,In_356,In_368);
or U2299 (N_2299,In_107,In_567);
or U2300 (N_2300,In_319,In_329);
nor U2301 (N_2301,In_476,In_550);
xor U2302 (N_2302,In_668,In_583);
nor U2303 (N_2303,In_465,In_748);
nor U2304 (N_2304,In_275,In_258);
xor U2305 (N_2305,In_358,In_727);
xnor U2306 (N_2306,In_245,In_89);
and U2307 (N_2307,In_587,In_249);
and U2308 (N_2308,In_697,In_219);
xor U2309 (N_2309,In_659,In_371);
and U2310 (N_2310,In_251,In_612);
nor U2311 (N_2311,In_65,In_53);
nand U2312 (N_2312,In_315,In_586);
xnor U2313 (N_2313,In_49,In_108);
nand U2314 (N_2314,In_185,In_193);
xor U2315 (N_2315,In_660,In_697);
xnor U2316 (N_2316,In_204,In_301);
nor U2317 (N_2317,In_588,In_564);
xor U2318 (N_2318,In_382,In_737);
and U2319 (N_2319,In_56,In_493);
and U2320 (N_2320,In_612,In_59);
nor U2321 (N_2321,In_571,In_252);
or U2322 (N_2322,In_70,In_340);
and U2323 (N_2323,In_741,In_656);
xor U2324 (N_2324,In_237,In_500);
and U2325 (N_2325,In_32,In_727);
nor U2326 (N_2326,In_431,In_180);
nand U2327 (N_2327,In_587,In_490);
nor U2328 (N_2328,In_304,In_414);
nand U2329 (N_2329,In_304,In_530);
or U2330 (N_2330,In_316,In_490);
nor U2331 (N_2331,In_650,In_205);
xor U2332 (N_2332,In_129,In_9);
xnor U2333 (N_2333,In_163,In_207);
and U2334 (N_2334,In_171,In_185);
and U2335 (N_2335,In_230,In_102);
nor U2336 (N_2336,In_678,In_694);
xnor U2337 (N_2337,In_424,In_265);
nand U2338 (N_2338,In_234,In_631);
nand U2339 (N_2339,In_658,In_355);
nand U2340 (N_2340,In_729,In_687);
or U2341 (N_2341,In_41,In_459);
xor U2342 (N_2342,In_660,In_306);
nand U2343 (N_2343,In_676,In_546);
xor U2344 (N_2344,In_326,In_239);
xnor U2345 (N_2345,In_287,In_1);
nor U2346 (N_2346,In_489,In_257);
nor U2347 (N_2347,In_223,In_553);
nor U2348 (N_2348,In_549,In_18);
or U2349 (N_2349,In_446,In_22);
nor U2350 (N_2350,In_553,In_358);
xor U2351 (N_2351,In_699,In_24);
or U2352 (N_2352,In_193,In_141);
and U2353 (N_2353,In_463,In_439);
or U2354 (N_2354,In_100,In_307);
nand U2355 (N_2355,In_474,In_146);
nor U2356 (N_2356,In_380,In_668);
nand U2357 (N_2357,In_64,In_35);
nand U2358 (N_2358,In_192,In_325);
xor U2359 (N_2359,In_192,In_641);
or U2360 (N_2360,In_115,In_256);
or U2361 (N_2361,In_124,In_725);
or U2362 (N_2362,In_347,In_678);
and U2363 (N_2363,In_115,In_485);
and U2364 (N_2364,In_530,In_648);
xnor U2365 (N_2365,In_48,In_733);
xnor U2366 (N_2366,In_518,In_696);
nand U2367 (N_2367,In_643,In_673);
and U2368 (N_2368,In_617,In_118);
or U2369 (N_2369,In_18,In_639);
xor U2370 (N_2370,In_559,In_420);
and U2371 (N_2371,In_338,In_122);
or U2372 (N_2372,In_594,In_269);
or U2373 (N_2373,In_129,In_19);
xnor U2374 (N_2374,In_625,In_27);
nor U2375 (N_2375,In_141,In_142);
nor U2376 (N_2376,In_498,In_320);
nand U2377 (N_2377,In_132,In_401);
or U2378 (N_2378,In_260,In_116);
xnor U2379 (N_2379,In_320,In_415);
or U2380 (N_2380,In_462,In_52);
xor U2381 (N_2381,In_699,In_437);
xnor U2382 (N_2382,In_276,In_225);
or U2383 (N_2383,In_246,In_2);
or U2384 (N_2384,In_609,In_497);
nand U2385 (N_2385,In_410,In_300);
and U2386 (N_2386,In_644,In_292);
xor U2387 (N_2387,In_679,In_268);
or U2388 (N_2388,In_521,In_563);
nand U2389 (N_2389,In_611,In_619);
nand U2390 (N_2390,In_350,In_609);
xnor U2391 (N_2391,In_698,In_241);
and U2392 (N_2392,In_292,In_192);
xnor U2393 (N_2393,In_544,In_293);
and U2394 (N_2394,In_294,In_411);
xor U2395 (N_2395,In_332,In_553);
xor U2396 (N_2396,In_681,In_351);
xor U2397 (N_2397,In_431,In_280);
nand U2398 (N_2398,In_537,In_70);
nor U2399 (N_2399,In_279,In_95);
nand U2400 (N_2400,In_648,In_727);
nor U2401 (N_2401,In_180,In_147);
nand U2402 (N_2402,In_474,In_111);
or U2403 (N_2403,In_664,In_667);
and U2404 (N_2404,In_598,In_626);
nand U2405 (N_2405,In_401,In_3);
nand U2406 (N_2406,In_378,In_129);
or U2407 (N_2407,In_116,In_224);
xnor U2408 (N_2408,In_5,In_666);
xnor U2409 (N_2409,In_511,In_710);
nand U2410 (N_2410,In_433,In_183);
nand U2411 (N_2411,In_660,In_313);
and U2412 (N_2412,In_323,In_261);
or U2413 (N_2413,In_745,In_237);
nor U2414 (N_2414,In_609,In_624);
nand U2415 (N_2415,In_54,In_310);
nand U2416 (N_2416,In_242,In_316);
and U2417 (N_2417,In_270,In_212);
nand U2418 (N_2418,In_357,In_276);
nand U2419 (N_2419,In_643,In_578);
and U2420 (N_2420,In_429,In_567);
xor U2421 (N_2421,In_678,In_379);
and U2422 (N_2422,In_420,In_594);
nor U2423 (N_2423,In_372,In_350);
or U2424 (N_2424,In_746,In_684);
xnor U2425 (N_2425,In_606,In_568);
nor U2426 (N_2426,In_334,In_157);
nor U2427 (N_2427,In_696,In_99);
or U2428 (N_2428,In_333,In_686);
xor U2429 (N_2429,In_398,In_361);
and U2430 (N_2430,In_715,In_377);
or U2431 (N_2431,In_439,In_298);
xor U2432 (N_2432,In_693,In_305);
or U2433 (N_2433,In_545,In_729);
xor U2434 (N_2434,In_290,In_510);
nand U2435 (N_2435,In_296,In_398);
xnor U2436 (N_2436,In_63,In_305);
and U2437 (N_2437,In_349,In_33);
or U2438 (N_2438,In_465,In_578);
and U2439 (N_2439,In_157,In_711);
and U2440 (N_2440,In_375,In_109);
nor U2441 (N_2441,In_548,In_159);
or U2442 (N_2442,In_647,In_481);
nor U2443 (N_2443,In_492,In_622);
and U2444 (N_2444,In_397,In_744);
or U2445 (N_2445,In_149,In_93);
xnor U2446 (N_2446,In_105,In_104);
or U2447 (N_2447,In_649,In_726);
nor U2448 (N_2448,In_342,In_488);
nor U2449 (N_2449,In_187,In_670);
and U2450 (N_2450,In_519,In_226);
and U2451 (N_2451,In_624,In_745);
xor U2452 (N_2452,In_441,In_421);
xnor U2453 (N_2453,In_115,In_471);
nand U2454 (N_2454,In_162,In_531);
xor U2455 (N_2455,In_447,In_576);
nor U2456 (N_2456,In_103,In_311);
nor U2457 (N_2457,In_191,In_445);
xor U2458 (N_2458,In_469,In_509);
nor U2459 (N_2459,In_614,In_385);
nor U2460 (N_2460,In_328,In_571);
and U2461 (N_2461,In_359,In_161);
nand U2462 (N_2462,In_691,In_544);
nor U2463 (N_2463,In_643,In_138);
or U2464 (N_2464,In_281,In_555);
nor U2465 (N_2465,In_573,In_374);
and U2466 (N_2466,In_490,In_11);
nor U2467 (N_2467,In_503,In_318);
nor U2468 (N_2468,In_206,In_499);
or U2469 (N_2469,In_278,In_479);
nor U2470 (N_2470,In_742,In_723);
xnor U2471 (N_2471,In_286,In_477);
nand U2472 (N_2472,In_371,In_247);
and U2473 (N_2473,In_743,In_307);
xnor U2474 (N_2474,In_409,In_297);
nand U2475 (N_2475,In_420,In_164);
nor U2476 (N_2476,In_66,In_351);
or U2477 (N_2477,In_242,In_561);
xor U2478 (N_2478,In_468,In_669);
nand U2479 (N_2479,In_337,In_65);
and U2480 (N_2480,In_130,In_345);
nand U2481 (N_2481,In_129,In_204);
nor U2482 (N_2482,In_367,In_117);
nand U2483 (N_2483,In_713,In_142);
nor U2484 (N_2484,In_414,In_641);
or U2485 (N_2485,In_538,In_724);
and U2486 (N_2486,In_259,In_726);
nand U2487 (N_2487,In_606,In_70);
nand U2488 (N_2488,In_170,In_639);
or U2489 (N_2489,In_528,In_704);
nor U2490 (N_2490,In_607,In_317);
or U2491 (N_2491,In_648,In_89);
xor U2492 (N_2492,In_263,In_403);
nand U2493 (N_2493,In_300,In_273);
nand U2494 (N_2494,In_720,In_494);
and U2495 (N_2495,In_626,In_625);
xor U2496 (N_2496,In_163,In_743);
xnor U2497 (N_2497,In_298,In_599);
and U2498 (N_2498,In_450,In_249);
or U2499 (N_2499,In_14,In_506);
or U2500 (N_2500,N_205,N_463);
or U2501 (N_2501,N_2425,N_1015);
or U2502 (N_2502,N_506,N_1975);
nor U2503 (N_2503,N_951,N_2449);
nand U2504 (N_2504,N_257,N_1246);
nand U2505 (N_2505,N_1502,N_2032);
xnor U2506 (N_2506,N_1083,N_1326);
and U2507 (N_2507,N_805,N_2233);
or U2508 (N_2508,N_2268,N_2237);
xor U2509 (N_2509,N_2080,N_813);
or U2510 (N_2510,N_1214,N_1271);
xor U2511 (N_2511,N_1794,N_661);
or U2512 (N_2512,N_258,N_1430);
xnor U2513 (N_2513,N_266,N_1432);
and U2514 (N_2514,N_1236,N_2314);
or U2515 (N_2515,N_1132,N_260);
nor U2516 (N_2516,N_161,N_64);
nor U2517 (N_2517,N_1796,N_1808);
or U2518 (N_2518,N_2374,N_1810);
xnor U2519 (N_2519,N_134,N_628);
xnor U2520 (N_2520,N_2120,N_838);
or U2521 (N_2521,N_1103,N_809);
and U2522 (N_2522,N_837,N_1688);
xor U2523 (N_2523,N_897,N_2059);
nor U2524 (N_2524,N_436,N_2036);
nor U2525 (N_2525,N_1397,N_2236);
and U2526 (N_2526,N_711,N_712);
xnor U2527 (N_2527,N_1092,N_1524);
xor U2528 (N_2528,N_2345,N_1857);
and U2529 (N_2529,N_1408,N_355);
and U2530 (N_2530,N_1405,N_138);
and U2531 (N_2531,N_1251,N_1517);
or U2532 (N_2532,N_1584,N_2416);
and U2533 (N_2533,N_753,N_2037);
xnor U2534 (N_2534,N_1485,N_887);
xnor U2535 (N_2535,N_1240,N_1967);
and U2536 (N_2536,N_1247,N_88);
and U2537 (N_2537,N_1242,N_2018);
nor U2538 (N_2538,N_1275,N_214);
nand U2539 (N_2539,N_328,N_1686);
or U2540 (N_2540,N_386,N_1495);
nor U2541 (N_2541,N_2039,N_2265);
nor U2542 (N_2542,N_2246,N_2296);
nor U2543 (N_2543,N_426,N_2348);
or U2544 (N_2544,N_1995,N_1518);
xor U2545 (N_2545,N_1964,N_1202);
nor U2546 (N_2546,N_700,N_473);
nand U2547 (N_2547,N_2317,N_1358);
xnor U2548 (N_2548,N_1321,N_2002);
nor U2549 (N_2549,N_1258,N_2440);
xnor U2550 (N_2550,N_1336,N_1488);
and U2551 (N_2551,N_1943,N_2000);
or U2552 (N_2552,N_1555,N_2377);
nor U2553 (N_2553,N_513,N_804);
nor U2554 (N_2554,N_2009,N_1694);
xnor U2555 (N_2555,N_1442,N_1290);
xor U2556 (N_2556,N_2321,N_1261);
nand U2557 (N_2557,N_2382,N_1632);
nand U2558 (N_2558,N_167,N_1297);
nor U2559 (N_2559,N_1532,N_768);
xor U2560 (N_2560,N_878,N_752);
and U2561 (N_2561,N_1210,N_1974);
nand U2562 (N_2562,N_259,N_141);
and U2563 (N_2563,N_2480,N_115);
nor U2564 (N_2564,N_2151,N_940);
nand U2565 (N_2565,N_502,N_806);
or U2566 (N_2566,N_2094,N_2179);
nand U2567 (N_2567,N_1328,N_1918);
xor U2568 (N_2568,N_1234,N_2160);
or U2569 (N_2569,N_1171,N_545);
xnor U2570 (N_2570,N_1831,N_943);
or U2571 (N_2571,N_2101,N_316);
nor U2572 (N_2572,N_2444,N_1424);
or U2573 (N_2573,N_1604,N_2158);
and U2574 (N_2574,N_1152,N_31);
xor U2575 (N_2575,N_2327,N_1071);
nand U2576 (N_2576,N_566,N_2066);
and U2577 (N_2577,N_779,N_1159);
and U2578 (N_2578,N_1802,N_1534);
nor U2579 (N_2579,N_717,N_187);
nand U2580 (N_2580,N_1611,N_1480);
nand U2581 (N_2581,N_223,N_1203);
xnor U2582 (N_2582,N_1392,N_1365);
or U2583 (N_2583,N_583,N_1007);
and U2584 (N_2584,N_915,N_2182);
and U2585 (N_2585,N_2109,N_1226);
or U2586 (N_2586,N_1853,N_2283);
and U2587 (N_2587,N_1340,N_1763);
xor U2588 (N_2588,N_740,N_1823);
nand U2589 (N_2589,N_830,N_609);
nand U2590 (N_2590,N_2213,N_1175);
and U2591 (N_2591,N_902,N_1441);
nor U2592 (N_2592,N_1695,N_345);
or U2593 (N_2593,N_1923,N_1603);
and U2594 (N_2594,N_2287,N_1661);
nor U2595 (N_2595,N_1474,N_1313);
xor U2596 (N_2596,N_1533,N_1186);
xnor U2597 (N_2597,N_771,N_2183);
xnor U2598 (N_2598,N_234,N_862);
nand U2599 (N_2599,N_974,N_1988);
nand U2600 (N_2600,N_523,N_298);
nand U2601 (N_2601,N_587,N_2168);
nand U2602 (N_2602,N_2142,N_2291);
nor U2603 (N_2603,N_1099,N_1043);
xnor U2604 (N_2604,N_856,N_667);
xor U2605 (N_2605,N_2255,N_2324);
nor U2606 (N_2606,N_430,N_332);
and U2607 (N_2607,N_783,N_567);
or U2608 (N_2608,N_1178,N_1068);
nand U2609 (N_2609,N_612,N_1700);
xor U2610 (N_2610,N_2430,N_901);
or U2611 (N_2611,N_1253,N_1384);
and U2612 (N_2612,N_1765,N_2251);
xor U2613 (N_2613,N_906,N_263);
nor U2614 (N_2614,N_122,N_826);
xor U2615 (N_2615,N_908,N_1299);
and U2616 (N_2616,N_329,N_701);
xnor U2617 (N_2617,N_1526,N_1703);
nand U2618 (N_2618,N_1754,N_1149);
xor U2619 (N_2619,N_624,N_1566);
nor U2620 (N_2620,N_1863,N_1956);
or U2621 (N_2621,N_2074,N_1548);
and U2622 (N_2622,N_836,N_2034);
and U2623 (N_2623,N_1933,N_2081);
or U2624 (N_2624,N_1032,N_2078);
xor U2625 (N_2625,N_2300,N_285);
nand U2626 (N_2626,N_993,N_603);
and U2627 (N_2627,N_1057,N_320);
and U2628 (N_2628,N_829,N_1744);
xor U2629 (N_2629,N_2279,N_1322);
xnor U2630 (N_2630,N_621,N_1865);
or U2631 (N_2631,N_2343,N_989);
nand U2632 (N_2632,N_588,N_44);
nor U2633 (N_2633,N_103,N_1293);
or U2634 (N_2634,N_2202,N_2150);
or U2635 (N_2635,N_1239,N_1279);
nor U2636 (N_2636,N_772,N_1282);
nand U2637 (N_2637,N_1066,N_198);
xnor U2638 (N_2638,N_77,N_1618);
nor U2639 (N_2639,N_118,N_876);
xnor U2640 (N_2640,N_1002,N_322);
xor U2641 (N_2641,N_406,N_2022);
or U2642 (N_2642,N_1138,N_1133);
nand U2643 (N_2643,N_337,N_1675);
nand U2644 (N_2644,N_1158,N_135);
nand U2645 (N_2645,N_1077,N_496);
or U2646 (N_2646,N_1067,N_623);
and U2647 (N_2647,N_1445,N_1745);
nand U2648 (N_2648,N_1304,N_2230);
and U2649 (N_2649,N_1512,N_1394);
and U2650 (N_2650,N_1949,N_1909);
nand U2651 (N_2651,N_154,N_1821);
nor U2652 (N_2652,N_1306,N_1217);
xor U2653 (N_2653,N_1115,N_2460);
nand U2654 (N_2654,N_670,N_2218);
nor U2655 (N_2655,N_2466,N_1131);
and U2656 (N_2656,N_379,N_1705);
or U2657 (N_2657,N_2139,N_1998);
or U2658 (N_2658,N_1013,N_2055);
or U2659 (N_2659,N_1916,N_2006);
and U2660 (N_2660,N_1697,N_1283);
nor U2661 (N_2661,N_921,N_340);
nand U2662 (N_2662,N_2176,N_268);
nand U2663 (N_2663,N_1870,N_1843);
nor U2664 (N_2664,N_339,N_1845);
nor U2665 (N_2665,N_808,N_2163);
nor U2666 (N_2666,N_1539,N_1560);
nand U2667 (N_2667,N_1504,N_534);
nor U2668 (N_2668,N_1717,N_1999);
or U2669 (N_2669,N_1937,N_1893);
nand U2670 (N_2670,N_499,N_326);
and U2671 (N_2671,N_1649,N_2359);
or U2672 (N_2672,N_390,N_2389);
nor U2673 (N_2673,N_1569,N_476);
or U2674 (N_2674,N_650,N_801);
nor U2675 (N_2675,N_1453,N_1090);
xor U2676 (N_2676,N_272,N_1088);
and U2677 (N_2677,N_501,N_422);
or U2678 (N_2678,N_1227,N_1761);
nor U2679 (N_2679,N_1087,N_536);
nand U2680 (N_2680,N_869,N_371);
or U2681 (N_2681,N_1721,N_2464);
nor U2682 (N_2682,N_1713,N_792);
xor U2683 (N_2683,N_917,N_803);
nor U2684 (N_2684,N_1318,N_858);
or U2685 (N_2685,N_59,N_241);
or U2686 (N_2686,N_762,N_2095);
and U2687 (N_2687,N_248,N_996);
xnor U2688 (N_2688,N_1116,N_1683);
nand U2689 (N_2689,N_1873,N_2068);
nor U2690 (N_2690,N_444,N_2244);
and U2691 (N_2691,N_2154,N_627);
xnor U2692 (N_2692,N_967,N_2405);
or U2693 (N_2693,N_1574,N_2308);
nand U2694 (N_2694,N_739,N_796);
or U2695 (N_2695,N_295,N_675);
xnor U2696 (N_2696,N_1855,N_1038);
nor U2697 (N_2697,N_445,N_486);
or U2698 (N_2698,N_954,N_278);
or U2699 (N_2699,N_1028,N_579);
nand U2700 (N_2700,N_1140,N_2446);
xor U2701 (N_2701,N_1693,N_480);
or U2702 (N_2702,N_417,N_1259);
xor U2703 (N_2703,N_286,N_1463);
nor U2704 (N_2704,N_53,N_991);
xnor U2705 (N_2705,N_2498,N_133);
nor U2706 (N_2706,N_1357,N_817);
and U2707 (N_2707,N_393,N_911);
or U2708 (N_2708,N_2043,N_1961);
xnor U2709 (N_2709,N_547,N_302);
xor U2710 (N_2710,N_1847,N_2025);
or U2711 (N_2711,N_2350,N_2414);
or U2712 (N_2712,N_2275,N_116);
and U2713 (N_2713,N_960,N_2058);
nor U2714 (N_2714,N_565,N_128);
nor U2715 (N_2715,N_194,N_2253);
and U2716 (N_2716,N_1570,N_57);
xor U2717 (N_2717,N_2393,N_1323);
or U2718 (N_2718,N_1784,N_375);
or U2719 (N_2719,N_798,N_963);
nand U2720 (N_2720,N_1698,N_1558);
xor U2721 (N_2721,N_2017,N_2028);
xnor U2722 (N_2722,N_443,N_104);
nand U2723 (N_2723,N_1750,N_489);
or U2724 (N_2724,N_529,N_97);
nand U2725 (N_2725,N_446,N_2269);
and U2726 (N_2726,N_2372,N_1730);
and U2727 (N_2727,N_1617,N_331);
and U2728 (N_2728,N_2422,N_1912);
xnor U2729 (N_2729,N_1380,N_719);
nand U2730 (N_2730,N_1471,N_2014);
nor U2731 (N_2731,N_2482,N_671);
nand U2732 (N_2732,N_582,N_1628);
and U2733 (N_2733,N_117,N_1148);
or U2734 (N_2734,N_1968,N_625);
xnor U2735 (N_2735,N_26,N_1469);
nand U2736 (N_2736,N_904,N_2323);
nand U2737 (N_2737,N_747,N_1913);
or U2738 (N_2738,N_742,N_1440);
nand U2739 (N_2739,N_1451,N_1378);
or U2740 (N_2740,N_2299,N_1482);
or U2741 (N_2741,N_702,N_1598);
or U2742 (N_2742,N_127,N_1861);
nand U2743 (N_2743,N_950,N_1003);
xnor U2744 (N_2744,N_418,N_2271);
or U2745 (N_2745,N_82,N_2152);
and U2746 (N_2746,N_1696,N_2220);
or U2747 (N_2747,N_1352,N_644);
xor U2748 (N_2748,N_325,N_1298);
nor U2749 (N_2749,N_151,N_1609);
or U2750 (N_2750,N_2329,N_2319);
nand U2751 (N_2751,N_1256,N_1731);
and U2752 (N_2752,N_290,N_2231);
and U2753 (N_2753,N_1477,N_1742);
xor U2754 (N_2754,N_107,N_2326);
nand U2755 (N_2755,N_598,N_2143);
nor U2756 (N_2756,N_593,N_1161);
nand U2757 (N_2757,N_1751,N_584);
and U2758 (N_2758,N_188,N_2064);
nor U2759 (N_2759,N_1108,N_1221);
or U2760 (N_2760,N_1264,N_96);
nor U2761 (N_2761,N_1971,N_1804);
or U2762 (N_2762,N_1546,N_1056);
nand U2763 (N_2763,N_370,N_1228);
nor U2764 (N_2764,N_518,N_1385);
and U2765 (N_2765,N_984,N_2428);
and U2766 (N_2766,N_1535,N_990);
and U2767 (N_2767,N_1634,N_2146);
nor U2768 (N_2768,N_2257,N_1136);
or U2769 (N_2769,N_1982,N_1173);
nor U2770 (N_2770,N_2342,N_1355);
nand U2771 (N_2771,N_452,N_427);
nor U2772 (N_2772,N_2167,N_2290);
nor U2773 (N_2773,N_1719,N_300);
or U2774 (N_2774,N_432,N_1780);
or U2775 (N_2775,N_799,N_1208);
nand U2776 (N_2776,N_985,N_571);
nor U2777 (N_2777,N_586,N_1935);
nand U2778 (N_2778,N_13,N_1194);
nand U2779 (N_2779,N_1523,N_425);
nor U2780 (N_2780,N_2131,N_1229);
and U2781 (N_2781,N_932,N_338);
xnor U2782 (N_2782,N_438,N_217);
xor U2783 (N_2783,N_468,N_165);
and U2784 (N_2784,N_453,N_1541);
nor U2785 (N_2785,N_2091,N_2189);
xor U2786 (N_2786,N_1302,N_1439);
or U2787 (N_2787,N_1881,N_1147);
xor U2788 (N_2788,N_1244,N_2070);
and U2789 (N_2789,N_1008,N_200);
or U2790 (N_2790,N_2277,N_1320);
xnor U2791 (N_2791,N_1950,N_544);
nor U2792 (N_2792,N_674,N_916);
nor U2793 (N_2793,N_1364,N_1372);
nor U2794 (N_2794,N_196,N_0);
or U2795 (N_2795,N_868,N_872);
or U2796 (N_2796,N_1543,N_317);
or U2797 (N_2797,N_287,N_666);
and U2798 (N_2798,N_1417,N_305);
nor U2799 (N_2799,N_292,N_1074);
xnor U2800 (N_2800,N_464,N_765);
nand U2801 (N_2801,N_413,N_1325);
nor U2802 (N_2802,N_1537,N_824);
nor U2803 (N_2803,N_2129,N_2354);
nand U2804 (N_2804,N_1309,N_114);
nor U2805 (N_2805,N_2483,N_1830);
and U2806 (N_2806,N_1054,N_981);
nor U2807 (N_2807,N_1638,N_716);
nand U2808 (N_2808,N_227,N_404);
nand U2809 (N_2809,N_730,N_1684);
or U2810 (N_2810,N_1010,N_1866);
and U2811 (N_2811,N_2,N_270);
xor U2812 (N_2812,N_2463,N_1273);
nand U2813 (N_2813,N_39,N_1120);
xor U2814 (N_2814,N_2478,N_1576);
nor U2815 (N_2815,N_1567,N_2267);
nor U2816 (N_2816,N_1407,N_2234);
or U2817 (N_2817,N_1809,N_140);
nand U2818 (N_2818,N_508,N_655);
nor U2819 (N_2819,N_1666,N_934);
nand U2820 (N_2820,N_601,N_1930);
nand U2821 (N_2821,N_2219,N_1165);
xnor U2822 (N_2822,N_2339,N_2235);
and U2823 (N_2823,N_1653,N_247);
and U2824 (N_2824,N_2188,N_166);
xor U2825 (N_2825,N_2357,N_1792);
nor U2826 (N_2826,N_1948,N_2045);
or U2827 (N_2827,N_1016,N_1265);
nand U2828 (N_2828,N_1749,N_2026);
xnor U2829 (N_2829,N_1207,N_213);
or U2830 (N_2830,N_1959,N_168);
nand U2831 (N_2831,N_540,N_2431);
and U2832 (N_2832,N_462,N_857);
nand U2833 (N_2833,N_1800,N_683);
or U2834 (N_2834,N_189,N_3);
nor U2835 (N_2835,N_2228,N_1599);
nor U2836 (N_2836,N_705,N_2020);
nand U2837 (N_2837,N_1970,N_521);
nor U2838 (N_2838,N_1704,N_387);
xor U2839 (N_2839,N_2015,N_959);
nor U2840 (N_2840,N_423,N_1072);
xnor U2841 (N_2841,N_1076,N_848);
and U2842 (N_2842,N_1732,N_1414);
and U2843 (N_2843,N_220,N_561);
and U2844 (N_2844,N_1435,N_1891);
or U2845 (N_2845,N_591,N_169);
or U2846 (N_2846,N_931,N_111);
nor U2847 (N_2847,N_715,N_131);
or U2848 (N_2848,N_132,N_1627);
or U2849 (N_2849,N_2148,N_2097);
and U2850 (N_2850,N_2285,N_1009);
and U2851 (N_2851,N_2470,N_86);
nand U2852 (N_2852,N_1728,N_539);
xor U2853 (N_2853,N_1768,N_232);
or U2854 (N_2854,N_459,N_863);
nand U2855 (N_2855,N_71,N_2266);
or U2856 (N_2856,N_1044,N_573);
nand U2857 (N_2857,N_2104,N_126);
nor U2858 (N_2858,N_2400,N_431);
nand U2859 (N_2859,N_1213,N_987);
xor U2860 (N_2860,N_669,N_2388);
nor U2861 (N_2861,N_2102,N_219);
nand U2862 (N_2862,N_1678,N_146);
nand U2863 (N_2863,N_727,N_1349);
xnor U2864 (N_2864,N_821,N_2494);
or U2865 (N_2865,N_871,N_528);
and U2866 (N_2866,N_697,N_1978);
and U2867 (N_2867,N_2209,N_654);
nor U2868 (N_2868,N_574,N_2312);
and U2869 (N_2869,N_2136,N_1053);
or U2870 (N_2870,N_2325,N_91);
nand U2871 (N_2871,N_36,N_1733);
or U2872 (N_2872,N_1390,N_1984);
xor U2873 (N_2873,N_2053,N_410);
or U2874 (N_2874,N_9,N_2174);
xor U2875 (N_2875,N_1775,N_875);
or U2876 (N_2876,N_657,N_1692);
and U2877 (N_2877,N_517,N_708);
nor U2878 (N_2878,N_277,N_2210);
nor U2879 (N_2879,N_2226,N_2457);
or U2880 (N_2880,N_211,N_1616);
nor U2881 (N_2881,N_1086,N_581);
xnor U2882 (N_2882,N_1075,N_244);
or U2883 (N_2883,N_228,N_1021);
nand U2884 (N_2884,N_1464,N_296);
nor U2885 (N_2885,N_1035,N_592);
xnor U2886 (N_2886,N_399,N_267);
nor U2887 (N_2887,N_1001,N_2001);
nand U2888 (N_2888,N_1123,N_392);
xor U2889 (N_2889,N_877,N_1945);
nand U2890 (N_2890,N_29,N_2208);
nand U2891 (N_2891,N_844,N_294);
and U2892 (N_2892,N_2216,N_1623);
nor U2893 (N_2893,N_870,N_206);
nand U2894 (N_2894,N_1516,N_1494);
nor U2895 (N_2895,N_5,N_1644);
nor U2896 (N_2896,N_2083,N_2309);
or U2897 (N_2897,N_1219,N_1735);
or U2898 (N_2898,N_2011,N_1972);
or U2899 (N_2899,N_2054,N_957);
xor U2900 (N_2900,N_1037,N_1192);
or U2901 (N_2901,N_156,N_1177);
nand U2902 (N_2902,N_2248,N_845);
xnor U2903 (N_2903,N_1846,N_2086);
nor U2904 (N_2904,N_2007,N_45);
or U2905 (N_2905,N_1312,N_110);
nand U2906 (N_2906,N_568,N_1932);
and U2907 (N_2907,N_2302,N_2351);
xor U2908 (N_2908,N_1838,N_1509);
nand U2909 (N_2909,N_458,N_2286);
nor U2910 (N_2910,N_1726,N_1174);
or U2911 (N_2911,N_1478,N_1278);
nand U2912 (N_2912,N_420,N_315);
xor U2913 (N_2913,N_2481,N_600);
nand U2914 (N_2914,N_2445,N_1180);
nor U2915 (N_2915,N_812,N_354);
xor U2916 (N_2916,N_1844,N_2225);
and U2917 (N_2917,N_790,N_49);
or U2918 (N_2918,N_2295,N_2227);
xnor U2919 (N_2919,N_2200,N_109);
and U2920 (N_2920,N_1391,N_1927);
nand U2921 (N_2921,N_505,N_1791);
or U2922 (N_2922,N_614,N_11);
or U2923 (N_2923,N_2370,N_709);
xor U2924 (N_2924,N_1455,N_1936);
and U2925 (N_2925,N_1760,N_572);
nand U2926 (N_2926,N_1906,N_769);
xor U2927 (N_2927,N_1739,N_488);
or U2928 (N_2928,N_347,N_1877);
or U2929 (N_2929,N_925,N_274);
and U2930 (N_2930,N_186,N_1597);
and U2931 (N_2931,N_42,N_1350);
nand U2932 (N_2932,N_652,N_734);
xnor U2933 (N_2933,N_1505,N_1206);
nand U2934 (N_2934,N_1456,N_1540);
or U2935 (N_2935,N_1851,N_2077);
xnor U2936 (N_2936,N_2206,N_958);
and U2937 (N_2937,N_2371,N_550);
nor U2938 (N_2938,N_460,N_465);
xnor U2939 (N_2939,N_1588,N_2363);
xor U2940 (N_2940,N_1641,N_466);
or U2941 (N_2941,N_1875,N_2030);
or U2942 (N_2942,N_1647,N_2443);
xor U2943 (N_2943,N_949,N_634);
and U2944 (N_2944,N_1303,N_1420);
nand U2945 (N_2945,N_98,N_1864);
xor U2946 (N_2946,N_733,N_2468);
nor U2947 (N_2947,N_1155,N_690);
and U2948 (N_2948,N_2128,N_659);
nand U2949 (N_2949,N_2474,N_2171);
xor U2950 (N_2950,N_1341,N_474);
nor U2951 (N_2951,N_2069,N_2184);
nor U2952 (N_2952,N_1366,N_2010);
nand U2953 (N_2953,N_2019,N_997);
xnor U2954 (N_2954,N_866,N_181);
and U2955 (N_2955,N_419,N_1926);
and U2956 (N_2956,N_2418,N_2385);
or U2957 (N_2957,N_699,N_815);
xor U2958 (N_2958,N_1807,N_2156);
xnor U2959 (N_2959,N_1167,N_1834);
xor U2960 (N_2960,N_335,N_264);
or U2961 (N_2961,N_1687,N_72);
and U2962 (N_2962,N_374,N_756);
xnor U2963 (N_2963,N_865,N_1189);
and U2964 (N_2964,N_2082,N_1940);
or U2965 (N_2965,N_1911,N_253);
nand U2966 (N_2966,N_2356,N_2462);
nand U2967 (N_2967,N_507,N_1752);
nand U2968 (N_2968,N_2197,N_284);
or U2969 (N_2969,N_2132,N_84);
xor U2970 (N_2970,N_47,N_1595);
nor U2971 (N_2971,N_421,N_986);
nand U2972 (N_2972,N_819,N_391);
and U2973 (N_2973,N_2258,N_785);
nand U2974 (N_2974,N_1708,N_555);
nor U2975 (N_2975,N_2281,N_1779);
nand U2976 (N_2976,N_318,N_1626);
nand U2977 (N_2977,N_1753,N_1811);
xnor U2978 (N_2978,N_1610,N_106);
or U2979 (N_2979,N_495,N_814);
xnor U2980 (N_2980,N_2448,N_1650);
nor U2981 (N_2981,N_23,N_2432);
nor U2982 (N_2982,N_520,N_2297);
xor U2983 (N_2983,N_2346,N_1362);
or U2984 (N_2984,N_2461,N_2135);
and U2985 (N_2985,N_924,N_1827);
xor U2986 (N_2986,N_1413,N_1166);
or U2987 (N_2987,N_913,N_1605);
nand U2988 (N_2988,N_807,N_909);
xnor U2989 (N_2989,N_1337,N_2065);
or U2990 (N_2990,N_1113,N_1139);
xnor U2991 (N_2991,N_889,N_15);
or U2992 (N_2992,N_1724,N_784);
or U2993 (N_2993,N_1024,N_1699);
nor U2994 (N_2994,N_1818,N_1338);
or U2995 (N_2995,N_1596,N_144);
nand U2996 (N_2996,N_635,N_560);
and U2997 (N_2997,N_490,N_1826);
nor U2998 (N_2998,N_1023,N_2399);
or U2999 (N_2999,N_2276,N_618);
nor U3000 (N_3000,N_1983,N_32);
or U3001 (N_3001,N_388,N_2384);
nand U3002 (N_3002,N_2090,N_689);
nor U3003 (N_3003,N_642,N_491);
and U3004 (N_3004,N_864,N_22);
nor U3005 (N_3005,N_789,N_524);
or U3006 (N_3006,N_1682,N_885);
and U3007 (N_3007,N_447,N_786);
nand U3008 (N_3008,N_309,N_2075);
and U3009 (N_3009,N_1117,N_541);
xor U3010 (N_3010,N_1901,N_1373);
nand U3011 (N_3011,N_2201,N_710);
xnor U3012 (N_3012,N_1151,N_841);
or U3013 (N_3013,N_240,N_1689);
xor U3014 (N_3014,N_823,N_1050);
nor U3015 (N_3015,N_1335,N_946);
nand U3016 (N_3016,N_532,N_262);
xor U3017 (N_3017,N_319,N_556);
nor U3018 (N_3018,N_1510,N_2263);
or U3019 (N_3019,N_1575,N_1677);
and U3020 (N_3020,N_1363,N_2403);
nor U3021 (N_3021,N_794,N_980);
nand U3022 (N_3022,N_1,N_2144);
or U3023 (N_3023,N_1272,N_2240);
or U3024 (N_3024,N_1890,N_846);
nand U3025 (N_3025,N_160,N_1100);
and U3026 (N_3026,N_2159,N_936);
or U3027 (N_3027,N_191,N_1182);
nor U3028 (N_3028,N_2330,N_361);
or U3029 (N_3029,N_2434,N_7);
and U3030 (N_3030,N_2447,N_1486);
xnor U3031 (N_3031,N_414,N_1419);
and U3032 (N_3032,N_1059,N_698);
xor U3033 (N_3033,N_707,N_2191);
xor U3034 (N_3034,N_362,N_879);
xnor U3035 (N_3035,N_1819,N_1393);
or U3036 (N_3036,N_1594,N_349);
nor U3037 (N_3037,N_2114,N_1070);
or U3038 (N_3038,N_1564,N_1590);
and U3039 (N_3039,N_433,N_2076);
nand U3040 (N_3040,N_793,N_619);
nor U3041 (N_3041,N_1063,N_1416);
nor U3042 (N_3042,N_1468,N_2041);
and U3043 (N_3043,N_1448,N_363);
xor U3044 (N_3044,N_1888,N_17);
nand U3045 (N_3045,N_939,N_158);
nor U3046 (N_3046,N_2004,N_1897);
and U3047 (N_3047,N_1327,N_691);
nor U3048 (N_3048,N_1230,N_333);
nor U3049 (N_3049,N_1048,N_1577);
xor U3050 (N_3050,N_2273,N_441);
nor U3051 (N_3051,N_1406,N_757);
xor U3052 (N_3052,N_791,N_364);
nand U3053 (N_3053,N_2366,N_239);
xnor U3054 (N_3054,N_995,N_34);
xnor U3055 (N_3055,N_1061,N_961);
nand U3056 (N_3056,N_1981,N_1859);
and U3057 (N_3057,N_471,N_979);
nand U3058 (N_3058,N_1118,N_604);
and U3059 (N_3059,N_663,N_2365);
nor U3060 (N_3060,N_2316,N_2223);
nand U3061 (N_3061,N_1033,N_1172);
xor U3062 (N_3062,N_2085,N_2173);
and U3063 (N_3063,N_1058,N_2270);
and U3064 (N_3064,N_152,N_1012);
or U3065 (N_3065,N_1497,N_365);
or U3066 (N_3066,N_323,N_1799);
nand U3067 (N_3067,N_101,N_2107);
xor U3068 (N_3068,N_2288,N_2016);
and U3069 (N_3069,N_2278,N_2435);
and U3070 (N_3070,N_2452,N_776);
or U3071 (N_3071,N_313,N_637);
or U3072 (N_3072,N_162,N_975);
nor U3073 (N_3073,N_487,N_2125);
and U3074 (N_3074,N_2047,N_1347);
and U3075 (N_3075,N_74,N_437);
nand U3076 (N_3076,N_229,N_1842);
nor U3077 (N_3077,N_2353,N_610);
nand U3078 (N_3078,N_1311,N_1245);
nand U3079 (N_3079,N_1646,N_512);
xor U3080 (N_3080,N_2048,N_2386);
or U3081 (N_3081,N_1925,N_732);
nor U3082 (N_3082,N_2005,N_1243);
and U3083 (N_3083,N_2496,N_155);
xnor U3084 (N_3084,N_79,N_777);
or U3085 (N_3085,N_770,N_542);
nand U3086 (N_3086,N_575,N_937);
xor U3087 (N_3087,N_1601,N_2040);
nand U3088 (N_3088,N_816,N_1344);
xor U3089 (N_3089,N_1840,N_1465);
nand U3090 (N_3090,N_2238,N_1931);
nand U3091 (N_3091,N_773,N_1762);
and U3092 (N_3092,N_1665,N_631);
and U3093 (N_3093,N_926,N_321);
nand U3094 (N_3094,N_1288,N_381);
nor U3095 (N_3095,N_207,N_1736);
nor U3096 (N_3096,N_65,N_1195);
nor U3097 (N_3097,N_1091,N_1691);
nor U3098 (N_3098,N_530,N_327);
nand U3099 (N_3099,N_1645,N_2499);
and U3100 (N_3100,N_1289,N_2488);
nand U3101 (N_3101,N_647,N_2190);
or U3102 (N_3102,N_1484,N_454);
nand U3103 (N_3103,N_119,N_1374);
xnor U3104 (N_3104,N_2476,N_1892);
xor U3105 (N_3105,N_440,N_1503);
nor U3106 (N_3106,N_2172,N_210);
xor U3107 (N_3107,N_143,N_748);
or U3108 (N_3108,N_197,N_1281);
nor U3109 (N_3109,N_2127,N_2390);
nor U3110 (N_3110,N_1353,N_787);
nor U3111 (N_3111,N_1314,N_781);
or U3112 (N_3112,N_2100,N_1046);
xor U3113 (N_3113,N_2196,N_484);
nor U3114 (N_3114,N_149,N_763);
or U3115 (N_3115,N_1499,N_833);
or U3116 (N_3116,N_2408,N_1268);
and U3117 (N_3117,N_1443,N_1462);
xnor U3118 (N_3118,N_1181,N_673);
and U3119 (N_3119,N_470,N_1829);
nor U3120 (N_3120,N_2178,N_835);
nor U3121 (N_3121,N_73,N_843);
xnor U3122 (N_3122,N_2426,N_171);
and U3123 (N_3123,N_595,N_68);
nor U3124 (N_3124,N_2315,N_1630);
nand U3125 (N_3125,N_706,N_2479);
nor U3126 (N_3126,N_1361,N_1446);
nand U3127 (N_3127,N_976,N_85);
nor U3128 (N_3128,N_2331,N_2232);
and U3129 (N_3129,N_2318,N_1073);
or U3130 (N_3130,N_1233,N_378);
nor U3131 (N_3131,N_2046,N_1052);
nor U3132 (N_3132,N_1629,N_1637);
nor U3133 (N_3133,N_972,N_2310);
nor U3134 (N_3134,N_1212,N_1806);
xor U3135 (N_3135,N_577,N_8);
or U3136 (N_3136,N_212,N_246);
and U3137 (N_3137,N_2456,N_2412);
nand U3138 (N_3138,N_324,N_563);
and U3139 (N_3139,N_183,N_968);
nand U3140 (N_3140,N_994,N_766);
and U3141 (N_3141,N_1801,N_43);
and U3142 (N_3142,N_1770,N_827);
or U3143 (N_3143,N_788,N_2130);
xnor U3144 (N_3144,N_121,N_1269);
nand U3145 (N_3145,N_383,N_1942);
and U3146 (N_3146,N_139,N_1421);
nor U3147 (N_3147,N_176,N_2421);
and U3148 (N_3148,N_1785,N_2212);
or U3149 (N_3149,N_467,N_30);
xor U3150 (N_3150,N_1979,N_1204);
and U3151 (N_3151,N_1527,N_948);
and U3152 (N_3152,N_1871,N_2469);
xor U3153 (N_3153,N_645,N_173);
and U3154 (N_3154,N_888,N_1218);
and U3155 (N_3155,N_2376,N_1817);
or U3156 (N_3156,N_28,N_224);
nor U3157 (N_3157,N_1833,N_2272);
or U3158 (N_3158,N_456,N_1232);
xnor U3159 (N_3159,N_2379,N_1924);
xnor U3160 (N_3160,N_2161,N_596);
or U3161 (N_3161,N_21,N_774);
nor U3162 (N_3162,N_608,N_651);
and U3163 (N_3163,N_1126,N_123);
xnor U3164 (N_3164,N_60,N_660);
and U3165 (N_3165,N_546,N_1257);
or U3166 (N_3166,N_589,N_1422);
nand U3167 (N_3167,N_1520,N_1119);
nand U3168 (N_3168,N_1386,N_2061);
nor U3169 (N_3169,N_1447,N_576);
or U3170 (N_3170,N_1919,N_243);
nor U3171 (N_3171,N_150,N_92);
xnor U3172 (N_3172,N_731,N_102);
nor U3173 (N_3173,N_1199,N_2192);
nand U3174 (N_3174,N_1428,N_1907);
nand U3175 (N_3175,N_2305,N_1345);
nand U3176 (N_3176,N_1587,N_356);
nand U3177 (N_3177,N_983,N_83);
or U3178 (N_3178,N_1461,N_1874);
nor U3179 (N_3179,N_1738,N_1938);
or U3180 (N_3180,N_1294,N_1492);
xnor U3181 (N_3181,N_2341,N_1069);
or U3182 (N_3182,N_1702,N_2073);
nand U3183 (N_3183,N_942,N_1019);
xor U3184 (N_3184,N_1388,N_2205);
or U3185 (N_3185,N_1778,N_686);
or U3186 (N_3186,N_1459,N_511);
and U3187 (N_3187,N_38,N_498);
xnor U3188 (N_3188,N_80,N_1989);
nand U3189 (N_3189,N_854,N_632);
nand U3190 (N_3190,N_164,N_2254);
nand U3191 (N_3191,N_1029,N_2355);
and U3192 (N_3192,N_1107,N_1343);
nor U3193 (N_3193,N_1782,N_352);
xnor U3194 (N_3194,N_382,N_1669);
or U3195 (N_3195,N_557,N_1714);
nor U3196 (N_3196,N_1183,N_1163);
or U3197 (N_3197,N_605,N_1460);
and U3198 (N_3198,N_722,N_1582);
and U3199 (N_3199,N_1157,N_1895);
and U3200 (N_3200,N_1403,N_395);
or U3201 (N_3201,N_2368,N_1903);
and U3202 (N_3202,N_69,N_416);
xor U3203 (N_3203,N_75,N_1593);
xor U3204 (N_3204,N_1156,N_1454);
or U3205 (N_3205,N_1319,N_1790);
xor U3206 (N_3206,N_1720,N_682);
and U3207 (N_3207,N_231,N_1191);
and U3208 (N_3208,N_2207,N_2454);
nand U3209 (N_3209,N_1795,N_99);
nor U3210 (N_3210,N_629,N_1489);
and U3211 (N_3211,N_235,N_1685);
nand U3212 (N_3212,N_558,N_2092);
nor U3213 (N_3213,N_527,N_2242);
and U3214 (N_3214,N_1614,N_475);
nor U3215 (N_3215,N_282,N_884);
or U3216 (N_3216,N_1193,N_1774);
xor U3217 (N_3217,N_831,N_1164);
nand U3218 (N_3218,N_1565,N_504);
nand U3219 (N_3219,N_2088,N_163);
nand U3220 (N_3220,N_1064,N_2035);
nand U3221 (N_3221,N_2038,N_2162);
xor U3222 (N_3222,N_680,N_694);
or U3223 (N_3223,N_1315,N_2352);
nor U3224 (N_3224,N_1973,N_2079);
and U3225 (N_3225,N_1370,N_1121);
or U3226 (N_3226,N_1030,N_2252);
or U3227 (N_3227,N_1060,N_688);
and U3228 (N_3228,N_2335,N_1955);
nor U3229 (N_3229,N_1572,N_1332);
nor U3230 (N_3230,N_81,N_1094);
nor U3231 (N_3231,N_125,N_2198);
nand U3232 (N_3232,N_736,N_658);
xor U3233 (N_3233,N_1082,N_1723);
or U3234 (N_3234,N_455,N_802);
nor U3235 (N_3235,N_428,N_1025);
nor U3236 (N_3236,N_1889,N_2241);
nand U3237 (N_3237,N_1885,N_613);
nand U3238 (N_3238,N_892,N_1986);
nand U3239 (N_3239,N_1145,N_254);
nor U3240 (N_3240,N_2401,N_912);
nor U3241 (N_3241,N_1093,N_1493);
or U3242 (N_3242,N_1743,N_1777);
nor U3243 (N_3243,N_1410,N_2413);
xor U3244 (N_3244,N_195,N_2419);
nand U3245 (N_3245,N_1789,N_226);
nand U3246 (N_3246,N_1854,N_2221);
nor U3247 (N_3247,N_2124,N_2391);
nand U3248 (N_3248,N_1433,N_403);
or U3249 (N_3249,N_2067,N_497);
xnor U3250 (N_3250,N_343,N_1561);
nand U3251 (N_3251,N_537,N_602);
xor U3252 (N_3252,N_1285,N_18);
nor U3253 (N_3253,N_822,N_2071);
nand U3254 (N_3254,N_2155,N_251);
and U3255 (N_3255,N_1701,N_1787);
xnor U3256 (N_3256,N_1852,N_755);
xnor U3257 (N_3257,N_1559,N_180);
and U3258 (N_3258,N_2362,N_873);
xor U3259 (N_3259,N_2157,N_590);
or U3260 (N_3260,N_1198,N_1080);
and U3261 (N_3261,N_2298,N_1143);
and U3262 (N_3262,N_1620,N_1880);
xor U3263 (N_3263,N_914,N_1624);
and U3264 (N_3264,N_1987,N_636);
and U3265 (N_3265,N_750,N_1263);
and U3266 (N_3266,N_360,N_2367);
and U3267 (N_3267,N_1102,N_941);
or U3268 (N_3268,N_2439,N_2304);
and U3269 (N_3269,N_2387,N_1856);
or U3270 (N_3270,N_2438,N_2186);
nand U3271 (N_3271,N_1813,N_170);
or U3272 (N_3272,N_2098,N_735);
xor U3273 (N_3273,N_510,N_2119);
nor U3274 (N_3274,N_66,N_1142);
and U3275 (N_3275,N_1224,N_130);
nand U3276 (N_3276,N_903,N_1905);
xor U3277 (N_3277,N_724,N_721);
and U3278 (N_3278,N_737,N_1690);
nor U3279 (N_3279,N_1452,N_1412);
nand U3280 (N_3280,N_1946,N_2475);
xnor U3281 (N_3281,N_2057,N_311);
and U3282 (N_3282,N_63,N_2484);
nor U3283 (N_3283,N_2093,N_377);
xnor U3284 (N_3284,N_1579,N_12);
xor U3285 (N_3285,N_500,N_1150);
and U3286 (N_3286,N_1681,N_1169);
or U3287 (N_3287,N_1026,N_56);
nand U3288 (N_3288,N_1976,N_1953);
or U3289 (N_3289,N_1729,N_2117);
or U3290 (N_3290,N_2072,N_1887);
or U3291 (N_3291,N_1608,N_373);
nor U3292 (N_3292,N_955,N_641);
or U3293 (N_3293,N_185,N_1920);
nand U3294 (N_3294,N_1934,N_1651);
xnor U3295 (N_3295,N_1398,N_2433);
nand U3296 (N_3296,N_1635,N_1928);
and U3297 (N_3297,N_1798,N_2050);
nor U3298 (N_3298,N_1078,N_969);
or U3299 (N_3299,N_1766,N_1400);
nand U3300 (N_3300,N_782,N_2441);
nor U3301 (N_3301,N_424,N_384);
nor U3302 (N_3302,N_2215,N_1711);
or U3303 (N_3303,N_1545,N_336);
or U3304 (N_3304,N_2087,N_1444);
or U3305 (N_3305,N_1367,N_1980);
and U3306 (N_3306,N_1065,N_2165);
nor U3307 (N_3307,N_929,N_1184);
nor U3308 (N_3308,N_2292,N_2149);
and U3309 (N_3309,N_2264,N_1308);
and U3310 (N_3310,N_1185,N_2332);
and U3311 (N_3311,N_1958,N_2099);
nor U3312 (N_3312,N_1960,N_1307);
or U3313 (N_3313,N_606,N_1671);
nand U3314 (N_3314,N_2261,N_664);
and U3315 (N_3315,N_376,N_1216);
nand U3316 (N_3316,N_745,N_2259);
or U3317 (N_3317,N_2204,N_744);
or U3318 (N_3318,N_1127,N_2492);
xor U3319 (N_3319,N_1759,N_1904);
nor U3320 (N_3320,N_535,N_1529);
xnor U3321 (N_3321,N_299,N_894);
nor U3322 (N_3322,N_1868,N_2424);
nor U3323 (N_3323,N_2320,N_714);
nor U3324 (N_3324,N_2364,N_1330);
and U3325 (N_3325,N_1110,N_389);
nand U3326 (N_3326,N_1097,N_1125);
nor U3327 (N_3327,N_1188,N_687);
and U3328 (N_3328,N_1144,N_357);
xor U3329 (N_3329,N_1501,N_216);
xnor U3330 (N_3330,N_1354,N_1654);
nand U3331 (N_3331,N_2063,N_304);
xnor U3332 (N_3332,N_1962,N_1295);
xnor U3333 (N_3333,N_1710,N_1600);
xnor U3334 (N_3334,N_95,N_1020);
xnor U3335 (N_3335,N_482,N_1371);
or U3336 (N_3336,N_2280,N_678);
or U3337 (N_3337,N_570,N_1467);
nor U3338 (N_3338,N_2153,N_2423);
nand U3339 (N_3339,N_893,N_509);
nand U3340 (N_3340,N_385,N_1041);
or U3341 (N_3341,N_283,N_867);
xor U3342 (N_3342,N_1602,N_896);
nor U3343 (N_3343,N_108,N_334);
and U3344 (N_3344,N_580,N_1209);
xor U3345 (N_3345,N_2096,N_478);
and U3346 (N_3346,N_2203,N_1674);
nand U3347 (N_3347,N_633,N_368);
and U3348 (N_3348,N_1815,N_1615);
xor U3349 (N_3349,N_597,N_1036);
xnor U3350 (N_3350,N_1146,N_1472);
xor U3351 (N_3351,N_208,N_192);
nand U3352 (N_3352,N_1200,N_2211);
nor U3353 (N_3353,N_2450,N_1490);
nor U3354 (N_3354,N_184,N_1639);
xnor U3355 (N_3355,N_1583,N_1652);
nand U3356 (N_3356,N_1111,N_1475);
xnor U3357 (N_3357,N_148,N_2338);
or U3358 (N_3358,N_905,N_780);
or U3359 (N_3359,N_221,N_933);
nand U3360 (N_3360,N_1130,N_910);
nand U3361 (N_3361,N_61,N_684);
nand U3362 (N_3362,N_1382,N_1122);
nor U3363 (N_3363,N_2337,N_758);
nor U3364 (N_3364,N_1018,N_1470);
nand U3365 (N_3365,N_526,N_1860);
and U3366 (N_3366,N_1262,N_2031);
or U3367 (N_3367,N_551,N_1376);
nor U3368 (N_3368,N_306,N_2361);
and U3369 (N_3369,N_1356,N_1722);
or U3370 (N_3370,N_2486,N_1137);
and U3371 (N_3371,N_1160,N_449);
nor U3372 (N_3372,N_1222,N_1515);
nor U3373 (N_3373,N_898,N_2108);
nand U3374 (N_3374,N_2133,N_1828);
nand U3375 (N_3375,N_1797,N_358);
and U3376 (N_3376,N_725,N_639);
nand U3377 (N_3377,N_1519,N_767);
or U3378 (N_3378,N_2180,N_964);
xnor U3379 (N_3379,N_1746,N_1633);
nor U3380 (N_3380,N_1487,N_1377);
and U3381 (N_3381,N_1425,N_1922);
and U3382 (N_3382,N_380,N_988);
or U3383 (N_3383,N_723,N_51);
xnor U3384 (N_3384,N_1334,N_2177);
nand U3385 (N_3385,N_1747,N_2347);
and U3386 (N_3386,N_245,N_1929);
nor U3387 (N_3387,N_297,N_2369);
nor U3388 (N_3388,N_553,N_1917);
or U3389 (N_3389,N_1254,N_70);
or U3390 (N_3390,N_2459,N_1951);
xor U3391 (N_3391,N_519,N_1712);
nand U3392 (N_3392,N_1153,N_202);
nor U3393 (N_3393,N_1957,N_1941);
or U3394 (N_3394,N_851,N_493);
nand U3395 (N_3395,N_54,N_157);
xor U3396 (N_3396,N_1022,N_1047);
or U3397 (N_3397,N_1231,N_2473);
and U3398 (N_3398,N_648,N_2358);
and U3399 (N_3399,N_346,N_351);
xor U3400 (N_3400,N_1437,N_1301);
and U3401 (N_3401,N_1837,N_825);
or U3402 (N_3402,N_649,N_741);
and U3403 (N_3403,N_754,N_52);
xor U3404 (N_3404,N_656,N_2411);
xnor U3405 (N_3405,N_1011,N_397);
nor U3406 (N_3406,N_1538,N_2407);
and U3407 (N_3407,N_1284,N_2137);
nor U3408 (N_3408,N_1977,N_2111);
nand U3409 (N_3409,N_2383,N_288);
and U3410 (N_3410,N_1824,N_190);
nand U3411 (N_3411,N_2214,N_1277);
xnor U3412 (N_3412,N_1648,N_1112);
nor U3413 (N_3413,N_2453,N_1662);
and U3414 (N_3414,N_2282,N_457);
or U3415 (N_3415,N_672,N_2427);
nor U3416 (N_3416,N_2301,N_531);
or U3417 (N_3417,N_638,N_2012);
and U3418 (N_3418,N_847,N_415);
nand U3419 (N_3419,N_1346,N_795);
nand U3420 (N_3420,N_2322,N_469);
nor U3421 (N_3421,N_2060,N_1513);
xor U3422 (N_3422,N_2378,N_859);
and U3423 (N_3423,N_492,N_35);
xor U3424 (N_3424,N_2455,N_1005);
and U3425 (N_3425,N_1803,N_273);
nor U3426 (N_3426,N_956,N_1415);
xor U3427 (N_3427,N_842,N_124);
nor U3428 (N_3428,N_1716,N_2489);
nor U3429 (N_3429,N_16,N_1436);
xor U3430 (N_3430,N_1994,N_2467);
nor U3431 (N_3431,N_1359,N_749);
and U3432 (N_3432,N_922,N_907);
xnor U3433 (N_3433,N_2195,N_665);
or U3434 (N_3434,N_1396,N_1522);
or U3435 (N_3435,N_1966,N_2169);
xnor U3436 (N_3436,N_1939,N_900);
nor U3437 (N_3437,N_626,N_2293);
or U3438 (N_3438,N_172,N_1664);
xor U3439 (N_3439,N_1902,N_249);
and U3440 (N_3440,N_236,N_1771);
or U3441 (N_3441,N_2138,N_2493);
or U3442 (N_3442,N_62,N_928);
nand U3443 (N_3443,N_2487,N_1547);
or U3444 (N_3444,N_1899,N_2084);
nand U3445 (N_3445,N_882,N_2110);
xnor U3446 (N_3446,N_1141,N_1793);
nor U3447 (N_3447,N_451,N_2497);
nor U3448 (N_3448,N_2126,N_2033);
nand U3449 (N_3449,N_1580,N_1429);
nand U3450 (N_3450,N_1551,N_1249);
or U3451 (N_3451,N_1619,N_1014);
xor U3452 (N_3452,N_1368,N_308);
nor U3453 (N_3453,N_1098,N_58);
or U3454 (N_3454,N_728,N_890);
or U3455 (N_3455,N_562,N_1287);
nor U3456 (N_3456,N_1755,N_1549);
and U3457 (N_3457,N_1305,N_2429);
xnor U3458 (N_3458,N_1270,N_1168);
or U3459 (N_3459,N_1727,N_2344);
xnor U3460 (N_3460,N_1858,N_938);
nor U3461 (N_3461,N_2260,N_797);
or U3462 (N_3462,N_348,N_1589);
xor U3463 (N_3463,N_177,N_2420);
nor U3464 (N_3464,N_2336,N_1869);
nand U3465 (N_3465,N_1573,N_1772);
or U3466 (N_3466,N_1051,N_1814);
nand U3467 (N_3467,N_930,N_2164);
nor U3468 (N_3468,N_199,N_372);
xor U3469 (N_3469,N_1707,N_105);
nor U3470 (N_3470,N_971,N_696);
nand U3471 (N_3471,N_2217,N_1506);
nor U3472 (N_3472,N_461,N_516);
and U3473 (N_3473,N_2417,N_1104);
nand U3474 (N_3474,N_695,N_242);
or U3475 (N_3475,N_1411,N_142);
xor U3476 (N_3476,N_450,N_40);
nor U3477 (N_3477,N_2465,N_1331);
nand U3478 (N_3478,N_1769,N_2307);
and U3479 (N_3479,N_448,N_27);
xor U3480 (N_3480,N_800,N_1276);
nor U3481 (N_3481,N_1900,N_1552);
xor U3482 (N_3482,N_1211,N_2451);
nor U3483 (N_3483,N_1525,N_1220);
and U3484 (N_3484,N_1530,N_100);
nor U3485 (N_3485,N_2056,N_1741);
and U3486 (N_3486,N_120,N_1135);
nor U3487 (N_3487,N_434,N_1196);
nand U3488 (N_3488,N_1867,N_1379);
xor U3489 (N_3489,N_1607,N_1556);
nand U3490 (N_3490,N_1563,N_408);
nor U3491 (N_3491,N_2245,N_713);
xnor U3492 (N_3492,N_1329,N_1248);
and U3493 (N_3493,N_668,N_1310);
xnor U3494 (N_3494,N_874,N_2089);
nor U3495 (N_3495,N_1521,N_1848);
nand U3496 (N_3496,N_301,N_1387);
nor U3497 (N_3497,N_41,N_2027);
and U3498 (N_3498,N_1625,N_1773);
nor U3499 (N_3499,N_525,N_87);
nor U3500 (N_3500,N_1621,N_1636);
xnor U3501 (N_3501,N_2406,N_1450);
and U3502 (N_3502,N_1658,N_136);
and U3503 (N_3503,N_1915,N_400);
nor U3504 (N_3504,N_1176,N_1381);
or U3505 (N_3505,N_147,N_407);
or U3506 (N_3506,N_2397,N_1586);
or U3507 (N_3507,N_2243,N_2112);
or U3508 (N_3508,N_76,N_1748);
and U3509 (N_3509,N_2194,N_1954);
nor U3510 (N_3510,N_662,N_1673);
nor U3511 (N_3511,N_1267,N_2436);
xor U3512 (N_3512,N_2185,N_398);
and U3513 (N_3513,N_1017,N_2284);
nand U3514 (N_3514,N_1300,N_1894);
or U3515 (N_3515,N_1260,N_1483);
nand U3516 (N_3516,N_2289,N_834);
xor U3517 (N_3517,N_1786,N_359);
nor U3518 (N_3518,N_307,N_1812);
nand U3519 (N_3519,N_1544,N_850);
nand U3520 (N_3520,N_1585,N_1715);
xnor U3521 (N_3521,N_2049,N_676);
xnor U3522 (N_3522,N_2147,N_1511);
nand U3523 (N_3523,N_503,N_2392);
or U3524 (N_3524,N_1034,N_37);
nor U3525 (N_3525,N_2349,N_927);
nand U3526 (N_3526,N_2274,N_1339);
xnor U3527 (N_3527,N_1223,N_761);
xnor U3528 (N_3528,N_2381,N_978);
nor U3529 (N_3529,N_554,N_1878);
nor U3530 (N_3530,N_25,N_1241);
nand U3531 (N_3531,N_1369,N_1776);
xnor U3532 (N_3532,N_1402,N_1952);
or U3533 (N_3533,N_2193,N_2115);
nor U3534 (N_3534,N_1095,N_367);
or U3535 (N_3535,N_2181,N_1498);
or U3536 (N_3536,N_1031,N_1317);
and U3537 (N_3537,N_760,N_435);
or U3538 (N_3538,N_1758,N_685);
nand U3539 (N_3539,N_238,N_1606);
nor U3540 (N_3540,N_1383,N_693);
nor U3541 (N_3541,N_2360,N_2409);
and U3542 (N_3542,N_2123,N_1805);
xnor U3543 (N_3543,N_1360,N_1187);
xnor U3544 (N_3544,N_1291,N_230);
and U3545 (N_3545,N_153,N_2042);
nor U3546 (N_3546,N_1883,N_6);
and U3547 (N_3547,N_1418,N_947);
nor U3548 (N_3548,N_1081,N_2415);
or U3549 (N_3549,N_2262,N_1993);
nand U3550 (N_3550,N_2306,N_237);
or U3551 (N_3551,N_992,N_179);
xnor U3552 (N_3552,N_718,N_564);
nand U3553 (N_3553,N_569,N_2170);
nor U3554 (N_3554,N_679,N_1657);
or U3555 (N_3555,N_2380,N_552);
nand U3556 (N_3556,N_94,N_2485);
xnor U3557 (N_3557,N_962,N_1458);
nor U3558 (N_3558,N_477,N_1101);
nor U3559 (N_3559,N_1514,N_1062);
or U3560 (N_3560,N_1536,N_982);
nor U3561 (N_3561,N_514,N_953);
or U3562 (N_3562,N_920,N_1201);
nand U3563 (N_3563,N_860,N_2116);
or U3564 (N_3564,N_1841,N_1886);
and U3565 (N_3565,N_396,N_1114);
nor U3566 (N_3566,N_1676,N_1027);
and U3567 (N_3567,N_218,N_48);
xnor U3568 (N_3568,N_2051,N_1040);
and U3569 (N_3569,N_2249,N_952);
nor U3570 (N_3570,N_543,N_1423);
xnor U3571 (N_3571,N_442,N_33);
and U3572 (N_3572,N_1409,N_966);
and U3573 (N_3573,N_923,N_549);
and U3574 (N_3574,N_818,N_2008);
or U3575 (N_3575,N_67,N_1896);
and U3576 (N_3576,N_895,N_1996);
and U3577 (N_3577,N_1124,N_585);
nand U3578 (N_3578,N_2491,N_1820);
nor U3579 (N_3579,N_14,N_1947);
or U3580 (N_3580,N_840,N_269);
and U3581 (N_3581,N_2442,N_2121);
nand U3582 (N_3582,N_1255,N_10);
nor U3583 (N_3583,N_405,N_1000);
or U3584 (N_3584,N_1500,N_919);
nor U3585 (N_3585,N_233,N_89);
or U3586 (N_3586,N_1944,N_1109);
nor U3587 (N_3587,N_1908,N_1039);
or U3588 (N_3588,N_1457,N_1507);
nor U3589 (N_3589,N_1985,N_1292);
or U3590 (N_3590,N_1849,N_222);
nor U3591 (N_3591,N_90,N_1106);
nand U3592 (N_3592,N_193,N_1342);
nor U3593 (N_3593,N_1992,N_1084);
nor U3594 (N_3594,N_751,N_1479);
nor U3595 (N_3595,N_2303,N_1718);
and U3596 (N_3596,N_832,N_1554);
and U3597 (N_3597,N_620,N_883);
and U3598 (N_3598,N_1434,N_2106);
nor U3599 (N_3599,N_965,N_1481);
xnor U3600 (N_3600,N_1835,N_113);
nand U3601 (N_3601,N_255,N_738);
nor U3602 (N_3602,N_726,N_1613);
nand U3603 (N_3603,N_559,N_2145);
nand U3604 (N_3604,N_1581,N_1333);
or U3605 (N_3605,N_1914,N_2404);
and U3606 (N_3606,N_2118,N_1496);
nor U3607 (N_3607,N_1725,N_1348);
xor U3608 (N_3608,N_112,N_1542);
nor U3609 (N_3609,N_2472,N_2333);
nand U3610 (N_3610,N_1839,N_2105);
or U3611 (N_3611,N_2140,N_1179);
or U3612 (N_3612,N_225,N_1438);
xnor U3613 (N_3613,N_1473,N_280);
xor U3614 (N_3614,N_853,N_4);
xor U3615 (N_3615,N_402,N_999);
nand U3616 (N_3616,N_256,N_20);
xnor U3617 (N_3617,N_409,N_2313);
xor U3618 (N_3618,N_1045,N_1643);
or U3619 (N_3619,N_2328,N_1642);
nand U3620 (N_3620,N_1764,N_1286);
nand U3621 (N_3621,N_279,N_1997);
xor U3622 (N_3622,N_1190,N_973);
or U3623 (N_3623,N_1631,N_729);
xnor U3624 (N_3624,N_175,N_1266);
nand U3625 (N_3625,N_2395,N_314);
nand U3626 (N_3626,N_1324,N_1862);
xnor U3627 (N_3627,N_1571,N_1667);
xnor U3628 (N_3628,N_828,N_2062);
nor U3629 (N_3629,N_703,N_515);
and U3630 (N_3630,N_1612,N_353);
xnor U3631 (N_3631,N_1668,N_342);
xnor U3632 (N_3632,N_861,N_2113);
or U3633 (N_3633,N_1670,N_2239);
nand U3634 (N_3634,N_2490,N_2229);
nor U3635 (N_3635,N_439,N_1660);
and U3636 (N_3636,N_1659,N_1898);
nor U3637 (N_3637,N_50,N_1788);
nand U3638 (N_3638,N_1531,N_886);
and U3639 (N_3639,N_704,N_646);
or U3640 (N_3640,N_764,N_1963);
nand U3641 (N_3641,N_681,N_970);
xor U3642 (N_3642,N_1399,N_1427);
and U3643 (N_3643,N_1351,N_1882);
or U3644 (N_3644,N_607,N_1553);
xor U3645 (N_3645,N_1557,N_616);
nor U3646 (N_3646,N_1965,N_261);
xnor U3647 (N_3647,N_1876,N_174);
and U3648 (N_3648,N_481,N_2199);
and U3649 (N_3649,N_293,N_880);
or U3650 (N_3650,N_2013,N_2003);
or U3651 (N_3651,N_1757,N_1042);
and U3652 (N_3652,N_341,N_1562);
and U3653 (N_3653,N_1401,N_129);
and U3654 (N_3654,N_1990,N_1822);
xor U3655 (N_3655,N_1431,N_2477);
nor U3656 (N_3656,N_1663,N_2224);
xor U3657 (N_3657,N_533,N_2103);
nand U3658 (N_3658,N_1205,N_271);
xor U3659 (N_3659,N_1134,N_1491);
nor U3660 (N_3660,N_201,N_1089);
and U3661 (N_3661,N_344,N_1578);
nand U3662 (N_3662,N_615,N_1672);
xnor U3663 (N_3663,N_1128,N_810);
xnor U3664 (N_3664,N_1466,N_55);
or U3665 (N_3665,N_281,N_1709);
nand U3666 (N_3666,N_303,N_899);
xor U3667 (N_3667,N_159,N_78);
or U3668 (N_3668,N_1426,N_1225);
nor U3669 (N_3669,N_2402,N_182);
nor U3670 (N_3670,N_918,N_178);
or U3671 (N_3671,N_1640,N_1085);
or U3672 (N_3672,N_366,N_1274);
and U3673 (N_3673,N_2458,N_2471);
nand U3674 (N_3674,N_1706,N_548);
and U3675 (N_3675,N_411,N_1655);
or U3676 (N_3676,N_137,N_945);
nand U3677 (N_3677,N_2334,N_1591);
xnor U3678 (N_3678,N_2052,N_2141);
nand U3679 (N_3679,N_483,N_204);
nor U3680 (N_3680,N_594,N_820);
nand U3681 (N_3681,N_881,N_252);
nand U3682 (N_3682,N_412,N_250);
nor U3683 (N_3683,N_2398,N_935);
or U3684 (N_3684,N_2311,N_485);
and U3685 (N_3685,N_1816,N_2340);
and U3686 (N_3686,N_479,N_472);
xnor U3687 (N_3687,N_1170,N_93);
xnor U3688 (N_3688,N_720,N_775);
nand U3689 (N_3689,N_2410,N_1004);
xnor U3690 (N_3690,N_1737,N_1825);
nand U3691 (N_3691,N_1476,N_1850);
and U3692 (N_3692,N_599,N_839);
nor U3693 (N_3693,N_1781,N_1235);
or U3694 (N_3694,N_891,N_289);
nor U3695 (N_3695,N_2294,N_24);
and U3696 (N_3696,N_653,N_630);
and U3697 (N_3697,N_1879,N_145);
xor U3698 (N_3698,N_1836,N_1096);
xnor U3699 (N_3699,N_2166,N_617);
nand U3700 (N_3700,N_1783,N_369);
or U3701 (N_3701,N_640,N_1550);
and U3702 (N_3702,N_1154,N_2394);
nand U3703 (N_3703,N_1316,N_19);
and U3704 (N_3704,N_522,N_276);
nor U3705 (N_3705,N_1105,N_2024);
nand U3706 (N_3706,N_849,N_2373);
nor U3707 (N_3707,N_2044,N_611);
and U3708 (N_3708,N_2247,N_1680);
nand U3709 (N_3709,N_622,N_1756);
nand U3710 (N_3710,N_46,N_209);
nand U3711 (N_3711,N_401,N_1740);
or U3712 (N_3712,N_2187,N_746);
or U3713 (N_3713,N_1884,N_1237);
nand U3714 (N_3714,N_778,N_1049);
xor U3715 (N_3715,N_692,N_1375);
nand U3716 (N_3716,N_1250,N_855);
or U3717 (N_3717,N_677,N_743);
nand U3718 (N_3718,N_1238,N_291);
nand U3719 (N_3719,N_1734,N_1055);
xnor U3720 (N_3720,N_394,N_1079);
nor U3721 (N_3721,N_1129,N_643);
and U3722 (N_3722,N_1528,N_811);
nand U3723 (N_3723,N_2122,N_203);
nand U3724 (N_3724,N_1872,N_1991);
nand U3725 (N_3725,N_275,N_1395);
nand U3726 (N_3726,N_1296,N_1404);
nor U3727 (N_3727,N_2437,N_429);
xnor U3728 (N_3728,N_578,N_538);
and U3729 (N_3729,N_312,N_1280);
and U3730 (N_3730,N_759,N_1592);
or U3731 (N_3731,N_1910,N_494);
or U3732 (N_3732,N_330,N_998);
nor U3733 (N_3733,N_1389,N_2256);
or U3734 (N_3734,N_2021,N_215);
and U3735 (N_3735,N_1832,N_1252);
nor U3736 (N_3736,N_2396,N_977);
xor U3737 (N_3737,N_2222,N_1215);
nor U3738 (N_3738,N_2250,N_1508);
nand U3739 (N_3739,N_2375,N_310);
xor U3740 (N_3740,N_1622,N_852);
and U3741 (N_3741,N_1679,N_1656);
xnor U3742 (N_3742,N_2029,N_265);
and U3743 (N_3743,N_2023,N_350);
nor U3744 (N_3744,N_1449,N_1921);
xor U3745 (N_3745,N_1006,N_2134);
nor U3746 (N_3746,N_2495,N_1767);
and U3747 (N_3747,N_944,N_1568);
nand U3748 (N_3748,N_2175,N_1162);
nor U3749 (N_3749,N_1969,N_1197);
or U3750 (N_3750,N_1220,N_2027);
and U3751 (N_3751,N_161,N_2247);
xor U3752 (N_3752,N_312,N_232);
nand U3753 (N_3753,N_18,N_639);
and U3754 (N_3754,N_1482,N_2037);
or U3755 (N_3755,N_1871,N_523);
nor U3756 (N_3756,N_100,N_281);
nor U3757 (N_3757,N_1067,N_684);
and U3758 (N_3758,N_646,N_492);
xor U3759 (N_3759,N_2334,N_2343);
nor U3760 (N_3760,N_1692,N_932);
nor U3761 (N_3761,N_610,N_36);
or U3762 (N_3762,N_741,N_488);
nand U3763 (N_3763,N_1527,N_947);
and U3764 (N_3764,N_1305,N_1623);
xnor U3765 (N_3765,N_1594,N_1878);
and U3766 (N_3766,N_1914,N_476);
and U3767 (N_3767,N_1225,N_1688);
nor U3768 (N_3768,N_920,N_39);
and U3769 (N_3769,N_1641,N_1406);
nor U3770 (N_3770,N_859,N_359);
nand U3771 (N_3771,N_1910,N_2138);
xnor U3772 (N_3772,N_1436,N_1201);
and U3773 (N_3773,N_1931,N_2196);
nand U3774 (N_3774,N_33,N_2224);
nor U3775 (N_3775,N_337,N_165);
xnor U3776 (N_3776,N_52,N_54);
xor U3777 (N_3777,N_2068,N_310);
or U3778 (N_3778,N_332,N_1593);
xor U3779 (N_3779,N_212,N_1546);
or U3780 (N_3780,N_2267,N_233);
nand U3781 (N_3781,N_1920,N_100);
and U3782 (N_3782,N_638,N_1930);
or U3783 (N_3783,N_833,N_1291);
xor U3784 (N_3784,N_2121,N_519);
and U3785 (N_3785,N_1790,N_2244);
and U3786 (N_3786,N_2082,N_1050);
nand U3787 (N_3787,N_1663,N_884);
xnor U3788 (N_3788,N_436,N_653);
nand U3789 (N_3789,N_1518,N_1057);
nor U3790 (N_3790,N_2240,N_1778);
nand U3791 (N_3791,N_1403,N_768);
nand U3792 (N_3792,N_325,N_621);
nand U3793 (N_3793,N_2140,N_670);
nor U3794 (N_3794,N_841,N_1576);
xor U3795 (N_3795,N_2201,N_1441);
nor U3796 (N_3796,N_786,N_2403);
nor U3797 (N_3797,N_1305,N_1401);
xor U3798 (N_3798,N_134,N_1562);
or U3799 (N_3799,N_50,N_855);
xnor U3800 (N_3800,N_2149,N_1560);
or U3801 (N_3801,N_498,N_2419);
nor U3802 (N_3802,N_880,N_712);
nor U3803 (N_3803,N_451,N_1374);
and U3804 (N_3804,N_2442,N_1952);
nor U3805 (N_3805,N_1841,N_2023);
or U3806 (N_3806,N_950,N_1440);
nand U3807 (N_3807,N_2470,N_572);
xnor U3808 (N_3808,N_1118,N_1074);
nor U3809 (N_3809,N_1848,N_922);
nand U3810 (N_3810,N_1469,N_387);
and U3811 (N_3811,N_418,N_503);
xor U3812 (N_3812,N_425,N_72);
nor U3813 (N_3813,N_1086,N_810);
and U3814 (N_3814,N_1867,N_2493);
xnor U3815 (N_3815,N_1712,N_1565);
nor U3816 (N_3816,N_458,N_2435);
xnor U3817 (N_3817,N_2332,N_27);
and U3818 (N_3818,N_1253,N_810);
or U3819 (N_3819,N_1245,N_108);
nor U3820 (N_3820,N_945,N_630);
or U3821 (N_3821,N_305,N_797);
nand U3822 (N_3822,N_2497,N_2216);
or U3823 (N_3823,N_1394,N_2447);
nand U3824 (N_3824,N_248,N_895);
or U3825 (N_3825,N_462,N_800);
xor U3826 (N_3826,N_647,N_661);
nor U3827 (N_3827,N_914,N_1779);
or U3828 (N_3828,N_1337,N_550);
and U3829 (N_3829,N_674,N_909);
nand U3830 (N_3830,N_1013,N_459);
nand U3831 (N_3831,N_366,N_2204);
and U3832 (N_3832,N_1456,N_2097);
nor U3833 (N_3833,N_2018,N_2380);
nor U3834 (N_3834,N_1500,N_1170);
xor U3835 (N_3835,N_1879,N_2222);
and U3836 (N_3836,N_1451,N_1164);
nor U3837 (N_3837,N_2181,N_1572);
and U3838 (N_3838,N_52,N_518);
or U3839 (N_3839,N_742,N_958);
nor U3840 (N_3840,N_1138,N_1541);
and U3841 (N_3841,N_1829,N_682);
or U3842 (N_3842,N_229,N_941);
nor U3843 (N_3843,N_1209,N_684);
xnor U3844 (N_3844,N_423,N_267);
nand U3845 (N_3845,N_213,N_1013);
or U3846 (N_3846,N_108,N_1586);
xnor U3847 (N_3847,N_1270,N_23);
xor U3848 (N_3848,N_1584,N_1310);
and U3849 (N_3849,N_1172,N_1749);
and U3850 (N_3850,N_976,N_959);
xnor U3851 (N_3851,N_300,N_1775);
or U3852 (N_3852,N_1810,N_568);
or U3853 (N_3853,N_2390,N_1834);
nor U3854 (N_3854,N_671,N_2367);
xnor U3855 (N_3855,N_766,N_576);
and U3856 (N_3856,N_1069,N_1055);
nand U3857 (N_3857,N_302,N_467);
xor U3858 (N_3858,N_523,N_645);
and U3859 (N_3859,N_1724,N_1087);
and U3860 (N_3860,N_531,N_1539);
and U3861 (N_3861,N_1117,N_2376);
xor U3862 (N_3862,N_67,N_1659);
or U3863 (N_3863,N_323,N_1175);
and U3864 (N_3864,N_2137,N_436);
or U3865 (N_3865,N_340,N_294);
and U3866 (N_3866,N_728,N_2026);
xor U3867 (N_3867,N_2458,N_1150);
nor U3868 (N_3868,N_1000,N_367);
nor U3869 (N_3869,N_1027,N_1520);
and U3870 (N_3870,N_1498,N_766);
and U3871 (N_3871,N_444,N_2139);
and U3872 (N_3872,N_305,N_1268);
and U3873 (N_3873,N_1911,N_2196);
xor U3874 (N_3874,N_1548,N_768);
xor U3875 (N_3875,N_1322,N_541);
and U3876 (N_3876,N_2156,N_673);
or U3877 (N_3877,N_1474,N_1689);
nor U3878 (N_3878,N_1347,N_695);
nand U3879 (N_3879,N_2182,N_2490);
nor U3880 (N_3880,N_1700,N_1204);
nor U3881 (N_3881,N_1413,N_1205);
nor U3882 (N_3882,N_2496,N_1719);
nor U3883 (N_3883,N_2382,N_1483);
nor U3884 (N_3884,N_470,N_1585);
nor U3885 (N_3885,N_685,N_1642);
or U3886 (N_3886,N_2310,N_523);
xnor U3887 (N_3887,N_1838,N_775);
or U3888 (N_3888,N_1469,N_1600);
nor U3889 (N_3889,N_324,N_583);
and U3890 (N_3890,N_831,N_522);
and U3891 (N_3891,N_1617,N_2262);
or U3892 (N_3892,N_1933,N_52);
and U3893 (N_3893,N_1403,N_922);
or U3894 (N_3894,N_805,N_2077);
or U3895 (N_3895,N_1889,N_996);
xor U3896 (N_3896,N_2002,N_1634);
xor U3897 (N_3897,N_275,N_1337);
or U3898 (N_3898,N_858,N_2181);
nand U3899 (N_3899,N_51,N_1945);
and U3900 (N_3900,N_1015,N_1327);
xor U3901 (N_3901,N_1611,N_1599);
xnor U3902 (N_3902,N_1019,N_801);
and U3903 (N_3903,N_1986,N_54);
nand U3904 (N_3904,N_366,N_1246);
xnor U3905 (N_3905,N_1998,N_1571);
and U3906 (N_3906,N_511,N_24);
or U3907 (N_3907,N_1289,N_2030);
nor U3908 (N_3908,N_1067,N_176);
xnor U3909 (N_3909,N_603,N_2239);
or U3910 (N_3910,N_2195,N_426);
or U3911 (N_3911,N_974,N_2152);
and U3912 (N_3912,N_640,N_218);
or U3913 (N_3913,N_2091,N_1745);
or U3914 (N_3914,N_670,N_1762);
nor U3915 (N_3915,N_37,N_2149);
and U3916 (N_3916,N_2116,N_424);
nor U3917 (N_3917,N_1156,N_1509);
nand U3918 (N_3918,N_201,N_29);
nor U3919 (N_3919,N_894,N_1818);
or U3920 (N_3920,N_1602,N_697);
and U3921 (N_3921,N_109,N_549);
nand U3922 (N_3922,N_1851,N_1153);
and U3923 (N_3923,N_437,N_266);
and U3924 (N_3924,N_1534,N_2072);
xnor U3925 (N_3925,N_1907,N_1426);
nand U3926 (N_3926,N_567,N_679);
xor U3927 (N_3927,N_490,N_1716);
nor U3928 (N_3928,N_1492,N_488);
nand U3929 (N_3929,N_1894,N_1757);
xnor U3930 (N_3930,N_95,N_2394);
nor U3931 (N_3931,N_1465,N_45);
and U3932 (N_3932,N_1236,N_798);
or U3933 (N_3933,N_1383,N_2184);
nor U3934 (N_3934,N_1723,N_1480);
or U3935 (N_3935,N_1519,N_1087);
nand U3936 (N_3936,N_348,N_391);
or U3937 (N_3937,N_1313,N_1116);
nand U3938 (N_3938,N_2137,N_2464);
nand U3939 (N_3939,N_1637,N_2422);
nand U3940 (N_3940,N_987,N_2137);
xor U3941 (N_3941,N_775,N_1266);
nand U3942 (N_3942,N_2049,N_1566);
nand U3943 (N_3943,N_998,N_1654);
nand U3944 (N_3944,N_1882,N_566);
or U3945 (N_3945,N_1011,N_1815);
xnor U3946 (N_3946,N_480,N_1885);
xor U3947 (N_3947,N_1296,N_2064);
nand U3948 (N_3948,N_1610,N_531);
xor U3949 (N_3949,N_729,N_231);
and U3950 (N_3950,N_2368,N_1416);
nor U3951 (N_3951,N_1165,N_2204);
nand U3952 (N_3952,N_370,N_1579);
nor U3953 (N_3953,N_1402,N_1549);
nand U3954 (N_3954,N_965,N_985);
nand U3955 (N_3955,N_2031,N_2117);
and U3956 (N_3956,N_8,N_1964);
xor U3957 (N_3957,N_2000,N_209);
xnor U3958 (N_3958,N_923,N_1532);
xnor U3959 (N_3959,N_1223,N_1339);
or U3960 (N_3960,N_555,N_1893);
and U3961 (N_3961,N_294,N_651);
nand U3962 (N_3962,N_802,N_2289);
or U3963 (N_3963,N_247,N_997);
nor U3964 (N_3964,N_2080,N_1970);
xor U3965 (N_3965,N_299,N_565);
nand U3966 (N_3966,N_2363,N_1658);
nor U3967 (N_3967,N_1039,N_92);
and U3968 (N_3968,N_502,N_616);
nor U3969 (N_3969,N_2064,N_2180);
nand U3970 (N_3970,N_1796,N_1389);
nand U3971 (N_3971,N_2293,N_2263);
or U3972 (N_3972,N_925,N_2334);
or U3973 (N_3973,N_115,N_1241);
xnor U3974 (N_3974,N_2298,N_596);
xnor U3975 (N_3975,N_1027,N_2312);
nor U3976 (N_3976,N_238,N_1875);
nand U3977 (N_3977,N_2350,N_679);
nor U3978 (N_3978,N_1476,N_1677);
nor U3979 (N_3979,N_561,N_812);
nor U3980 (N_3980,N_1616,N_2436);
and U3981 (N_3981,N_9,N_2342);
xnor U3982 (N_3982,N_1190,N_434);
nand U3983 (N_3983,N_462,N_950);
or U3984 (N_3984,N_986,N_2190);
or U3985 (N_3985,N_2240,N_1327);
nand U3986 (N_3986,N_1460,N_1398);
and U3987 (N_3987,N_680,N_558);
nand U3988 (N_3988,N_1433,N_1364);
nand U3989 (N_3989,N_293,N_496);
xor U3990 (N_3990,N_656,N_1823);
and U3991 (N_3991,N_147,N_1597);
xnor U3992 (N_3992,N_2261,N_2270);
xnor U3993 (N_3993,N_1386,N_1206);
and U3994 (N_3994,N_1847,N_201);
nor U3995 (N_3995,N_726,N_211);
and U3996 (N_3996,N_391,N_59);
xor U3997 (N_3997,N_1292,N_1522);
nor U3998 (N_3998,N_1063,N_463);
nand U3999 (N_3999,N_895,N_1545);
and U4000 (N_4000,N_397,N_877);
and U4001 (N_4001,N_2368,N_212);
nand U4002 (N_4002,N_67,N_1948);
nand U4003 (N_4003,N_431,N_1353);
and U4004 (N_4004,N_1524,N_763);
or U4005 (N_4005,N_1929,N_240);
nor U4006 (N_4006,N_1557,N_53);
xor U4007 (N_4007,N_1896,N_2106);
and U4008 (N_4008,N_1441,N_1943);
nor U4009 (N_4009,N_356,N_179);
or U4010 (N_4010,N_2402,N_2267);
or U4011 (N_4011,N_2125,N_671);
xnor U4012 (N_4012,N_825,N_1860);
nand U4013 (N_4013,N_1323,N_2096);
nand U4014 (N_4014,N_1546,N_516);
xnor U4015 (N_4015,N_1380,N_1504);
nand U4016 (N_4016,N_443,N_2115);
nor U4017 (N_4017,N_862,N_502);
nand U4018 (N_4018,N_395,N_1225);
nor U4019 (N_4019,N_2453,N_420);
and U4020 (N_4020,N_120,N_1401);
nand U4021 (N_4021,N_224,N_383);
and U4022 (N_4022,N_529,N_176);
xnor U4023 (N_4023,N_2457,N_1094);
xnor U4024 (N_4024,N_2444,N_2225);
xor U4025 (N_4025,N_2132,N_1053);
or U4026 (N_4026,N_297,N_549);
xor U4027 (N_4027,N_1081,N_524);
and U4028 (N_4028,N_2034,N_153);
or U4029 (N_4029,N_1443,N_1918);
or U4030 (N_4030,N_130,N_2347);
nor U4031 (N_4031,N_942,N_2344);
nor U4032 (N_4032,N_1952,N_1810);
nand U4033 (N_4033,N_1519,N_1234);
xnor U4034 (N_4034,N_1514,N_1314);
or U4035 (N_4035,N_2429,N_1962);
xnor U4036 (N_4036,N_1610,N_748);
xor U4037 (N_4037,N_303,N_1323);
xnor U4038 (N_4038,N_189,N_1716);
nand U4039 (N_4039,N_369,N_2251);
nand U4040 (N_4040,N_1388,N_695);
nand U4041 (N_4041,N_278,N_2080);
nor U4042 (N_4042,N_42,N_62);
nor U4043 (N_4043,N_872,N_1642);
nor U4044 (N_4044,N_987,N_2094);
and U4045 (N_4045,N_701,N_1006);
xor U4046 (N_4046,N_1873,N_2200);
xor U4047 (N_4047,N_1136,N_158);
xor U4048 (N_4048,N_565,N_635);
nand U4049 (N_4049,N_1478,N_2183);
and U4050 (N_4050,N_1896,N_1436);
nor U4051 (N_4051,N_2478,N_760);
nor U4052 (N_4052,N_1751,N_552);
xnor U4053 (N_4053,N_1763,N_2114);
xor U4054 (N_4054,N_1934,N_1723);
or U4055 (N_4055,N_66,N_1016);
nand U4056 (N_4056,N_1401,N_1897);
and U4057 (N_4057,N_1941,N_2392);
nor U4058 (N_4058,N_1798,N_1245);
and U4059 (N_4059,N_159,N_584);
or U4060 (N_4060,N_172,N_432);
or U4061 (N_4061,N_209,N_478);
xnor U4062 (N_4062,N_46,N_1621);
and U4063 (N_4063,N_1226,N_492);
nor U4064 (N_4064,N_725,N_1705);
and U4065 (N_4065,N_759,N_777);
or U4066 (N_4066,N_23,N_596);
xnor U4067 (N_4067,N_469,N_217);
xnor U4068 (N_4068,N_112,N_913);
or U4069 (N_4069,N_839,N_2371);
nand U4070 (N_4070,N_1001,N_2244);
nand U4071 (N_4071,N_122,N_385);
and U4072 (N_4072,N_598,N_984);
nand U4073 (N_4073,N_1730,N_326);
and U4074 (N_4074,N_734,N_952);
nor U4075 (N_4075,N_624,N_3);
xnor U4076 (N_4076,N_1996,N_1258);
and U4077 (N_4077,N_573,N_1428);
nand U4078 (N_4078,N_153,N_2045);
or U4079 (N_4079,N_1271,N_1535);
or U4080 (N_4080,N_463,N_1562);
and U4081 (N_4081,N_484,N_1858);
or U4082 (N_4082,N_205,N_820);
xor U4083 (N_4083,N_913,N_2063);
nand U4084 (N_4084,N_2086,N_1358);
xor U4085 (N_4085,N_1651,N_2470);
or U4086 (N_4086,N_1819,N_198);
nand U4087 (N_4087,N_911,N_1574);
xnor U4088 (N_4088,N_2330,N_2184);
nand U4089 (N_4089,N_1083,N_1392);
or U4090 (N_4090,N_2437,N_2367);
or U4091 (N_4091,N_1400,N_1359);
xnor U4092 (N_4092,N_185,N_2445);
nor U4093 (N_4093,N_1350,N_1000);
xnor U4094 (N_4094,N_1691,N_2429);
and U4095 (N_4095,N_2312,N_465);
nand U4096 (N_4096,N_1726,N_148);
nor U4097 (N_4097,N_2001,N_575);
and U4098 (N_4098,N_2258,N_1583);
nor U4099 (N_4099,N_965,N_2048);
xor U4100 (N_4100,N_924,N_2271);
nor U4101 (N_4101,N_411,N_571);
xnor U4102 (N_4102,N_658,N_467);
nand U4103 (N_4103,N_471,N_2078);
xnor U4104 (N_4104,N_502,N_822);
xor U4105 (N_4105,N_1326,N_1702);
or U4106 (N_4106,N_906,N_801);
or U4107 (N_4107,N_717,N_1269);
or U4108 (N_4108,N_2283,N_2340);
xnor U4109 (N_4109,N_1801,N_405);
and U4110 (N_4110,N_332,N_532);
nand U4111 (N_4111,N_542,N_2283);
and U4112 (N_4112,N_1452,N_1428);
and U4113 (N_4113,N_31,N_143);
or U4114 (N_4114,N_2243,N_1184);
and U4115 (N_4115,N_647,N_796);
nand U4116 (N_4116,N_1556,N_1087);
nand U4117 (N_4117,N_1142,N_738);
nand U4118 (N_4118,N_1189,N_777);
or U4119 (N_4119,N_1811,N_595);
nand U4120 (N_4120,N_219,N_1492);
or U4121 (N_4121,N_1430,N_193);
or U4122 (N_4122,N_495,N_1687);
nor U4123 (N_4123,N_1015,N_535);
and U4124 (N_4124,N_1152,N_1779);
and U4125 (N_4125,N_182,N_30);
nand U4126 (N_4126,N_291,N_305);
nand U4127 (N_4127,N_1935,N_2043);
and U4128 (N_4128,N_516,N_1241);
xnor U4129 (N_4129,N_30,N_2456);
nor U4130 (N_4130,N_2450,N_471);
or U4131 (N_4131,N_1987,N_418);
and U4132 (N_4132,N_1615,N_1022);
nand U4133 (N_4133,N_1139,N_1093);
xnor U4134 (N_4134,N_1412,N_1572);
or U4135 (N_4135,N_1745,N_291);
nor U4136 (N_4136,N_380,N_513);
xor U4137 (N_4137,N_1485,N_2265);
or U4138 (N_4138,N_2378,N_553);
nor U4139 (N_4139,N_2015,N_1242);
and U4140 (N_4140,N_1444,N_2200);
xor U4141 (N_4141,N_2346,N_447);
xor U4142 (N_4142,N_1506,N_1003);
nor U4143 (N_4143,N_1114,N_452);
xor U4144 (N_4144,N_2387,N_1221);
and U4145 (N_4145,N_2167,N_602);
nor U4146 (N_4146,N_2026,N_1550);
nand U4147 (N_4147,N_845,N_783);
nand U4148 (N_4148,N_54,N_2044);
xor U4149 (N_4149,N_1122,N_1456);
and U4150 (N_4150,N_1215,N_468);
nor U4151 (N_4151,N_2290,N_73);
or U4152 (N_4152,N_1244,N_1392);
nand U4153 (N_4153,N_386,N_1337);
or U4154 (N_4154,N_1096,N_896);
or U4155 (N_4155,N_2200,N_1462);
nand U4156 (N_4156,N_2145,N_125);
nand U4157 (N_4157,N_2357,N_364);
and U4158 (N_4158,N_809,N_1187);
and U4159 (N_4159,N_1992,N_1337);
and U4160 (N_4160,N_2066,N_760);
nand U4161 (N_4161,N_1482,N_28);
nor U4162 (N_4162,N_2208,N_1425);
or U4163 (N_4163,N_2242,N_1384);
xnor U4164 (N_4164,N_430,N_2205);
nand U4165 (N_4165,N_649,N_2293);
or U4166 (N_4166,N_1309,N_153);
and U4167 (N_4167,N_371,N_174);
or U4168 (N_4168,N_1208,N_1129);
and U4169 (N_4169,N_500,N_2082);
nand U4170 (N_4170,N_268,N_1514);
nand U4171 (N_4171,N_1990,N_249);
nand U4172 (N_4172,N_1652,N_944);
and U4173 (N_4173,N_1584,N_1036);
or U4174 (N_4174,N_1343,N_2014);
nor U4175 (N_4175,N_203,N_762);
nor U4176 (N_4176,N_21,N_2452);
or U4177 (N_4177,N_1282,N_1852);
nand U4178 (N_4178,N_2396,N_1405);
and U4179 (N_4179,N_175,N_260);
and U4180 (N_4180,N_56,N_679);
xor U4181 (N_4181,N_479,N_1735);
nand U4182 (N_4182,N_338,N_229);
or U4183 (N_4183,N_992,N_1269);
and U4184 (N_4184,N_698,N_2343);
and U4185 (N_4185,N_590,N_2406);
nor U4186 (N_4186,N_1749,N_749);
or U4187 (N_4187,N_1199,N_603);
and U4188 (N_4188,N_1805,N_1403);
or U4189 (N_4189,N_1122,N_617);
nor U4190 (N_4190,N_244,N_1009);
nand U4191 (N_4191,N_2403,N_394);
nor U4192 (N_4192,N_913,N_566);
nand U4193 (N_4193,N_100,N_1854);
nor U4194 (N_4194,N_2287,N_1028);
nor U4195 (N_4195,N_770,N_181);
nand U4196 (N_4196,N_955,N_531);
and U4197 (N_4197,N_2402,N_2485);
nand U4198 (N_4198,N_232,N_811);
nand U4199 (N_4199,N_1057,N_316);
or U4200 (N_4200,N_852,N_842);
and U4201 (N_4201,N_1734,N_604);
or U4202 (N_4202,N_249,N_1260);
and U4203 (N_4203,N_19,N_1655);
or U4204 (N_4204,N_2410,N_1551);
or U4205 (N_4205,N_1102,N_935);
nand U4206 (N_4206,N_2283,N_985);
or U4207 (N_4207,N_2378,N_1709);
nand U4208 (N_4208,N_969,N_2388);
xor U4209 (N_4209,N_1646,N_1788);
xnor U4210 (N_4210,N_1413,N_256);
and U4211 (N_4211,N_105,N_1469);
and U4212 (N_4212,N_1792,N_332);
nor U4213 (N_4213,N_226,N_2371);
and U4214 (N_4214,N_265,N_1628);
nand U4215 (N_4215,N_124,N_1687);
and U4216 (N_4216,N_2414,N_1713);
xnor U4217 (N_4217,N_366,N_1275);
or U4218 (N_4218,N_1420,N_1249);
nand U4219 (N_4219,N_293,N_2455);
and U4220 (N_4220,N_2427,N_1454);
and U4221 (N_4221,N_483,N_1835);
nor U4222 (N_4222,N_596,N_1631);
nor U4223 (N_4223,N_1851,N_1784);
nor U4224 (N_4224,N_1971,N_2027);
nor U4225 (N_4225,N_1044,N_620);
xnor U4226 (N_4226,N_372,N_868);
nand U4227 (N_4227,N_1448,N_150);
or U4228 (N_4228,N_1881,N_1546);
and U4229 (N_4229,N_2295,N_2203);
xnor U4230 (N_4230,N_1722,N_1559);
nand U4231 (N_4231,N_354,N_2360);
or U4232 (N_4232,N_770,N_1839);
xnor U4233 (N_4233,N_2493,N_877);
nor U4234 (N_4234,N_784,N_97);
and U4235 (N_4235,N_294,N_887);
nor U4236 (N_4236,N_26,N_2260);
and U4237 (N_4237,N_1812,N_2231);
nand U4238 (N_4238,N_2462,N_1425);
or U4239 (N_4239,N_2460,N_216);
nand U4240 (N_4240,N_580,N_2182);
nor U4241 (N_4241,N_673,N_1688);
xor U4242 (N_4242,N_289,N_1938);
xnor U4243 (N_4243,N_1506,N_2312);
xor U4244 (N_4244,N_1521,N_445);
xnor U4245 (N_4245,N_1510,N_1809);
and U4246 (N_4246,N_47,N_1281);
xor U4247 (N_4247,N_2431,N_276);
and U4248 (N_4248,N_1754,N_1425);
nor U4249 (N_4249,N_199,N_1709);
and U4250 (N_4250,N_1201,N_1166);
and U4251 (N_4251,N_2321,N_244);
or U4252 (N_4252,N_789,N_2118);
and U4253 (N_4253,N_1377,N_491);
xnor U4254 (N_4254,N_175,N_2121);
xor U4255 (N_4255,N_1967,N_1711);
or U4256 (N_4256,N_649,N_2305);
xor U4257 (N_4257,N_1692,N_2051);
and U4258 (N_4258,N_2040,N_776);
nand U4259 (N_4259,N_1169,N_397);
and U4260 (N_4260,N_1786,N_857);
nand U4261 (N_4261,N_509,N_1887);
nand U4262 (N_4262,N_251,N_1818);
and U4263 (N_4263,N_83,N_649);
nand U4264 (N_4264,N_1359,N_1543);
or U4265 (N_4265,N_341,N_226);
or U4266 (N_4266,N_222,N_246);
xor U4267 (N_4267,N_9,N_1278);
and U4268 (N_4268,N_99,N_2231);
or U4269 (N_4269,N_1536,N_1532);
xnor U4270 (N_4270,N_282,N_1084);
nor U4271 (N_4271,N_1948,N_30);
and U4272 (N_4272,N_554,N_948);
or U4273 (N_4273,N_137,N_9);
nand U4274 (N_4274,N_1604,N_544);
xor U4275 (N_4275,N_369,N_1041);
or U4276 (N_4276,N_103,N_336);
nand U4277 (N_4277,N_637,N_2343);
or U4278 (N_4278,N_1224,N_61);
xor U4279 (N_4279,N_2072,N_367);
and U4280 (N_4280,N_1181,N_547);
and U4281 (N_4281,N_2377,N_290);
nor U4282 (N_4282,N_1147,N_1936);
or U4283 (N_4283,N_1252,N_1382);
nor U4284 (N_4284,N_2151,N_190);
and U4285 (N_4285,N_644,N_208);
nand U4286 (N_4286,N_1084,N_2306);
and U4287 (N_4287,N_1374,N_76);
xnor U4288 (N_4288,N_1035,N_415);
or U4289 (N_4289,N_2148,N_346);
nor U4290 (N_4290,N_2489,N_488);
or U4291 (N_4291,N_1668,N_2357);
xor U4292 (N_4292,N_514,N_93);
or U4293 (N_4293,N_1089,N_1355);
and U4294 (N_4294,N_1301,N_1565);
nor U4295 (N_4295,N_2470,N_1873);
and U4296 (N_4296,N_713,N_958);
xnor U4297 (N_4297,N_693,N_258);
nand U4298 (N_4298,N_1655,N_550);
or U4299 (N_4299,N_1976,N_2177);
nand U4300 (N_4300,N_217,N_2127);
nor U4301 (N_4301,N_2119,N_2373);
and U4302 (N_4302,N_1452,N_204);
or U4303 (N_4303,N_1599,N_2178);
xor U4304 (N_4304,N_2198,N_2405);
xor U4305 (N_4305,N_1825,N_1730);
and U4306 (N_4306,N_441,N_1801);
nor U4307 (N_4307,N_733,N_1850);
xor U4308 (N_4308,N_769,N_1249);
and U4309 (N_4309,N_2441,N_1758);
or U4310 (N_4310,N_1038,N_1802);
and U4311 (N_4311,N_1225,N_2404);
xnor U4312 (N_4312,N_1692,N_499);
and U4313 (N_4313,N_1841,N_1506);
xor U4314 (N_4314,N_419,N_790);
nand U4315 (N_4315,N_2186,N_2234);
and U4316 (N_4316,N_520,N_1279);
nand U4317 (N_4317,N_1186,N_676);
xor U4318 (N_4318,N_555,N_837);
or U4319 (N_4319,N_1144,N_441);
and U4320 (N_4320,N_2293,N_1153);
nor U4321 (N_4321,N_492,N_2374);
nor U4322 (N_4322,N_318,N_1105);
xor U4323 (N_4323,N_1850,N_333);
and U4324 (N_4324,N_963,N_639);
or U4325 (N_4325,N_2377,N_1547);
or U4326 (N_4326,N_1249,N_584);
nand U4327 (N_4327,N_113,N_811);
and U4328 (N_4328,N_820,N_202);
xnor U4329 (N_4329,N_124,N_925);
nor U4330 (N_4330,N_1605,N_305);
and U4331 (N_4331,N_2119,N_522);
nor U4332 (N_4332,N_2364,N_161);
xnor U4333 (N_4333,N_922,N_1158);
nor U4334 (N_4334,N_36,N_1486);
or U4335 (N_4335,N_173,N_1629);
nor U4336 (N_4336,N_82,N_1086);
nor U4337 (N_4337,N_2216,N_922);
xnor U4338 (N_4338,N_1245,N_522);
or U4339 (N_4339,N_438,N_633);
or U4340 (N_4340,N_77,N_1286);
nor U4341 (N_4341,N_1271,N_873);
xor U4342 (N_4342,N_1353,N_103);
nor U4343 (N_4343,N_1656,N_2184);
or U4344 (N_4344,N_1635,N_405);
xnor U4345 (N_4345,N_1108,N_310);
xor U4346 (N_4346,N_2441,N_772);
nor U4347 (N_4347,N_47,N_1179);
or U4348 (N_4348,N_1165,N_1615);
xor U4349 (N_4349,N_625,N_1248);
nor U4350 (N_4350,N_1572,N_2334);
nand U4351 (N_4351,N_2118,N_1219);
and U4352 (N_4352,N_257,N_956);
nor U4353 (N_4353,N_713,N_414);
xor U4354 (N_4354,N_1267,N_1268);
xor U4355 (N_4355,N_1133,N_736);
xnor U4356 (N_4356,N_638,N_1549);
xnor U4357 (N_4357,N_178,N_2306);
or U4358 (N_4358,N_1219,N_956);
nor U4359 (N_4359,N_793,N_1540);
nand U4360 (N_4360,N_1677,N_623);
or U4361 (N_4361,N_1869,N_987);
and U4362 (N_4362,N_1157,N_273);
nand U4363 (N_4363,N_550,N_2136);
or U4364 (N_4364,N_1019,N_1926);
xnor U4365 (N_4365,N_1727,N_1648);
xnor U4366 (N_4366,N_1143,N_100);
nand U4367 (N_4367,N_1575,N_76);
or U4368 (N_4368,N_2315,N_1785);
xnor U4369 (N_4369,N_2010,N_770);
xor U4370 (N_4370,N_314,N_1687);
nand U4371 (N_4371,N_1660,N_545);
nand U4372 (N_4372,N_1416,N_218);
nor U4373 (N_4373,N_1331,N_639);
and U4374 (N_4374,N_228,N_1077);
nand U4375 (N_4375,N_742,N_398);
nor U4376 (N_4376,N_777,N_1714);
nand U4377 (N_4377,N_584,N_675);
and U4378 (N_4378,N_137,N_1262);
or U4379 (N_4379,N_1505,N_227);
or U4380 (N_4380,N_2174,N_857);
and U4381 (N_4381,N_1479,N_104);
and U4382 (N_4382,N_208,N_1793);
and U4383 (N_4383,N_1068,N_2401);
or U4384 (N_4384,N_1420,N_608);
nand U4385 (N_4385,N_495,N_1374);
nor U4386 (N_4386,N_1167,N_1854);
nand U4387 (N_4387,N_1725,N_590);
or U4388 (N_4388,N_347,N_1024);
nand U4389 (N_4389,N_1415,N_1177);
and U4390 (N_4390,N_522,N_1575);
xor U4391 (N_4391,N_595,N_1828);
and U4392 (N_4392,N_129,N_62);
nand U4393 (N_4393,N_799,N_377);
nor U4394 (N_4394,N_878,N_2461);
or U4395 (N_4395,N_1904,N_275);
nand U4396 (N_4396,N_1960,N_2476);
nor U4397 (N_4397,N_1384,N_165);
or U4398 (N_4398,N_175,N_21);
nand U4399 (N_4399,N_94,N_2100);
or U4400 (N_4400,N_1159,N_2231);
or U4401 (N_4401,N_2341,N_952);
nand U4402 (N_4402,N_1016,N_2424);
xnor U4403 (N_4403,N_1375,N_1528);
xnor U4404 (N_4404,N_1867,N_693);
xnor U4405 (N_4405,N_2380,N_2100);
xnor U4406 (N_4406,N_354,N_1371);
or U4407 (N_4407,N_157,N_14);
and U4408 (N_4408,N_1872,N_897);
nand U4409 (N_4409,N_196,N_1146);
nor U4410 (N_4410,N_338,N_1002);
nand U4411 (N_4411,N_485,N_2131);
nand U4412 (N_4412,N_2227,N_181);
and U4413 (N_4413,N_2356,N_476);
and U4414 (N_4414,N_752,N_773);
and U4415 (N_4415,N_2325,N_2099);
nor U4416 (N_4416,N_305,N_691);
nand U4417 (N_4417,N_732,N_2167);
nor U4418 (N_4418,N_1596,N_1593);
or U4419 (N_4419,N_266,N_2400);
nand U4420 (N_4420,N_264,N_2202);
nand U4421 (N_4421,N_932,N_345);
xor U4422 (N_4422,N_2219,N_577);
nor U4423 (N_4423,N_171,N_1119);
and U4424 (N_4424,N_2474,N_482);
or U4425 (N_4425,N_1323,N_27);
xnor U4426 (N_4426,N_1422,N_902);
nand U4427 (N_4427,N_1668,N_1004);
nand U4428 (N_4428,N_1539,N_748);
or U4429 (N_4429,N_2440,N_166);
nor U4430 (N_4430,N_826,N_947);
or U4431 (N_4431,N_568,N_2152);
or U4432 (N_4432,N_1876,N_638);
or U4433 (N_4433,N_309,N_1733);
or U4434 (N_4434,N_1990,N_742);
or U4435 (N_4435,N_1468,N_221);
nor U4436 (N_4436,N_1385,N_949);
xor U4437 (N_4437,N_1378,N_249);
and U4438 (N_4438,N_1455,N_499);
nand U4439 (N_4439,N_672,N_332);
xor U4440 (N_4440,N_1254,N_1200);
nand U4441 (N_4441,N_1539,N_1567);
nor U4442 (N_4442,N_1600,N_1505);
nor U4443 (N_4443,N_2134,N_1457);
or U4444 (N_4444,N_814,N_1543);
and U4445 (N_4445,N_243,N_304);
nand U4446 (N_4446,N_1380,N_1903);
nand U4447 (N_4447,N_2071,N_645);
nand U4448 (N_4448,N_2110,N_2471);
or U4449 (N_4449,N_1063,N_1172);
xor U4450 (N_4450,N_2467,N_882);
or U4451 (N_4451,N_695,N_813);
xor U4452 (N_4452,N_1942,N_1775);
nor U4453 (N_4453,N_1484,N_811);
or U4454 (N_4454,N_1025,N_174);
and U4455 (N_4455,N_1725,N_1298);
and U4456 (N_4456,N_678,N_474);
and U4457 (N_4457,N_1784,N_507);
nor U4458 (N_4458,N_1555,N_1307);
and U4459 (N_4459,N_505,N_2147);
xnor U4460 (N_4460,N_1256,N_1752);
nor U4461 (N_4461,N_1765,N_2064);
nor U4462 (N_4462,N_1586,N_1715);
or U4463 (N_4463,N_918,N_2165);
nand U4464 (N_4464,N_524,N_1679);
or U4465 (N_4465,N_70,N_987);
nor U4466 (N_4466,N_8,N_1098);
or U4467 (N_4467,N_2020,N_407);
xnor U4468 (N_4468,N_1123,N_502);
and U4469 (N_4469,N_1747,N_1780);
and U4470 (N_4470,N_176,N_1074);
and U4471 (N_4471,N_5,N_2061);
nor U4472 (N_4472,N_271,N_80);
and U4473 (N_4473,N_2085,N_1799);
nor U4474 (N_4474,N_1220,N_45);
or U4475 (N_4475,N_1008,N_1291);
nand U4476 (N_4476,N_2444,N_1732);
and U4477 (N_4477,N_545,N_118);
nor U4478 (N_4478,N_1133,N_1155);
nor U4479 (N_4479,N_79,N_1854);
nor U4480 (N_4480,N_1290,N_1200);
or U4481 (N_4481,N_852,N_1864);
or U4482 (N_4482,N_315,N_1502);
nor U4483 (N_4483,N_2238,N_678);
nand U4484 (N_4484,N_583,N_1030);
nor U4485 (N_4485,N_1486,N_121);
nor U4486 (N_4486,N_1835,N_1903);
nor U4487 (N_4487,N_1514,N_1998);
and U4488 (N_4488,N_1197,N_967);
and U4489 (N_4489,N_2084,N_967);
or U4490 (N_4490,N_2154,N_322);
nand U4491 (N_4491,N_1056,N_2262);
nand U4492 (N_4492,N_2338,N_2482);
xnor U4493 (N_4493,N_595,N_1009);
or U4494 (N_4494,N_757,N_648);
nand U4495 (N_4495,N_1650,N_441);
nand U4496 (N_4496,N_2451,N_1966);
and U4497 (N_4497,N_524,N_1380);
nor U4498 (N_4498,N_847,N_798);
and U4499 (N_4499,N_2495,N_148);
xor U4500 (N_4500,N_171,N_37);
nand U4501 (N_4501,N_2344,N_194);
nand U4502 (N_4502,N_415,N_687);
nor U4503 (N_4503,N_1656,N_1543);
and U4504 (N_4504,N_1982,N_316);
or U4505 (N_4505,N_1091,N_2079);
nand U4506 (N_4506,N_1765,N_374);
nor U4507 (N_4507,N_2022,N_991);
and U4508 (N_4508,N_673,N_184);
nand U4509 (N_4509,N_863,N_2323);
or U4510 (N_4510,N_2101,N_800);
nor U4511 (N_4511,N_553,N_177);
nand U4512 (N_4512,N_1695,N_1311);
nor U4513 (N_4513,N_1246,N_2309);
nor U4514 (N_4514,N_1220,N_924);
nor U4515 (N_4515,N_407,N_539);
nor U4516 (N_4516,N_1397,N_2349);
nand U4517 (N_4517,N_1063,N_838);
xor U4518 (N_4518,N_1740,N_1818);
nand U4519 (N_4519,N_55,N_1610);
nand U4520 (N_4520,N_1477,N_455);
xor U4521 (N_4521,N_2069,N_1379);
nor U4522 (N_4522,N_872,N_486);
nor U4523 (N_4523,N_186,N_2362);
nand U4524 (N_4524,N_218,N_1194);
nor U4525 (N_4525,N_65,N_784);
xor U4526 (N_4526,N_2258,N_272);
xnor U4527 (N_4527,N_1817,N_88);
or U4528 (N_4528,N_1731,N_289);
nor U4529 (N_4529,N_2115,N_738);
xor U4530 (N_4530,N_2086,N_1944);
and U4531 (N_4531,N_548,N_846);
and U4532 (N_4532,N_2431,N_1426);
nor U4533 (N_4533,N_1024,N_493);
or U4534 (N_4534,N_529,N_1169);
nor U4535 (N_4535,N_325,N_1482);
or U4536 (N_4536,N_1913,N_979);
nand U4537 (N_4537,N_2485,N_249);
and U4538 (N_4538,N_1068,N_1270);
and U4539 (N_4539,N_277,N_1469);
and U4540 (N_4540,N_2293,N_1756);
xor U4541 (N_4541,N_89,N_1081);
nand U4542 (N_4542,N_466,N_350);
or U4543 (N_4543,N_1701,N_981);
and U4544 (N_4544,N_2442,N_594);
and U4545 (N_4545,N_540,N_1932);
or U4546 (N_4546,N_338,N_1381);
nand U4547 (N_4547,N_2346,N_2224);
xnor U4548 (N_4548,N_1491,N_650);
and U4549 (N_4549,N_2250,N_1612);
or U4550 (N_4550,N_830,N_1589);
xnor U4551 (N_4551,N_2097,N_1166);
nand U4552 (N_4552,N_1775,N_2406);
or U4553 (N_4553,N_2228,N_315);
nor U4554 (N_4554,N_1264,N_2458);
nand U4555 (N_4555,N_2423,N_790);
or U4556 (N_4556,N_798,N_448);
xor U4557 (N_4557,N_1640,N_2217);
or U4558 (N_4558,N_1940,N_2474);
and U4559 (N_4559,N_1777,N_639);
or U4560 (N_4560,N_906,N_2046);
xnor U4561 (N_4561,N_1635,N_1874);
nor U4562 (N_4562,N_678,N_506);
and U4563 (N_4563,N_2476,N_570);
nor U4564 (N_4564,N_1228,N_447);
nand U4565 (N_4565,N_2164,N_1296);
and U4566 (N_4566,N_238,N_1488);
xnor U4567 (N_4567,N_1047,N_11);
nand U4568 (N_4568,N_2011,N_1267);
nand U4569 (N_4569,N_264,N_67);
or U4570 (N_4570,N_1424,N_360);
or U4571 (N_4571,N_2281,N_586);
nand U4572 (N_4572,N_2457,N_1261);
nor U4573 (N_4573,N_1267,N_677);
nor U4574 (N_4574,N_842,N_702);
nand U4575 (N_4575,N_382,N_1251);
nand U4576 (N_4576,N_1199,N_2353);
nor U4577 (N_4577,N_1154,N_1411);
nand U4578 (N_4578,N_741,N_2195);
nor U4579 (N_4579,N_1825,N_131);
nor U4580 (N_4580,N_2458,N_1320);
xor U4581 (N_4581,N_2422,N_313);
xor U4582 (N_4582,N_1417,N_849);
and U4583 (N_4583,N_2485,N_1414);
or U4584 (N_4584,N_1088,N_23);
xnor U4585 (N_4585,N_1853,N_1319);
and U4586 (N_4586,N_935,N_2401);
nand U4587 (N_4587,N_380,N_1611);
xor U4588 (N_4588,N_175,N_992);
and U4589 (N_4589,N_995,N_2215);
or U4590 (N_4590,N_2364,N_863);
or U4591 (N_4591,N_140,N_641);
nand U4592 (N_4592,N_2281,N_61);
nor U4593 (N_4593,N_696,N_577);
or U4594 (N_4594,N_2496,N_690);
and U4595 (N_4595,N_258,N_2470);
xnor U4596 (N_4596,N_2163,N_1533);
xnor U4597 (N_4597,N_1247,N_959);
or U4598 (N_4598,N_1543,N_2054);
or U4599 (N_4599,N_1670,N_2479);
nand U4600 (N_4600,N_1320,N_2049);
xor U4601 (N_4601,N_1903,N_1984);
or U4602 (N_4602,N_1897,N_1943);
nand U4603 (N_4603,N_1656,N_1989);
nand U4604 (N_4604,N_932,N_1768);
xor U4605 (N_4605,N_2433,N_942);
nor U4606 (N_4606,N_496,N_1894);
nor U4607 (N_4607,N_1870,N_1120);
nor U4608 (N_4608,N_57,N_722);
nand U4609 (N_4609,N_994,N_2450);
xnor U4610 (N_4610,N_1431,N_929);
or U4611 (N_4611,N_1871,N_1592);
nor U4612 (N_4612,N_780,N_589);
nor U4613 (N_4613,N_1094,N_1831);
xor U4614 (N_4614,N_1126,N_740);
and U4615 (N_4615,N_97,N_136);
or U4616 (N_4616,N_239,N_1335);
xor U4617 (N_4617,N_1517,N_1756);
nand U4618 (N_4618,N_541,N_138);
nor U4619 (N_4619,N_417,N_1232);
nand U4620 (N_4620,N_229,N_1100);
nand U4621 (N_4621,N_66,N_75);
nor U4622 (N_4622,N_520,N_1314);
and U4623 (N_4623,N_371,N_237);
xor U4624 (N_4624,N_1301,N_267);
nand U4625 (N_4625,N_88,N_2422);
xnor U4626 (N_4626,N_1812,N_1128);
nor U4627 (N_4627,N_5,N_1356);
nor U4628 (N_4628,N_2464,N_1835);
or U4629 (N_4629,N_1967,N_2215);
or U4630 (N_4630,N_831,N_2402);
or U4631 (N_4631,N_2476,N_2106);
or U4632 (N_4632,N_356,N_2394);
nor U4633 (N_4633,N_2265,N_802);
xnor U4634 (N_4634,N_27,N_1511);
and U4635 (N_4635,N_370,N_2036);
nor U4636 (N_4636,N_1212,N_1236);
nand U4637 (N_4637,N_504,N_31);
nand U4638 (N_4638,N_2239,N_1957);
or U4639 (N_4639,N_2265,N_1807);
nand U4640 (N_4640,N_997,N_2255);
nor U4641 (N_4641,N_525,N_1995);
and U4642 (N_4642,N_901,N_1708);
nand U4643 (N_4643,N_313,N_971);
nand U4644 (N_4644,N_2239,N_2381);
nor U4645 (N_4645,N_488,N_1172);
or U4646 (N_4646,N_1357,N_362);
or U4647 (N_4647,N_91,N_2088);
xnor U4648 (N_4648,N_785,N_416);
nand U4649 (N_4649,N_491,N_2068);
xnor U4650 (N_4650,N_613,N_528);
and U4651 (N_4651,N_430,N_2496);
xor U4652 (N_4652,N_23,N_104);
xor U4653 (N_4653,N_2348,N_756);
or U4654 (N_4654,N_1605,N_55);
or U4655 (N_4655,N_2141,N_1826);
nor U4656 (N_4656,N_1787,N_1034);
and U4657 (N_4657,N_481,N_761);
nor U4658 (N_4658,N_1339,N_139);
nand U4659 (N_4659,N_1507,N_1862);
xnor U4660 (N_4660,N_1042,N_2109);
or U4661 (N_4661,N_510,N_530);
or U4662 (N_4662,N_1767,N_1331);
nor U4663 (N_4663,N_1722,N_1652);
and U4664 (N_4664,N_2248,N_260);
xor U4665 (N_4665,N_1656,N_645);
xnor U4666 (N_4666,N_209,N_2291);
xor U4667 (N_4667,N_983,N_404);
and U4668 (N_4668,N_1782,N_703);
nor U4669 (N_4669,N_2265,N_1033);
or U4670 (N_4670,N_358,N_192);
and U4671 (N_4671,N_2162,N_557);
nor U4672 (N_4672,N_1329,N_2324);
xnor U4673 (N_4673,N_630,N_717);
nand U4674 (N_4674,N_1785,N_386);
xor U4675 (N_4675,N_607,N_1544);
xnor U4676 (N_4676,N_2329,N_260);
or U4677 (N_4677,N_1691,N_882);
nand U4678 (N_4678,N_2320,N_1367);
or U4679 (N_4679,N_1006,N_1575);
xor U4680 (N_4680,N_410,N_920);
nor U4681 (N_4681,N_584,N_1005);
xor U4682 (N_4682,N_1146,N_1701);
and U4683 (N_4683,N_1015,N_1035);
nor U4684 (N_4684,N_893,N_2267);
nand U4685 (N_4685,N_992,N_2316);
and U4686 (N_4686,N_1617,N_1543);
nor U4687 (N_4687,N_1411,N_1005);
nor U4688 (N_4688,N_2084,N_990);
or U4689 (N_4689,N_76,N_238);
nand U4690 (N_4690,N_1500,N_452);
and U4691 (N_4691,N_1913,N_876);
and U4692 (N_4692,N_174,N_10);
xnor U4693 (N_4693,N_609,N_610);
xnor U4694 (N_4694,N_1565,N_1035);
xor U4695 (N_4695,N_1990,N_1885);
and U4696 (N_4696,N_2292,N_2264);
xnor U4697 (N_4697,N_2311,N_880);
xnor U4698 (N_4698,N_2393,N_911);
xor U4699 (N_4699,N_614,N_113);
xor U4700 (N_4700,N_84,N_95);
and U4701 (N_4701,N_580,N_1628);
or U4702 (N_4702,N_449,N_2247);
nand U4703 (N_4703,N_2175,N_434);
nand U4704 (N_4704,N_1771,N_938);
and U4705 (N_4705,N_2275,N_207);
nand U4706 (N_4706,N_1600,N_681);
nor U4707 (N_4707,N_350,N_1223);
or U4708 (N_4708,N_1754,N_2102);
or U4709 (N_4709,N_2325,N_442);
nand U4710 (N_4710,N_2171,N_1590);
and U4711 (N_4711,N_830,N_1804);
xnor U4712 (N_4712,N_1578,N_983);
or U4713 (N_4713,N_2359,N_2224);
or U4714 (N_4714,N_2274,N_2165);
or U4715 (N_4715,N_1934,N_308);
nor U4716 (N_4716,N_229,N_1694);
nand U4717 (N_4717,N_2257,N_122);
or U4718 (N_4718,N_67,N_875);
nor U4719 (N_4719,N_668,N_2261);
nor U4720 (N_4720,N_274,N_1716);
and U4721 (N_4721,N_2028,N_603);
or U4722 (N_4722,N_740,N_2274);
and U4723 (N_4723,N_2066,N_2156);
and U4724 (N_4724,N_1666,N_1224);
and U4725 (N_4725,N_2086,N_1876);
nor U4726 (N_4726,N_966,N_89);
and U4727 (N_4727,N_2171,N_1178);
and U4728 (N_4728,N_1187,N_1782);
nor U4729 (N_4729,N_2402,N_991);
xor U4730 (N_4730,N_1544,N_530);
nand U4731 (N_4731,N_2485,N_1853);
and U4732 (N_4732,N_2139,N_1315);
nand U4733 (N_4733,N_1614,N_35);
or U4734 (N_4734,N_1616,N_2438);
nand U4735 (N_4735,N_1772,N_2293);
and U4736 (N_4736,N_2191,N_2164);
and U4737 (N_4737,N_116,N_1028);
or U4738 (N_4738,N_1085,N_1555);
xnor U4739 (N_4739,N_321,N_1932);
nor U4740 (N_4740,N_1004,N_263);
and U4741 (N_4741,N_2287,N_159);
and U4742 (N_4742,N_1334,N_2217);
nor U4743 (N_4743,N_52,N_2257);
or U4744 (N_4744,N_1191,N_525);
or U4745 (N_4745,N_1987,N_1614);
nor U4746 (N_4746,N_1762,N_983);
nor U4747 (N_4747,N_2115,N_933);
or U4748 (N_4748,N_263,N_2415);
and U4749 (N_4749,N_1266,N_322);
and U4750 (N_4750,N_1034,N_1496);
and U4751 (N_4751,N_1562,N_655);
nor U4752 (N_4752,N_2481,N_832);
nor U4753 (N_4753,N_1295,N_959);
and U4754 (N_4754,N_1172,N_923);
and U4755 (N_4755,N_152,N_2058);
or U4756 (N_4756,N_561,N_2318);
nor U4757 (N_4757,N_1571,N_297);
nor U4758 (N_4758,N_608,N_2145);
xor U4759 (N_4759,N_119,N_1474);
or U4760 (N_4760,N_1213,N_1479);
nor U4761 (N_4761,N_2106,N_1883);
or U4762 (N_4762,N_2170,N_1629);
or U4763 (N_4763,N_1830,N_2231);
nand U4764 (N_4764,N_1560,N_181);
xor U4765 (N_4765,N_445,N_993);
xor U4766 (N_4766,N_927,N_167);
and U4767 (N_4767,N_2482,N_1596);
nand U4768 (N_4768,N_777,N_1965);
nor U4769 (N_4769,N_775,N_511);
nand U4770 (N_4770,N_349,N_2015);
xnor U4771 (N_4771,N_806,N_1161);
nor U4772 (N_4772,N_918,N_2316);
nand U4773 (N_4773,N_2071,N_1791);
and U4774 (N_4774,N_332,N_805);
or U4775 (N_4775,N_1588,N_786);
nand U4776 (N_4776,N_390,N_715);
xor U4777 (N_4777,N_2013,N_1727);
and U4778 (N_4778,N_904,N_2184);
nand U4779 (N_4779,N_1040,N_1919);
or U4780 (N_4780,N_1535,N_878);
xnor U4781 (N_4781,N_337,N_1647);
or U4782 (N_4782,N_2484,N_887);
and U4783 (N_4783,N_409,N_1092);
or U4784 (N_4784,N_2319,N_1902);
nand U4785 (N_4785,N_636,N_1688);
or U4786 (N_4786,N_2412,N_2138);
nor U4787 (N_4787,N_336,N_1267);
and U4788 (N_4788,N_653,N_484);
xnor U4789 (N_4789,N_2431,N_2372);
nand U4790 (N_4790,N_1611,N_1330);
nor U4791 (N_4791,N_775,N_2451);
or U4792 (N_4792,N_352,N_608);
xnor U4793 (N_4793,N_755,N_1038);
or U4794 (N_4794,N_695,N_714);
nand U4795 (N_4795,N_1032,N_536);
nor U4796 (N_4796,N_1640,N_1634);
or U4797 (N_4797,N_2106,N_699);
and U4798 (N_4798,N_1982,N_1077);
nor U4799 (N_4799,N_1817,N_1780);
xor U4800 (N_4800,N_618,N_1033);
or U4801 (N_4801,N_1915,N_1351);
nor U4802 (N_4802,N_2093,N_2339);
xnor U4803 (N_4803,N_1498,N_38);
and U4804 (N_4804,N_1604,N_904);
nor U4805 (N_4805,N_2335,N_1388);
nand U4806 (N_4806,N_126,N_2024);
nor U4807 (N_4807,N_1459,N_2140);
or U4808 (N_4808,N_1613,N_2290);
xnor U4809 (N_4809,N_2345,N_1245);
or U4810 (N_4810,N_1146,N_185);
and U4811 (N_4811,N_170,N_919);
nand U4812 (N_4812,N_948,N_216);
xor U4813 (N_4813,N_919,N_912);
nand U4814 (N_4814,N_752,N_2387);
or U4815 (N_4815,N_1882,N_57);
nor U4816 (N_4816,N_1359,N_1399);
and U4817 (N_4817,N_1135,N_603);
nor U4818 (N_4818,N_209,N_255);
xnor U4819 (N_4819,N_2207,N_241);
or U4820 (N_4820,N_127,N_1938);
xnor U4821 (N_4821,N_573,N_2213);
and U4822 (N_4822,N_927,N_47);
or U4823 (N_4823,N_1027,N_1610);
xnor U4824 (N_4824,N_1165,N_402);
nand U4825 (N_4825,N_1535,N_917);
or U4826 (N_4826,N_1926,N_525);
xnor U4827 (N_4827,N_1776,N_813);
or U4828 (N_4828,N_2283,N_1979);
or U4829 (N_4829,N_435,N_1517);
or U4830 (N_4830,N_2464,N_699);
nand U4831 (N_4831,N_1440,N_1991);
nor U4832 (N_4832,N_138,N_30);
or U4833 (N_4833,N_1005,N_1130);
and U4834 (N_4834,N_1967,N_292);
or U4835 (N_4835,N_1627,N_583);
xnor U4836 (N_4836,N_549,N_2029);
nand U4837 (N_4837,N_574,N_425);
xor U4838 (N_4838,N_1123,N_1943);
or U4839 (N_4839,N_2096,N_2144);
nor U4840 (N_4840,N_2206,N_2235);
xnor U4841 (N_4841,N_799,N_848);
and U4842 (N_4842,N_1020,N_1818);
and U4843 (N_4843,N_967,N_282);
nor U4844 (N_4844,N_1494,N_2218);
and U4845 (N_4845,N_958,N_426);
and U4846 (N_4846,N_319,N_1794);
xnor U4847 (N_4847,N_1237,N_837);
and U4848 (N_4848,N_111,N_343);
xor U4849 (N_4849,N_276,N_1126);
nand U4850 (N_4850,N_1434,N_945);
nor U4851 (N_4851,N_276,N_1068);
and U4852 (N_4852,N_2034,N_1544);
xor U4853 (N_4853,N_530,N_706);
and U4854 (N_4854,N_1713,N_1406);
nor U4855 (N_4855,N_1659,N_493);
or U4856 (N_4856,N_572,N_2157);
nor U4857 (N_4857,N_850,N_14);
and U4858 (N_4858,N_1594,N_356);
nor U4859 (N_4859,N_911,N_1744);
nand U4860 (N_4860,N_398,N_1855);
nor U4861 (N_4861,N_1131,N_1418);
xor U4862 (N_4862,N_2459,N_2187);
nand U4863 (N_4863,N_148,N_156);
xnor U4864 (N_4864,N_554,N_2164);
and U4865 (N_4865,N_252,N_2320);
or U4866 (N_4866,N_910,N_1801);
nand U4867 (N_4867,N_1547,N_2033);
xor U4868 (N_4868,N_741,N_1437);
xnor U4869 (N_4869,N_220,N_261);
or U4870 (N_4870,N_26,N_2351);
nand U4871 (N_4871,N_1237,N_981);
nand U4872 (N_4872,N_1815,N_1319);
or U4873 (N_4873,N_460,N_773);
nand U4874 (N_4874,N_2267,N_158);
nand U4875 (N_4875,N_1808,N_236);
or U4876 (N_4876,N_1712,N_2381);
and U4877 (N_4877,N_1393,N_1956);
nand U4878 (N_4878,N_1452,N_1478);
xor U4879 (N_4879,N_2266,N_1465);
nor U4880 (N_4880,N_2072,N_448);
or U4881 (N_4881,N_2323,N_1590);
nand U4882 (N_4882,N_2232,N_1506);
xnor U4883 (N_4883,N_2407,N_167);
and U4884 (N_4884,N_84,N_1297);
and U4885 (N_4885,N_1780,N_1894);
nand U4886 (N_4886,N_226,N_1444);
or U4887 (N_4887,N_875,N_912);
nor U4888 (N_4888,N_151,N_1064);
or U4889 (N_4889,N_1128,N_1126);
xor U4890 (N_4890,N_901,N_2494);
or U4891 (N_4891,N_1788,N_2165);
nor U4892 (N_4892,N_198,N_273);
nand U4893 (N_4893,N_1990,N_1282);
or U4894 (N_4894,N_1337,N_75);
xnor U4895 (N_4895,N_541,N_2225);
nor U4896 (N_4896,N_1614,N_92);
xor U4897 (N_4897,N_278,N_1189);
and U4898 (N_4898,N_1617,N_1094);
or U4899 (N_4899,N_2316,N_2383);
nand U4900 (N_4900,N_396,N_945);
nor U4901 (N_4901,N_1346,N_1190);
and U4902 (N_4902,N_476,N_413);
or U4903 (N_4903,N_941,N_969);
and U4904 (N_4904,N_1067,N_1890);
and U4905 (N_4905,N_717,N_2214);
and U4906 (N_4906,N_1647,N_1347);
and U4907 (N_4907,N_167,N_573);
or U4908 (N_4908,N_1549,N_1259);
and U4909 (N_4909,N_2081,N_1359);
and U4910 (N_4910,N_2135,N_1381);
nand U4911 (N_4911,N_220,N_2238);
nor U4912 (N_4912,N_549,N_2312);
xor U4913 (N_4913,N_1626,N_997);
xnor U4914 (N_4914,N_2335,N_1565);
nand U4915 (N_4915,N_1582,N_2292);
or U4916 (N_4916,N_755,N_98);
or U4917 (N_4917,N_615,N_1197);
xor U4918 (N_4918,N_1903,N_509);
nand U4919 (N_4919,N_556,N_773);
nand U4920 (N_4920,N_2417,N_664);
xnor U4921 (N_4921,N_820,N_2479);
xnor U4922 (N_4922,N_2022,N_983);
and U4923 (N_4923,N_907,N_609);
nor U4924 (N_4924,N_2313,N_641);
xnor U4925 (N_4925,N_1800,N_1909);
nand U4926 (N_4926,N_783,N_1746);
nor U4927 (N_4927,N_850,N_2328);
nand U4928 (N_4928,N_540,N_497);
or U4929 (N_4929,N_1615,N_1203);
nand U4930 (N_4930,N_749,N_1433);
and U4931 (N_4931,N_2040,N_1181);
or U4932 (N_4932,N_2313,N_539);
nand U4933 (N_4933,N_552,N_1336);
and U4934 (N_4934,N_1702,N_2462);
and U4935 (N_4935,N_1837,N_2002);
or U4936 (N_4936,N_2101,N_1053);
or U4937 (N_4937,N_2380,N_983);
nor U4938 (N_4938,N_913,N_1781);
xnor U4939 (N_4939,N_876,N_301);
and U4940 (N_4940,N_735,N_1546);
nand U4941 (N_4941,N_2303,N_424);
and U4942 (N_4942,N_1097,N_1584);
nor U4943 (N_4943,N_1580,N_1010);
nand U4944 (N_4944,N_1299,N_1238);
nand U4945 (N_4945,N_485,N_2152);
nor U4946 (N_4946,N_1857,N_909);
and U4947 (N_4947,N_896,N_1030);
or U4948 (N_4948,N_2197,N_260);
nor U4949 (N_4949,N_2175,N_1381);
or U4950 (N_4950,N_1424,N_1092);
and U4951 (N_4951,N_1391,N_738);
nand U4952 (N_4952,N_2211,N_572);
and U4953 (N_4953,N_1789,N_618);
nand U4954 (N_4954,N_1903,N_299);
nand U4955 (N_4955,N_1952,N_2374);
or U4956 (N_4956,N_1112,N_1238);
xnor U4957 (N_4957,N_1003,N_1191);
nand U4958 (N_4958,N_1382,N_1034);
and U4959 (N_4959,N_639,N_314);
nor U4960 (N_4960,N_138,N_668);
xnor U4961 (N_4961,N_717,N_1512);
xnor U4962 (N_4962,N_532,N_1175);
nor U4963 (N_4963,N_723,N_920);
nand U4964 (N_4964,N_1600,N_259);
nand U4965 (N_4965,N_1208,N_1217);
and U4966 (N_4966,N_263,N_705);
or U4967 (N_4967,N_1710,N_1031);
xor U4968 (N_4968,N_1693,N_1965);
xor U4969 (N_4969,N_1348,N_1681);
xor U4970 (N_4970,N_1446,N_414);
xor U4971 (N_4971,N_310,N_435);
nor U4972 (N_4972,N_278,N_1993);
nand U4973 (N_4973,N_379,N_650);
nor U4974 (N_4974,N_2303,N_1188);
and U4975 (N_4975,N_1580,N_446);
and U4976 (N_4976,N_1936,N_2466);
xnor U4977 (N_4977,N_289,N_399);
xor U4978 (N_4978,N_848,N_1576);
nand U4979 (N_4979,N_235,N_2050);
nand U4980 (N_4980,N_2130,N_1427);
and U4981 (N_4981,N_1819,N_1425);
or U4982 (N_4982,N_1300,N_1742);
nand U4983 (N_4983,N_1321,N_739);
nand U4984 (N_4984,N_1235,N_1554);
nor U4985 (N_4985,N_328,N_1726);
or U4986 (N_4986,N_289,N_927);
or U4987 (N_4987,N_717,N_392);
xor U4988 (N_4988,N_1811,N_857);
xnor U4989 (N_4989,N_381,N_2327);
nor U4990 (N_4990,N_2496,N_1528);
or U4991 (N_4991,N_2371,N_258);
nor U4992 (N_4992,N_2345,N_1035);
and U4993 (N_4993,N_124,N_1317);
nor U4994 (N_4994,N_2044,N_1404);
nor U4995 (N_4995,N_160,N_1165);
and U4996 (N_4996,N_2274,N_1601);
and U4997 (N_4997,N_476,N_2082);
or U4998 (N_4998,N_1244,N_1939);
nor U4999 (N_4999,N_177,N_2294);
nor UO_0 (O_0,N_3075,N_4788);
or UO_1 (O_1,N_3606,N_4255);
nand UO_2 (O_2,N_4451,N_3714);
nand UO_3 (O_3,N_3574,N_4698);
xnor UO_4 (O_4,N_2523,N_4626);
nand UO_5 (O_5,N_3206,N_3937);
xnor UO_6 (O_6,N_4340,N_3820);
xnor UO_7 (O_7,N_2900,N_3215);
or UO_8 (O_8,N_3487,N_3744);
xor UO_9 (O_9,N_3725,N_4143);
xor UO_10 (O_10,N_3842,N_4251);
xor UO_11 (O_11,N_3561,N_4252);
nor UO_12 (O_12,N_4199,N_3021);
or UO_13 (O_13,N_4138,N_2667);
and UO_14 (O_14,N_2829,N_4690);
or UO_15 (O_15,N_3609,N_4605);
nor UO_16 (O_16,N_4769,N_4249);
nand UO_17 (O_17,N_2584,N_3961);
and UO_18 (O_18,N_2526,N_3197);
nand UO_19 (O_19,N_3862,N_3988);
nor UO_20 (O_20,N_4184,N_4342);
nor UO_21 (O_21,N_3575,N_3421);
nor UO_22 (O_22,N_4446,N_4073);
xnor UO_23 (O_23,N_3173,N_3560);
or UO_24 (O_24,N_4011,N_4445);
nand UO_25 (O_25,N_2565,N_4993);
nor UO_26 (O_26,N_3357,N_4645);
nor UO_27 (O_27,N_4860,N_3145);
or UO_28 (O_28,N_4204,N_3439);
nand UO_29 (O_29,N_3216,N_3517);
or UO_30 (O_30,N_3117,N_3464);
nor UO_31 (O_31,N_3412,N_2623);
xor UO_32 (O_32,N_4044,N_2692);
and UO_33 (O_33,N_3044,N_3001);
nand UO_34 (O_34,N_2820,N_4966);
nand UO_35 (O_35,N_3223,N_3522);
nand UO_36 (O_36,N_4875,N_2703);
nand UO_37 (O_37,N_2574,N_3070);
nor UO_38 (O_38,N_3892,N_2772);
xor UO_39 (O_39,N_4236,N_4990);
xnor UO_40 (O_40,N_4114,N_3022);
nand UO_41 (O_41,N_4090,N_4594);
or UO_42 (O_42,N_4646,N_4331);
xnor UO_43 (O_43,N_3932,N_2676);
or UO_44 (O_44,N_4045,N_3824);
xnor UO_45 (O_45,N_3454,N_3297);
and UO_46 (O_46,N_3653,N_3495);
or UO_47 (O_47,N_4816,N_3855);
or UO_48 (O_48,N_3181,N_4317);
xnor UO_49 (O_49,N_2952,N_4714);
nand UO_50 (O_50,N_4740,N_4739);
or UO_51 (O_51,N_4152,N_3761);
or UO_52 (O_52,N_2789,N_4492);
nand UO_53 (O_53,N_4001,N_3423);
nor UO_54 (O_54,N_2970,N_3898);
or UO_55 (O_55,N_4093,N_3141);
and UO_56 (O_56,N_4444,N_4115);
nor UO_57 (O_57,N_4868,N_3968);
or UO_58 (O_58,N_4402,N_3016);
and UO_59 (O_59,N_2766,N_3447);
xor UO_60 (O_60,N_3983,N_3453);
or UO_61 (O_61,N_3243,N_4633);
nand UO_62 (O_62,N_3912,N_4725);
nor UO_63 (O_63,N_2817,N_2519);
nor UO_64 (O_64,N_4949,N_4774);
xnor UO_65 (O_65,N_4453,N_3493);
nand UO_66 (O_66,N_3072,N_4231);
nand UO_67 (O_67,N_4787,N_3036);
nand UO_68 (O_68,N_4829,N_4542);
nor UO_69 (O_69,N_3459,N_2979);
xor UO_70 (O_70,N_4107,N_3797);
or UO_71 (O_71,N_2943,N_2804);
and UO_72 (O_72,N_3269,N_4103);
nor UO_73 (O_73,N_4910,N_4510);
xor UO_74 (O_74,N_4549,N_4395);
or UO_75 (O_75,N_4535,N_3395);
nor UO_76 (O_76,N_2514,N_3446);
nand UO_77 (O_77,N_3033,N_4610);
nor UO_78 (O_78,N_4474,N_4709);
and UO_79 (O_79,N_4847,N_3093);
or UO_80 (O_80,N_3681,N_3712);
nor UO_81 (O_81,N_3994,N_3853);
or UO_82 (O_82,N_4345,N_4560);
nand UO_83 (O_83,N_3596,N_4675);
nor UO_84 (O_84,N_3953,N_3232);
and UO_85 (O_85,N_2516,N_2744);
and UO_86 (O_86,N_4614,N_4408);
or UO_87 (O_87,N_4593,N_4040);
xor UO_88 (O_88,N_4768,N_4659);
nand UO_89 (O_89,N_4384,N_2544);
nor UO_90 (O_90,N_4872,N_2524);
nand UO_91 (O_91,N_3276,N_4590);
or UO_92 (O_92,N_3875,N_3006);
nand UO_93 (O_93,N_3941,N_3967);
and UO_94 (O_94,N_4671,N_4952);
or UO_95 (O_95,N_3474,N_3477);
xnor UO_96 (O_96,N_3335,N_4425);
and UO_97 (O_97,N_3844,N_3390);
xor UO_98 (O_98,N_4578,N_2760);
nor UO_99 (O_99,N_3231,N_3150);
xor UO_100 (O_100,N_2893,N_4338);
and UO_101 (O_101,N_4664,N_2951);
and UO_102 (O_102,N_3905,N_4328);
nand UO_103 (O_103,N_4796,N_2803);
nor UO_104 (O_104,N_2662,N_3951);
or UO_105 (O_105,N_3865,N_4435);
nor UO_106 (O_106,N_3724,N_2721);
nand UO_107 (O_107,N_4630,N_3624);
and UO_108 (O_108,N_4381,N_4814);
and UO_109 (O_109,N_3255,N_3848);
nor UO_110 (O_110,N_4760,N_2773);
and UO_111 (O_111,N_2700,N_4106);
xor UO_112 (O_112,N_2694,N_3656);
and UO_113 (O_113,N_4117,N_2749);
and UO_114 (O_114,N_2794,N_4971);
nor UO_115 (O_115,N_4771,N_3564);
nor UO_116 (O_116,N_4520,N_3299);
xor UO_117 (O_117,N_4521,N_3312);
and UO_118 (O_118,N_3202,N_4853);
and UO_119 (O_119,N_4612,N_2786);
nor UO_120 (O_120,N_4185,N_3555);
and UO_121 (O_121,N_3236,N_4906);
xor UO_122 (O_122,N_3726,N_4758);
nor UO_123 (O_123,N_4780,N_4817);
nor UO_124 (O_124,N_2816,N_3540);
xnor UO_125 (O_125,N_4992,N_4364);
xor UO_126 (O_126,N_3113,N_3414);
nor UO_127 (O_127,N_3040,N_3282);
xnor UO_128 (O_128,N_4471,N_4122);
nand UO_129 (O_129,N_4812,N_3644);
and UO_130 (O_130,N_4757,N_3880);
nor UO_131 (O_131,N_4259,N_4449);
nor UO_132 (O_132,N_4438,N_3711);
and UO_133 (O_133,N_4233,N_4287);
or UO_134 (O_134,N_3514,N_3370);
or UO_135 (O_135,N_2799,N_2857);
nand UO_136 (O_136,N_3752,N_3211);
nand UO_137 (O_137,N_3557,N_3305);
nand UO_138 (O_138,N_3743,N_4443);
nor UO_139 (O_139,N_3501,N_3252);
and UO_140 (O_140,N_4433,N_4583);
and UO_141 (O_141,N_3497,N_3319);
nor UO_142 (O_142,N_2784,N_4892);
and UO_143 (O_143,N_2964,N_4657);
or UO_144 (O_144,N_3998,N_4466);
nand UO_145 (O_145,N_3971,N_3729);
nand UO_146 (O_146,N_3738,N_3472);
nand UO_147 (O_147,N_3207,N_4689);
or UO_148 (O_148,N_2652,N_3697);
xor UO_149 (O_149,N_3693,N_3654);
xnor UO_150 (O_150,N_4918,N_2935);
and UO_151 (O_151,N_3627,N_3253);
xor UO_152 (O_152,N_2678,N_4953);
xnor UO_153 (O_153,N_4129,N_4455);
xor UO_154 (O_154,N_2824,N_4546);
nor UO_155 (O_155,N_4468,N_4691);
or UO_156 (O_156,N_4300,N_3595);
or UO_157 (O_157,N_2896,N_2758);
and UO_158 (O_158,N_3879,N_3131);
nor UO_159 (O_159,N_4382,N_4726);
nor UO_160 (O_160,N_4065,N_4619);
or UO_161 (O_161,N_3935,N_4254);
nand UO_162 (O_162,N_2539,N_3676);
or UO_163 (O_163,N_4522,N_2780);
nand UO_164 (O_164,N_4724,N_3339);
nor UO_165 (O_165,N_3062,N_2973);
nand UO_166 (O_166,N_3023,N_3334);
or UO_167 (O_167,N_3315,N_4037);
or UO_168 (O_168,N_4149,N_3435);
and UO_169 (O_169,N_4688,N_4750);
nand UO_170 (O_170,N_2620,N_3102);
xnor UO_171 (O_171,N_3132,N_4431);
and UO_172 (O_172,N_4810,N_4119);
nor UO_173 (O_173,N_4801,N_4068);
or UO_174 (O_174,N_4261,N_3838);
xor UO_175 (O_175,N_4987,N_4576);
or UO_176 (O_176,N_4540,N_3521);
nand UO_177 (O_177,N_2836,N_3224);
or UO_178 (O_178,N_3764,N_2564);
nand UO_179 (O_179,N_4208,N_2895);
xnor UO_180 (O_180,N_3283,N_3810);
xor UO_181 (O_181,N_3632,N_3544);
and UO_182 (O_182,N_4034,N_2507);
or UO_183 (O_183,N_3385,N_4859);
and UO_184 (O_184,N_3746,N_4609);
xnor UO_185 (O_185,N_4125,N_4092);
nor UO_186 (O_186,N_4809,N_4452);
and UO_187 (O_187,N_4672,N_3767);
and UO_188 (O_188,N_3826,N_4416);
xor UO_189 (O_189,N_4245,N_3946);
nand UO_190 (O_190,N_4584,N_3220);
and UO_191 (O_191,N_4955,N_4228);
or UO_192 (O_192,N_2959,N_2569);
and UO_193 (O_193,N_3986,N_4643);
and UO_194 (O_194,N_2971,N_3333);
xnor UO_195 (O_195,N_4469,N_4807);
xnor UO_196 (O_196,N_3415,N_4215);
and UO_197 (O_197,N_4891,N_4734);
nand UO_198 (O_198,N_3913,N_3230);
nor UO_199 (O_199,N_3786,N_2510);
nand UO_200 (O_200,N_2728,N_4286);
nand UO_201 (O_201,N_2580,N_4298);
and UO_202 (O_202,N_4173,N_4465);
or UO_203 (O_203,N_4116,N_4080);
and UO_204 (O_204,N_2955,N_2697);
nand UO_205 (O_205,N_3164,N_3389);
nor UO_206 (O_206,N_4505,N_4694);
or UO_207 (O_207,N_2977,N_3944);
and UO_208 (O_208,N_3804,N_4457);
nand UO_209 (O_209,N_4196,N_2621);
nand UO_210 (O_210,N_3188,N_2683);
or UO_211 (O_211,N_2878,N_4927);
or UO_212 (O_212,N_4289,N_3558);
or UO_213 (O_213,N_2792,N_3985);
nand UO_214 (O_214,N_3060,N_4862);
and UO_215 (O_215,N_3802,N_4487);
and UO_216 (O_216,N_4700,N_4258);
nand UO_217 (O_217,N_3134,N_4961);
nor UO_218 (O_218,N_3193,N_2534);
nand UO_219 (O_219,N_3448,N_4648);
xor UO_220 (O_220,N_4494,N_3925);
nor UO_221 (O_221,N_2762,N_2778);
or UO_222 (O_222,N_3248,N_4800);
nor UO_223 (O_223,N_4618,N_3148);
or UO_224 (O_224,N_3272,N_4797);
and UO_225 (O_225,N_4368,N_3121);
xnor UO_226 (O_226,N_2592,N_4180);
xnor UO_227 (O_227,N_2619,N_2546);
or UO_228 (O_228,N_4840,N_3929);
xor UO_229 (O_229,N_2549,N_3887);
nor UO_230 (O_230,N_3634,N_4450);
nand UO_231 (O_231,N_4363,N_4415);
and UO_232 (O_232,N_3700,N_4615);
and UO_233 (O_233,N_4305,N_4101);
and UO_234 (O_234,N_4386,N_3041);
and UO_235 (O_235,N_4625,N_2587);
and UO_236 (O_236,N_4747,N_4385);
xor UO_237 (O_237,N_2897,N_4137);
nand UO_238 (O_238,N_4569,N_3024);
or UO_239 (O_239,N_2688,N_4403);
nand UO_240 (O_240,N_3531,N_4670);
xor UO_241 (O_241,N_3200,N_3535);
xor UO_242 (O_242,N_4226,N_3155);
nand UO_243 (O_243,N_3168,N_4970);
nand UO_244 (O_244,N_2894,N_3111);
or UO_245 (O_245,N_2888,N_4727);
or UO_246 (O_246,N_3837,N_4655);
nor UO_247 (O_247,N_4572,N_3313);
and UO_248 (O_248,N_3884,N_3516);
nor UO_249 (O_249,N_3287,N_4097);
nand UO_250 (O_250,N_4607,N_4956);
nor UO_251 (O_251,N_3427,N_3227);
nor UO_252 (O_252,N_2990,N_3602);
nor UO_253 (O_253,N_2764,N_2869);
and UO_254 (O_254,N_2718,N_2814);
xor UO_255 (O_255,N_3359,N_3499);
and UO_256 (O_256,N_4805,N_4361);
or UO_257 (O_257,N_3717,N_3590);
and UO_258 (O_258,N_3130,N_3162);
and UO_259 (O_259,N_3769,N_2846);
and UO_260 (O_260,N_2547,N_4429);
nand UO_261 (O_261,N_2598,N_2594);
xnor UO_262 (O_262,N_4530,N_2616);
nand UO_263 (O_263,N_4472,N_3601);
nand UO_264 (O_264,N_4157,N_3568);
or UO_265 (O_265,N_4644,N_4491);
or UO_266 (O_266,N_3151,N_4876);
xor UO_267 (O_267,N_3103,N_3662);
nand UO_268 (O_268,N_2914,N_4055);
nor UO_269 (O_269,N_4335,N_4321);
nand UO_270 (O_270,N_2679,N_4477);
or UO_271 (O_271,N_4874,N_2756);
nand UO_272 (O_272,N_4753,N_3303);
or UO_273 (O_273,N_2681,N_3950);
nand UO_274 (O_274,N_4209,N_2622);
nand UO_275 (O_275,N_4454,N_4111);
xnor UO_276 (O_276,N_3629,N_3807);
xor UO_277 (O_277,N_2719,N_3734);
and UO_278 (O_278,N_4815,N_4203);
nor UO_279 (O_279,N_4667,N_4509);
xor UO_280 (O_280,N_4878,N_4102);
nand UO_281 (O_281,N_3233,N_4207);
nand UO_282 (O_282,N_4350,N_4846);
and UO_283 (O_283,N_4634,N_4580);
nor UO_284 (O_284,N_3736,N_3663);
and UO_285 (O_285,N_4064,N_4166);
xnor UO_286 (O_286,N_4686,N_4851);
or UO_287 (O_287,N_3413,N_3776);
nand UO_288 (O_288,N_3751,N_4617);
nor UO_289 (O_289,N_2635,N_4084);
or UO_290 (O_290,N_3133,N_3543);
xor UO_291 (O_291,N_4311,N_4399);
xnor UO_292 (O_292,N_4366,N_4436);
or UO_293 (O_293,N_4271,N_4665);
nand UO_294 (O_294,N_3294,N_3592);
xor UO_295 (O_295,N_4030,N_4274);
or UO_296 (O_296,N_4272,N_3684);
xnor UO_297 (O_297,N_2506,N_4857);
nor UO_298 (O_298,N_4718,N_4723);
and UO_299 (O_299,N_3019,N_2847);
nor UO_300 (O_300,N_4935,N_3980);
xnor UO_301 (O_301,N_3043,N_3559);
xnor UO_302 (O_302,N_3818,N_3649);
xor UO_303 (O_303,N_4419,N_3660);
and UO_304 (O_304,N_3931,N_4072);
and UO_305 (O_305,N_3638,N_3537);
xor UO_306 (O_306,N_2796,N_4417);
and UO_307 (O_307,N_3302,N_2709);
and UO_308 (O_308,N_4219,N_4778);
xnor UO_309 (O_309,N_3722,N_4934);
nor UO_310 (O_310,N_4375,N_4925);
xnor UO_311 (O_311,N_2558,N_3452);
nand UO_312 (O_312,N_3934,N_3977);
xor UO_313 (O_313,N_3301,N_2873);
nor UO_314 (O_314,N_2832,N_4748);
nor UO_315 (O_315,N_4039,N_3280);
or UO_316 (O_316,N_4291,N_3954);
nor UO_317 (O_317,N_3106,N_2736);
or UO_318 (O_318,N_2603,N_3507);
xnor UO_319 (O_319,N_4803,N_3431);
nor UO_320 (O_320,N_3571,N_4060);
nor UO_321 (O_321,N_3254,N_3035);
nand UO_322 (O_322,N_4848,N_3127);
and UO_323 (O_323,N_2752,N_2704);
xor UO_324 (O_324,N_4029,N_4647);
or UO_325 (O_325,N_2757,N_4901);
nand UO_326 (O_326,N_4460,N_3694);
nand UO_327 (O_327,N_3871,N_4292);
or UO_328 (O_328,N_4432,N_4380);
nor UO_329 (O_329,N_3456,N_3484);
xnor UO_330 (O_330,N_4257,N_4200);
nand UO_331 (O_331,N_3351,N_4722);
or UO_332 (O_332,N_3311,N_3896);
nor UO_333 (O_333,N_2909,N_4058);
nand UO_334 (O_334,N_4567,N_4599);
nand UO_335 (O_335,N_2653,N_3204);
and UO_336 (O_336,N_3608,N_3066);
nor UO_337 (O_337,N_4652,N_3483);
nand UO_338 (O_338,N_2663,N_3161);
nand UO_339 (O_339,N_2673,N_2930);
nand UO_340 (O_340,N_3042,N_3976);
xor UO_341 (O_341,N_3088,N_3870);
or UO_342 (O_342,N_4178,N_4110);
nor UO_343 (O_343,N_4879,N_3402);
xor UO_344 (O_344,N_4418,N_2822);
nor UO_345 (O_345,N_2657,N_4049);
nor UO_346 (O_346,N_4754,N_3081);
xnor UO_347 (O_347,N_3646,N_4944);
or UO_348 (O_348,N_2919,N_3829);
xnor UO_349 (O_349,N_3083,N_3281);
and UO_350 (O_350,N_2726,N_2785);
nand UO_351 (O_351,N_4159,N_3182);
nor UO_352 (O_352,N_3471,N_4370);
nor UO_353 (O_353,N_4025,N_3636);
nand UO_354 (O_354,N_3674,N_3605);
nand UO_355 (O_355,N_4931,N_2889);
nand UO_356 (O_356,N_2642,N_3398);
or UO_357 (O_357,N_3065,N_3631);
xnor UO_358 (O_358,N_3271,N_3296);
xor UO_359 (O_359,N_2972,N_4921);
and UO_360 (O_360,N_3610,N_3554);
nand UO_361 (O_361,N_3475,N_3523);
nor UO_362 (O_362,N_3773,N_4631);
nand UO_363 (O_363,N_4692,N_4928);
xor UO_364 (O_364,N_2597,N_4010);
xnor UO_365 (O_365,N_4140,N_3519);
nand UO_366 (O_366,N_2761,N_2633);
xnor UO_367 (O_367,N_3965,N_4193);
or UO_368 (O_368,N_3856,N_4556);
and UO_369 (O_369,N_4824,N_3054);
nand UO_370 (O_370,N_4083,N_3715);
or UO_371 (O_371,N_3777,N_2969);
xnor UO_372 (O_372,N_3110,N_2831);
nand UO_373 (O_373,N_3910,N_2685);
or UO_374 (O_374,N_2614,N_2800);
xor UO_375 (O_375,N_4705,N_4728);
and UO_376 (O_376,N_3430,N_3857);
and UO_377 (O_377,N_2573,N_2818);
nand UO_378 (O_378,N_3118,N_4820);
and UO_379 (O_379,N_4483,N_3026);
xor UO_380 (O_380,N_4248,N_4206);
and UO_381 (O_381,N_2963,N_3418);
nor UO_382 (O_382,N_3583,N_3970);
and UO_383 (O_383,N_4427,N_4070);
or UO_384 (O_384,N_3494,N_2730);
nor UO_385 (O_385,N_4337,N_4962);
nor UO_386 (O_386,N_4608,N_4917);
and UO_387 (O_387,N_2566,N_3048);
or UO_388 (O_388,N_2948,N_3208);
nand UO_389 (O_389,N_3160,N_4877);
nand UO_390 (O_390,N_4371,N_3146);
or UO_391 (O_391,N_4676,N_4770);
and UO_392 (O_392,N_4174,N_4085);
nor UO_393 (O_393,N_3092,N_4972);
nand UO_394 (O_394,N_2981,N_3174);
xor UO_395 (O_395,N_3341,N_4864);
xor UO_396 (O_396,N_2947,N_3222);
nor UO_397 (O_397,N_4920,N_3432);
nand UO_398 (O_398,N_4202,N_4679);
xor UO_399 (O_399,N_3455,N_4653);
xnor UO_400 (O_400,N_2689,N_4589);
or UO_401 (O_401,N_3262,N_2654);
and UO_402 (O_402,N_3831,N_2841);
nand UO_403 (O_403,N_2520,N_4464);
and UO_404 (O_404,N_3920,N_2611);
nand UO_405 (O_405,N_4210,N_3539);
nor UO_406 (O_406,N_2682,N_3598);
nand UO_407 (O_407,N_3013,N_3635);
and UO_408 (O_408,N_3765,N_3030);
or UO_409 (O_409,N_2581,N_3264);
or UO_410 (O_410,N_3235,N_4393);
and UO_411 (O_411,N_2837,N_2779);
nor UO_412 (O_412,N_2880,N_4963);
and UO_413 (O_413,N_4318,N_2849);
and UO_414 (O_414,N_4006,N_4514);
or UO_415 (O_415,N_3307,N_4982);
nand UO_416 (O_416,N_4825,N_4332);
or UO_417 (O_417,N_4169,N_4516);
nor UO_418 (O_418,N_2590,N_3260);
or UO_419 (O_419,N_3485,N_3138);
nand UO_420 (O_420,N_4792,N_3467);
nand UO_421 (O_421,N_3668,N_3076);
and UO_422 (O_422,N_4673,N_3273);
and UO_423 (O_423,N_3794,N_3811);
nor UO_424 (O_424,N_3960,N_4168);
xor UO_425 (O_425,N_4260,N_3234);
and UO_426 (O_426,N_2739,N_2797);
nor UO_427 (O_427,N_2727,N_3000);
xnor UO_428 (O_428,N_2567,N_4685);
nand UO_429 (O_429,N_4124,N_4881);
nor UO_430 (O_430,N_3336,N_4738);
xor UO_431 (O_431,N_3330,N_4497);
and UO_432 (O_432,N_2670,N_4627);
and UO_433 (O_433,N_4564,N_4818);
xnor UO_434 (O_434,N_3721,N_3100);
and UO_435 (O_435,N_2552,N_2529);
or UO_436 (O_436,N_2957,N_4089);
or UO_437 (O_437,N_3259,N_3520);
nand UO_438 (O_438,N_4232,N_2860);
or UO_439 (O_439,N_3194,N_3274);
xor UO_440 (O_440,N_3828,N_3108);
xor UO_441 (O_441,N_4496,N_3250);
or UO_442 (O_442,N_4978,N_2562);
or UO_443 (O_443,N_4784,N_4005);
xor UO_444 (O_444,N_3545,N_2596);
nand UO_445 (O_445,N_3144,N_3219);
or UO_446 (O_446,N_4945,N_3442);
nor UO_447 (O_447,N_3067,N_4057);
nor UO_448 (O_448,N_3177,N_2706);
or UO_449 (O_449,N_4563,N_4896);
nor UO_450 (O_450,N_4933,N_3257);
nor UO_451 (O_451,N_4442,N_4802);
nor UO_452 (O_452,N_2807,N_3926);
xor UO_453 (O_453,N_2759,N_3153);
or UO_454 (O_454,N_3665,N_4941);
xnor UO_455 (O_455,N_4264,N_2821);
nor UO_456 (O_456,N_3614,N_3321);
or UO_457 (O_457,N_3628,N_3462);
xnor UO_458 (O_458,N_4682,N_4900);
and UO_459 (O_459,N_4638,N_3101);
nand UO_460 (O_460,N_3068,N_2533);
or UO_461 (O_461,N_2863,N_4181);
and UO_462 (O_462,N_3969,N_3286);
xnor UO_463 (O_463,N_3139,N_4146);
nor UO_464 (O_464,N_3845,N_4782);
or UO_465 (O_465,N_3476,N_2643);
and UO_466 (O_466,N_2665,N_3217);
and UO_467 (O_467,N_4324,N_3504);
or UO_468 (O_468,N_4369,N_4737);
xnor UO_469 (O_469,N_4234,N_2638);
or UO_470 (O_470,N_2608,N_4789);
xor UO_471 (O_471,N_2532,N_3686);
nor UO_472 (O_472,N_4479,N_3409);
and UO_473 (O_473,N_4275,N_3914);
and UO_474 (O_474,N_3899,N_4639);
nand UO_475 (O_475,N_3817,N_3513);
or UO_476 (O_476,N_3778,N_2782);
or UO_477 (O_477,N_4214,N_4358);
and UO_478 (O_478,N_3534,N_4536);
xnor UO_479 (O_479,N_4973,N_3733);
xor UO_480 (O_480,N_2815,N_3186);
and UO_481 (O_481,N_4319,N_2656);
or UO_482 (O_482,N_4155,N_4046);
or UO_483 (O_483,N_4575,N_4091);
xnor UO_484 (O_484,N_4574,N_3866);
and UO_485 (O_485,N_2712,N_2672);
nand UO_486 (O_486,N_3801,N_3371);
nor UO_487 (O_487,N_4280,N_4515);
nand UO_488 (O_488,N_3849,N_4136);
nand UO_489 (O_489,N_3099,N_3261);
nand UO_490 (O_490,N_3340,N_3683);
xnor UO_491 (O_491,N_3049,N_3071);
nand UO_492 (O_492,N_4392,N_2879);
xnor UO_493 (O_493,N_3393,N_2984);
or UO_494 (O_494,N_3372,N_3548);
and UO_495 (O_495,N_2504,N_2699);
nor UO_496 (O_496,N_4602,N_3238);
nor UO_497 (O_497,N_4462,N_3361);
nor UO_498 (O_498,N_2858,N_2588);
and UO_499 (O_499,N_3401,N_2639);
xor UO_500 (O_500,N_2572,N_2791);
and UO_501 (O_501,N_4282,N_2626);
xnor UO_502 (O_502,N_4861,N_4975);
or UO_503 (O_503,N_3529,N_3938);
nand UO_504 (O_504,N_4870,N_4511);
and UO_505 (O_505,N_3057,N_4858);
nand UO_506 (O_506,N_4325,N_3184);
nor UO_507 (O_507,N_4669,N_4745);
and UO_508 (O_508,N_2917,N_3648);
nor UO_509 (O_509,N_4704,N_4054);
or UO_510 (O_510,N_4668,N_4243);
nand UO_511 (O_511,N_2578,N_4710);
nor UO_512 (O_512,N_3643,N_3196);
xnor UO_513 (O_513,N_4528,N_3840);
or UO_514 (O_514,N_2659,N_3858);
nand UO_515 (O_515,N_2605,N_4606);
or UO_516 (O_516,N_2735,N_4314);
or UO_517 (O_517,N_3527,N_2945);
xnor UO_518 (O_518,N_3061,N_4702);
xor UO_519 (O_519,N_4316,N_4736);
nor UO_520 (O_520,N_4297,N_2925);
or UO_521 (O_521,N_4804,N_2913);
nand UO_522 (O_522,N_4327,N_3928);
nor UO_523 (O_523,N_4843,N_4360);
nor UO_524 (O_524,N_3874,N_4067);
nand UO_525 (O_525,N_3830,N_4811);
xor UO_526 (O_526,N_4059,N_3748);
nand UO_527 (O_527,N_3891,N_4222);
or UO_528 (O_528,N_2859,N_4827);
or UO_529 (O_529,N_4288,N_2810);
nand UO_530 (O_530,N_3422,N_4842);
xor UO_531 (O_531,N_4148,N_3839);
nand UO_532 (O_532,N_4886,N_3058);
or UO_533 (O_533,N_3268,N_3482);
or UO_534 (O_534,N_4926,N_2805);
or UO_535 (O_535,N_4167,N_3291);
or UO_536 (O_536,N_4499,N_2850);
nand UO_537 (O_537,N_3256,N_4751);
or UO_538 (O_538,N_3416,N_3466);
or UO_539 (O_539,N_4600,N_3380);
and UO_540 (O_540,N_4629,N_3353);
and UO_541 (O_541,N_3984,N_4562);
nand UO_542 (O_542,N_4018,N_4586);
xor UO_543 (O_543,N_4703,N_3356);
xor UO_544 (O_544,N_3433,N_4041);
and UO_545 (O_545,N_3642,N_2733);
and UO_546 (O_546,N_4731,N_3673);
nor UO_547 (O_547,N_4439,N_4063);
nand UO_548 (O_548,N_3753,N_3933);
or UO_549 (O_549,N_3974,N_2905);
xor UO_550 (O_550,N_3591,N_3179);
and UO_551 (O_551,N_4687,N_2753);
xor UO_552 (O_552,N_3798,N_2691);
nand UO_553 (O_553,N_4795,N_2751);
and UO_554 (O_554,N_3854,N_4490);
or UO_555 (O_555,N_3549,N_3097);
nor UO_556 (O_556,N_2891,N_4969);
and UO_557 (O_557,N_3275,N_3708);
or UO_558 (O_558,N_3212,N_4635);
or UO_559 (O_559,N_4377,N_4262);
nand UO_560 (O_560,N_3792,N_3713);
nor UO_561 (O_561,N_4929,N_4441);
nor UO_562 (O_562,N_3157,N_4762);
and UO_563 (O_563,N_4729,N_2874);
or UO_564 (O_564,N_4047,N_2649);
nand UO_565 (O_565,N_3667,N_3739);
nor UO_566 (O_566,N_3623,N_2513);
xor UO_567 (O_567,N_2828,N_3515);
nand UO_568 (O_568,N_3137,N_2934);
nor UO_569 (O_569,N_3705,N_4850);
or UO_570 (O_570,N_4218,N_4043);
nand UO_571 (O_571,N_4430,N_4538);
and UO_572 (O_572,N_2845,N_4595);
nand UO_573 (O_573,N_2711,N_3465);
xor UO_574 (O_574,N_4518,N_3428);
nand UO_575 (O_575,N_3658,N_4551);
nand UO_576 (O_576,N_3890,N_3285);
nor UO_577 (O_577,N_3688,N_4032);
nor UO_578 (O_578,N_4713,N_2798);
or UO_579 (O_579,N_3142,N_4960);
or UO_580 (O_580,N_4151,N_4502);
nand UO_581 (O_581,N_4683,N_3009);
and UO_582 (O_582,N_3695,N_3813);
or UO_583 (O_583,N_3868,N_4017);
xnor UO_584 (O_584,N_4002,N_2903);
and UO_585 (O_585,N_3553,N_4663);
or UO_586 (O_586,N_2515,N_3822);
or UO_587 (O_587,N_3199,N_3295);
xor UO_588 (O_588,N_3135,N_2577);
xnor UO_589 (O_589,N_4374,N_3239);
or UO_590 (O_590,N_4882,N_3124);
and UO_591 (O_591,N_3298,N_4706);
and UO_592 (O_592,N_3784,N_3109);
xor UO_593 (O_593,N_4553,N_4897);
and UO_594 (O_594,N_3923,N_3795);
nor UO_595 (O_595,N_3463,N_2992);
xnor UO_596 (O_596,N_3940,N_4008);
or UO_597 (O_597,N_3791,N_4622);
xnor UO_598 (O_598,N_4699,N_3265);
and UO_599 (O_599,N_3429,N_2615);
nand UO_600 (O_600,N_2553,N_3038);
nand UO_601 (O_601,N_3749,N_2644);
nor UO_602 (O_602,N_3567,N_4440);
and UO_603 (O_603,N_4182,N_4221);
and UO_604 (O_604,N_4603,N_4164);
and UO_605 (O_605,N_4968,N_3706);
xor UO_606 (O_606,N_4779,N_3956);
xnor UO_607 (O_607,N_2531,N_3616);
nand UO_608 (O_608,N_3129,N_3763);
xor UO_609 (O_609,N_4720,N_2543);
and UO_610 (O_610,N_3012,N_3664);
nor UO_611 (O_611,N_3119,N_3737);
or UO_612 (O_612,N_3927,N_4397);
and UO_613 (O_613,N_3819,N_3716);
nor UO_614 (O_614,N_4937,N_3091);
xor UO_615 (O_615,N_2865,N_3834);
and UO_616 (O_616,N_2559,N_4570);
nand UO_617 (O_617,N_3641,N_3964);
nor UO_618 (O_618,N_3140,N_3185);
nor UO_619 (O_619,N_4190,N_3996);
and UO_620 (O_620,N_4623,N_2839);
nand UO_621 (O_621,N_3350,N_4118);
and UO_622 (O_622,N_4548,N_3279);
or UO_623 (O_623,N_2500,N_3888);
or UO_624 (O_624,N_4004,N_2996);
and UO_625 (O_625,N_2993,N_3966);
xor UO_626 (O_626,N_3637,N_4947);
and UO_627 (O_627,N_3190,N_4893);
nor UO_628 (O_628,N_3228,N_4696);
nor UO_629 (O_629,N_4566,N_3895);
and UO_630 (O_630,N_3440,N_2870);
or UO_631 (O_631,N_3930,N_3143);
and UO_632 (O_632,N_4458,N_2904);
nand UO_633 (O_633,N_4156,N_4224);
or UO_634 (O_634,N_4504,N_3374);
nand UO_635 (O_635,N_4565,N_2939);
nand UO_636 (O_636,N_3538,N_4398);
or UO_637 (O_637,N_4898,N_3704);
and UO_638 (O_638,N_4579,N_4326);
nor UO_639 (O_639,N_4105,N_4428);
or UO_640 (O_640,N_2687,N_4832);
nand UO_641 (O_641,N_4899,N_4349);
or UO_642 (O_642,N_4989,N_2617);
nor UO_643 (O_643,N_4033,N_4790);
nor UO_644 (O_644,N_2702,N_2582);
or UO_645 (O_645,N_2801,N_4640);
xor UO_646 (O_646,N_3187,N_3490);
or UO_647 (O_647,N_2901,N_2509);
nor UO_648 (O_648,N_3251,N_4031);
and UO_649 (O_649,N_4957,N_3392);
nand UO_650 (O_650,N_3774,N_2554);
xnor UO_651 (O_651,N_2548,N_4674);
or UO_652 (O_652,N_2740,N_3963);
nor UO_653 (O_653,N_4601,N_3354);
xnor UO_654 (O_654,N_4844,N_4170);
xor UO_655 (O_655,N_4744,N_2601);
xnor UO_656 (O_656,N_4558,N_2982);
and UO_657 (O_657,N_3909,N_3051);
nor UO_658 (O_658,N_3098,N_4229);
xnor UO_659 (O_659,N_3288,N_3921);
nand UO_660 (O_660,N_4940,N_2690);
xnor UO_661 (O_661,N_2787,N_3876);
xor UO_662 (O_662,N_4281,N_4604);
and UO_663 (O_663,N_4016,N_3126);
nand UO_664 (O_664,N_4096,N_4913);
and UO_665 (O_665,N_3346,N_2771);
nor UO_666 (O_666,N_3419,N_4488);
xnor UO_667 (O_667,N_4109,N_2852);
nand UO_668 (O_668,N_4480,N_4946);
and UO_669 (O_669,N_3572,N_4035);
nand UO_670 (O_670,N_3982,N_2628);
nor UO_671 (O_671,N_3159,N_3955);
nand UO_672 (O_672,N_2827,N_3017);
nor UO_673 (O_673,N_2695,N_3620);
or UO_674 (O_674,N_3018,N_4009);
nor UO_675 (O_675,N_2907,N_4422);
and UO_676 (O_676,N_3981,N_2540);
nor UO_677 (O_677,N_3344,N_3502);
and UO_678 (O_678,N_3011,N_3814);
nand UO_679 (O_679,N_2809,N_4711);
nand UO_680 (O_680,N_4680,N_4310);
nand UO_681 (O_681,N_3936,N_4112);
and UO_682 (O_682,N_4050,N_3293);
nand UO_683 (O_683,N_3210,N_4141);
and UO_684 (O_684,N_2501,N_3468);
and UO_685 (O_685,N_3503,N_4015);
and UO_686 (O_686,N_4077,N_2842);
and UO_687 (O_687,N_3029,N_4773);
and UO_688 (O_688,N_4086,N_3613);
nand UO_689 (O_689,N_3473,N_2707);
nor UO_690 (O_690,N_3821,N_3405);
and UO_691 (O_691,N_2851,N_3883);
and UO_692 (O_692,N_4819,N_2968);
xor UO_693 (O_693,N_4923,N_4995);
nor UO_694 (O_694,N_4552,N_4852);
nor UO_695 (O_695,N_4823,N_4007);
or UO_696 (O_696,N_4598,N_2974);
or UO_697 (O_697,N_2755,N_2898);
nor UO_698 (O_698,N_4786,N_3805);
and UO_699 (O_699,N_3787,N_3806);
nor UO_700 (O_700,N_3424,N_3457);
and UO_701 (O_701,N_4708,N_4075);
nor UO_702 (O_702,N_3165,N_3562);
and UO_703 (O_703,N_4561,N_4056);
or UO_704 (O_704,N_4493,N_4139);
or UO_705 (O_705,N_3850,N_2882);
nor UO_706 (O_706,N_2586,N_4977);
nor UO_707 (O_707,N_4543,N_4628);
or UO_708 (O_708,N_2502,N_3292);
nand UO_709 (O_709,N_4717,N_2825);
nor UO_710 (O_710,N_2966,N_4756);
nor UO_711 (O_711,N_4904,N_3323);
and UO_712 (O_712,N_2527,N_3176);
or UO_713 (O_713,N_2717,N_3317);
or UO_714 (O_714,N_2997,N_3582);
nand UO_715 (O_715,N_4133,N_4693);
nor UO_716 (O_716,N_4997,N_2908);
nand UO_717 (O_717,N_3833,N_2640);
and UO_718 (O_718,N_2868,N_3799);
nor UO_719 (O_719,N_2980,N_3218);
or UO_720 (O_720,N_4299,N_3979);
and UO_721 (O_721,N_3768,N_3566);
xor UO_722 (O_722,N_4295,N_3444);
nand UO_723 (O_723,N_3727,N_4434);
nand UO_724 (O_724,N_2871,N_4591);
xnor UO_725 (O_725,N_3163,N_4405);
xor UO_726 (O_726,N_3420,N_3718);
or UO_727 (O_727,N_4241,N_2867);
xor UO_728 (O_728,N_2579,N_3373);
and UO_729 (O_729,N_3358,N_4636);
nand UO_730 (O_730,N_4830,N_3263);
and UO_731 (O_731,N_3593,N_4186);
xor UO_732 (O_732,N_4592,N_4132);
xnor UO_733 (O_733,N_3078,N_3364);
nor UO_734 (O_734,N_4213,N_3191);
or UO_735 (O_735,N_3995,N_3436);
and UO_736 (O_736,N_2790,N_4263);
nand UO_737 (O_737,N_4347,N_4983);
or UO_738 (O_738,N_3785,N_4550);
or UO_739 (O_739,N_3491,N_2720);
xor UO_740 (O_740,N_4269,N_4423);
xnor UO_741 (O_741,N_4539,N_3766);
and UO_742 (O_742,N_3115,N_4735);
nor UO_743 (O_743,N_3355,N_3481);
or UO_744 (O_744,N_3363,N_4835);
and UO_745 (O_745,N_4354,N_3478);
and UO_746 (O_746,N_3028,N_3975);
and UO_747 (O_747,N_4759,N_3114);
nor UO_748 (O_748,N_3388,N_3122);
or UO_749 (O_749,N_3589,N_3325);
xnor UO_750 (O_750,N_3958,N_4367);
nand UO_751 (O_751,N_4942,N_3809);
nand UO_752 (O_752,N_3770,N_4279);
and UO_753 (O_753,N_4656,N_3679);
nand UO_754 (O_754,N_4994,N_4188);
or UO_755 (O_755,N_2632,N_4066);
or UO_756 (O_756,N_2668,N_2961);
nor UO_757 (O_757,N_3087,N_2606);
nor UO_758 (O_758,N_4894,N_4273);
and UO_759 (O_759,N_3803,N_4806);
xnor UO_760 (O_760,N_4359,N_3597);
xnor UO_761 (O_761,N_3972,N_4312);
and UO_762 (O_762,N_2899,N_4355);
and UO_763 (O_763,N_3916,N_4225);
and UO_764 (O_764,N_2834,N_4329);
xnor UO_765 (O_765,N_4456,N_4678);
xnor UO_766 (O_766,N_3586,N_3090);
or UO_767 (O_767,N_2994,N_4484);
xor UO_768 (O_768,N_2946,N_3897);
and UO_769 (O_769,N_2910,N_4179);
xnor UO_770 (O_770,N_2517,N_4763);
xnor UO_771 (O_771,N_3408,N_3835);
nand UO_772 (O_772,N_2811,N_4684);
xnor UO_773 (O_773,N_3506,N_3327);
nor UO_774 (O_774,N_3991,N_4743);
and UO_775 (O_775,N_3989,N_3707);
xor UO_776 (O_776,N_3594,N_2918);
nor UO_777 (O_777,N_3069,N_2557);
and UO_778 (O_778,N_3460,N_2560);
nand UO_779 (O_779,N_3245,N_3924);
nor UO_780 (O_780,N_2928,N_2571);
or UO_781 (O_781,N_2956,N_2844);
or UO_782 (O_782,N_4414,N_4379);
nand UO_783 (O_783,N_4421,N_2570);
nand UO_784 (O_784,N_2921,N_3214);
or UO_785 (O_785,N_3861,N_3320);
nor UO_786 (O_786,N_2677,N_3528);
nand UO_787 (O_787,N_4144,N_4936);
nor UO_788 (O_788,N_3630,N_4478);
nand UO_789 (O_789,N_2823,N_3488);
or UO_790 (O_790,N_2607,N_2535);
or UO_791 (O_791,N_2645,N_4476);
or UO_792 (O_792,N_3331,N_3911);
xor UO_793 (O_793,N_3692,N_2724);
or UO_794 (O_794,N_3815,N_3348);
or UO_795 (O_795,N_2604,N_3047);
xor UO_796 (O_796,N_4905,N_3689);
and UO_797 (O_797,N_2876,N_2583);
or UO_798 (O_798,N_4154,N_2561);
nor UO_799 (O_799,N_2987,N_3943);
or UO_800 (O_800,N_2862,N_2866);
xnor UO_801 (O_801,N_2833,N_4967);
and UO_802 (O_802,N_4544,N_4776);
xor UO_803 (O_803,N_3192,N_3085);
and UO_804 (O_804,N_4557,N_4062);
nor UO_805 (O_805,N_3394,N_4194);
and UO_806 (O_806,N_3270,N_3687);
nor UO_807 (O_807,N_2568,N_4895);
nor UO_808 (O_808,N_3580,N_4412);
or UO_809 (O_809,N_3867,N_3949);
and UO_810 (O_810,N_2658,N_4301);
nand UO_811 (O_811,N_3180,N_3149);
nand UO_812 (O_812,N_4176,N_4396);
and UO_813 (O_813,N_2734,N_3244);
xor UO_814 (O_814,N_4069,N_3780);
nor UO_815 (O_815,N_3709,N_2806);
nand UO_816 (O_816,N_3702,N_3640);
nor UO_817 (O_817,N_2556,N_4650);
and UO_818 (O_818,N_3378,N_4372);
or UO_819 (O_819,N_4526,N_3237);
nand UO_820 (O_820,N_3847,N_4306);
nand UO_821 (O_821,N_4315,N_4352);
or UO_822 (O_822,N_4869,N_3366);
and UO_823 (O_823,N_4485,N_3500);
nand UO_824 (O_824,N_4517,N_3247);
nand UO_825 (O_825,N_3079,N_2953);
nor UO_826 (O_826,N_4270,N_4265);
and UO_827 (O_827,N_3962,N_2793);
and UO_828 (O_828,N_4986,N_4741);
and UO_829 (O_829,N_2741,N_2813);
nand UO_830 (O_830,N_2634,N_3685);
or UO_831 (O_831,N_3750,N_4042);
and UO_832 (O_832,N_2714,N_4411);
and UO_833 (O_833,N_4277,N_4715);
or UO_834 (O_834,N_4903,N_3014);
nor UO_835 (O_835,N_4304,N_3306);
nand UO_836 (O_836,N_2788,N_3277);
and UO_837 (O_837,N_4681,N_3489);
nand UO_838 (O_838,N_3377,N_4914);
xor UO_839 (O_839,N_4268,N_3945);
nor UO_840 (O_840,N_2763,N_3783);
or UO_841 (O_841,N_3578,N_4353);
and UO_842 (O_842,N_2991,N_3703);
nand UO_843 (O_843,N_4390,N_4473);
nand UO_844 (O_844,N_3556,N_3198);
nor UO_845 (O_845,N_4712,N_2713);
xnor UO_846 (O_846,N_4613,N_3672);
or UO_847 (O_847,N_3304,N_3008);
xnor UO_848 (O_848,N_4013,N_2927);
and UO_849 (O_849,N_3904,N_2902);
and UO_850 (O_850,N_4524,N_4662);
nor UO_851 (O_851,N_2999,N_2912);
and UO_852 (O_852,N_4003,N_4021);
xnor UO_853 (O_853,N_2525,N_4401);
or UO_854 (O_854,N_3386,N_3397);
nand UO_855 (O_855,N_2536,N_4732);
nor UO_856 (O_856,N_3221,N_2765);
nand UO_857 (O_857,N_3915,N_3579);
or UO_858 (O_858,N_3360,N_3877);
or UO_859 (O_859,N_3367,N_3015);
or UO_860 (O_860,N_4250,N_3379);
nor UO_861 (O_861,N_4908,N_4641);
or UO_862 (O_862,N_2542,N_2660);
and UO_863 (O_863,N_4822,N_2732);
nor UO_864 (O_864,N_4746,N_4223);
nand UO_865 (O_865,N_4285,N_4996);
and UO_866 (O_866,N_3169,N_3639);
nand UO_867 (O_867,N_3205,N_3178);
xor UO_868 (O_868,N_4527,N_2669);
and UO_869 (O_869,N_3469,N_4362);
nor UO_870 (O_870,N_2637,N_4854);
nand UO_871 (O_871,N_3587,N_4012);
and UO_872 (O_872,N_4799,N_4242);
xor UO_873 (O_873,N_4742,N_3872);
nand UO_874 (O_874,N_2965,N_4357);
and UO_875 (O_875,N_3757,N_2674);
xnor UO_876 (O_876,N_4525,N_3524);
nor UO_877 (O_877,N_3939,N_4120);
or UO_878 (O_878,N_3010,N_3326);
nor UO_879 (O_879,N_4642,N_2743);
and UO_880 (O_880,N_3992,N_3059);
nand UO_881 (O_881,N_2768,N_3762);
xor UO_882 (O_882,N_4883,N_4849);
or UO_883 (O_883,N_3678,N_4088);
or UO_884 (O_884,N_4695,N_2655);
nor UO_885 (O_885,N_3903,N_2975);
or UO_886 (O_886,N_2593,N_3690);
xor UO_887 (O_887,N_2664,N_3050);
nor UO_888 (O_888,N_2819,N_4577);
nand UO_889 (O_889,N_2872,N_2708);
or UO_890 (O_890,N_3852,N_2595);
nand UO_891 (O_891,N_2591,N_2958);
or UO_892 (O_892,N_3758,N_4621);
nor UO_893 (O_893,N_3461,N_4061);
nor UO_894 (O_894,N_2933,N_3438);
or UO_895 (O_895,N_3034,N_4661);
xor UO_896 (O_896,N_4887,N_4828);
and UO_897 (O_897,N_2738,N_3175);
or UO_898 (O_898,N_3284,N_3183);
or UO_899 (O_899,N_4666,N_2754);
nor UO_900 (O_900,N_3063,N_3136);
xor UO_901 (O_901,N_4051,N_3343);
xnor UO_902 (O_902,N_4130,N_2563);
nand UO_903 (O_903,N_2962,N_3599);
nor UO_904 (O_904,N_2890,N_4303);
nor UO_905 (O_905,N_4394,N_3661);
and UO_906 (O_906,N_3719,N_3445);
and UO_907 (O_907,N_4534,N_2613);
xor UO_908 (O_908,N_3404,N_2864);
nand UO_909 (O_909,N_3226,N_2774);
and UO_910 (O_910,N_3647,N_4976);
nand UO_911 (O_911,N_4426,N_3781);
nor UO_912 (O_912,N_4943,N_3007);
nand UO_913 (O_913,N_3604,N_4293);
or UO_914 (O_914,N_3039,N_2989);
and UO_915 (O_915,N_3365,N_4197);
nand UO_916 (O_916,N_3701,N_3449);
xor UO_917 (O_917,N_4240,N_2518);
xnor UO_918 (O_918,N_3864,N_4147);
nand UO_919 (O_919,N_4348,N_3045);
and UO_920 (O_920,N_3004,N_3615);
and UO_921 (O_921,N_4158,N_4244);
nor UO_922 (O_922,N_2978,N_3387);
xor UO_923 (O_923,N_4902,N_3249);
or UO_924 (O_924,N_4701,N_2775);
nand UO_925 (O_925,N_3760,N_4023);
nor UO_926 (O_926,N_4036,N_4529);
nor UO_927 (O_927,N_2995,N_4865);
xnor UO_928 (O_928,N_4596,N_3278);
xnor UO_929 (O_929,N_2745,N_3152);
and UO_930 (O_930,N_3005,N_4341);
and UO_931 (O_931,N_4654,N_4356);
and UO_932 (O_932,N_4113,N_4932);
or UO_933 (O_933,N_4128,N_2856);
nand UO_934 (O_934,N_3906,N_4247);
and UO_935 (O_935,N_2722,N_4930);
or UO_936 (O_936,N_3793,N_2835);
nand UO_937 (O_937,N_3973,N_3550);
nor UO_938 (O_938,N_3172,N_4559);
nor UO_939 (O_939,N_3720,N_3246);
xor UO_940 (O_940,N_2967,N_2843);
and UO_941 (O_941,N_4512,N_3789);
nand UO_942 (O_942,N_2600,N_2630);
or UO_943 (O_943,N_3542,N_3573);
nor UO_944 (O_944,N_4573,N_2648);
nand UO_945 (O_945,N_3376,N_4475);
xor UO_946 (O_946,N_2576,N_4205);
xnor UO_947 (O_947,N_4246,N_3403);
nand UO_948 (O_948,N_4330,N_4082);
and UO_949 (O_949,N_2808,N_4276);
nor UO_950 (O_950,N_2861,N_4313);
and UO_951 (O_951,N_4922,N_2929);
nor UO_952 (O_952,N_4766,N_3584);
or UO_953 (O_953,N_2906,N_4237);
nor UO_954 (O_954,N_2651,N_2589);
nor UO_955 (O_955,N_2886,N_3352);
and UO_956 (O_956,N_2511,N_4024);
nand UO_957 (O_957,N_4841,N_3508);
and UO_958 (O_958,N_3443,N_3745);
nor UO_959 (O_959,N_2624,N_4302);
nor UO_960 (O_960,N_4239,N_4028);
and UO_961 (O_961,N_4238,N_4964);
and UO_962 (O_962,N_3893,N_2920);
nor UO_963 (O_963,N_3655,N_3565);
or UO_964 (O_964,N_2631,N_3046);
or UO_965 (O_965,N_4845,N_3056);
or UO_966 (O_966,N_3611,N_4296);
nor UO_967 (O_967,N_3779,N_4838);
or UO_968 (O_968,N_2922,N_4938);
nor UO_969 (O_969,N_3096,N_4919);
xnor UO_970 (O_970,N_3052,N_2781);
nand UO_971 (O_971,N_3997,N_3347);
or UO_972 (O_972,N_2641,N_4404);
nor UO_973 (O_973,N_4547,N_4507);
nand UO_974 (O_974,N_3771,N_2505);
or UO_975 (O_975,N_2941,N_4649);
xor UO_976 (O_976,N_2538,N_3095);
or UO_977 (O_977,N_4014,N_4278);
nor UO_978 (O_978,N_4624,N_2885);
and UO_979 (O_979,N_3987,N_4500);
and UO_980 (O_980,N_4409,N_3328);
or UO_981 (O_981,N_3345,N_4160);
nand UO_982 (O_982,N_3116,N_4123);
or UO_983 (O_983,N_3959,N_3577);
nand UO_984 (O_984,N_2853,N_4984);
or UO_985 (O_985,N_4834,N_4022);
or UO_986 (O_986,N_4351,N_2612);
xnor UO_987 (O_987,N_3003,N_3128);
xor UO_988 (O_988,N_3496,N_4410);
and UO_989 (O_989,N_4611,N_3645);
nand UO_990 (O_990,N_3800,N_3213);
or UO_991 (O_991,N_3399,N_4855);
and UO_992 (O_992,N_4052,N_3878);
nand UO_993 (O_993,N_3978,N_4098);
or UO_994 (O_994,N_4495,N_3450);
or UO_995 (O_995,N_2671,N_4376);
xnor UO_996 (O_996,N_4198,N_4388);
and UO_997 (O_997,N_4467,N_4153);
xor UO_998 (O_998,N_2776,N_3342);
nand UO_999 (O_999,N_4470,N_2705);
endmodule