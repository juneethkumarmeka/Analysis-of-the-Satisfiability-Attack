module basic_1000_10000_1500_5_levels_5xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nand U0 (N_0,In_794,In_278);
nor U1 (N_1,In_270,In_660);
or U2 (N_2,In_966,In_213);
nand U3 (N_3,In_439,In_42);
or U4 (N_4,In_547,In_591);
or U5 (N_5,In_40,In_463);
xnor U6 (N_6,In_623,In_344);
and U7 (N_7,In_609,In_723);
or U8 (N_8,In_722,In_556);
nand U9 (N_9,In_783,In_269);
nor U10 (N_10,In_995,In_90);
or U11 (N_11,In_369,In_301);
xnor U12 (N_12,In_837,In_186);
and U13 (N_13,In_587,In_230);
or U14 (N_14,In_629,In_529);
nand U15 (N_15,In_41,In_784);
nor U16 (N_16,In_858,In_296);
nand U17 (N_17,In_956,In_645);
or U18 (N_18,In_236,In_251);
nor U19 (N_19,In_974,In_504);
or U20 (N_20,In_949,In_738);
nor U21 (N_21,In_265,In_245);
or U22 (N_22,In_436,In_212);
nor U23 (N_23,In_688,In_55);
nand U24 (N_24,In_701,In_778);
nor U25 (N_25,In_300,In_295);
nand U26 (N_26,In_482,In_345);
nor U27 (N_27,In_443,In_33);
nand U28 (N_28,In_707,In_259);
and U29 (N_29,In_50,In_942);
and U30 (N_30,In_963,In_53);
xnor U31 (N_31,In_390,In_503);
nand U32 (N_32,In_931,In_351);
and U33 (N_33,In_462,In_170);
xor U34 (N_34,In_861,In_367);
nor U35 (N_35,In_842,In_135);
nand U36 (N_36,In_145,In_530);
or U37 (N_37,In_908,In_128);
or U38 (N_38,In_820,In_646);
nand U39 (N_39,In_275,In_161);
and U40 (N_40,In_194,In_287);
nand U41 (N_41,In_119,In_324);
and U42 (N_42,In_959,In_8);
or U43 (N_43,In_468,In_284);
nor U44 (N_44,In_435,In_457);
nand U45 (N_45,In_467,In_495);
or U46 (N_46,In_860,In_661);
or U47 (N_47,In_444,In_699);
nor U48 (N_48,In_322,In_597);
or U49 (N_49,In_334,In_249);
nor U50 (N_50,In_555,In_39);
nand U51 (N_51,In_593,In_473);
nand U52 (N_52,In_440,In_990);
or U53 (N_53,In_834,In_674);
xnor U54 (N_54,In_852,In_305);
nor U55 (N_55,In_209,In_810);
or U56 (N_56,In_365,In_184);
nor U57 (N_57,In_805,In_283);
and U58 (N_58,In_200,In_940);
nand U59 (N_59,In_747,In_330);
nor U60 (N_60,In_299,In_698);
and U61 (N_61,In_453,In_592);
nand U62 (N_62,In_204,In_628);
or U63 (N_63,In_341,In_233);
nor U64 (N_64,In_665,In_74);
nand U65 (N_65,In_621,In_590);
xnor U66 (N_66,In_420,In_122);
or U67 (N_67,In_835,In_441);
and U68 (N_68,In_166,In_653);
nor U69 (N_69,In_957,In_915);
or U70 (N_70,In_932,In_767);
or U71 (N_71,In_411,In_370);
and U72 (N_72,In_573,In_791);
nor U73 (N_73,In_340,In_45);
nand U74 (N_74,In_325,In_154);
nand U75 (N_75,In_558,In_920);
nor U76 (N_76,In_906,In_356);
nand U77 (N_77,In_313,In_884);
and U78 (N_78,In_537,In_950);
or U79 (N_79,In_17,In_790);
or U80 (N_80,In_712,In_536);
nor U81 (N_81,In_160,In_126);
nand U82 (N_82,In_903,In_879);
nor U83 (N_83,In_943,In_508);
nor U84 (N_84,In_402,In_358);
or U85 (N_85,In_152,In_760);
and U86 (N_86,In_512,In_899);
and U87 (N_87,In_538,In_190);
nor U88 (N_88,In_663,In_877);
and U89 (N_89,In_523,In_916);
and U90 (N_90,In_181,In_434);
or U91 (N_91,In_706,In_695);
or U92 (N_92,In_228,In_44);
nor U93 (N_93,In_531,In_427);
nor U94 (N_94,In_612,In_570);
or U95 (N_95,In_187,In_148);
nor U96 (N_96,In_757,In_242);
or U97 (N_97,In_286,In_828);
or U98 (N_98,In_195,In_282);
nor U99 (N_99,In_853,In_486);
nand U100 (N_100,In_261,In_851);
nor U101 (N_101,In_733,In_718);
nor U102 (N_102,In_132,In_541);
nand U103 (N_103,In_11,In_927);
or U104 (N_104,In_566,In_934);
and U105 (N_105,In_26,In_203);
nand U106 (N_106,In_938,In_456);
xnor U107 (N_107,In_856,In_936);
nand U108 (N_108,In_481,In_437);
or U109 (N_109,In_979,In_379);
and U110 (N_110,In_821,In_23);
nor U111 (N_111,In_826,In_27);
nor U112 (N_112,In_548,In_73);
nor U113 (N_113,In_37,In_475);
and U114 (N_114,In_543,In_279);
or U115 (N_115,In_1,In_825);
nor U116 (N_116,In_378,In_954);
nand U117 (N_117,In_280,In_546);
or U118 (N_118,In_363,In_110);
and U119 (N_119,In_227,In_525);
or U120 (N_120,In_338,In_897);
or U121 (N_121,In_400,In_193);
or U122 (N_122,In_180,In_923);
and U123 (N_123,In_297,In_347);
xnor U124 (N_124,In_422,In_844);
nand U125 (N_125,In_572,In_424);
nand U126 (N_126,In_32,In_409);
nor U127 (N_127,In_106,In_635);
nor U128 (N_128,In_291,In_658);
and U129 (N_129,In_501,In_214);
nand U130 (N_130,In_637,In_650);
nor U131 (N_131,In_211,In_777);
nand U132 (N_132,In_649,In_492);
nor U133 (N_133,In_999,In_490);
or U134 (N_134,In_735,In_670);
and U135 (N_135,In_127,In_406);
or U136 (N_136,In_859,In_375);
or U137 (N_137,In_780,In_891);
and U138 (N_138,In_306,In_361);
nand U139 (N_139,In_144,In_739);
or U140 (N_140,In_5,In_312);
nor U141 (N_141,In_65,In_937);
nand U142 (N_142,In_4,In_332);
or U143 (N_143,In_318,In_407);
nor U144 (N_144,In_958,In_466);
and U145 (N_145,In_813,In_841);
or U146 (N_146,In_253,In_880);
xor U147 (N_147,In_857,In_385);
nand U148 (N_148,In_526,In_307);
and U149 (N_149,In_395,In_292);
nor U150 (N_150,In_303,In_30);
xnor U151 (N_151,In_798,In_410);
or U152 (N_152,In_199,In_125);
nand U153 (N_153,In_578,In_745);
nand U154 (N_154,In_15,In_24);
xnor U155 (N_155,In_641,In_973);
or U156 (N_156,In_19,In_913);
xor U157 (N_157,In_716,In_383);
nor U158 (N_158,In_532,In_129);
nor U159 (N_159,In_54,In_631);
nand U160 (N_160,In_517,In_964);
nand U161 (N_161,In_445,In_933);
xnor U162 (N_162,In_61,In_878);
xor U163 (N_163,In_626,In_876);
and U164 (N_164,In_470,In_601);
nor U165 (N_165,In_732,In_364);
or U166 (N_166,In_192,In_3);
nand U167 (N_167,In_171,In_756);
and U168 (N_168,In_946,In_510);
and U169 (N_169,In_677,In_764);
or U170 (N_170,In_373,In_978);
and U171 (N_171,In_662,In_316);
and U172 (N_172,In_634,In_48);
and U173 (N_173,In_173,In_429);
nand U174 (N_174,In_75,In_667);
nand U175 (N_175,In_803,In_331);
nor U176 (N_176,In_93,In_70);
and U177 (N_177,In_516,In_359);
nor U178 (N_178,In_730,In_524);
nand U179 (N_179,In_206,In_518);
and U180 (N_180,In_225,In_560);
or U181 (N_181,In_57,In_666);
xnor U182 (N_182,In_496,In_918);
nor U183 (N_183,In_86,In_682);
nand U184 (N_184,In_99,In_602);
or U185 (N_185,In_31,In_46);
xor U186 (N_186,In_981,In_174);
nor U187 (N_187,In_534,In_172);
or U188 (N_188,In_52,In_874);
or U189 (N_189,In_800,In_575);
nand U190 (N_190,In_72,In_396);
and U191 (N_191,In_116,In_519);
nand U192 (N_192,In_766,In_246);
or U193 (N_193,In_360,In_502);
nor U194 (N_194,In_36,In_819);
or U195 (N_195,In_189,In_799);
and U196 (N_196,In_98,In_727);
nor U197 (N_197,In_792,In_627);
nand U198 (N_198,In_43,In_260);
or U199 (N_199,In_115,In_124);
and U200 (N_200,In_498,In_238);
xnor U201 (N_201,In_845,In_684);
and U202 (N_202,In_149,In_117);
nand U203 (N_203,In_185,In_740);
and U204 (N_204,In_571,In_673);
and U205 (N_205,In_337,In_693);
or U206 (N_206,In_352,In_714);
xnor U207 (N_207,In_690,In_277);
or U208 (N_208,In_644,In_162);
or U209 (N_209,In_522,In_461);
or U210 (N_210,In_909,In_892);
nand U211 (N_211,In_281,In_977);
nor U212 (N_212,In_133,In_768);
nor U213 (N_213,In_619,In_630);
nor U214 (N_214,In_136,In_59);
and U215 (N_215,In_394,In_500);
xnor U216 (N_216,In_219,In_382);
or U217 (N_217,In_729,In_980);
nand U218 (N_218,In_22,In_568);
xor U219 (N_219,In_140,In_655);
and U220 (N_220,In_247,In_314);
xnor U221 (N_221,In_355,In_472);
nand U222 (N_222,In_158,In_167);
nand U223 (N_223,In_561,In_875);
and U224 (N_224,In_871,In_838);
and U225 (N_225,In_450,In_188);
xnor U226 (N_226,In_986,In_762);
and U227 (N_227,In_16,In_432);
xor U228 (N_228,In_624,In_459);
nand U229 (N_229,In_890,In_335);
nor U230 (N_230,In_131,In_881);
nand U231 (N_231,In_2,In_51);
and U232 (N_232,In_721,In_528);
xor U233 (N_233,In_812,In_428);
and U234 (N_234,In_430,In_786);
or U235 (N_235,In_847,In_917);
and U236 (N_236,In_970,In_987);
nand U237 (N_237,In_616,In_288);
and U238 (N_238,In_659,In_357);
or U239 (N_239,In_539,In_506);
and U240 (N_240,In_807,In_788);
nand U241 (N_241,In_863,In_685);
nor U242 (N_242,In_885,In_368);
nand U243 (N_243,In_580,In_678);
or U244 (N_244,In_703,In_687);
and U245 (N_245,In_267,In_754);
and U246 (N_246,In_843,In_511);
nor U247 (N_247,In_273,In_285);
nor U248 (N_248,In_614,In_12);
or U249 (N_249,In_244,In_697);
nand U250 (N_250,In_551,In_968);
nand U251 (N_251,In_224,In_120);
and U252 (N_252,In_143,In_66);
nand U253 (N_253,In_736,In_724);
nand U254 (N_254,In_0,In_452);
nand U255 (N_255,In_535,In_507);
or U256 (N_256,In_464,In_728);
and U257 (N_257,In_67,In_380);
and U258 (N_258,In_71,In_309);
nand U259 (N_259,In_175,In_681);
or U260 (N_260,In_376,In_311);
nand U261 (N_261,In_618,In_771);
or U262 (N_262,In_711,In_971);
or U263 (N_263,In_588,In_342);
nor U264 (N_264,In_317,In_493);
and U265 (N_265,In_617,In_554);
nand U266 (N_266,In_773,In_708);
or U267 (N_267,In_755,In_221);
or U268 (N_268,In_328,In_272);
nand U269 (N_269,In_371,In_802);
nand U270 (N_270,In_888,In_914);
and U271 (N_271,In_290,In_945);
nand U272 (N_272,In_700,In_622);
nand U273 (N_273,In_640,In_239);
nor U274 (N_274,In_992,In_176);
or U275 (N_275,In_7,In_202);
nor U276 (N_276,In_408,In_669);
xnor U277 (N_277,In_56,In_607);
nand U278 (N_278,In_717,In_421);
nor U279 (N_279,In_222,In_625);
nand U280 (N_280,In_82,In_743);
nor U281 (N_281,In_632,In_392);
and U282 (N_282,In_961,In_919);
xor U283 (N_283,In_901,In_60);
nor U284 (N_284,In_169,In_121);
and U285 (N_285,In_513,In_95);
nor U286 (N_286,In_20,In_836);
or U287 (N_287,In_268,In_550);
and U288 (N_288,In_731,In_595);
nand U289 (N_289,In_78,In_774);
or U290 (N_290,In_865,In_654);
and U291 (N_291,In_354,In_178);
or U292 (N_292,In_586,In_704);
or U293 (N_293,In_226,In_509);
or U294 (N_294,In_930,In_737);
nand U295 (N_295,In_479,In_478);
nor U296 (N_296,In_862,In_208);
or U297 (N_297,In_254,In_753);
and U298 (N_298,In_846,In_983);
xnor U299 (N_299,In_585,In_955);
nand U300 (N_300,In_248,In_92);
or U301 (N_301,In_237,In_257);
or U302 (N_302,In_112,In_336);
or U303 (N_303,In_982,In_793);
nand U304 (N_304,In_579,In_480);
nand U305 (N_305,In_997,In_989);
or U306 (N_306,In_164,In_994);
and U307 (N_307,In_266,In_751);
nor U308 (N_308,In_157,In_89);
xor U309 (N_309,In_883,In_76);
or U310 (N_310,In_900,In_540);
nor U311 (N_311,In_811,In_928);
or U312 (N_312,In_346,In_873);
or U313 (N_313,In_894,In_474);
or U314 (N_314,In_196,In_118);
nor U315 (N_315,In_107,In_868);
or U316 (N_316,In_683,In_458);
or U317 (N_317,In_608,In_403);
nand U318 (N_318,In_469,In_386);
xnor U319 (N_319,In_97,In_159);
or U320 (N_320,In_201,In_77);
and U321 (N_321,In_829,In_652);
nand U322 (N_322,In_62,In_460);
or U323 (N_323,In_720,In_414);
xor U324 (N_324,In_809,In_141);
nor U325 (N_325,In_271,In_326);
or U326 (N_326,In_867,In_818);
nor U327 (N_327,In_263,In_638);
nand U328 (N_328,In_972,In_866);
or U329 (N_329,In_898,In_234);
xor U330 (N_330,In_744,In_565);
nand U331 (N_331,In_611,In_869);
nor U332 (N_332,In_220,In_569);
nand U333 (N_333,In_719,In_433);
or U334 (N_334,In_374,In_343);
and U335 (N_335,In_6,In_848);
or U336 (N_336,In_262,In_451);
and U337 (N_337,In_413,In_941);
nand U338 (N_338,In_864,In_553);
or U339 (N_339,In_431,In_715);
nand U340 (N_340,In_679,In_151);
or U341 (N_341,In_921,In_320);
nor U342 (N_342,In_146,In_80);
nand U343 (N_343,In_250,In_574);
xor U344 (N_344,In_58,In_564);
and U345 (N_345,In_710,In_103);
or U346 (N_346,In_804,In_763);
and U347 (N_347,In_870,In_223);
nor U348 (N_348,In_929,In_832);
or U349 (N_349,In_258,In_521);
and U350 (N_350,In_438,In_68);
or U351 (N_351,In_139,In_984);
nand U352 (N_352,In_398,In_599);
nor U353 (N_353,In_922,In_642);
nand U354 (N_354,In_150,In_217);
or U355 (N_355,In_18,In_533);
xnor U356 (N_356,In_63,In_339);
nand U357 (N_357,In_746,In_415);
nand U358 (N_358,In_134,In_887);
nor U359 (N_359,In_814,In_750);
nor U360 (N_360,In_9,In_494);
nand U361 (N_361,In_321,In_520);
xor U362 (N_362,In_713,In_976);
and U363 (N_363,In_417,In_606);
nand U364 (N_364,In_589,In_726);
nand U365 (N_365,In_489,In_581);
and U366 (N_366,In_680,In_404);
xnor U367 (N_367,In_372,In_64);
nor U368 (N_368,In_749,In_775);
nand U369 (N_369,In_948,In_13);
and U370 (N_370,In_84,In_21);
or U371 (N_371,In_675,In_975);
nor U372 (N_372,In_100,In_425);
nand U373 (N_373,In_232,In_85);
and U374 (N_374,In_639,In_985);
or U375 (N_375,In_882,In_557);
or U376 (N_376,In_387,In_109);
or U377 (N_377,In_789,In_787);
xor U378 (N_378,In_991,In_229);
or U379 (N_379,In_418,In_889);
nand U380 (N_380,In_902,In_758);
or U381 (N_381,In_765,In_672);
and U382 (N_382,In_643,In_240);
nand U383 (N_383,In_939,In_734);
and U384 (N_384,In_177,In_183);
and U385 (N_385,In_455,In_327);
or U386 (N_386,In_515,In_702);
or U387 (N_387,In_967,In_742);
and U388 (N_388,In_349,In_584);
or U389 (N_389,In_147,In_831);
nand U390 (N_390,In_231,In_497);
nor U391 (N_391,In_308,In_822);
and U392 (N_392,In_477,In_505);
or U393 (N_393,In_514,In_393);
nor U394 (N_394,In_633,In_485);
nand U395 (N_395,In_153,In_850);
xnor U396 (N_396,In_49,In_544);
or U397 (N_397,In_454,In_542);
nand U398 (N_398,In_353,In_319);
nand U399 (N_399,In_123,In_839);
and U400 (N_400,In_657,In_849);
or U401 (N_401,In_34,In_648);
or U402 (N_402,In_582,In_96);
nor U403 (N_403,In_419,In_333);
xor U404 (N_404,In_401,In_910);
or U405 (N_405,In_855,In_668);
nand U406 (N_406,In_600,In_748);
or U407 (N_407,In_692,In_442);
or U408 (N_408,In_576,In_694);
nand U409 (N_409,In_613,In_397);
nor U410 (N_410,In_276,In_953);
nand U411 (N_411,In_28,In_491);
nor U412 (N_412,In_210,In_993);
nor U413 (N_413,In_782,In_562);
xor U414 (N_414,In_448,In_113);
xor U415 (N_415,In_725,In_384);
and U416 (N_416,In_111,In_907);
nand U417 (N_417,In_952,In_545);
nor U418 (N_418,In_91,In_926);
and U419 (N_419,In_636,In_476);
nand U420 (N_420,In_197,In_83);
or U421 (N_421,In_304,In_664);
nor U422 (N_422,In_252,In_423);
nand U423 (N_423,In_761,In_274);
nor U424 (N_424,In_366,In_484);
and U425 (N_425,In_559,In_815);
or U426 (N_426,In_905,In_465);
nand U427 (N_427,In_323,In_998);
xnor U428 (N_428,In_389,In_895);
nor U429 (N_429,In_264,In_168);
nor U430 (N_430,In_329,In_620);
nor U431 (N_431,In_785,In_965);
nor U432 (N_432,In_302,In_951);
or U433 (N_433,In_88,In_38);
and U434 (N_434,In_647,In_362);
nor U435 (N_435,In_691,In_912);
nor U436 (N_436,In_594,In_577);
nor U437 (N_437,In_935,In_310);
or U438 (N_438,In_947,In_205);
xor U439 (N_439,In_25,In_709);
nand U440 (N_440,In_808,In_610);
and U441 (N_441,In_824,In_893);
nand U442 (N_442,In_769,In_705);
or U443 (N_443,In_69,In_488);
or U444 (N_444,In_911,In_255);
nor U445 (N_445,In_741,In_872);
nor U446 (N_446,In_549,In_138);
or U447 (N_447,In_904,In_686);
and U448 (N_448,In_759,In_182);
nand U449 (N_449,In_416,In_105);
nor U450 (N_450,In_471,In_35);
xor U451 (N_451,In_806,In_886);
xnor U452 (N_452,In_216,In_776);
nand U453 (N_453,In_47,In_10);
and U454 (N_454,In_483,In_527);
nand U455 (N_455,In_405,In_81);
nand U456 (N_456,In_924,In_962);
and U457 (N_457,In_207,In_108);
and U458 (N_458,In_823,In_101);
and U459 (N_459,In_315,In_615);
or U460 (N_460,In_796,In_388);
nand U461 (N_461,In_137,In_689);
and U462 (N_462,In_426,In_142);
nor U463 (N_463,In_598,In_583);
nor U464 (N_464,In_391,In_779);
nand U465 (N_465,In_960,In_833);
and U466 (N_466,In_348,In_29);
nor U467 (N_467,In_988,In_114);
nand U468 (N_468,In_198,In_399);
nand U469 (N_469,In_840,In_381);
or U470 (N_470,In_487,In_696);
or U471 (N_471,In_289,In_801);
or U472 (N_472,In_179,In_94);
nor U473 (N_473,In_651,In_218);
or U474 (N_474,In_155,In_603);
nand U475 (N_475,In_567,In_795);
nand U476 (N_476,In_944,In_350);
nor U477 (N_477,In_156,In_676);
nand U478 (N_478,In_797,In_563);
or U479 (N_479,In_235,In_449);
and U480 (N_480,In_14,In_854);
or U481 (N_481,In_604,In_996);
nor U482 (N_482,In_605,In_241);
or U483 (N_483,In_830,In_104);
xnor U484 (N_484,In_447,In_896);
and U485 (N_485,In_130,In_191);
and U486 (N_486,In_816,In_770);
or U487 (N_487,In_165,In_671);
or U488 (N_488,In_552,In_298);
nor U489 (N_489,In_925,In_772);
or U490 (N_490,In_87,In_969);
or U491 (N_491,In_781,In_243);
and U492 (N_492,In_256,In_827);
or U493 (N_493,In_79,In_215);
or U494 (N_494,In_163,In_499);
and U495 (N_495,In_446,In_294);
or U496 (N_496,In_817,In_412);
and U497 (N_497,In_752,In_596);
nand U498 (N_498,In_293,In_102);
nand U499 (N_499,In_377,In_656);
and U500 (N_500,In_528,In_31);
nand U501 (N_501,In_372,In_553);
nor U502 (N_502,In_908,In_112);
and U503 (N_503,In_879,In_120);
nor U504 (N_504,In_767,In_130);
nor U505 (N_505,In_157,In_730);
or U506 (N_506,In_348,In_253);
and U507 (N_507,In_298,In_261);
xor U508 (N_508,In_979,In_273);
nand U509 (N_509,In_775,In_738);
and U510 (N_510,In_389,In_637);
or U511 (N_511,In_157,In_23);
nand U512 (N_512,In_182,In_401);
nor U513 (N_513,In_559,In_199);
nand U514 (N_514,In_120,In_619);
nand U515 (N_515,In_701,In_206);
nor U516 (N_516,In_445,In_343);
and U517 (N_517,In_453,In_88);
nand U518 (N_518,In_328,In_719);
nor U519 (N_519,In_344,In_170);
nand U520 (N_520,In_661,In_53);
nand U521 (N_521,In_458,In_925);
nor U522 (N_522,In_447,In_686);
xor U523 (N_523,In_538,In_966);
nor U524 (N_524,In_793,In_152);
nand U525 (N_525,In_367,In_15);
nor U526 (N_526,In_837,In_617);
and U527 (N_527,In_824,In_654);
and U528 (N_528,In_151,In_858);
xor U529 (N_529,In_232,In_32);
or U530 (N_530,In_199,In_3);
nor U531 (N_531,In_950,In_592);
nand U532 (N_532,In_322,In_280);
or U533 (N_533,In_603,In_103);
or U534 (N_534,In_198,In_514);
nand U535 (N_535,In_448,In_484);
and U536 (N_536,In_47,In_972);
and U537 (N_537,In_497,In_655);
nand U538 (N_538,In_818,In_383);
nor U539 (N_539,In_645,In_293);
nor U540 (N_540,In_92,In_961);
nor U541 (N_541,In_484,In_417);
nor U542 (N_542,In_716,In_252);
and U543 (N_543,In_303,In_368);
or U544 (N_544,In_571,In_796);
or U545 (N_545,In_225,In_374);
or U546 (N_546,In_101,In_701);
xnor U547 (N_547,In_449,In_313);
nand U548 (N_548,In_255,In_126);
nor U549 (N_549,In_751,In_633);
and U550 (N_550,In_314,In_575);
or U551 (N_551,In_3,In_215);
and U552 (N_552,In_887,In_372);
nand U553 (N_553,In_321,In_311);
and U554 (N_554,In_629,In_896);
or U555 (N_555,In_911,In_725);
xor U556 (N_556,In_288,In_672);
and U557 (N_557,In_279,In_405);
nand U558 (N_558,In_593,In_994);
nor U559 (N_559,In_569,In_262);
and U560 (N_560,In_368,In_134);
nor U561 (N_561,In_786,In_126);
or U562 (N_562,In_287,In_361);
or U563 (N_563,In_491,In_5);
or U564 (N_564,In_740,In_913);
and U565 (N_565,In_495,In_441);
nor U566 (N_566,In_364,In_91);
nor U567 (N_567,In_95,In_38);
or U568 (N_568,In_848,In_463);
nand U569 (N_569,In_419,In_759);
nand U570 (N_570,In_356,In_232);
and U571 (N_571,In_493,In_614);
nor U572 (N_572,In_250,In_510);
and U573 (N_573,In_299,In_781);
xor U574 (N_574,In_517,In_762);
xor U575 (N_575,In_684,In_436);
or U576 (N_576,In_433,In_373);
and U577 (N_577,In_338,In_909);
and U578 (N_578,In_836,In_778);
nor U579 (N_579,In_739,In_44);
xnor U580 (N_580,In_170,In_666);
nand U581 (N_581,In_911,In_835);
nand U582 (N_582,In_449,In_180);
or U583 (N_583,In_74,In_914);
and U584 (N_584,In_1,In_68);
xor U585 (N_585,In_768,In_837);
or U586 (N_586,In_800,In_127);
nor U587 (N_587,In_187,In_337);
or U588 (N_588,In_340,In_677);
nand U589 (N_589,In_445,In_433);
and U590 (N_590,In_675,In_879);
and U591 (N_591,In_609,In_923);
xnor U592 (N_592,In_873,In_575);
nand U593 (N_593,In_818,In_304);
or U594 (N_594,In_992,In_417);
nor U595 (N_595,In_691,In_169);
nand U596 (N_596,In_54,In_179);
nand U597 (N_597,In_355,In_17);
or U598 (N_598,In_887,In_62);
nor U599 (N_599,In_214,In_724);
nand U600 (N_600,In_890,In_121);
nand U601 (N_601,In_769,In_539);
nand U602 (N_602,In_844,In_400);
xor U603 (N_603,In_959,In_629);
or U604 (N_604,In_882,In_747);
or U605 (N_605,In_580,In_203);
or U606 (N_606,In_495,In_119);
and U607 (N_607,In_631,In_175);
and U608 (N_608,In_320,In_448);
and U609 (N_609,In_109,In_726);
nand U610 (N_610,In_478,In_888);
and U611 (N_611,In_817,In_291);
and U612 (N_612,In_691,In_239);
nor U613 (N_613,In_793,In_30);
xor U614 (N_614,In_98,In_657);
nor U615 (N_615,In_540,In_999);
and U616 (N_616,In_377,In_940);
or U617 (N_617,In_267,In_446);
xor U618 (N_618,In_799,In_289);
nor U619 (N_619,In_726,In_27);
nand U620 (N_620,In_115,In_559);
or U621 (N_621,In_295,In_346);
and U622 (N_622,In_356,In_734);
nor U623 (N_623,In_177,In_901);
and U624 (N_624,In_614,In_577);
nand U625 (N_625,In_677,In_426);
or U626 (N_626,In_152,In_156);
xor U627 (N_627,In_33,In_289);
and U628 (N_628,In_942,In_870);
and U629 (N_629,In_927,In_500);
nand U630 (N_630,In_412,In_660);
nand U631 (N_631,In_472,In_516);
nand U632 (N_632,In_602,In_573);
nor U633 (N_633,In_757,In_530);
nand U634 (N_634,In_162,In_824);
or U635 (N_635,In_68,In_751);
or U636 (N_636,In_945,In_434);
and U637 (N_637,In_141,In_113);
or U638 (N_638,In_536,In_191);
and U639 (N_639,In_503,In_941);
or U640 (N_640,In_122,In_920);
and U641 (N_641,In_434,In_130);
and U642 (N_642,In_486,In_623);
xnor U643 (N_643,In_330,In_324);
and U644 (N_644,In_394,In_469);
nor U645 (N_645,In_135,In_629);
xor U646 (N_646,In_991,In_714);
nor U647 (N_647,In_742,In_792);
or U648 (N_648,In_455,In_143);
and U649 (N_649,In_834,In_359);
nand U650 (N_650,In_786,In_509);
or U651 (N_651,In_783,In_460);
nor U652 (N_652,In_128,In_367);
nor U653 (N_653,In_391,In_25);
nor U654 (N_654,In_953,In_873);
and U655 (N_655,In_691,In_847);
nor U656 (N_656,In_789,In_485);
xor U657 (N_657,In_647,In_980);
and U658 (N_658,In_821,In_12);
nand U659 (N_659,In_852,In_302);
and U660 (N_660,In_612,In_562);
or U661 (N_661,In_564,In_913);
or U662 (N_662,In_894,In_782);
and U663 (N_663,In_759,In_148);
nand U664 (N_664,In_714,In_433);
nor U665 (N_665,In_231,In_54);
nor U666 (N_666,In_15,In_214);
or U667 (N_667,In_905,In_637);
xor U668 (N_668,In_382,In_259);
xor U669 (N_669,In_92,In_144);
nand U670 (N_670,In_152,In_661);
nand U671 (N_671,In_686,In_337);
and U672 (N_672,In_442,In_852);
or U673 (N_673,In_806,In_167);
and U674 (N_674,In_623,In_657);
xnor U675 (N_675,In_102,In_554);
and U676 (N_676,In_914,In_468);
nor U677 (N_677,In_53,In_757);
or U678 (N_678,In_599,In_571);
xnor U679 (N_679,In_668,In_353);
or U680 (N_680,In_183,In_499);
nand U681 (N_681,In_947,In_397);
or U682 (N_682,In_52,In_557);
or U683 (N_683,In_262,In_489);
or U684 (N_684,In_281,In_584);
xnor U685 (N_685,In_260,In_492);
nor U686 (N_686,In_225,In_52);
and U687 (N_687,In_549,In_593);
or U688 (N_688,In_424,In_628);
nor U689 (N_689,In_178,In_696);
and U690 (N_690,In_198,In_497);
nand U691 (N_691,In_986,In_880);
and U692 (N_692,In_551,In_171);
and U693 (N_693,In_691,In_926);
nor U694 (N_694,In_75,In_763);
and U695 (N_695,In_378,In_105);
xnor U696 (N_696,In_915,In_661);
and U697 (N_697,In_48,In_396);
or U698 (N_698,In_136,In_242);
xnor U699 (N_699,In_806,In_972);
and U700 (N_700,In_553,In_276);
and U701 (N_701,In_570,In_286);
nand U702 (N_702,In_848,In_879);
and U703 (N_703,In_987,In_258);
and U704 (N_704,In_506,In_889);
nor U705 (N_705,In_992,In_116);
nor U706 (N_706,In_284,In_65);
nor U707 (N_707,In_400,In_267);
nand U708 (N_708,In_228,In_249);
nand U709 (N_709,In_842,In_496);
nand U710 (N_710,In_940,In_637);
or U711 (N_711,In_679,In_127);
or U712 (N_712,In_691,In_918);
or U713 (N_713,In_273,In_213);
xnor U714 (N_714,In_49,In_78);
and U715 (N_715,In_215,In_885);
xnor U716 (N_716,In_996,In_696);
nand U717 (N_717,In_496,In_725);
and U718 (N_718,In_592,In_58);
nor U719 (N_719,In_64,In_940);
and U720 (N_720,In_839,In_974);
nor U721 (N_721,In_366,In_501);
nor U722 (N_722,In_811,In_431);
nor U723 (N_723,In_700,In_630);
or U724 (N_724,In_427,In_158);
xnor U725 (N_725,In_696,In_568);
and U726 (N_726,In_932,In_293);
or U727 (N_727,In_771,In_153);
and U728 (N_728,In_814,In_622);
nand U729 (N_729,In_555,In_298);
and U730 (N_730,In_446,In_461);
nor U731 (N_731,In_382,In_14);
or U732 (N_732,In_593,In_929);
nor U733 (N_733,In_842,In_775);
or U734 (N_734,In_226,In_10);
nor U735 (N_735,In_707,In_321);
nor U736 (N_736,In_860,In_807);
or U737 (N_737,In_63,In_876);
or U738 (N_738,In_326,In_142);
nor U739 (N_739,In_239,In_497);
nor U740 (N_740,In_409,In_472);
nor U741 (N_741,In_695,In_205);
or U742 (N_742,In_663,In_856);
nand U743 (N_743,In_943,In_689);
or U744 (N_744,In_885,In_209);
xnor U745 (N_745,In_718,In_385);
xnor U746 (N_746,In_784,In_543);
and U747 (N_747,In_416,In_612);
xnor U748 (N_748,In_712,In_160);
nand U749 (N_749,In_249,In_452);
nand U750 (N_750,In_378,In_609);
nand U751 (N_751,In_320,In_180);
nand U752 (N_752,In_6,In_505);
nor U753 (N_753,In_531,In_23);
xor U754 (N_754,In_397,In_49);
or U755 (N_755,In_620,In_447);
or U756 (N_756,In_682,In_338);
nor U757 (N_757,In_163,In_115);
and U758 (N_758,In_241,In_509);
nor U759 (N_759,In_298,In_68);
or U760 (N_760,In_950,In_813);
nor U761 (N_761,In_667,In_623);
or U762 (N_762,In_432,In_87);
or U763 (N_763,In_672,In_724);
nand U764 (N_764,In_768,In_428);
nor U765 (N_765,In_232,In_309);
nor U766 (N_766,In_653,In_793);
or U767 (N_767,In_592,In_539);
or U768 (N_768,In_955,In_266);
xnor U769 (N_769,In_985,In_396);
and U770 (N_770,In_898,In_452);
xnor U771 (N_771,In_61,In_675);
xor U772 (N_772,In_761,In_44);
and U773 (N_773,In_146,In_322);
xnor U774 (N_774,In_152,In_375);
nor U775 (N_775,In_696,In_675);
or U776 (N_776,In_928,In_335);
or U777 (N_777,In_418,In_35);
xnor U778 (N_778,In_677,In_493);
nand U779 (N_779,In_406,In_574);
nand U780 (N_780,In_556,In_706);
or U781 (N_781,In_782,In_968);
or U782 (N_782,In_794,In_826);
nand U783 (N_783,In_131,In_139);
or U784 (N_784,In_15,In_705);
and U785 (N_785,In_226,In_515);
nor U786 (N_786,In_608,In_227);
and U787 (N_787,In_49,In_413);
xor U788 (N_788,In_63,In_929);
or U789 (N_789,In_474,In_93);
and U790 (N_790,In_998,In_852);
nand U791 (N_791,In_58,In_534);
or U792 (N_792,In_922,In_312);
xnor U793 (N_793,In_229,In_750);
nor U794 (N_794,In_444,In_284);
and U795 (N_795,In_288,In_296);
xnor U796 (N_796,In_122,In_108);
nand U797 (N_797,In_171,In_768);
or U798 (N_798,In_173,In_537);
nand U799 (N_799,In_947,In_769);
nor U800 (N_800,In_384,In_197);
or U801 (N_801,In_740,In_288);
or U802 (N_802,In_249,In_612);
and U803 (N_803,In_545,In_977);
or U804 (N_804,In_662,In_253);
and U805 (N_805,In_206,In_461);
xor U806 (N_806,In_704,In_47);
nand U807 (N_807,In_920,In_131);
nand U808 (N_808,In_796,In_766);
nand U809 (N_809,In_951,In_772);
or U810 (N_810,In_737,In_560);
or U811 (N_811,In_749,In_993);
nand U812 (N_812,In_636,In_673);
nor U813 (N_813,In_61,In_454);
and U814 (N_814,In_392,In_875);
or U815 (N_815,In_19,In_410);
and U816 (N_816,In_489,In_525);
and U817 (N_817,In_505,In_676);
nand U818 (N_818,In_648,In_285);
or U819 (N_819,In_835,In_567);
nor U820 (N_820,In_388,In_842);
or U821 (N_821,In_467,In_899);
nor U822 (N_822,In_28,In_889);
nand U823 (N_823,In_265,In_295);
and U824 (N_824,In_815,In_607);
nand U825 (N_825,In_645,In_275);
nor U826 (N_826,In_697,In_962);
xor U827 (N_827,In_541,In_334);
nand U828 (N_828,In_317,In_221);
nor U829 (N_829,In_735,In_10);
nor U830 (N_830,In_287,In_228);
nor U831 (N_831,In_241,In_623);
nor U832 (N_832,In_210,In_337);
nand U833 (N_833,In_174,In_366);
or U834 (N_834,In_797,In_14);
nand U835 (N_835,In_928,In_589);
or U836 (N_836,In_395,In_130);
and U837 (N_837,In_172,In_995);
or U838 (N_838,In_454,In_596);
nand U839 (N_839,In_961,In_891);
and U840 (N_840,In_156,In_276);
or U841 (N_841,In_80,In_929);
or U842 (N_842,In_309,In_484);
nor U843 (N_843,In_328,In_60);
nand U844 (N_844,In_543,In_863);
nand U845 (N_845,In_981,In_383);
xnor U846 (N_846,In_904,In_788);
nand U847 (N_847,In_597,In_688);
or U848 (N_848,In_186,In_472);
nand U849 (N_849,In_959,In_670);
nand U850 (N_850,In_913,In_279);
or U851 (N_851,In_846,In_839);
or U852 (N_852,In_701,In_45);
nand U853 (N_853,In_210,In_320);
nor U854 (N_854,In_381,In_366);
nand U855 (N_855,In_62,In_255);
and U856 (N_856,In_261,In_653);
or U857 (N_857,In_417,In_734);
nor U858 (N_858,In_888,In_462);
and U859 (N_859,In_932,In_613);
nor U860 (N_860,In_96,In_342);
nor U861 (N_861,In_767,In_629);
xnor U862 (N_862,In_979,In_274);
nor U863 (N_863,In_903,In_428);
nand U864 (N_864,In_970,In_371);
or U865 (N_865,In_696,In_8);
nand U866 (N_866,In_887,In_643);
xor U867 (N_867,In_603,In_732);
xnor U868 (N_868,In_497,In_869);
and U869 (N_869,In_271,In_25);
nand U870 (N_870,In_812,In_592);
and U871 (N_871,In_313,In_534);
xor U872 (N_872,In_31,In_552);
and U873 (N_873,In_575,In_948);
nand U874 (N_874,In_870,In_627);
or U875 (N_875,In_59,In_558);
or U876 (N_876,In_215,In_52);
nand U877 (N_877,In_237,In_282);
or U878 (N_878,In_371,In_139);
nand U879 (N_879,In_936,In_476);
and U880 (N_880,In_943,In_763);
nor U881 (N_881,In_34,In_356);
nor U882 (N_882,In_520,In_581);
or U883 (N_883,In_914,In_432);
or U884 (N_884,In_607,In_590);
nand U885 (N_885,In_929,In_808);
xor U886 (N_886,In_280,In_691);
and U887 (N_887,In_629,In_806);
nand U888 (N_888,In_843,In_112);
or U889 (N_889,In_359,In_32);
nor U890 (N_890,In_366,In_765);
nor U891 (N_891,In_290,In_122);
and U892 (N_892,In_454,In_706);
or U893 (N_893,In_126,In_372);
nand U894 (N_894,In_984,In_369);
or U895 (N_895,In_875,In_312);
and U896 (N_896,In_299,In_203);
nor U897 (N_897,In_59,In_113);
nand U898 (N_898,In_0,In_913);
and U899 (N_899,In_162,In_430);
nand U900 (N_900,In_255,In_103);
and U901 (N_901,In_930,In_712);
xor U902 (N_902,In_233,In_581);
xnor U903 (N_903,In_322,In_37);
or U904 (N_904,In_900,In_887);
or U905 (N_905,In_21,In_463);
nand U906 (N_906,In_46,In_732);
and U907 (N_907,In_752,In_569);
or U908 (N_908,In_398,In_914);
and U909 (N_909,In_498,In_927);
and U910 (N_910,In_160,In_53);
nand U911 (N_911,In_14,In_955);
nand U912 (N_912,In_623,In_961);
nand U913 (N_913,In_453,In_665);
nand U914 (N_914,In_236,In_155);
nand U915 (N_915,In_654,In_849);
or U916 (N_916,In_152,In_179);
nand U917 (N_917,In_712,In_974);
and U918 (N_918,In_847,In_668);
xor U919 (N_919,In_653,In_569);
nor U920 (N_920,In_767,In_84);
and U921 (N_921,In_246,In_181);
xnor U922 (N_922,In_564,In_165);
or U923 (N_923,In_660,In_478);
nor U924 (N_924,In_212,In_124);
or U925 (N_925,In_206,In_205);
nor U926 (N_926,In_527,In_826);
nand U927 (N_927,In_853,In_284);
xor U928 (N_928,In_632,In_661);
and U929 (N_929,In_134,In_778);
xnor U930 (N_930,In_734,In_535);
or U931 (N_931,In_15,In_657);
or U932 (N_932,In_2,In_346);
or U933 (N_933,In_289,In_598);
nand U934 (N_934,In_239,In_228);
and U935 (N_935,In_474,In_393);
nor U936 (N_936,In_850,In_47);
nand U937 (N_937,In_527,In_441);
nor U938 (N_938,In_292,In_124);
nand U939 (N_939,In_936,In_960);
nand U940 (N_940,In_833,In_425);
nor U941 (N_941,In_617,In_183);
nand U942 (N_942,In_575,In_712);
or U943 (N_943,In_816,In_359);
or U944 (N_944,In_53,In_81);
nand U945 (N_945,In_699,In_379);
and U946 (N_946,In_407,In_527);
and U947 (N_947,In_232,In_794);
or U948 (N_948,In_100,In_663);
nand U949 (N_949,In_704,In_935);
or U950 (N_950,In_876,In_718);
or U951 (N_951,In_594,In_699);
and U952 (N_952,In_71,In_127);
and U953 (N_953,In_725,In_900);
or U954 (N_954,In_101,In_486);
nand U955 (N_955,In_776,In_783);
xor U956 (N_956,In_476,In_488);
or U957 (N_957,In_814,In_751);
nand U958 (N_958,In_93,In_33);
and U959 (N_959,In_959,In_412);
nor U960 (N_960,In_345,In_60);
or U961 (N_961,In_492,In_799);
xnor U962 (N_962,In_983,In_900);
xnor U963 (N_963,In_284,In_100);
nand U964 (N_964,In_398,In_34);
or U965 (N_965,In_676,In_699);
nor U966 (N_966,In_801,In_426);
nand U967 (N_967,In_465,In_293);
nor U968 (N_968,In_981,In_16);
nand U969 (N_969,In_429,In_402);
nand U970 (N_970,In_45,In_654);
nor U971 (N_971,In_352,In_422);
xnor U972 (N_972,In_385,In_732);
or U973 (N_973,In_103,In_247);
and U974 (N_974,In_633,In_35);
or U975 (N_975,In_27,In_729);
nand U976 (N_976,In_181,In_326);
xnor U977 (N_977,In_929,In_290);
and U978 (N_978,In_781,In_577);
nor U979 (N_979,In_87,In_779);
or U980 (N_980,In_195,In_324);
nand U981 (N_981,In_569,In_580);
or U982 (N_982,In_633,In_170);
nand U983 (N_983,In_843,In_58);
or U984 (N_984,In_80,In_809);
nor U985 (N_985,In_50,In_140);
nand U986 (N_986,In_168,In_654);
nand U987 (N_987,In_546,In_445);
nor U988 (N_988,In_19,In_198);
xor U989 (N_989,In_115,In_682);
nor U990 (N_990,In_299,In_624);
nand U991 (N_991,In_184,In_134);
nand U992 (N_992,In_943,In_757);
and U993 (N_993,In_121,In_173);
nor U994 (N_994,In_899,In_0);
and U995 (N_995,In_110,In_50);
or U996 (N_996,In_184,In_842);
or U997 (N_997,In_312,In_739);
nand U998 (N_998,In_303,In_37);
nand U999 (N_999,In_52,In_572);
nor U1000 (N_1000,In_451,In_746);
or U1001 (N_1001,In_192,In_289);
and U1002 (N_1002,In_866,In_310);
and U1003 (N_1003,In_521,In_613);
nand U1004 (N_1004,In_814,In_233);
nand U1005 (N_1005,In_314,In_533);
nand U1006 (N_1006,In_463,In_371);
and U1007 (N_1007,In_950,In_15);
nor U1008 (N_1008,In_374,In_200);
and U1009 (N_1009,In_94,In_434);
nor U1010 (N_1010,In_173,In_435);
nor U1011 (N_1011,In_436,In_728);
and U1012 (N_1012,In_131,In_404);
and U1013 (N_1013,In_407,In_862);
nor U1014 (N_1014,In_706,In_95);
or U1015 (N_1015,In_140,In_761);
and U1016 (N_1016,In_625,In_632);
nor U1017 (N_1017,In_73,In_435);
nor U1018 (N_1018,In_973,In_981);
nand U1019 (N_1019,In_140,In_211);
nand U1020 (N_1020,In_293,In_5);
or U1021 (N_1021,In_125,In_919);
or U1022 (N_1022,In_55,In_383);
and U1023 (N_1023,In_789,In_562);
and U1024 (N_1024,In_847,In_164);
or U1025 (N_1025,In_922,In_858);
or U1026 (N_1026,In_23,In_871);
nand U1027 (N_1027,In_759,In_259);
nand U1028 (N_1028,In_138,In_953);
or U1029 (N_1029,In_374,In_264);
and U1030 (N_1030,In_587,In_933);
xnor U1031 (N_1031,In_932,In_511);
nand U1032 (N_1032,In_780,In_69);
or U1033 (N_1033,In_456,In_230);
nand U1034 (N_1034,In_635,In_623);
nand U1035 (N_1035,In_478,In_589);
or U1036 (N_1036,In_120,In_495);
nor U1037 (N_1037,In_395,In_366);
xor U1038 (N_1038,In_301,In_857);
nand U1039 (N_1039,In_286,In_306);
or U1040 (N_1040,In_217,In_651);
or U1041 (N_1041,In_434,In_296);
and U1042 (N_1042,In_268,In_453);
and U1043 (N_1043,In_188,In_235);
xor U1044 (N_1044,In_903,In_833);
nor U1045 (N_1045,In_422,In_500);
nand U1046 (N_1046,In_643,In_548);
nand U1047 (N_1047,In_8,In_382);
nand U1048 (N_1048,In_487,In_939);
or U1049 (N_1049,In_481,In_313);
nand U1050 (N_1050,In_332,In_904);
and U1051 (N_1051,In_688,In_878);
nor U1052 (N_1052,In_540,In_103);
or U1053 (N_1053,In_865,In_954);
nand U1054 (N_1054,In_753,In_429);
xor U1055 (N_1055,In_630,In_674);
nand U1056 (N_1056,In_586,In_557);
or U1057 (N_1057,In_743,In_703);
nor U1058 (N_1058,In_104,In_158);
nor U1059 (N_1059,In_56,In_681);
nor U1060 (N_1060,In_535,In_930);
nor U1061 (N_1061,In_995,In_348);
nand U1062 (N_1062,In_380,In_486);
nand U1063 (N_1063,In_778,In_556);
xor U1064 (N_1064,In_113,In_550);
nor U1065 (N_1065,In_577,In_423);
nand U1066 (N_1066,In_935,In_228);
nor U1067 (N_1067,In_666,In_845);
or U1068 (N_1068,In_817,In_889);
nand U1069 (N_1069,In_868,In_199);
and U1070 (N_1070,In_343,In_567);
nand U1071 (N_1071,In_982,In_145);
or U1072 (N_1072,In_646,In_821);
and U1073 (N_1073,In_461,In_780);
nand U1074 (N_1074,In_242,In_348);
nor U1075 (N_1075,In_390,In_628);
nor U1076 (N_1076,In_452,In_295);
or U1077 (N_1077,In_50,In_931);
nor U1078 (N_1078,In_653,In_1);
nand U1079 (N_1079,In_307,In_932);
or U1080 (N_1080,In_295,In_987);
and U1081 (N_1081,In_771,In_64);
or U1082 (N_1082,In_699,In_300);
nand U1083 (N_1083,In_696,In_627);
or U1084 (N_1084,In_315,In_850);
and U1085 (N_1085,In_741,In_745);
nor U1086 (N_1086,In_425,In_495);
nor U1087 (N_1087,In_452,In_311);
or U1088 (N_1088,In_689,In_391);
or U1089 (N_1089,In_913,In_657);
and U1090 (N_1090,In_263,In_734);
nor U1091 (N_1091,In_403,In_777);
nand U1092 (N_1092,In_404,In_246);
and U1093 (N_1093,In_534,In_583);
nor U1094 (N_1094,In_548,In_81);
nand U1095 (N_1095,In_645,In_376);
xnor U1096 (N_1096,In_537,In_819);
nor U1097 (N_1097,In_877,In_292);
or U1098 (N_1098,In_74,In_984);
nand U1099 (N_1099,In_254,In_713);
nand U1100 (N_1100,In_178,In_375);
nand U1101 (N_1101,In_946,In_870);
or U1102 (N_1102,In_675,In_972);
or U1103 (N_1103,In_647,In_519);
nor U1104 (N_1104,In_283,In_816);
nor U1105 (N_1105,In_401,In_954);
nand U1106 (N_1106,In_288,In_381);
nor U1107 (N_1107,In_283,In_786);
nand U1108 (N_1108,In_74,In_61);
and U1109 (N_1109,In_289,In_458);
nand U1110 (N_1110,In_314,In_857);
or U1111 (N_1111,In_753,In_252);
nor U1112 (N_1112,In_752,In_43);
or U1113 (N_1113,In_555,In_161);
nor U1114 (N_1114,In_391,In_530);
nor U1115 (N_1115,In_250,In_851);
or U1116 (N_1116,In_864,In_783);
xor U1117 (N_1117,In_219,In_896);
nor U1118 (N_1118,In_253,In_401);
xor U1119 (N_1119,In_680,In_322);
nor U1120 (N_1120,In_438,In_708);
and U1121 (N_1121,In_258,In_830);
and U1122 (N_1122,In_959,In_923);
nand U1123 (N_1123,In_363,In_204);
and U1124 (N_1124,In_931,In_822);
and U1125 (N_1125,In_60,In_50);
xnor U1126 (N_1126,In_158,In_351);
xor U1127 (N_1127,In_893,In_593);
nor U1128 (N_1128,In_634,In_321);
nand U1129 (N_1129,In_345,In_923);
or U1130 (N_1130,In_875,In_247);
nand U1131 (N_1131,In_434,In_139);
or U1132 (N_1132,In_256,In_940);
and U1133 (N_1133,In_123,In_66);
and U1134 (N_1134,In_490,In_985);
and U1135 (N_1135,In_191,In_48);
nand U1136 (N_1136,In_712,In_507);
nor U1137 (N_1137,In_756,In_436);
nand U1138 (N_1138,In_557,In_393);
nand U1139 (N_1139,In_605,In_773);
or U1140 (N_1140,In_814,In_546);
and U1141 (N_1141,In_278,In_185);
or U1142 (N_1142,In_645,In_660);
or U1143 (N_1143,In_843,In_695);
or U1144 (N_1144,In_213,In_243);
or U1145 (N_1145,In_65,In_136);
nor U1146 (N_1146,In_329,In_386);
nor U1147 (N_1147,In_933,In_997);
nor U1148 (N_1148,In_221,In_859);
nand U1149 (N_1149,In_896,In_618);
and U1150 (N_1150,In_555,In_146);
nor U1151 (N_1151,In_826,In_114);
and U1152 (N_1152,In_574,In_447);
nor U1153 (N_1153,In_228,In_331);
nor U1154 (N_1154,In_53,In_990);
or U1155 (N_1155,In_82,In_721);
nand U1156 (N_1156,In_753,In_968);
and U1157 (N_1157,In_663,In_993);
and U1158 (N_1158,In_209,In_774);
and U1159 (N_1159,In_45,In_181);
nand U1160 (N_1160,In_614,In_572);
or U1161 (N_1161,In_879,In_453);
and U1162 (N_1162,In_330,In_749);
nand U1163 (N_1163,In_943,In_932);
xnor U1164 (N_1164,In_816,In_476);
nand U1165 (N_1165,In_424,In_889);
or U1166 (N_1166,In_990,In_589);
and U1167 (N_1167,In_530,In_713);
and U1168 (N_1168,In_63,In_543);
nand U1169 (N_1169,In_570,In_639);
xnor U1170 (N_1170,In_931,In_607);
nand U1171 (N_1171,In_167,In_183);
nand U1172 (N_1172,In_12,In_975);
nor U1173 (N_1173,In_870,In_593);
nor U1174 (N_1174,In_903,In_479);
and U1175 (N_1175,In_728,In_940);
nor U1176 (N_1176,In_805,In_122);
xnor U1177 (N_1177,In_527,In_828);
or U1178 (N_1178,In_243,In_773);
nand U1179 (N_1179,In_298,In_916);
and U1180 (N_1180,In_578,In_77);
and U1181 (N_1181,In_443,In_75);
and U1182 (N_1182,In_25,In_852);
xor U1183 (N_1183,In_609,In_828);
and U1184 (N_1184,In_674,In_67);
xor U1185 (N_1185,In_637,In_796);
nand U1186 (N_1186,In_72,In_719);
or U1187 (N_1187,In_629,In_692);
nand U1188 (N_1188,In_346,In_953);
or U1189 (N_1189,In_912,In_162);
and U1190 (N_1190,In_809,In_520);
nand U1191 (N_1191,In_583,In_777);
or U1192 (N_1192,In_641,In_951);
and U1193 (N_1193,In_308,In_759);
nand U1194 (N_1194,In_344,In_27);
and U1195 (N_1195,In_288,In_716);
nand U1196 (N_1196,In_84,In_41);
or U1197 (N_1197,In_253,In_324);
and U1198 (N_1198,In_293,In_951);
and U1199 (N_1199,In_941,In_648);
nand U1200 (N_1200,In_390,In_229);
xor U1201 (N_1201,In_412,In_622);
or U1202 (N_1202,In_702,In_974);
xnor U1203 (N_1203,In_299,In_278);
nand U1204 (N_1204,In_163,In_591);
nor U1205 (N_1205,In_556,In_226);
xnor U1206 (N_1206,In_274,In_27);
nor U1207 (N_1207,In_296,In_181);
nand U1208 (N_1208,In_441,In_437);
nand U1209 (N_1209,In_569,In_675);
and U1210 (N_1210,In_625,In_997);
xnor U1211 (N_1211,In_649,In_904);
nor U1212 (N_1212,In_615,In_726);
nor U1213 (N_1213,In_526,In_879);
nor U1214 (N_1214,In_688,In_444);
nand U1215 (N_1215,In_252,In_374);
xor U1216 (N_1216,In_834,In_68);
nor U1217 (N_1217,In_9,In_937);
and U1218 (N_1218,In_884,In_346);
and U1219 (N_1219,In_8,In_436);
xnor U1220 (N_1220,In_877,In_372);
or U1221 (N_1221,In_985,In_909);
nor U1222 (N_1222,In_424,In_354);
xnor U1223 (N_1223,In_331,In_2);
nand U1224 (N_1224,In_604,In_192);
nand U1225 (N_1225,In_745,In_402);
xnor U1226 (N_1226,In_849,In_243);
or U1227 (N_1227,In_774,In_696);
and U1228 (N_1228,In_919,In_366);
or U1229 (N_1229,In_541,In_401);
or U1230 (N_1230,In_533,In_938);
and U1231 (N_1231,In_145,In_238);
xor U1232 (N_1232,In_266,In_538);
and U1233 (N_1233,In_779,In_250);
or U1234 (N_1234,In_713,In_235);
or U1235 (N_1235,In_774,In_640);
and U1236 (N_1236,In_404,In_523);
nand U1237 (N_1237,In_150,In_932);
and U1238 (N_1238,In_307,In_340);
nand U1239 (N_1239,In_451,In_412);
nor U1240 (N_1240,In_244,In_421);
nand U1241 (N_1241,In_907,In_366);
or U1242 (N_1242,In_981,In_742);
nand U1243 (N_1243,In_874,In_545);
xor U1244 (N_1244,In_260,In_952);
nand U1245 (N_1245,In_277,In_175);
nand U1246 (N_1246,In_995,In_132);
and U1247 (N_1247,In_998,In_584);
nor U1248 (N_1248,In_525,In_518);
nand U1249 (N_1249,In_347,In_168);
or U1250 (N_1250,In_758,In_887);
and U1251 (N_1251,In_934,In_863);
or U1252 (N_1252,In_248,In_463);
xor U1253 (N_1253,In_720,In_826);
nand U1254 (N_1254,In_841,In_96);
and U1255 (N_1255,In_47,In_597);
nor U1256 (N_1256,In_93,In_693);
and U1257 (N_1257,In_315,In_622);
nand U1258 (N_1258,In_273,In_105);
nand U1259 (N_1259,In_422,In_162);
xor U1260 (N_1260,In_244,In_948);
nand U1261 (N_1261,In_899,In_963);
nor U1262 (N_1262,In_283,In_853);
nor U1263 (N_1263,In_997,In_448);
and U1264 (N_1264,In_96,In_163);
nand U1265 (N_1265,In_377,In_81);
nand U1266 (N_1266,In_119,In_743);
xor U1267 (N_1267,In_752,In_241);
and U1268 (N_1268,In_222,In_5);
and U1269 (N_1269,In_572,In_146);
or U1270 (N_1270,In_772,In_679);
nand U1271 (N_1271,In_130,In_822);
nor U1272 (N_1272,In_18,In_12);
and U1273 (N_1273,In_791,In_705);
nor U1274 (N_1274,In_464,In_804);
or U1275 (N_1275,In_646,In_566);
xnor U1276 (N_1276,In_894,In_944);
nand U1277 (N_1277,In_318,In_888);
or U1278 (N_1278,In_985,In_300);
nor U1279 (N_1279,In_580,In_745);
nor U1280 (N_1280,In_548,In_728);
nor U1281 (N_1281,In_6,In_388);
or U1282 (N_1282,In_31,In_846);
nand U1283 (N_1283,In_291,In_272);
nand U1284 (N_1284,In_232,In_839);
nand U1285 (N_1285,In_737,In_306);
or U1286 (N_1286,In_99,In_717);
or U1287 (N_1287,In_636,In_870);
or U1288 (N_1288,In_569,In_674);
or U1289 (N_1289,In_168,In_12);
or U1290 (N_1290,In_68,In_575);
xnor U1291 (N_1291,In_564,In_444);
nand U1292 (N_1292,In_96,In_579);
xor U1293 (N_1293,In_88,In_505);
nor U1294 (N_1294,In_434,In_83);
nor U1295 (N_1295,In_452,In_886);
nand U1296 (N_1296,In_103,In_237);
nor U1297 (N_1297,In_121,In_458);
or U1298 (N_1298,In_38,In_392);
nand U1299 (N_1299,In_650,In_514);
or U1300 (N_1300,In_672,In_757);
and U1301 (N_1301,In_561,In_402);
or U1302 (N_1302,In_397,In_976);
xnor U1303 (N_1303,In_686,In_440);
nor U1304 (N_1304,In_113,In_157);
nand U1305 (N_1305,In_974,In_580);
nand U1306 (N_1306,In_680,In_146);
nand U1307 (N_1307,In_502,In_694);
and U1308 (N_1308,In_727,In_2);
or U1309 (N_1309,In_611,In_433);
nand U1310 (N_1310,In_992,In_38);
nand U1311 (N_1311,In_309,In_210);
xnor U1312 (N_1312,In_157,In_309);
or U1313 (N_1313,In_97,In_283);
nor U1314 (N_1314,In_783,In_292);
and U1315 (N_1315,In_544,In_343);
and U1316 (N_1316,In_795,In_130);
nor U1317 (N_1317,In_501,In_47);
and U1318 (N_1318,In_595,In_382);
nor U1319 (N_1319,In_419,In_760);
or U1320 (N_1320,In_879,In_485);
xor U1321 (N_1321,In_314,In_783);
and U1322 (N_1322,In_57,In_239);
or U1323 (N_1323,In_205,In_138);
and U1324 (N_1324,In_653,In_534);
nand U1325 (N_1325,In_838,In_687);
or U1326 (N_1326,In_752,In_630);
nor U1327 (N_1327,In_771,In_769);
or U1328 (N_1328,In_698,In_689);
or U1329 (N_1329,In_604,In_645);
nand U1330 (N_1330,In_827,In_201);
and U1331 (N_1331,In_304,In_808);
or U1332 (N_1332,In_160,In_521);
nor U1333 (N_1333,In_365,In_234);
and U1334 (N_1334,In_742,In_335);
nand U1335 (N_1335,In_575,In_807);
nor U1336 (N_1336,In_720,In_148);
and U1337 (N_1337,In_127,In_762);
nand U1338 (N_1338,In_705,In_471);
and U1339 (N_1339,In_315,In_528);
nand U1340 (N_1340,In_288,In_221);
or U1341 (N_1341,In_91,In_331);
nand U1342 (N_1342,In_347,In_760);
nor U1343 (N_1343,In_791,In_641);
nand U1344 (N_1344,In_284,In_854);
nand U1345 (N_1345,In_385,In_703);
and U1346 (N_1346,In_16,In_578);
nand U1347 (N_1347,In_351,In_86);
and U1348 (N_1348,In_825,In_666);
nor U1349 (N_1349,In_816,In_761);
or U1350 (N_1350,In_453,In_617);
and U1351 (N_1351,In_424,In_774);
nor U1352 (N_1352,In_843,In_937);
nand U1353 (N_1353,In_840,In_855);
xnor U1354 (N_1354,In_657,In_404);
xor U1355 (N_1355,In_207,In_59);
nor U1356 (N_1356,In_523,In_700);
and U1357 (N_1357,In_340,In_42);
nand U1358 (N_1358,In_99,In_340);
nor U1359 (N_1359,In_813,In_685);
nor U1360 (N_1360,In_985,In_754);
or U1361 (N_1361,In_932,In_275);
and U1362 (N_1362,In_422,In_384);
or U1363 (N_1363,In_80,In_391);
nor U1364 (N_1364,In_368,In_480);
and U1365 (N_1365,In_324,In_511);
and U1366 (N_1366,In_675,In_489);
and U1367 (N_1367,In_249,In_395);
and U1368 (N_1368,In_896,In_641);
nor U1369 (N_1369,In_570,In_206);
nor U1370 (N_1370,In_909,In_135);
nand U1371 (N_1371,In_498,In_534);
xor U1372 (N_1372,In_182,In_399);
nor U1373 (N_1373,In_838,In_891);
or U1374 (N_1374,In_265,In_872);
nand U1375 (N_1375,In_580,In_698);
and U1376 (N_1376,In_497,In_915);
nand U1377 (N_1377,In_880,In_272);
or U1378 (N_1378,In_574,In_104);
nor U1379 (N_1379,In_287,In_588);
or U1380 (N_1380,In_434,In_159);
nand U1381 (N_1381,In_896,In_178);
or U1382 (N_1382,In_708,In_544);
nor U1383 (N_1383,In_691,In_52);
nand U1384 (N_1384,In_656,In_799);
or U1385 (N_1385,In_884,In_700);
or U1386 (N_1386,In_274,In_74);
nand U1387 (N_1387,In_839,In_622);
xor U1388 (N_1388,In_254,In_530);
nand U1389 (N_1389,In_968,In_874);
and U1390 (N_1390,In_751,In_747);
nor U1391 (N_1391,In_283,In_683);
nor U1392 (N_1392,In_151,In_780);
nor U1393 (N_1393,In_514,In_105);
nand U1394 (N_1394,In_965,In_420);
xor U1395 (N_1395,In_567,In_910);
and U1396 (N_1396,In_76,In_752);
nand U1397 (N_1397,In_411,In_408);
and U1398 (N_1398,In_227,In_18);
nand U1399 (N_1399,In_478,In_908);
xor U1400 (N_1400,In_250,In_975);
nor U1401 (N_1401,In_96,In_816);
nand U1402 (N_1402,In_403,In_470);
and U1403 (N_1403,In_104,In_828);
or U1404 (N_1404,In_147,In_275);
or U1405 (N_1405,In_403,In_533);
nand U1406 (N_1406,In_947,In_268);
nor U1407 (N_1407,In_864,In_155);
or U1408 (N_1408,In_714,In_961);
xnor U1409 (N_1409,In_84,In_967);
nor U1410 (N_1410,In_218,In_387);
nor U1411 (N_1411,In_673,In_356);
nor U1412 (N_1412,In_329,In_364);
or U1413 (N_1413,In_744,In_626);
nand U1414 (N_1414,In_948,In_306);
nand U1415 (N_1415,In_963,In_876);
or U1416 (N_1416,In_706,In_426);
or U1417 (N_1417,In_589,In_911);
nor U1418 (N_1418,In_699,In_408);
nor U1419 (N_1419,In_34,In_270);
nand U1420 (N_1420,In_920,In_89);
xnor U1421 (N_1421,In_409,In_371);
or U1422 (N_1422,In_938,In_541);
or U1423 (N_1423,In_840,In_145);
nand U1424 (N_1424,In_755,In_903);
or U1425 (N_1425,In_665,In_293);
nand U1426 (N_1426,In_460,In_163);
nand U1427 (N_1427,In_460,In_87);
and U1428 (N_1428,In_794,In_844);
nor U1429 (N_1429,In_419,In_613);
nand U1430 (N_1430,In_928,In_981);
and U1431 (N_1431,In_522,In_914);
or U1432 (N_1432,In_41,In_68);
and U1433 (N_1433,In_972,In_338);
and U1434 (N_1434,In_798,In_287);
and U1435 (N_1435,In_673,In_485);
or U1436 (N_1436,In_758,In_74);
xor U1437 (N_1437,In_303,In_426);
or U1438 (N_1438,In_432,In_602);
or U1439 (N_1439,In_314,In_553);
or U1440 (N_1440,In_867,In_273);
nor U1441 (N_1441,In_965,In_818);
or U1442 (N_1442,In_284,In_338);
nor U1443 (N_1443,In_939,In_539);
nor U1444 (N_1444,In_671,In_522);
xor U1445 (N_1445,In_243,In_780);
nor U1446 (N_1446,In_124,In_114);
and U1447 (N_1447,In_149,In_418);
nor U1448 (N_1448,In_853,In_130);
and U1449 (N_1449,In_773,In_813);
or U1450 (N_1450,In_522,In_42);
xnor U1451 (N_1451,In_901,In_449);
xnor U1452 (N_1452,In_806,In_803);
nand U1453 (N_1453,In_916,In_469);
xor U1454 (N_1454,In_201,In_499);
nand U1455 (N_1455,In_640,In_929);
and U1456 (N_1456,In_697,In_593);
nor U1457 (N_1457,In_414,In_168);
and U1458 (N_1458,In_57,In_85);
and U1459 (N_1459,In_928,In_478);
nor U1460 (N_1460,In_909,In_518);
or U1461 (N_1461,In_887,In_438);
xor U1462 (N_1462,In_586,In_737);
xnor U1463 (N_1463,In_483,In_245);
and U1464 (N_1464,In_588,In_550);
nand U1465 (N_1465,In_603,In_847);
nor U1466 (N_1466,In_522,In_792);
or U1467 (N_1467,In_30,In_968);
nand U1468 (N_1468,In_398,In_649);
and U1469 (N_1469,In_141,In_710);
or U1470 (N_1470,In_592,In_946);
nor U1471 (N_1471,In_101,In_946);
and U1472 (N_1472,In_757,In_799);
nand U1473 (N_1473,In_939,In_304);
nor U1474 (N_1474,In_816,In_624);
or U1475 (N_1475,In_630,In_35);
nor U1476 (N_1476,In_158,In_716);
or U1477 (N_1477,In_460,In_593);
nand U1478 (N_1478,In_604,In_390);
or U1479 (N_1479,In_841,In_45);
nor U1480 (N_1480,In_960,In_347);
nand U1481 (N_1481,In_796,In_332);
and U1482 (N_1482,In_27,In_11);
nand U1483 (N_1483,In_384,In_988);
nor U1484 (N_1484,In_213,In_279);
nor U1485 (N_1485,In_626,In_348);
xnor U1486 (N_1486,In_960,In_403);
or U1487 (N_1487,In_15,In_565);
nand U1488 (N_1488,In_845,In_180);
and U1489 (N_1489,In_557,In_397);
xor U1490 (N_1490,In_853,In_145);
xnor U1491 (N_1491,In_354,In_840);
and U1492 (N_1492,In_710,In_609);
nand U1493 (N_1493,In_413,In_434);
and U1494 (N_1494,In_4,In_739);
and U1495 (N_1495,In_682,In_229);
xnor U1496 (N_1496,In_145,In_279);
xnor U1497 (N_1497,In_425,In_700);
nor U1498 (N_1498,In_741,In_992);
and U1499 (N_1499,In_989,In_964);
and U1500 (N_1500,In_556,In_487);
nand U1501 (N_1501,In_292,In_73);
nand U1502 (N_1502,In_720,In_711);
or U1503 (N_1503,In_617,In_352);
and U1504 (N_1504,In_392,In_645);
and U1505 (N_1505,In_598,In_904);
or U1506 (N_1506,In_352,In_780);
or U1507 (N_1507,In_474,In_780);
and U1508 (N_1508,In_110,In_484);
or U1509 (N_1509,In_32,In_439);
nor U1510 (N_1510,In_996,In_816);
nand U1511 (N_1511,In_265,In_20);
or U1512 (N_1512,In_821,In_512);
nand U1513 (N_1513,In_84,In_962);
and U1514 (N_1514,In_919,In_727);
nand U1515 (N_1515,In_662,In_525);
and U1516 (N_1516,In_624,In_55);
or U1517 (N_1517,In_494,In_537);
nand U1518 (N_1518,In_273,In_717);
nand U1519 (N_1519,In_367,In_645);
nand U1520 (N_1520,In_803,In_644);
nand U1521 (N_1521,In_728,In_751);
and U1522 (N_1522,In_652,In_710);
nand U1523 (N_1523,In_67,In_945);
nor U1524 (N_1524,In_414,In_338);
nand U1525 (N_1525,In_534,In_667);
nand U1526 (N_1526,In_570,In_10);
and U1527 (N_1527,In_886,In_998);
or U1528 (N_1528,In_540,In_973);
nand U1529 (N_1529,In_19,In_698);
nand U1530 (N_1530,In_623,In_605);
or U1531 (N_1531,In_488,In_757);
or U1532 (N_1532,In_958,In_549);
nand U1533 (N_1533,In_626,In_975);
nor U1534 (N_1534,In_921,In_557);
nand U1535 (N_1535,In_225,In_379);
and U1536 (N_1536,In_463,In_278);
nor U1537 (N_1537,In_974,In_109);
or U1538 (N_1538,In_491,In_604);
or U1539 (N_1539,In_856,In_169);
nand U1540 (N_1540,In_515,In_495);
and U1541 (N_1541,In_824,In_773);
and U1542 (N_1542,In_619,In_550);
or U1543 (N_1543,In_414,In_46);
or U1544 (N_1544,In_445,In_690);
or U1545 (N_1545,In_811,In_207);
and U1546 (N_1546,In_638,In_726);
or U1547 (N_1547,In_431,In_173);
and U1548 (N_1548,In_303,In_672);
and U1549 (N_1549,In_272,In_423);
nor U1550 (N_1550,In_547,In_17);
xor U1551 (N_1551,In_109,In_475);
and U1552 (N_1552,In_56,In_334);
xnor U1553 (N_1553,In_253,In_49);
and U1554 (N_1554,In_863,In_115);
and U1555 (N_1555,In_654,In_539);
or U1556 (N_1556,In_150,In_608);
xnor U1557 (N_1557,In_803,In_426);
nand U1558 (N_1558,In_335,In_72);
or U1559 (N_1559,In_724,In_968);
xor U1560 (N_1560,In_262,In_989);
and U1561 (N_1561,In_72,In_110);
nor U1562 (N_1562,In_757,In_287);
nor U1563 (N_1563,In_239,In_512);
and U1564 (N_1564,In_2,In_157);
or U1565 (N_1565,In_499,In_650);
and U1566 (N_1566,In_785,In_860);
or U1567 (N_1567,In_589,In_569);
or U1568 (N_1568,In_527,In_671);
and U1569 (N_1569,In_417,In_906);
and U1570 (N_1570,In_56,In_31);
or U1571 (N_1571,In_966,In_801);
or U1572 (N_1572,In_919,In_69);
or U1573 (N_1573,In_341,In_450);
nor U1574 (N_1574,In_360,In_944);
or U1575 (N_1575,In_25,In_73);
and U1576 (N_1576,In_890,In_728);
nor U1577 (N_1577,In_262,In_425);
nand U1578 (N_1578,In_587,In_85);
or U1579 (N_1579,In_659,In_354);
and U1580 (N_1580,In_220,In_818);
xnor U1581 (N_1581,In_959,In_708);
or U1582 (N_1582,In_17,In_733);
nand U1583 (N_1583,In_615,In_805);
or U1584 (N_1584,In_997,In_560);
and U1585 (N_1585,In_679,In_136);
xor U1586 (N_1586,In_694,In_86);
and U1587 (N_1587,In_491,In_355);
nor U1588 (N_1588,In_161,In_193);
and U1589 (N_1589,In_797,In_879);
nand U1590 (N_1590,In_604,In_567);
nand U1591 (N_1591,In_429,In_690);
xnor U1592 (N_1592,In_504,In_947);
nor U1593 (N_1593,In_711,In_434);
and U1594 (N_1594,In_867,In_627);
and U1595 (N_1595,In_818,In_577);
or U1596 (N_1596,In_935,In_973);
nand U1597 (N_1597,In_404,In_612);
and U1598 (N_1598,In_246,In_163);
or U1599 (N_1599,In_23,In_877);
nor U1600 (N_1600,In_404,In_446);
and U1601 (N_1601,In_938,In_768);
and U1602 (N_1602,In_122,In_976);
or U1603 (N_1603,In_251,In_626);
nand U1604 (N_1604,In_796,In_93);
or U1605 (N_1605,In_520,In_773);
xor U1606 (N_1606,In_3,In_581);
and U1607 (N_1607,In_154,In_237);
nand U1608 (N_1608,In_672,In_563);
or U1609 (N_1609,In_556,In_667);
and U1610 (N_1610,In_527,In_657);
nand U1611 (N_1611,In_738,In_674);
or U1612 (N_1612,In_644,In_934);
or U1613 (N_1613,In_616,In_570);
and U1614 (N_1614,In_820,In_344);
and U1615 (N_1615,In_237,In_478);
nand U1616 (N_1616,In_230,In_212);
nand U1617 (N_1617,In_241,In_394);
xnor U1618 (N_1618,In_502,In_421);
and U1619 (N_1619,In_80,In_632);
nor U1620 (N_1620,In_176,In_794);
xnor U1621 (N_1621,In_556,In_904);
and U1622 (N_1622,In_968,In_514);
or U1623 (N_1623,In_623,In_200);
and U1624 (N_1624,In_765,In_957);
nand U1625 (N_1625,In_741,In_42);
nor U1626 (N_1626,In_651,In_653);
or U1627 (N_1627,In_524,In_576);
or U1628 (N_1628,In_969,In_205);
or U1629 (N_1629,In_519,In_235);
or U1630 (N_1630,In_727,In_445);
and U1631 (N_1631,In_190,In_83);
and U1632 (N_1632,In_292,In_34);
or U1633 (N_1633,In_614,In_809);
nand U1634 (N_1634,In_511,In_596);
or U1635 (N_1635,In_880,In_879);
nor U1636 (N_1636,In_34,In_37);
or U1637 (N_1637,In_223,In_71);
nor U1638 (N_1638,In_229,In_552);
and U1639 (N_1639,In_231,In_228);
nand U1640 (N_1640,In_212,In_412);
or U1641 (N_1641,In_58,In_218);
nor U1642 (N_1642,In_534,In_704);
or U1643 (N_1643,In_660,In_816);
nand U1644 (N_1644,In_438,In_40);
nand U1645 (N_1645,In_417,In_22);
and U1646 (N_1646,In_284,In_983);
nand U1647 (N_1647,In_719,In_448);
xnor U1648 (N_1648,In_994,In_162);
nor U1649 (N_1649,In_684,In_447);
xor U1650 (N_1650,In_238,In_400);
xnor U1651 (N_1651,In_315,In_107);
or U1652 (N_1652,In_346,In_601);
or U1653 (N_1653,In_11,In_936);
nand U1654 (N_1654,In_735,In_925);
nor U1655 (N_1655,In_487,In_494);
or U1656 (N_1656,In_824,In_39);
nand U1657 (N_1657,In_379,In_566);
or U1658 (N_1658,In_78,In_948);
or U1659 (N_1659,In_26,In_104);
nand U1660 (N_1660,In_373,In_933);
or U1661 (N_1661,In_888,In_864);
nand U1662 (N_1662,In_876,In_156);
or U1663 (N_1663,In_271,In_987);
nand U1664 (N_1664,In_692,In_957);
and U1665 (N_1665,In_708,In_929);
nand U1666 (N_1666,In_408,In_768);
nor U1667 (N_1667,In_505,In_113);
nand U1668 (N_1668,In_738,In_704);
or U1669 (N_1669,In_646,In_193);
or U1670 (N_1670,In_687,In_237);
nor U1671 (N_1671,In_760,In_56);
and U1672 (N_1672,In_232,In_249);
or U1673 (N_1673,In_195,In_829);
nand U1674 (N_1674,In_125,In_551);
nand U1675 (N_1675,In_190,In_692);
nand U1676 (N_1676,In_485,In_759);
nand U1677 (N_1677,In_374,In_201);
nand U1678 (N_1678,In_320,In_105);
xnor U1679 (N_1679,In_277,In_987);
or U1680 (N_1680,In_588,In_385);
or U1681 (N_1681,In_845,In_776);
nand U1682 (N_1682,In_789,In_152);
or U1683 (N_1683,In_809,In_776);
and U1684 (N_1684,In_771,In_656);
or U1685 (N_1685,In_851,In_306);
nor U1686 (N_1686,In_875,In_835);
or U1687 (N_1687,In_772,In_394);
or U1688 (N_1688,In_731,In_856);
and U1689 (N_1689,In_95,In_685);
or U1690 (N_1690,In_91,In_374);
nor U1691 (N_1691,In_180,In_99);
or U1692 (N_1692,In_69,In_863);
nor U1693 (N_1693,In_143,In_530);
or U1694 (N_1694,In_710,In_713);
and U1695 (N_1695,In_972,In_198);
and U1696 (N_1696,In_170,In_877);
nor U1697 (N_1697,In_170,In_134);
nor U1698 (N_1698,In_485,In_224);
or U1699 (N_1699,In_994,In_300);
and U1700 (N_1700,In_92,In_70);
nand U1701 (N_1701,In_4,In_750);
nor U1702 (N_1702,In_739,In_736);
nor U1703 (N_1703,In_659,In_683);
xor U1704 (N_1704,In_768,In_329);
nand U1705 (N_1705,In_871,In_485);
or U1706 (N_1706,In_673,In_489);
and U1707 (N_1707,In_400,In_191);
nor U1708 (N_1708,In_705,In_629);
and U1709 (N_1709,In_367,In_642);
or U1710 (N_1710,In_375,In_169);
or U1711 (N_1711,In_420,In_410);
or U1712 (N_1712,In_743,In_570);
nand U1713 (N_1713,In_88,In_565);
nand U1714 (N_1714,In_455,In_850);
and U1715 (N_1715,In_213,In_365);
and U1716 (N_1716,In_127,In_995);
or U1717 (N_1717,In_275,In_250);
nand U1718 (N_1718,In_935,In_695);
nand U1719 (N_1719,In_247,In_95);
xnor U1720 (N_1720,In_442,In_658);
and U1721 (N_1721,In_985,In_698);
nand U1722 (N_1722,In_810,In_93);
nand U1723 (N_1723,In_296,In_427);
nand U1724 (N_1724,In_636,In_300);
nand U1725 (N_1725,In_252,In_15);
nor U1726 (N_1726,In_255,In_626);
nor U1727 (N_1727,In_747,In_138);
nand U1728 (N_1728,In_984,In_741);
and U1729 (N_1729,In_615,In_927);
or U1730 (N_1730,In_374,In_60);
or U1731 (N_1731,In_817,In_959);
nand U1732 (N_1732,In_915,In_421);
or U1733 (N_1733,In_781,In_832);
nand U1734 (N_1734,In_825,In_331);
and U1735 (N_1735,In_709,In_60);
nand U1736 (N_1736,In_946,In_153);
or U1737 (N_1737,In_958,In_510);
or U1738 (N_1738,In_159,In_824);
nor U1739 (N_1739,In_58,In_489);
and U1740 (N_1740,In_564,In_40);
and U1741 (N_1741,In_824,In_723);
or U1742 (N_1742,In_831,In_505);
and U1743 (N_1743,In_217,In_6);
xnor U1744 (N_1744,In_252,In_922);
nand U1745 (N_1745,In_973,In_316);
nand U1746 (N_1746,In_958,In_112);
nand U1747 (N_1747,In_190,In_625);
and U1748 (N_1748,In_150,In_352);
nor U1749 (N_1749,In_384,In_169);
nor U1750 (N_1750,In_246,In_11);
and U1751 (N_1751,In_513,In_992);
xor U1752 (N_1752,In_32,In_135);
nor U1753 (N_1753,In_664,In_869);
and U1754 (N_1754,In_459,In_619);
nor U1755 (N_1755,In_104,In_135);
nand U1756 (N_1756,In_583,In_971);
nand U1757 (N_1757,In_814,In_150);
nand U1758 (N_1758,In_252,In_530);
or U1759 (N_1759,In_576,In_370);
nand U1760 (N_1760,In_322,In_720);
nor U1761 (N_1761,In_285,In_561);
nor U1762 (N_1762,In_604,In_568);
or U1763 (N_1763,In_602,In_314);
nand U1764 (N_1764,In_170,In_445);
or U1765 (N_1765,In_831,In_704);
or U1766 (N_1766,In_89,In_313);
nor U1767 (N_1767,In_852,In_309);
and U1768 (N_1768,In_4,In_773);
or U1769 (N_1769,In_399,In_339);
or U1770 (N_1770,In_344,In_50);
nand U1771 (N_1771,In_888,In_919);
or U1772 (N_1772,In_20,In_951);
nand U1773 (N_1773,In_258,In_106);
nor U1774 (N_1774,In_567,In_476);
nor U1775 (N_1775,In_815,In_250);
or U1776 (N_1776,In_251,In_908);
or U1777 (N_1777,In_515,In_719);
nand U1778 (N_1778,In_51,In_402);
nand U1779 (N_1779,In_219,In_669);
and U1780 (N_1780,In_216,In_259);
nand U1781 (N_1781,In_881,In_751);
and U1782 (N_1782,In_664,In_476);
nand U1783 (N_1783,In_639,In_927);
nand U1784 (N_1784,In_971,In_530);
and U1785 (N_1785,In_132,In_999);
and U1786 (N_1786,In_532,In_140);
nand U1787 (N_1787,In_510,In_227);
xnor U1788 (N_1788,In_772,In_628);
nand U1789 (N_1789,In_403,In_352);
nand U1790 (N_1790,In_750,In_403);
nor U1791 (N_1791,In_983,In_975);
nand U1792 (N_1792,In_517,In_729);
and U1793 (N_1793,In_928,In_831);
nor U1794 (N_1794,In_6,In_27);
nor U1795 (N_1795,In_539,In_308);
xor U1796 (N_1796,In_554,In_176);
nand U1797 (N_1797,In_77,In_19);
or U1798 (N_1798,In_342,In_675);
and U1799 (N_1799,In_1,In_403);
or U1800 (N_1800,In_17,In_459);
nand U1801 (N_1801,In_585,In_36);
nor U1802 (N_1802,In_487,In_101);
nand U1803 (N_1803,In_946,In_179);
xnor U1804 (N_1804,In_162,In_594);
nand U1805 (N_1805,In_968,In_31);
nand U1806 (N_1806,In_913,In_178);
xor U1807 (N_1807,In_736,In_407);
and U1808 (N_1808,In_579,In_206);
nor U1809 (N_1809,In_808,In_935);
nor U1810 (N_1810,In_342,In_679);
or U1811 (N_1811,In_830,In_825);
and U1812 (N_1812,In_502,In_697);
and U1813 (N_1813,In_109,In_949);
nand U1814 (N_1814,In_457,In_884);
or U1815 (N_1815,In_680,In_806);
nor U1816 (N_1816,In_774,In_919);
and U1817 (N_1817,In_678,In_933);
or U1818 (N_1818,In_511,In_275);
or U1819 (N_1819,In_591,In_596);
and U1820 (N_1820,In_453,In_270);
and U1821 (N_1821,In_6,In_495);
or U1822 (N_1822,In_449,In_920);
or U1823 (N_1823,In_840,In_954);
nor U1824 (N_1824,In_382,In_789);
nor U1825 (N_1825,In_247,In_692);
and U1826 (N_1826,In_558,In_38);
nand U1827 (N_1827,In_186,In_752);
nand U1828 (N_1828,In_64,In_688);
or U1829 (N_1829,In_102,In_732);
and U1830 (N_1830,In_547,In_173);
nand U1831 (N_1831,In_849,In_13);
and U1832 (N_1832,In_294,In_810);
and U1833 (N_1833,In_379,In_372);
or U1834 (N_1834,In_155,In_993);
nor U1835 (N_1835,In_740,In_26);
and U1836 (N_1836,In_733,In_945);
or U1837 (N_1837,In_625,In_368);
or U1838 (N_1838,In_574,In_7);
or U1839 (N_1839,In_575,In_439);
xnor U1840 (N_1840,In_123,In_507);
nand U1841 (N_1841,In_981,In_66);
nand U1842 (N_1842,In_687,In_487);
nand U1843 (N_1843,In_373,In_372);
or U1844 (N_1844,In_680,In_338);
nor U1845 (N_1845,In_758,In_295);
nor U1846 (N_1846,In_163,In_130);
and U1847 (N_1847,In_792,In_152);
or U1848 (N_1848,In_626,In_716);
or U1849 (N_1849,In_625,In_443);
and U1850 (N_1850,In_902,In_212);
nor U1851 (N_1851,In_313,In_350);
nor U1852 (N_1852,In_107,In_269);
or U1853 (N_1853,In_215,In_163);
nor U1854 (N_1854,In_460,In_619);
and U1855 (N_1855,In_997,In_937);
nand U1856 (N_1856,In_271,In_334);
nor U1857 (N_1857,In_59,In_45);
or U1858 (N_1858,In_822,In_652);
nor U1859 (N_1859,In_288,In_304);
and U1860 (N_1860,In_417,In_508);
nor U1861 (N_1861,In_20,In_454);
nor U1862 (N_1862,In_193,In_918);
and U1863 (N_1863,In_175,In_31);
and U1864 (N_1864,In_365,In_494);
nand U1865 (N_1865,In_200,In_211);
nand U1866 (N_1866,In_396,In_253);
and U1867 (N_1867,In_387,In_266);
and U1868 (N_1868,In_445,In_166);
xnor U1869 (N_1869,In_285,In_726);
nand U1870 (N_1870,In_769,In_100);
or U1871 (N_1871,In_298,In_706);
and U1872 (N_1872,In_78,In_210);
or U1873 (N_1873,In_431,In_520);
and U1874 (N_1874,In_963,In_951);
nor U1875 (N_1875,In_536,In_437);
nand U1876 (N_1876,In_364,In_293);
nor U1877 (N_1877,In_253,In_328);
nor U1878 (N_1878,In_630,In_966);
and U1879 (N_1879,In_186,In_934);
or U1880 (N_1880,In_34,In_742);
or U1881 (N_1881,In_400,In_677);
nor U1882 (N_1882,In_232,In_409);
nor U1883 (N_1883,In_619,In_970);
nor U1884 (N_1884,In_226,In_657);
nor U1885 (N_1885,In_173,In_751);
or U1886 (N_1886,In_365,In_384);
and U1887 (N_1887,In_267,In_349);
nor U1888 (N_1888,In_906,In_814);
xnor U1889 (N_1889,In_353,In_297);
and U1890 (N_1890,In_951,In_864);
or U1891 (N_1891,In_344,In_922);
nand U1892 (N_1892,In_411,In_469);
nand U1893 (N_1893,In_864,In_381);
nand U1894 (N_1894,In_651,In_816);
nor U1895 (N_1895,In_62,In_904);
nor U1896 (N_1896,In_715,In_501);
nand U1897 (N_1897,In_27,In_560);
nor U1898 (N_1898,In_417,In_144);
nand U1899 (N_1899,In_928,In_482);
nand U1900 (N_1900,In_437,In_750);
and U1901 (N_1901,In_978,In_967);
nor U1902 (N_1902,In_334,In_554);
and U1903 (N_1903,In_325,In_188);
nand U1904 (N_1904,In_799,In_722);
nand U1905 (N_1905,In_917,In_426);
or U1906 (N_1906,In_237,In_320);
nand U1907 (N_1907,In_460,In_907);
nand U1908 (N_1908,In_815,In_134);
or U1909 (N_1909,In_461,In_644);
and U1910 (N_1910,In_556,In_305);
xnor U1911 (N_1911,In_56,In_130);
or U1912 (N_1912,In_920,In_318);
nor U1913 (N_1913,In_156,In_99);
nand U1914 (N_1914,In_629,In_725);
and U1915 (N_1915,In_77,In_598);
nand U1916 (N_1916,In_44,In_154);
nor U1917 (N_1917,In_639,In_856);
or U1918 (N_1918,In_397,In_369);
and U1919 (N_1919,In_376,In_329);
or U1920 (N_1920,In_615,In_733);
xor U1921 (N_1921,In_267,In_542);
and U1922 (N_1922,In_601,In_337);
xor U1923 (N_1923,In_810,In_387);
and U1924 (N_1924,In_567,In_807);
nor U1925 (N_1925,In_627,In_738);
nand U1926 (N_1926,In_233,In_531);
xnor U1927 (N_1927,In_229,In_592);
and U1928 (N_1928,In_894,In_714);
and U1929 (N_1929,In_493,In_825);
nand U1930 (N_1930,In_965,In_440);
and U1931 (N_1931,In_770,In_5);
xor U1932 (N_1932,In_0,In_494);
xnor U1933 (N_1933,In_96,In_36);
nand U1934 (N_1934,In_134,In_644);
and U1935 (N_1935,In_145,In_893);
nor U1936 (N_1936,In_447,In_415);
and U1937 (N_1937,In_920,In_610);
nand U1938 (N_1938,In_361,In_219);
nor U1939 (N_1939,In_908,In_120);
and U1940 (N_1940,In_509,In_583);
nand U1941 (N_1941,In_721,In_138);
nor U1942 (N_1942,In_540,In_132);
and U1943 (N_1943,In_908,In_879);
and U1944 (N_1944,In_425,In_868);
nand U1945 (N_1945,In_740,In_695);
or U1946 (N_1946,In_537,In_677);
nand U1947 (N_1947,In_705,In_618);
and U1948 (N_1948,In_821,In_621);
and U1949 (N_1949,In_516,In_736);
xnor U1950 (N_1950,In_233,In_731);
and U1951 (N_1951,In_349,In_521);
nand U1952 (N_1952,In_957,In_850);
nor U1953 (N_1953,In_820,In_355);
and U1954 (N_1954,In_595,In_889);
or U1955 (N_1955,In_425,In_295);
xor U1956 (N_1956,In_158,In_78);
nor U1957 (N_1957,In_686,In_187);
or U1958 (N_1958,In_138,In_873);
xnor U1959 (N_1959,In_759,In_279);
xor U1960 (N_1960,In_899,In_929);
xnor U1961 (N_1961,In_535,In_982);
nand U1962 (N_1962,In_68,In_944);
nor U1963 (N_1963,In_231,In_102);
and U1964 (N_1964,In_358,In_995);
nand U1965 (N_1965,In_814,In_149);
or U1966 (N_1966,In_516,In_463);
or U1967 (N_1967,In_878,In_919);
or U1968 (N_1968,In_441,In_608);
and U1969 (N_1969,In_422,In_338);
nand U1970 (N_1970,In_500,In_961);
nand U1971 (N_1971,In_912,In_667);
and U1972 (N_1972,In_230,In_698);
nand U1973 (N_1973,In_670,In_26);
and U1974 (N_1974,In_733,In_638);
or U1975 (N_1975,In_627,In_506);
xnor U1976 (N_1976,In_556,In_225);
nand U1977 (N_1977,In_518,In_964);
or U1978 (N_1978,In_397,In_494);
nand U1979 (N_1979,In_342,In_271);
and U1980 (N_1980,In_14,In_265);
nor U1981 (N_1981,In_978,In_462);
nor U1982 (N_1982,In_586,In_894);
or U1983 (N_1983,In_207,In_552);
or U1984 (N_1984,In_210,In_450);
or U1985 (N_1985,In_787,In_288);
and U1986 (N_1986,In_991,In_461);
nand U1987 (N_1987,In_3,In_685);
nand U1988 (N_1988,In_958,In_856);
nor U1989 (N_1989,In_938,In_39);
nor U1990 (N_1990,In_131,In_391);
and U1991 (N_1991,In_460,In_249);
nand U1992 (N_1992,In_632,In_329);
or U1993 (N_1993,In_843,In_784);
and U1994 (N_1994,In_923,In_328);
or U1995 (N_1995,In_586,In_590);
nand U1996 (N_1996,In_669,In_734);
or U1997 (N_1997,In_519,In_55);
and U1998 (N_1998,In_897,In_468);
nand U1999 (N_1999,In_182,In_408);
nor U2000 (N_2000,N_963,N_720);
nand U2001 (N_2001,N_100,N_1913);
and U2002 (N_2002,N_816,N_220);
nor U2003 (N_2003,N_543,N_245);
nand U2004 (N_2004,N_919,N_469);
nand U2005 (N_2005,N_897,N_1071);
and U2006 (N_2006,N_934,N_402);
nor U2007 (N_2007,N_1979,N_279);
nor U2008 (N_2008,N_1522,N_38);
or U2009 (N_2009,N_1353,N_1443);
nor U2010 (N_2010,N_1728,N_607);
nor U2011 (N_2011,N_216,N_1413);
nand U2012 (N_2012,N_567,N_909);
xnor U2013 (N_2013,N_954,N_1714);
nor U2014 (N_2014,N_535,N_95);
and U2015 (N_2015,N_1999,N_1405);
nor U2016 (N_2016,N_1208,N_1492);
and U2017 (N_2017,N_1193,N_1624);
or U2018 (N_2018,N_1472,N_1339);
nor U2019 (N_2019,N_508,N_692);
and U2020 (N_2020,N_1276,N_1816);
nor U2021 (N_2021,N_1115,N_233);
xnor U2022 (N_2022,N_1227,N_324);
and U2023 (N_2023,N_1506,N_1774);
nor U2024 (N_2024,N_1290,N_1588);
nand U2025 (N_2025,N_1474,N_772);
or U2026 (N_2026,N_1349,N_1994);
nor U2027 (N_2027,N_518,N_140);
nand U2028 (N_2028,N_864,N_568);
or U2029 (N_2029,N_178,N_1436);
nand U2030 (N_2030,N_1235,N_1579);
nand U2031 (N_2031,N_1259,N_494);
and U2032 (N_2032,N_612,N_1401);
xor U2033 (N_2033,N_1150,N_1245);
nor U2034 (N_2034,N_261,N_1059);
nor U2035 (N_2035,N_1511,N_775);
or U2036 (N_2036,N_387,N_268);
nor U2037 (N_2037,N_711,N_1817);
or U2038 (N_2038,N_1866,N_1283);
nor U2039 (N_2039,N_906,N_454);
or U2040 (N_2040,N_1786,N_1824);
nor U2041 (N_2041,N_724,N_1448);
nand U2042 (N_2042,N_1847,N_1111);
xor U2043 (N_2043,N_125,N_559);
nand U2044 (N_2044,N_786,N_1569);
nand U2045 (N_2045,N_93,N_1789);
and U2046 (N_2046,N_383,N_1654);
and U2047 (N_2047,N_825,N_422);
and U2048 (N_2048,N_1247,N_1814);
or U2049 (N_2049,N_1264,N_1546);
or U2050 (N_2050,N_1250,N_644);
or U2051 (N_2051,N_1981,N_332);
or U2052 (N_2052,N_530,N_1088);
nor U2053 (N_2053,N_845,N_1161);
nor U2054 (N_2054,N_1904,N_235);
nor U2055 (N_2055,N_427,N_69);
nor U2056 (N_2056,N_99,N_647);
nor U2057 (N_2057,N_153,N_605);
nand U2058 (N_2058,N_1215,N_476);
or U2059 (N_2059,N_232,N_707);
nor U2060 (N_2060,N_810,N_893);
or U2061 (N_2061,N_617,N_1122);
nand U2062 (N_2062,N_1151,N_289);
nand U2063 (N_2063,N_187,N_46);
and U2064 (N_2064,N_836,N_1384);
nand U2065 (N_2065,N_1284,N_507);
and U2066 (N_2066,N_1729,N_1836);
xor U2067 (N_2067,N_1554,N_1246);
and U2068 (N_2068,N_610,N_1281);
nor U2069 (N_2069,N_124,N_111);
nand U2070 (N_2070,N_453,N_765);
nand U2071 (N_2071,N_1336,N_251);
nand U2072 (N_2072,N_159,N_155);
xnor U2073 (N_2073,N_669,N_599);
nor U2074 (N_2074,N_393,N_467);
nand U2075 (N_2075,N_1528,N_286);
nand U2076 (N_2076,N_804,N_272);
xnor U2077 (N_2077,N_728,N_277);
nor U2078 (N_2078,N_598,N_1599);
and U2079 (N_2079,N_996,N_472);
nand U2080 (N_2080,N_754,N_204);
nand U2081 (N_2081,N_1343,N_106);
or U2082 (N_2082,N_1810,N_368);
or U2083 (N_2083,N_971,N_1975);
xnor U2084 (N_2084,N_1432,N_1854);
and U2085 (N_2085,N_1998,N_1333);
nand U2086 (N_2086,N_1147,N_1792);
and U2087 (N_2087,N_1177,N_426);
or U2088 (N_2088,N_215,N_759);
nand U2089 (N_2089,N_94,N_206);
nand U2090 (N_2090,N_1692,N_1076);
xor U2091 (N_2091,N_1602,N_705);
or U2092 (N_2092,N_616,N_1838);
nand U2093 (N_2093,N_1895,N_1565);
nor U2094 (N_2094,N_1100,N_1769);
and U2095 (N_2095,N_1548,N_384);
nor U2096 (N_2096,N_1342,N_1083);
nand U2097 (N_2097,N_869,N_1734);
xor U2098 (N_2098,N_562,N_1760);
or U2099 (N_2099,N_1559,N_645);
nor U2100 (N_2100,N_566,N_34);
or U2101 (N_2101,N_1470,N_366);
nor U2102 (N_2102,N_17,N_295);
nand U2103 (N_2103,N_1762,N_861);
or U2104 (N_2104,N_445,N_1633);
nand U2105 (N_2105,N_1656,N_1051);
or U2106 (N_2106,N_1042,N_1289);
nor U2107 (N_2107,N_1143,N_194);
nand U2108 (N_2108,N_1857,N_1431);
and U2109 (N_2109,N_1921,N_1253);
nand U2110 (N_2110,N_989,N_1267);
nor U2111 (N_2111,N_1035,N_1755);
and U2112 (N_2112,N_1219,N_633);
or U2113 (N_2113,N_1341,N_757);
and U2114 (N_2114,N_737,N_1204);
nand U2115 (N_2115,N_1038,N_1099);
nand U2116 (N_2116,N_351,N_579);
nor U2117 (N_2117,N_854,N_675);
and U2118 (N_2118,N_1382,N_965);
nor U2119 (N_2119,N_1784,N_385);
or U2120 (N_2120,N_1756,N_1152);
or U2121 (N_2121,N_490,N_142);
and U2122 (N_2122,N_358,N_1577);
nor U2123 (N_2123,N_666,N_1863);
or U2124 (N_2124,N_942,N_1323);
and U2125 (N_2125,N_1303,N_837);
xnor U2126 (N_2126,N_15,N_1305);
and U2127 (N_2127,N_872,N_503);
nand U2128 (N_2128,N_37,N_362);
xor U2129 (N_2129,N_1513,N_1710);
nand U2130 (N_2130,N_949,N_1301);
and U2131 (N_2131,N_1704,N_1918);
or U2132 (N_2132,N_483,N_850);
xor U2133 (N_2133,N_1618,N_1288);
nand U2134 (N_2134,N_1778,N_460);
nor U2135 (N_2135,N_554,N_1363);
nand U2136 (N_2136,N_284,N_326);
xor U2137 (N_2137,N_614,N_981);
nand U2138 (N_2138,N_1427,N_1055);
and U2139 (N_2139,N_556,N_1031);
and U2140 (N_2140,N_589,N_66);
and U2141 (N_2141,N_654,N_1648);
nor U2142 (N_2142,N_1881,N_308);
nand U2143 (N_2143,N_878,N_1074);
nor U2144 (N_2144,N_1039,N_678);
or U2145 (N_2145,N_998,N_1536);
and U2146 (N_2146,N_1945,N_832);
or U2147 (N_2147,N_306,N_1580);
or U2148 (N_2148,N_1291,N_1662);
nand U2149 (N_2149,N_1715,N_747);
and U2150 (N_2150,N_390,N_1309);
or U2151 (N_2151,N_214,N_1404);
nand U2152 (N_2152,N_528,N_197);
nor U2153 (N_2153,N_1829,N_1331);
and U2154 (N_2154,N_1397,N_1271);
xnor U2155 (N_2155,N_416,N_1986);
or U2156 (N_2156,N_855,N_565);
nor U2157 (N_2157,N_1210,N_994);
nand U2158 (N_2158,N_67,N_1899);
nor U2159 (N_2159,N_189,N_504);
or U2160 (N_2160,N_1661,N_269);
nand U2161 (N_2161,N_1324,N_320);
and U2162 (N_2162,N_1772,N_635);
and U2163 (N_2163,N_89,N_1007);
nand U2164 (N_2164,N_609,N_1665);
nand U2165 (N_2165,N_1096,N_1677);
xor U2166 (N_2166,N_1621,N_1860);
and U2167 (N_2167,N_1949,N_1399);
and U2168 (N_2168,N_1425,N_840);
nand U2169 (N_2169,N_1030,N_1721);
or U2170 (N_2170,N_1103,N_1357);
nand U2171 (N_2171,N_1400,N_1542);
and U2172 (N_2172,N_394,N_1930);
xnor U2173 (N_2173,N_896,N_780);
or U2174 (N_2174,N_951,N_450);
nor U2175 (N_2175,N_653,N_739);
and U2176 (N_2176,N_625,N_962);
nor U2177 (N_2177,N_1048,N_1943);
and U2178 (N_2178,N_770,N_755);
and U2179 (N_2179,N_409,N_285);
nor U2180 (N_2180,N_1089,N_1298);
or U2181 (N_2181,N_1642,N_1426);
and U2182 (N_2182,N_22,N_1851);
nor U2183 (N_2183,N_629,N_1780);
nand U2184 (N_2184,N_1178,N_1182);
nor U2185 (N_2185,N_1419,N_1138);
or U2186 (N_2186,N_1262,N_1980);
nand U2187 (N_2187,N_824,N_938);
or U2188 (N_2188,N_54,N_1002);
nand U2189 (N_2189,N_1718,N_1187);
and U2190 (N_2190,N_588,N_1174);
xnor U2191 (N_2191,N_844,N_813);
and U2192 (N_2192,N_1795,N_944);
xnor U2193 (N_2193,N_1025,N_334);
nand U2194 (N_2194,N_1575,N_240);
nor U2195 (N_2195,N_78,N_1175);
or U2196 (N_2196,N_929,N_234);
nor U2197 (N_2197,N_943,N_1909);
nand U2198 (N_2198,N_83,N_1682);
xnor U2199 (N_2199,N_908,N_369);
and U2200 (N_2200,N_16,N_948);
nor U2201 (N_2201,N_735,N_486);
nor U2202 (N_2202,N_1417,N_1626);
xnor U2203 (N_2203,N_355,N_1312);
and U2204 (N_2204,N_1666,N_1660);
nand U2205 (N_2205,N_659,N_712);
and U2206 (N_2206,N_241,N_1200);
or U2207 (N_2207,N_1763,N_1676);
or U2208 (N_2208,N_1509,N_413);
nand U2209 (N_2209,N_613,N_671);
nand U2210 (N_2210,N_313,N_1738);
or U2211 (N_2211,N_1912,N_680);
and U2212 (N_2212,N_1158,N_1359);
xnor U2213 (N_2213,N_151,N_1350);
nor U2214 (N_2214,N_801,N_1097);
or U2215 (N_2215,N_1672,N_1709);
and U2216 (N_2216,N_926,N_939);
and U2217 (N_2217,N_398,N_457);
and U2218 (N_2218,N_835,N_782);
and U2219 (N_2219,N_1233,N_1675);
and U2220 (N_2220,N_152,N_1519);
or U2221 (N_2221,N_164,N_59);
xnor U2222 (N_2222,N_1573,N_177);
or U2223 (N_2223,N_44,N_606);
nand U2224 (N_2224,N_418,N_1114);
or U2225 (N_2225,N_1646,N_1241);
or U2226 (N_2226,N_1344,N_491);
nor U2227 (N_2227,N_1917,N_231);
nand U2228 (N_2228,N_1809,N_170);
xor U2229 (N_2229,N_375,N_1387);
and U2230 (N_2230,N_1856,N_1320);
nand U2231 (N_2231,N_1547,N_1438);
or U2232 (N_2232,N_407,N_1455);
or U2233 (N_2233,N_371,N_1942);
or U2234 (N_2234,N_860,N_968);
nand U2235 (N_2235,N_715,N_1467);
nor U2236 (N_2236,N_716,N_1885);
nor U2237 (N_2237,N_363,N_335);
or U2238 (N_2238,N_1123,N_437);
nor U2239 (N_2239,N_501,N_668);
nor U2240 (N_2240,N_974,N_13);
nor U2241 (N_2241,N_560,N_1985);
and U2242 (N_2242,N_276,N_638);
nand U2243 (N_2243,N_1578,N_706);
and U2244 (N_2244,N_1477,N_496);
nor U2245 (N_2245,N_624,N_969);
nand U2246 (N_2246,N_96,N_336);
or U2247 (N_2247,N_1613,N_726);
nor U2248 (N_2248,N_547,N_783);
or U2249 (N_2249,N_1315,N_1663);
nand U2250 (N_2250,N_1012,N_1925);
nand U2251 (N_2251,N_1388,N_1976);
xor U2252 (N_2252,N_1832,N_18);
and U2253 (N_2253,N_350,N_1274);
nand U2254 (N_2254,N_1882,N_1328);
nor U2255 (N_2255,N_1517,N_555);
nor U2256 (N_2256,N_1104,N_834);
and U2257 (N_2257,N_907,N_1855);
and U2258 (N_2258,N_1804,N_756);
nand U2259 (N_2259,N_630,N_493);
nor U2260 (N_2260,N_1697,N_1695);
and U2261 (N_2261,N_1598,N_495);
nand U2262 (N_2262,N_760,N_1263);
or U2263 (N_2263,N_331,N_743);
and U2264 (N_2264,N_701,N_649);
or U2265 (N_2265,N_1272,N_24);
nand U2266 (N_2266,N_1524,N_1016);
nand U2267 (N_2267,N_56,N_1785);
nand U2268 (N_2268,N_451,N_98);
nand U2269 (N_2269,N_1040,N_1889);
xor U2270 (N_2270,N_474,N_797);
xor U2271 (N_2271,N_219,N_468);
or U2272 (N_2272,N_202,N_32);
and U2273 (N_2273,N_1282,N_1527);
nor U2274 (N_2274,N_281,N_438);
nor U2275 (N_2275,N_594,N_109);
nand U2276 (N_2276,N_168,N_563);
nor U2277 (N_2277,N_417,N_1671);
and U2278 (N_2278,N_1534,N_1045);
nor U2279 (N_2279,N_1017,N_456);
or U2280 (N_2280,N_820,N_403);
nor U2281 (N_2281,N_1947,N_329);
nand U2282 (N_2282,N_307,N_858);
and U2283 (N_2283,N_1205,N_992);
nand U2284 (N_2284,N_211,N_514);
or U2285 (N_2285,N_1368,N_785);
or U2286 (N_2286,N_1616,N_619);
xor U2287 (N_2287,N_1933,N_150);
nor U2288 (N_2288,N_767,N_356);
nor U2289 (N_2289,N_738,N_652);
nand U2290 (N_2290,N_461,N_972);
and U2291 (N_2291,N_1951,N_829);
xor U2292 (N_2292,N_120,N_805);
or U2293 (N_2293,N_1212,N_1098);
nor U2294 (N_2294,N_222,N_440);
or U2295 (N_2295,N_1422,N_1988);
nand U2296 (N_2296,N_1759,N_1993);
nor U2297 (N_2297,N_1195,N_1984);
and U2298 (N_2298,N_76,N_793);
or U2299 (N_2299,N_1188,N_255);
and U2300 (N_2300,N_1963,N_1903);
xnor U2301 (N_2301,N_1645,N_1068);
nor U2302 (N_2302,N_1418,N_297);
and U2303 (N_2303,N_626,N_1587);
or U2304 (N_2304,N_537,N_1242);
xnor U2305 (N_2305,N_1965,N_1620);
xor U2306 (N_2306,N_452,N_985);
nand U2307 (N_2307,N_1126,N_764);
or U2308 (N_2308,N_1139,N_1908);
nand U2309 (N_2309,N_1507,N_997);
and U2310 (N_2310,N_1297,N_1469);
or U2311 (N_2311,N_1629,N_1466);
nand U2312 (N_2312,N_1287,N_1699);
and U2313 (N_2313,N_280,N_1410);
and U2314 (N_2314,N_283,N_360);
and U2315 (N_2315,N_1162,N_627);
nor U2316 (N_2316,N_79,N_344);
and U2317 (N_2317,N_915,N_1346);
nor U2318 (N_2318,N_1337,N_1490);
and U2319 (N_2319,N_500,N_1430);
nand U2320 (N_2320,N_1192,N_1731);
or U2321 (N_2321,N_1664,N_1216);
and U2322 (N_2322,N_1801,N_795);
nand U2323 (N_2323,N_367,N_734);
and U2324 (N_2324,N_166,N_103);
nor U2325 (N_2325,N_488,N_1777);
nor U2326 (N_2326,N_621,N_830);
nand U2327 (N_2327,N_1906,N_538);
and U2328 (N_2328,N_1116,N_973);
nor U2329 (N_2329,N_1929,N_1468);
nand U2330 (N_2330,N_1000,N_1010);
or U2331 (N_2331,N_947,N_1080);
xor U2332 (N_2332,N_1920,N_1148);
nand U2333 (N_2333,N_1757,N_1574);
nand U2334 (N_2334,N_1510,N_148);
nor U2335 (N_2335,N_789,N_799);
nand U2336 (N_2336,N_26,N_304);
and U2337 (N_2337,N_798,N_61);
nor U2338 (N_2338,N_575,N_911);
and U2339 (N_2339,N_1354,N_1313);
or U2340 (N_2340,N_1926,N_1416);
or U2341 (N_2341,N_119,N_637);
and U2342 (N_2342,N_217,N_814);
nand U2343 (N_2343,N_122,N_173);
nor U2344 (N_2344,N_1694,N_1458);
and U2345 (N_2345,N_1739,N_784);
or U2346 (N_2346,N_851,N_1190);
and U2347 (N_2347,N_1722,N_1252);
nand U2348 (N_2348,N_646,N_116);
or U2349 (N_2349,N_193,N_1269);
or U2350 (N_2350,N_704,N_48);
and U2351 (N_2351,N_791,N_1257);
and U2352 (N_2352,N_1402,N_988);
and U2353 (N_2353,N_1968,N_90);
nor U2354 (N_2354,N_532,N_1171);
or U2355 (N_2355,N_144,N_986);
or U2356 (N_2356,N_875,N_198);
or U2357 (N_2357,N_960,N_1793);
and U2358 (N_2358,N_1799,N_1953);
or U2359 (N_2359,N_21,N_807);
or U2360 (N_2360,N_702,N_209);
nand U2361 (N_2361,N_1691,N_1717);
nand U2362 (N_2362,N_1060,N_60);
nand U2363 (N_2363,N_444,N_1159);
nor U2364 (N_2364,N_435,N_1132);
nand U2365 (N_2365,N_761,N_5);
nand U2366 (N_2366,N_913,N_1843);
or U2367 (N_2367,N_464,N_910);
and U2368 (N_2368,N_1770,N_91);
and U2369 (N_2369,N_343,N_1532);
or U2370 (N_2370,N_1120,N_1378);
and U2371 (N_2371,N_1916,N_293);
and U2372 (N_2372,N_1224,N_449);
and U2373 (N_2373,N_1766,N_1607);
xnor U2374 (N_2374,N_718,N_823);
or U2375 (N_2375,N_1592,N_516);
nand U2376 (N_2376,N_1,N_1658);
nor U2377 (N_2377,N_1142,N_1545);
and U2378 (N_2378,N_886,N_248);
or U2379 (N_2379,N_1499,N_1238);
nand U2380 (N_2380,N_1831,N_812);
nand U2381 (N_2381,N_1037,N_1849);
or U2382 (N_2382,N_361,N_1237);
xnor U2383 (N_2383,N_870,N_788);
nor U2384 (N_2384,N_689,N_327);
and U2385 (N_2385,N_1302,N_684);
nand U2386 (N_2386,N_1015,N_1608);
and U2387 (N_2387,N_157,N_790);
or U2388 (N_2388,N_657,N_572);
nor U2389 (N_2389,N_1390,N_587);
nand U2390 (N_2390,N_1915,N_1144);
or U2391 (N_2391,N_1779,N_1723);
or U2392 (N_2392,N_833,N_1669);
and U2393 (N_2393,N_1090,N_806);
xnor U2394 (N_2394,N_717,N_901);
nor U2395 (N_2395,N_544,N_1356);
or U2396 (N_2396,N_552,N_64);
xor U2397 (N_2397,N_1876,N_1463);
and U2398 (N_2398,N_731,N_1673);
or U2399 (N_2399,N_1459,N_68);
or U2400 (N_2400,N_1670,N_527);
nand U2401 (N_2401,N_1970,N_571);
nor U2402 (N_2402,N_1220,N_640);
nor U2403 (N_2403,N_341,N_1280);
nand U2404 (N_2404,N_639,N_397);
nor U2405 (N_2405,N_1110,N_1610);
or U2406 (N_2406,N_162,N_225);
or U2407 (N_2407,N_581,N_1892);
nand U2408 (N_2408,N_1612,N_1218);
or U2409 (N_2409,N_374,N_1582);
and U2410 (N_2410,N_1516,N_1605);
nand U2411 (N_2411,N_1166,N_838);
and U2412 (N_2412,N_1877,N_1823);
xnor U2413 (N_2413,N_936,N_1130);
or U2414 (N_2414,N_1299,N_1029);
nor U2415 (N_2415,N_1032,N_857);
and U2416 (N_2416,N_902,N_1541);
nor U2417 (N_2417,N_1950,N_1452);
or U2418 (N_2418,N_1421,N_1705);
nor U2419 (N_2419,N_47,N_1846);
and U2420 (N_2420,N_927,N_379);
nor U2421 (N_2421,N_459,N_686);
nand U2422 (N_2422,N_1072,N_378);
nand U2423 (N_2423,N_1084,N_773);
or U2424 (N_2424,N_1462,N_1322);
nand U2425 (N_2425,N_884,N_1194);
or U2426 (N_2426,N_443,N_388);
and U2427 (N_2427,N_874,N_1450);
xor U2428 (N_2428,N_411,N_867);
or U2429 (N_2429,N_466,N_428);
and U2430 (N_2430,N_597,N_564);
and U2431 (N_2431,N_1078,N_1085);
nor U2432 (N_2432,N_1494,N_966);
nor U2433 (N_2433,N_766,N_628);
and U2434 (N_2434,N_822,N_1479);
nand U2435 (N_2435,N_1690,N_97);
nand U2436 (N_2436,N_1758,N_1334);
nor U2437 (N_2437,N_608,N_710);
or U2438 (N_2438,N_1079,N_741);
nand U2439 (N_2439,N_11,N_184);
or U2440 (N_2440,N_1451,N_1744);
nand U2441 (N_2441,N_1934,N_1615);
or U2442 (N_2442,N_266,N_1749);
xor U2443 (N_2443,N_1603,N_1544);
nand U2444 (N_2444,N_1883,N_287);
nor U2445 (N_2445,N_1327,N_933);
and U2446 (N_2446,N_282,N_1800);
nor U2447 (N_2447,N_1797,N_1741);
or U2448 (N_2448,N_1498,N_1409);
or U2449 (N_2449,N_108,N_895);
nor U2450 (N_2450,N_1940,N_4);
nor U2451 (N_2451,N_243,N_238);
or U2452 (N_2452,N_688,N_1414);
nor U2453 (N_2453,N_742,N_322);
nor U2454 (N_2454,N_1674,N_1844);
or U2455 (N_2455,N_478,N_1812);
nor U2456 (N_2456,N_519,N_1249);
and U2457 (N_2457,N_1596,N_1875);
nor U2458 (N_2458,N_749,N_1131);
nor U2459 (N_2459,N_1884,N_1213);
nand U2460 (N_2460,N_138,N_1659);
nand U2461 (N_2461,N_310,N_1270);
or U2462 (N_2462,N_1295,N_1868);
nand U2463 (N_2463,N_311,N_1018);
nor U2464 (N_2464,N_1364,N_1394);
nand U2465 (N_2465,N_693,N_1650);
or U2466 (N_2466,N_1408,N_298);
or U2467 (N_2467,N_128,N_1733);
nand U2468 (N_2468,N_439,N_485);
nand U2469 (N_2469,N_1886,N_257);
or U2470 (N_2470,N_75,N_1708);
nor U2471 (N_2471,N_1021,N_1523);
nand U2472 (N_2472,N_1803,N_1564);
nand U2473 (N_2473,N_1525,N_685);
xnor U2474 (N_2474,N_1712,N_914);
and U2475 (N_2475,N_1611,N_1255);
nand U2476 (N_2476,N_406,N_1067);
nor U2477 (N_2477,N_1058,N_1375);
and U2478 (N_2478,N_903,N_299);
xor U2479 (N_2479,N_848,N_1526);
and U2480 (N_2480,N_1636,N_309);
nand U2481 (N_2481,N_1637,N_1179);
xnor U2482 (N_2482,N_62,N_1300);
xnor U2483 (N_2483,N_463,N_1181);
or U2484 (N_2484,N_553,N_1261);
xor U2485 (N_2485,N_736,N_1790);
nor U2486 (N_2486,N_1160,N_865);
nor U2487 (N_2487,N_1743,N_364);
or U2488 (N_2488,N_1737,N_447);
and U2489 (N_2489,N_1753,N_1732);
or U2490 (N_2490,N_224,N_1537);
xnor U2491 (N_2491,N_312,N_339);
nor U2492 (N_2492,N_1101,N_156);
nor U2493 (N_2493,N_1754,N_1638);
or U2494 (N_2494,N_540,N_1653);
nand U2495 (N_2495,N_1293,N_839);
nand U2496 (N_2496,N_1285,N_506);
and U2497 (N_2497,N_499,N_1093);
nor U2498 (N_2498,N_107,N_1563);
nor U2499 (N_2499,N_1614,N_1222);
nand U2500 (N_2500,N_1685,N_877);
and U2501 (N_2501,N_1202,N_1859);
nor U2502 (N_2502,N_419,N_1073);
xnor U2503 (N_2503,N_846,N_252);
and U2504 (N_2504,N_542,N_1497);
nand U2505 (N_2505,N_1374,N_725);
nor U2506 (N_2506,N_771,N_1726);
or U2507 (N_2507,N_1745,N_405);
and U2508 (N_2508,N_1825,N_497);
and U2509 (N_2509,N_681,N_796);
and U2510 (N_2510,N_1345,N_133);
nor U2511 (N_2511,N_180,N_1735);
and U2512 (N_2512,N_1657,N_585);
nand U2513 (N_2513,N_955,N_1369);
nor U2514 (N_2514,N_643,N_976);
and U2515 (N_2515,N_748,N_1229);
nor U2516 (N_2516,N_1113,N_964);
nor U2517 (N_2517,N_1361,N_525);
nand U2518 (N_2518,N_1681,N_891);
or U2519 (N_2519,N_561,N_1767);
xor U2520 (N_2520,N_86,N_1641);
nor U2521 (N_2521,N_1553,N_550);
and U2522 (N_2522,N_1938,N_27);
nor U2523 (N_2523,N_1446,N_249);
and U2524 (N_2524,N_410,N_1398);
and U2525 (N_2525,N_1716,N_223);
nand U2526 (N_2526,N_1063,N_925);
nand U2527 (N_2527,N_1678,N_1157);
or U2528 (N_2528,N_890,N_593);
nor U2529 (N_2529,N_642,N_1948);
nor U2530 (N_2530,N_36,N_213);
nor U2531 (N_2531,N_545,N_937);
nand U2532 (N_2532,N_1070,N_604);
nor U2533 (N_2533,N_1783,N_227);
and U2534 (N_2534,N_573,N_1260);
xor U2535 (N_2535,N_414,N_1955);
or U2536 (N_2536,N_421,N_892);
and U2537 (N_2537,N_977,N_1852);
nand U2538 (N_2538,N_104,N_1062);
and U2539 (N_2539,N_1258,N_1639);
nand U2540 (N_2540,N_1473,N_515);
nand U2541 (N_2541,N_191,N_359);
nand U2542 (N_2542,N_1619,N_1256);
nor U2543 (N_2543,N_382,N_665);
nor U2544 (N_2544,N_1504,N_112);
nor U2545 (N_2545,N_1061,N_1486);
or U2546 (N_2546,N_305,N_302);
nand U2547 (N_2547,N_1496,N_207);
and U2548 (N_2548,N_1987,N_487);
nand U2549 (N_2549,N_1075,N_1381);
and U2550 (N_2550,N_1962,N_531);
and U2551 (N_2551,N_1702,N_1403);
and U2552 (N_2552,N_576,N_650);
nand U2553 (N_2553,N_1643,N_446);
and U2554 (N_2554,N_602,N_1041);
or U2555 (N_2555,N_275,N_509);
xor U2556 (N_2556,N_1217,N_904);
and U2557 (N_2557,N_1457,N_990);
nand U2558 (N_2558,N_161,N_333);
or U2559 (N_2559,N_274,N_221);
nand U2560 (N_2560,N_77,N_74);
and U2561 (N_2561,N_1279,N_808);
and U2562 (N_2562,N_1982,N_620);
nor U2563 (N_2563,N_480,N_477);
nand U2564 (N_2564,N_84,N_1560);
nor U2565 (N_2565,N_113,N_1992);
and U2566 (N_2566,N_826,N_1232);
nor U2567 (N_2567,N_448,N_1453);
nand U2568 (N_2568,N_57,N_1440);
and U2569 (N_2569,N_774,N_1201);
or U2570 (N_2570,N_391,N_1266);
or U2571 (N_2571,N_165,N_174);
and U2572 (N_2572,N_1773,N_983);
or U2573 (N_2573,N_667,N_967);
nand U2574 (N_2574,N_697,N_863);
nor U2575 (N_2575,N_912,N_727);
and U2576 (N_2576,N_1449,N_1820);
nand U2577 (N_2577,N_1454,N_1197);
xor U2578 (N_2578,N_470,N_1698);
nor U2579 (N_2579,N_1841,N_1340);
nor U2580 (N_2580,N_167,N_534);
and U2581 (N_2581,N_1972,N_879);
and U2582 (N_2582,N_887,N_294);
xnor U2583 (N_2583,N_482,N_1064);
and U2584 (N_2584,N_1594,N_1781);
nor U2585 (N_2585,N_1765,N_924);
nand U2586 (N_2586,N_183,N_172);
or U2587 (N_2587,N_930,N_762);
and U2588 (N_2588,N_852,N_492);
or U2589 (N_2589,N_1046,N_1796);
nand U2590 (N_2590,N_1170,N_803);
nor U2591 (N_2591,N_1186,N_1049);
or U2592 (N_2592,N_586,N_337);
nor U2593 (N_2593,N_1826,N_952);
nand U2594 (N_2594,N_1990,N_536);
and U2595 (N_2595,N_479,N_1189);
and U2596 (N_2596,N_1835,N_1493);
nand U2597 (N_2597,N_458,N_549);
nor U2598 (N_2598,N_1693,N_303);
and U2599 (N_2599,N_1748,N_584);
nor U2600 (N_2600,N_154,N_228);
or U2601 (N_2601,N_751,N_205);
or U2602 (N_2602,N_300,N_1052);
xnor U2603 (N_2603,N_1811,N_1460);
or U2604 (N_2604,N_33,N_105);
nor U2605 (N_2605,N_1004,N_719);
and U2606 (N_2606,N_779,N_1609);
nand U2607 (N_2607,N_1332,N_296);
nor U2608 (N_2608,N_1989,N_1360);
xor U2609 (N_2609,N_1791,N_511);
xnor U2610 (N_2610,N_1156,N_1347);
or U2611 (N_2611,N_1680,N_1529);
nand U2612 (N_2612,N_1539,N_1538);
and U2613 (N_2613,N_1971,N_1869);
nand U2614 (N_2614,N_995,N_815);
nor U2615 (N_2615,N_674,N_1475);
and U2616 (N_2616,N_1583,N_1294);
nand U2617 (N_2617,N_1191,N_82);
nand U2618 (N_2618,N_389,N_1198);
nand U2619 (N_2619,N_853,N_1761);
xor U2620 (N_2620,N_1128,N_1923);
or U2621 (N_2621,N_1747,N_843);
nor U2622 (N_2622,N_827,N_1686);
nand U2623 (N_2623,N_777,N_1873);
and U2624 (N_2624,N_1306,N_818);
nand U2625 (N_2625,N_348,N_1874);
or U2626 (N_2626,N_1461,N_1065);
nand U2627 (N_2627,N_601,N_208);
or U2628 (N_2628,N_1069,N_1818);
or U2629 (N_2629,N_288,N_1481);
nor U2630 (N_2630,N_932,N_894);
nand U2631 (N_2631,N_1081,N_1689);
xor U2632 (N_2632,N_1406,N_1751);
nand U2633 (N_2633,N_661,N_1112);
nor U2634 (N_2634,N_979,N_920);
nand U2635 (N_2635,N_1286,N_1628);
and U2636 (N_2636,N_1632,N_250);
and U2637 (N_2637,N_1604,N_1173);
nor U2638 (N_2638,N_1815,N_65);
nand U2639 (N_2639,N_372,N_163);
and U2640 (N_2640,N_399,N_218);
and U2641 (N_2641,N_1314,N_970);
or U2642 (N_2642,N_45,N_123);
nand U2643 (N_2643,N_1169,N_1521);
xnor U2644 (N_2644,N_683,N_110);
and U2645 (N_2645,N_583,N_1488);
and U2646 (N_2646,N_740,N_141);
nor U2647 (N_2647,N_1531,N_1141);
and U2648 (N_2648,N_1711,N_1456);
and U2649 (N_2649,N_641,N_136);
and U2650 (N_2650,N_1372,N_1483);
and U2651 (N_2651,N_1435,N_1640);
nor U2652 (N_2652,N_1495,N_475);
nand U2653 (N_2653,N_1888,N_7);
or U2654 (N_2654,N_679,N_1006);
and U2655 (N_2655,N_1244,N_1750);
nor U2656 (N_2656,N_1106,N_430);
xor U2657 (N_2657,N_1377,N_1520);
or U2658 (N_2658,N_1225,N_101);
nor U2659 (N_2659,N_520,N_999);
nor U2660 (N_2660,N_632,N_158);
and U2661 (N_2661,N_744,N_1476);
or U2662 (N_2662,N_1556,N_946);
nand U2663 (N_2663,N_1830,N_1775);
or U2664 (N_2664,N_1533,N_1043);
nor U2665 (N_2665,N_866,N_396);
nor U2666 (N_2666,N_776,N_1420);
xnor U2667 (N_2667,N_1326,N_957);
or U2668 (N_2668,N_940,N_1960);
and U2669 (N_2669,N_841,N_1939);
and U2670 (N_2670,N_1897,N_1050);
nor U2671 (N_2671,N_600,N_1057);
or U2672 (N_2672,N_1558,N_1180);
nor U2673 (N_2673,N_1028,N_182);
and U2674 (N_2674,N_317,N_1688);
xor U2675 (N_2675,N_577,N_1231);
nor U2676 (N_2676,N_1027,N_1595);
and U2677 (N_2677,N_1995,N_1969);
xor U2678 (N_2678,N_1167,N_132);
nand U2679 (N_2679,N_1278,N_1606);
or U2680 (N_2680,N_1867,N_1958);
nor U2681 (N_2681,N_1308,N_687);
nand U2682 (N_2682,N_1683,N_1505);
and U2683 (N_2683,N_392,N_1207);
nand U2684 (N_2684,N_1713,N_88);
nor U2685 (N_2685,N_1019,N_1385);
or U2686 (N_2686,N_1827,N_1706);
nor U2687 (N_2687,N_254,N_696);
xor U2688 (N_2688,N_1184,N_1243);
nand U2689 (N_2689,N_982,N_1091);
nand U2690 (N_2690,N_1898,N_695);
and U2691 (N_2691,N_676,N_876);
or U2692 (N_2692,N_171,N_871);
or U2693 (N_2693,N_342,N_700);
xnor U2694 (N_2694,N_1822,N_636);
and U2695 (N_2695,N_1185,N_526);
and U2696 (N_2696,N_230,N_365);
xnor U2697 (N_2697,N_541,N_196);
xor U2698 (N_2698,N_1500,N_1922);
and U2699 (N_2699,N_1914,N_118);
nor U2700 (N_2700,N_1617,N_8);
and U2701 (N_2701,N_905,N_1226);
nor U2702 (N_2702,N_242,N_1865);
or U2703 (N_2703,N_1172,N_43);
and U2704 (N_2704,N_1667,N_201);
nand U2705 (N_2705,N_1833,N_993);
nor U2706 (N_2706,N_1155,N_1429);
and U2707 (N_2707,N_1808,N_1880);
or U2708 (N_2708,N_264,N_498);
and U2709 (N_2709,N_1586,N_1240);
nand U2710 (N_2710,N_134,N_1720);
nor U2711 (N_2711,N_1802,N_1597);
or U2712 (N_2712,N_787,N_87);
or U2713 (N_2713,N_425,N_1581);
xnor U2714 (N_2714,N_1296,N_1540);
or U2715 (N_2715,N_548,N_881);
or U2716 (N_2716,N_980,N_1991);
nor U2717 (N_2717,N_662,N_1746);
nand U2718 (N_2718,N_200,N_750);
or U2719 (N_2719,N_1623,N_1622);
nor U2720 (N_2720,N_253,N_146);
xor U2721 (N_2721,N_1214,N_1894);
nor U2722 (N_2722,N_1776,N_1135);
nor U2723 (N_2723,N_730,N_1118);
nor U2724 (N_2724,N_19,N_271);
nand U2725 (N_2725,N_433,N_1941);
nor U2726 (N_2726,N_373,N_1543);
nand U2727 (N_2727,N_135,N_918);
nand U2728 (N_2728,N_1557,N_239);
or U2729 (N_2729,N_935,N_1230);
or U2730 (N_2730,N_656,N_781);
or U2731 (N_2731,N_1902,N_984);
nor U2732 (N_2732,N_1491,N_1701);
nor U2733 (N_2733,N_1630,N_1358);
nand U2734 (N_2734,N_673,N_473);
and U2735 (N_2735,N_1502,N_1376);
nor U2736 (N_2736,N_592,N_1740);
xor U2737 (N_2737,N_1134,N_529);
nand U2738 (N_2738,N_899,N_524);
or U2739 (N_2739,N_1203,N_1329);
nand U2740 (N_2740,N_1465,N_51);
nor U2741 (N_2741,N_401,N_1514);
nand U2742 (N_2742,N_1066,N_1501);
nand U2743 (N_2743,N_1014,N_346);
and U2744 (N_2744,N_1555,N_1412);
or U2745 (N_2745,N_1095,N_1572);
xor U2746 (N_2746,N_663,N_1277);
or U2747 (N_2747,N_259,N_580);
nand U2748 (N_2748,N_20,N_63);
or U2749 (N_2749,N_1627,N_23);
or U2750 (N_2750,N_188,N_953);
nand U2751 (N_2751,N_1445,N_883);
nand U2752 (N_2752,N_130,N_1077);
or U2753 (N_2753,N_1023,N_574);
nand U2754 (N_2754,N_179,N_291);
nand U2755 (N_2755,N_591,N_691);
nand U2756 (N_2756,N_143,N_677);
or U2757 (N_2757,N_31,N_1129);
nor U2758 (N_2758,N_53,N_1821);
and U2759 (N_2759,N_328,N_352);
or U2760 (N_2760,N_1024,N_623);
nand U2761 (N_2761,N_578,N_347);
nand U2762 (N_2762,N_192,N_1444);
nor U2763 (N_2763,N_290,N_1551);
or U2764 (N_2764,N_1946,N_1983);
or U2765 (N_2765,N_1145,N_817);
and U2766 (N_2766,N_370,N_648);
nand U2767 (N_2767,N_1355,N_1001);
or U2768 (N_2768,N_1105,N_338);
xor U2769 (N_2769,N_978,N_1373);
xor U2770 (N_2770,N_1590,N_81);
nand U2771 (N_2771,N_1956,N_1787);
and U2772 (N_2772,N_729,N_203);
nor U2773 (N_2773,N_1959,N_703);
nor U2774 (N_2774,N_395,N_1600);
nand U2775 (N_2775,N_1996,N_1589);
nor U2776 (N_2776,N_682,N_1591);
xor U2777 (N_2777,N_190,N_1649);
or U2778 (N_2778,N_1878,N_1927);
nand U2779 (N_2779,N_1928,N_1317);
nor U2780 (N_2780,N_462,N_212);
and U2781 (N_2781,N_880,N_752);
nor U2782 (N_2782,N_28,N_733);
and U2783 (N_2783,N_273,N_690);
nor U2784 (N_2784,N_1011,N_408);
and U2785 (N_2785,N_1196,N_1900);
or U2786 (N_2786,N_1407,N_941);
nor U2787 (N_2787,N_354,N_1764);
nand U2788 (N_2788,N_1318,N_1005);
xnor U2789 (N_2789,N_1647,N_102);
nor U2790 (N_2790,N_278,N_267);
or U2791 (N_2791,N_570,N_1871);
or U2792 (N_2792,N_1352,N_956);
and U2793 (N_2793,N_1601,N_1396);
or U2794 (N_2794,N_800,N_634);
or U2795 (N_2795,N_1853,N_1367);
nand U2796 (N_2796,N_1768,N_1625);
and U2797 (N_2797,N_856,N_1858);
and U2798 (N_2798,N_664,N_847);
nor U2799 (N_2799,N_1009,N_1593);
or U2800 (N_2800,N_551,N_517);
nor U2801 (N_2801,N_386,N_1819);
and U2802 (N_2802,N_1634,N_169);
xor U2803 (N_2803,N_145,N_1165);
or U2804 (N_2804,N_1102,N_1932);
and U2805 (N_2805,N_185,N_1478);
or U2806 (N_2806,N_898,N_794);
nor U2807 (N_2807,N_1047,N_819);
and U2808 (N_2808,N_961,N_959);
nor U2809 (N_2809,N_247,N_714);
nand U2810 (N_2810,N_1428,N_1961);
or U2811 (N_2811,N_1316,N_1644);
or U2812 (N_2812,N_868,N_615);
nand U2813 (N_2813,N_1107,N_330);
nand U2814 (N_2814,N_1265,N_175);
nor U2815 (N_2815,N_237,N_484);
xnor U2816 (N_2816,N_1489,N_522);
nor U2817 (N_2817,N_1806,N_1441);
and U2818 (N_2818,N_1325,N_1870);
nor U2819 (N_2819,N_1805,N_831);
or U2820 (N_2820,N_1036,N_71);
nor U2821 (N_2821,N_1013,N_595);
or U2822 (N_2822,N_1026,N_1700);
nor U2823 (N_2823,N_1911,N_244);
or U2824 (N_2824,N_1108,N_723);
or U2825 (N_2825,N_1515,N_732);
and U2826 (N_2826,N_1254,N_1571);
or U2827 (N_2827,N_1321,N_1304);
nor U2828 (N_2828,N_127,N_1034);
nor U2829 (N_2829,N_849,N_928);
nand U2830 (N_2830,N_380,N_1366);
nand U2831 (N_2831,N_42,N_1168);
nand U2832 (N_2832,N_1905,N_1423);
nor U2833 (N_2833,N_828,N_931);
nand U2834 (N_2834,N_1395,N_1484);
or U2835 (N_2835,N_236,N_1974);
nor U2836 (N_2836,N_129,N_1480);
or U2837 (N_2837,N_1518,N_1228);
nand U2838 (N_2838,N_1471,N_1840);
and U2839 (N_2839,N_945,N_318);
xor U2840 (N_2840,N_1631,N_1437);
or U2841 (N_2841,N_1845,N_746);
nand U2842 (N_2842,N_25,N_1153);
nand U2843 (N_2843,N_1679,N_1392);
nor U2844 (N_2844,N_1655,N_922);
nor U2845 (N_2845,N_1003,N_139);
and U2846 (N_2846,N_1273,N_1464);
nand U2847 (N_2847,N_1053,N_1842);
or U2848 (N_2848,N_1149,N_1788);
xnor U2849 (N_2849,N_917,N_1771);
nor U2850 (N_2850,N_889,N_9);
and U2851 (N_2851,N_263,N_1236);
nand U2852 (N_2852,N_809,N_596);
or U2853 (N_2853,N_1997,N_1487);
nand U2854 (N_2854,N_160,N_1552);
nand U2855 (N_2855,N_1176,N_699);
and U2856 (N_2856,N_1183,N_80);
nand U2857 (N_2857,N_455,N_1872);
or U2858 (N_2858,N_270,N_55);
or U2859 (N_2859,N_1782,N_1535);
nand U2860 (N_2860,N_655,N_353);
or U2861 (N_2861,N_1954,N_1550);
nor U2862 (N_2862,N_1206,N_1901);
or U2863 (N_2863,N_1248,N_1937);
nor U2864 (N_2864,N_246,N_1127);
nor U2865 (N_2865,N_753,N_603);
nand U2866 (N_2866,N_1124,N_325);
nand U2867 (N_2867,N_558,N_1567);
and U2868 (N_2868,N_1379,N_1292);
or U2869 (N_2869,N_1087,N_1307);
nor U2870 (N_2870,N_1807,N_6);
nor U2871 (N_2871,N_1635,N_1687);
nor U2872 (N_2872,N_292,N_1424);
and U2873 (N_2873,N_1652,N_1879);
nand U2874 (N_2874,N_186,N_888);
and U2875 (N_2875,N_1752,N_1319);
nand U2876 (N_2876,N_1268,N_512);
nor U2877 (N_2877,N_92,N_950);
nand U2878 (N_2878,N_713,N_1957);
or U2879 (N_2879,N_1887,N_10);
nor U2880 (N_2880,N_1813,N_73);
and U2881 (N_2881,N_1117,N_1146);
xnor U2882 (N_2882,N_1086,N_1209);
nor U2883 (N_2883,N_226,N_489);
xor U2884 (N_2884,N_321,N_958);
nand U2885 (N_2885,N_1164,N_404);
nand U2886 (N_2886,N_436,N_30);
xor U2887 (N_2887,N_1140,N_1561);
nand U2888 (N_2888,N_1850,N_1977);
xor U2889 (N_2889,N_694,N_131);
nand U2890 (N_2890,N_1861,N_708);
or U2891 (N_2891,N_176,N_121);
and U2892 (N_2892,N_50,N_1562);
and U2893 (N_2893,N_377,N_1371);
nand U2894 (N_2894,N_0,N_1570);
nor U2895 (N_2895,N_1482,N_400);
nand U2896 (N_2896,N_1386,N_1211);
nor U2897 (N_2897,N_415,N_147);
nor U2898 (N_2898,N_441,N_1798);
or U2899 (N_2899,N_1896,N_1864);
and U2900 (N_2900,N_137,N_301);
nand U2901 (N_2901,N_1549,N_349);
nand U2902 (N_2902,N_1924,N_1365);
nor U2903 (N_2903,N_323,N_265);
and U2904 (N_2904,N_3,N_521);
xor U2905 (N_2905,N_758,N_873);
and U2906 (N_2906,N_1964,N_210);
nor U2907 (N_2907,N_442,N_546);
and U2908 (N_2908,N_1696,N_1447);
nor U2909 (N_2909,N_1839,N_1223);
nor U2910 (N_2910,N_721,N_29);
xnor U2911 (N_2911,N_1393,N_1837);
nor U2912 (N_2912,N_1893,N_357);
and U2913 (N_2913,N_631,N_582);
nand U2914 (N_2914,N_1736,N_1362);
nor U2915 (N_2915,N_1978,N_510);
nor U2916 (N_2916,N_114,N_1919);
nand U2917 (N_2917,N_778,N_1239);
or U2918 (N_2918,N_1330,N_1056);
nor U2919 (N_2919,N_1119,N_117);
or U2920 (N_2920,N_1503,N_698);
nor U2921 (N_2921,N_431,N_916);
or U2922 (N_2922,N_1022,N_502);
or U2923 (N_2923,N_229,N_72);
xor U2924 (N_2924,N_987,N_763);
and U2925 (N_2925,N_882,N_1154);
nor U2926 (N_2926,N_434,N_745);
or U2927 (N_2927,N_1221,N_1935);
nor U2928 (N_2928,N_1389,N_412);
or U2929 (N_2929,N_658,N_1275);
and U2930 (N_2930,N_1310,N_1251);
and U2931 (N_2931,N_1133,N_1568);
nand U2932 (N_2932,N_1730,N_651);
or U2933 (N_2933,N_523,N_1125);
nor U2934 (N_2934,N_1082,N_260);
nand U2935 (N_2935,N_1008,N_722);
and U2936 (N_2936,N_557,N_611);
nand U2937 (N_2937,N_429,N_1092);
nand U2938 (N_2938,N_1707,N_533);
nor U2939 (N_2939,N_1411,N_2);
nand U2940 (N_2940,N_340,N_1508);
nor U2941 (N_2941,N_1136,N_1651);
and U2942 (N_2942,N_149,N_1584);
and U2943 (N_2943,N_49,N_1512);
nor U2944 (N_2944,N_513,N_1944);
and U2945 (N_2945,N_85,N_921);
and U2946 (N_2946,N_1794,N_1485);
nand U2947 (N_2947,N_1725,N_590);
and U2948 (N_2948,N_1703,N_115);
and U2949 (N_2949,N_1137,N_39);
nor U2950 (N_2950,N_862,N_424);
or U2951 (N_2951,N_792,N_1907);
nand U2952 (N_2952,N_1727,N_1163);
xor U2953 (N_2953,N_1415,N_1890);
nand U2954 (N_2954,N_1054,N_432);
or U2955 (N_2955,N_539,N_672);
nor U2956 (N_2956,N_1121,N_1348);
or U2957 (N_2957,N_315,N_1439);
and U2958 (N_2958,N_1391,N_465);
nand U2959 (N_2959,N_900,N_420);
nand U2960 (N_2960,N_1383,N_345);
nor U2961 (N_2961,N_1434,N_1952);
or U2962 (N_2962,N_1966,N_885);
nor U2963 (N_2963,N_181,N_1931);
and U2964 (N_2964,N_256,N_1684);
and U2965 (N_2965,N_1234,N_1848);
or U2966 (N_2966,N_58,N_811);
and U2967 (N_2967,N_1585,N_1094);
nand U2968 (N_2968,N_1724,N_1380);
and U2969 (N_2969,N_1936,N_319);
nand U2970 (N_2970,N_1311,N_381);
or U2971 (N_2971,N_1566,N_1109);
nand U2972 (N_2972,N_709,N_1719);
or U2973 (N_2973,N_991,N_769);
nand U2974 (N_2974,N_52,N_670);
nand U2975 (N_2975,N_41,N_1020);
and U2976 (N_2976,N_505,N_314);
or U2977 (N_2977,N_1862,N_569);
or U2978 (N_2978,N_1530,N_1834);
or U2979 (N_2979,N_923,N_199);
or U2980 (N_2980,N_70,N_660);
and U2981 (N_2981,N_975,N_1828);
nand U2982 (N_2982,N_1338,N_12);
nand U2983 (N_2983,N_768,N_618);
xor U2984 (N_2984,N_842,N_1033);
nor U2985 (N_2985,N_1351,N_1370);
nor U2986 (N_2986,N_1442,N_316);
xnor U2987 (N_2987,N_126,N_821);
nand U2988 (N_2988,N_1668,N_1199);
nand U2989 (N_2989,N_1576,N_802);
nand U2990 (N_2990,N_423,N_622);
or U2991 (N_2991,N_35,N_1433);
nor U2992 (N_2992,N_1910,N_1044);
nor U2993 (N_2993,N_481,N_376);
nand U2994 (N_2994,N_471,N_1973);
nor U2995 (N_2995,N_195,N_859);
nor U2996 (N_2996,N_258,N_1742);
and U2997 (N_2997,N_1967,N_14);
nand U2998 (N_2998,N_262,N_1335);
nand U2999 (N_2999,N_40,N_1891);
nor U3000 (N_3000,N_405,N_1537);
nand U3001 (N_3001,N_927,N_1742);
xnor U3002 (N_3002,N_1444,N_1566);
and U3003 (N_3003,N_1130,N_10);
or U3004 (N_3004,N_55,N_750);
or U3005 (N_3005,N_1678,N_1765);
nand U3006 (N_3006,N_1883,N_1435);
or U3007 (N_3007,N_531,N_1773);
nand U3008 (N_3008,N_556,N_1384);
nand U3009 (N_3009,N_131,N_310);
nand U3010 (N_3010,N_1354,N_1276);
nand U3011 (N_3011,N_1065,N_176);
nand U3012 (N_3012,N_1129,N_1312);
or U3013 (N_3013,N_1983,N_1093);
nor U3014 (N_3014,N_1196,N_271);
xnor U3015 (N_3015,N_1702,N_1916);
or U3016 (N_3016,N_1290,N_1601);
or U3017 (N_3017,N_1633,N_1732);
nand U3018 (N_3018,N_321,N_422);
and U3019 (N_3019,N_1098,N_1377);
or U3020 (N_3020,N_1348,N_439);
and U3021 (N_3021,N_1668,N_594);
nand U3022 (N_3022,N_1724,N_1667);
or U3023 (N_3023,N_1628,N_419);
nand U3024 (N_3024,N_201,N_5);
nand U3025 (N_3025,N_56,N_1934);
or U3026 (N_3026,N_325,N_1120);
or U3027 (N_3027,N_149,N_1798);
or U3028 (N_3028,N_1032,N_609);
or U3029 (N_3029,N_1066,N_250);
nand U3030 (N_3030,N_499,N_1186);
and U3031 (N_3031,N_1190,N_1461);
nand U3032 (N_3032,N_725,N_1042);
and U3033 (N_3033,N_1584,N_1243);
and U3034 (N_3034,N_1147,N_1177);
xnor U3035 (N_3035,N_282,N_693);
nor U3036 (N_3036,N_1541,N_70);
and U3037 (N_3037,N_1911,N_77);
xnor U3038 (N_3038,N_163,N_1488);
or U3039 (N_3039,N_534,N_1562);
nand U3040 (N_3040,N_393,N_244);
nand U3041 (N_3041,N_5,N_1904);
and U3042 (N_3042,N_1677,N_1011);
nor U3043 (N_3043,N_6,N_1162);
or U3044 (N_3044,N_734,N_977);
or U3045 (N_3045,N_793,N_1389);
or U3046 (N_3046,N_384,N_373);
nor U3047 (N_3047,N_59,N_1023);
nor U3048 (N_3048,N_724,N_5);
xor U3049 (N_3049,N_836,N_1227);
xor U3050 (N_3050,N_32,N_618);
or U3051 (N_3051,N_868,N_1994);
nand U3052 (N_3052,N_862,N_963);
nor U3053 (N_3053,N_1834,N_210);
and U3054 (N_3054,N_882,N_1690);
nor U3055 (N_3055,N_153,N_1722);
or U3056 (N_3056,N_1904,N_1060);
or U3057 (N_3057,N_693,N_1973);
nor U3058 (N_3058,N_586,N_1251);
or U3059 (N_3059,N_1319,N_647);
nor U3060 (N_3060,N_1233,N_1879);
nand U3061 (N_3061,N_1927,N_715);
and U3062 (N_3062,N_1607,N_695);
xnor U3063 (N_3063,N_1294,N_1485);
nand U3064 (N_3064,N_1604,N_65);
and U3065 (N_3065,N_258,N_871);
or U3066 (N_3066,N_1361,N_1554);
nor U3067 (N_3067,N_73,N_1909);
nand U3068 (N_3068,N_52,N_131);
or U3069 (N_3069,N_322,N_285);
nor U3070 (N_3070,N_526,N_581);
nand U3071 (N_3071,N_1658,N_613);
nand U3072 (N_3072,N_601,N_1029);
nand U3073 (N_3073,N_1175,N_1767);
and U3074 (N_3074,N_1028,N_815);
nor U3075 (N_3075,N_707,N_757);
xnor U3076 (N_3076,N_1685,N_1030);
nand U3077 (N_3077,N_1222,N_135);
nand U3078 (N_3078,N_963,N_251);
nand U3079 (N_3079,N_1920,N_888);
or U3080 (N_3080,N_269,N_1711);
xnor U3081 (N_3081,N_31,N_925);
xnor U3082 (N_3082,N_492,N_53);
and U3083 (N_3083,N_37,N_1681);
nand U3084 (N_3084,N_419,N_630);
and U3085 (N_3085,N_1949,N_996);
and U3086 (N_3086,N_583,N_770);
and U3087 (N_3087,N_492,N_932);
xnor U3088 (N_3088,N_1936,N_1273);
xnor U3089 (N_3089,N_1786,N_409);
or U3090 (N_3090,N_1510,N_1375);
or U3091 (N_3091,N_308,N_1948);
or U3092 (N_3092,N_1004,N_1940);
nor U3093 (N_3093,N_1878,N_1657);
nand U3094 (N_3094,N_293,N_1268);
and U3095 (N_3095,N_293,N_1488);
nand U3096 (N_3096,N_1602,N_596);
xnor U3097 (N_3097,N_806,N_523);
or U3098 (N_3098,N_1236,N_573);
xnor U3099 (N_3099,N_1833,N_716);
nand U3100 (N_3100,N_792,N_1997);
nor U3101 (N_3101,N_1007,N_170);
and U3102 (N_3102,N_1190,N_895);
or U3103 (N_3103,N_100,N_986);
or U3104 (N_3104,N_563,N_496);
nand U3105 (N_3105,N_992,N_1130);
nor U3106 (N_3106,N_779,N_173);
and U3107 (N_3107,N_244,N_1161);
and U3108 (N_3108,N_607,N_1922);
nor U3109 (N_3109,N_463,N_1124);
nor U3110 (N_3110,N_204,N_970);
and U3111 (N_3111,N_1445,N_517);
xor U3112 (N_3112,N_1696,N_608);
or U3113 (N_3113,N_621,N_1789);
or U3114 (N_3114,N_1125,N_391);
nor U3115 (N_3115,N_1376,N_79);
nor U3116 (N_3116,N_1531,N_1791);
or U3117 (N_3117,N_63,N_1302);
nand U3118 (N_3118,N_1103,N_534);
and U3119 (N_3119,N_1441,N_1423);
nand U3120 (N_3120,N_1913,N_14);
nand U3121 (N_3121,N_253,N_942);
and U3122 (N_3122,N_212,N_1585);
nand U3123 (N_3123,N_482,N_1346);
nor U3124 (N_3124,N_957,N_1990);
nor U3125 (N_3125,N_788,N_1245);
or U3126 (N_3126,N_1825,N_1618);
xnor U3127 (N_3127,N_217,N_729);
nand U3128 (N_3128,N_855,N_96);
xnor U3129 (N_3129,N_77,N_549);
nor U3130 (N_3130,N_237,N_263);
nor U3131 (N_3131,N_535,N_818);
or U3132 (N_3132,N_537,N_1464);
and U3133 (N_3133,N_289,N_1682);
and U3134 (N_3134,N_1666,N_394);
or U3135 (N_3135,N_863,N_64);
or U3136 (N_3136,N_1535,N_1665);
nor U3137 (N_3137,N_468,N_1846);
nor U3138 (N_3138,N_213,N_780);
nor U3139 (N_3139,N_878,N_109);
or U3140 (N_3140,N_569,N_1827);
and U3141 (N_3141,N_1304,N_1174);
nor U3142 (N_3142,N_504,N_389);
and U3143 (N_3143,N_1347,N_664);
or U3144 (N_3144,N_797,N_1806);
nand U3145 (N_3145,N_14,N_1766);
and U3146 (N_3146,N_1237,N_548);
xor U3147 (N_3147,N_1563,N_1055);
nor U3148 (N_3148,N_1979,N_198);
nor U3149 (N_3149,N_1705,N_1033);
or U3150 (N_3150,N_311,N_1870);
or U3151 (N_3151,N_688,N_735);
or U3152 (N_3152,N_700,N_1111);
or U3153 (N_3153,N_1972,N_358);
and U3154 (N_3154,N_1188,N_1361);
nand U3155 (N_3155,N_1520,N_1669);
nor U3156 (N_3156,N_836,N_1677);
nand U3157 (N_3157,N_1349,N_1540);
xor U3158 (N_3158,N_33,N_606);
nor U3159 (N_3159,N_1905,N_1585);
nor U3160 (N_3160,N_1580,N_1824);
or U3161 (N_3161,N_1682,N_713);
xor U3162 (N_3162,N_1838,N_1397);
nand U3163 (N_3163,N_1352,N_1226);
or U3164 (N_3164,N_103,N_502);
and U3165 (N_3165,N_1439,N_795);
or U3166 (N_3166,N_42,N_1203);
nor U3167 (N_3167,N_1994,N_532);
and U3168 (N_3168,N_1117,N_977);
xor U3169 (N_3169,N_510,N_1917);
xor U3170 (N_3170,N_1994,N_959);
and U3171 (N_3171,N_1194,N_1297);
or U3172 (N_3172,N_450,N_65);
nor U3173 (N_3173,N_1857,N_1990);
or U3174 (N_3174,N_906,N_246);
and U3175 (N_3175,N_964,N_1424);
and U3176 (N_3176,N_71,N_1144);
or U3177 (N_3177,N_1222,N_1027);
xnor U3178 (N_3178,N_1701,N_1811);
or U3179 (N_3179,N_1416,N_1533);
nor U3180 (N_3180,N_512,N_114);
and U3181 (N_3181,N_1094,N_669);
or U3182 (N_3182,N_1859,N_343);
or U3183 (N_3183,N_1175,N_156);
nand U3184 (N_3184,N_7,N_1209);
xnor U3185 (N_3185,N_497,N_1208);
nand U3186 (N_3186,N_760,N_775);
nor U3187 (N_3187,N_1914,N_1626);
nand U3188 (N_3188,N_1335,N_1130);
xor U3189 (N_3189,N_1752,N_1244);
nor U3190 (N_3190,N_1541,N_1240);
and U3191 (N_3191,N_888,N_1612);
or U3192 (N_3192,N_771,N_122);
nand U3193 (N_3193,N_1141,N_1803);
or U3194 (N_3194,N_474,N_861);
or U3195 (N_3195,N_713,N_1350);
and U3196 (N_3196,N_1553,N_1081);
and U3197 (N_3197,N_1675,N_1291);
or U3198 (N_3198,N_1965,N_830);
and U3199 (N_3199,N_97,N_1452);
nand U3200 (N_3200,N_40,N_954);
or U3201 (N_3201,N_834,N_588);
nor U3202 (N_3202,N_1733,N_409);
nor U3203 (N_3203,N_650,N_1032);
xor U3204 (N_3204,N_1599,N_96);
or U3205 (N_3205,N_1157,N_1670);
or U3206 (N_3206,N_906,N_1561);
or U3207 (N_3207,N_25,N_1060);
and U3208 (N_3208,N_546,N_382);
xnor U3209 (N_3209,N_864,N_1030);
and U3210 (N_3210,N_247,N_1383);
and U3211 (N_3211,N_475,N_1740);
and U3212 (N_3212,N_244,N_511);
nand U3213 (N_3213,N_1700,N_1662);
or U3214 (N_3214,N_1661,N_1377);
xnor U3215 (N_3215,N_415,N_1470);
nor U3216 (N_3216,N_1789,N_1487);
nor U3217 (N_3217,N_1946,N_1762);
nand U3218 (N_3218,N_323,N_865);
xor U3219 (N_3219,N_159,N_359);
or U3220 (N_3220,N_1165,N_275);
nand U3221 (N_3221,N_113,N_396);
and U3222 (N_3222,N_1049,N_95);
xnor U3223 (N_3223,N_946,N_42);
nand U3224 (N_3224,N_998,N_830);
and U3225 (N_3225,N_1833,N_1609);
nor U3226 (N_3226,N_621,N_96);
xnor U3227 (N_3227,N_1093,N_641);
nor U3228 (N_3228,N_1527,N_1926);
and U3229 (N_3229,N_1420,N_105);
and U3230 (N_3230,N_369,N_81);
xor U3231 (N_3231,N_116,N_1493);
or U3232 (N_3232,N_367,N_1911);
or U3233 (N_3233,N_1803,N_758);
nand U3234 (N_3234,N_1953,N_1265);
or U3235 (N_3235,N_537,N_989);
or U3236 (N_3236,N_327,N_281);
nor U3237 (N_3237,N_476,N_1126);
xnor U3238 (N_3238,N_624,N_396);
nand U3239 (N_3239,N_556,N_292);
nor U3240 (N_3240,N_1244,N_1513);
nor U3241 (N_3241,N_594,N_1009);
nor U3242 (N_3242,N_54,N_611);
and U3243 (N_3243,N_301,N_1044);
or U3244 (N_3244,N_449,N_321);
nor U3245 (N_3245,N_610,N_1875);
nand U3246 (N_3246,N_1509,N_1859);
nand U3247 (N_3247,N_1484,N_1584);
and U3248 (N_3248,N_1136,N_1010);
nor U3249 (N_3249,N_1229,N_1182);
nor U3250 (N_3250,N_788,N_676);
or U3251 (N_3251,N_1804,N_1878);
and U3252 (N_3252,N_745,N_1175);
xor U3253 (N_3253,N_1169,N_175);
or U3254 (N_3254,N_1508,N_742);
nand U3255 (N_3255,N_930,N_285);
nor U3256 (N_3256,N_1745,N_1094);
nand U3257 (N_3257,N_544,N_851);
xor U3258 (N_3258,N_1574,N_203);
or U3259 (N_3259,N_467,N_219);
or U3260 (N_3260,N_435,N_53);
nor U3261 (N_3261,N_66,N_1178);
nand U3262 (N_3262,N_1362,N_1094);
and U3263 (N_3263,N_517,N_80);
nor U3264 (N_3264,N_1131,N_837);
xnor U3265 (N_3265,N_551,N_188);
and U3266 (N_3266,N_108,N_592);
or U3267 (N_3267,N_430,N_206);
or U3268 (N_3268,N_58,N_1266);
or U3269 (N_3269,N_197,N_984);
xnor U3270 (N_3270,N_396,N_1695);
nor U3271 (N_3271,N_448,N_9);
or U3272 (N_3272,N_1418,N_935);
or U3273 (N_3273,N_1286,N_635);
or U3274 (N_3274,N_378,N_1766);
and U3275 (N_3275,N_123,N_340);
or U3276 (N_3276,N_274,N_760);
or U3277 (N_3277,N_1142,N_1454);
or U3278 (N_3278,N_1168,N_865);
nand U3279 (N_3279,N_1005,N_659);
or U3280 (N_3280,N_788,N_1819);
nor U3281 (N_3281,N_1966,N_1697);
or U3282 (N_3282,N_1897,N_955);
nand U3283 (N_3283,N_1255,N_1897);
or U3284 (N_3284,N_1391,N_1349);
nand U3285 (N_3285,N_1443,N_526);
xor U3286 (N_3286,N_206,N_1599);
and U3287 (N_3287,N_581,N_353);
nand U3288 (N_3288,N_412,N_702);
and U3289 (N_3289,N_737,N_1371);
or U3290 (N_3290,N_711,N_849);
nor U3291 (N_3291,N_1887,N_1694);
or U3292 (N_3292,N_827,N_1790);
nor U3293 (N_3293,N_1128,N_1502);
nand U3294 (N_3294,N_422,N_735);
and U3295 (N_3295,N_864,N_1150);
nor U3296 (N_3296,N_220,N_832);
or U3297 (N_3297,N_1456,N_36);
nor U3298 (N_3298,N_792,N_217);
or U3299 (N_3299,N_1175,N_1894);
nand U3300 (N_3300,N_1723,N_1805);
and U3301 (N_3301,N_1316,N_1073);
or U3302 (N_3302,N_1042,N_514);
nor U3303 (N_3303,N_1834,N_206);
nand U3304 (N_3304,N_674,N_1890);
nor U3305 (N_3305,N_575,N_803);
and U3306 (N_3306,N_731,N_1133);
or U3307 (N_3307,N_935,N_1175);
nor U3308 (N_3308,N_756,N_416);
and U3309 (N_3309,N_579,N_1320);
or U3310 (N_3310,N_973,N_1384);
xnor U3311 (N_3311,N_772,N_1281);
nor U3312 (N_3312,N_17,N_26);
nand U3313 (N_3313,N_1200,N_1849);
nand U3314 (N_3314,N_612,N_493);
nand U3315 (N_3315,N_839,N_1472);
xor U3316 (N_3316,N_1940,N_440);
nor U3317 (N_3317,N_870,N_444);
and U3318 (N_3318,N_1389,N_1113);
nand U3319 (N_3319,N_1119,N_4);
or U3320 (N_3320,N_1029,N_709);
nor U3321 (N_3321,N_1853,N_1845);
nand U3322 (N_3322,N_1241,N_1455);
nand U3323 (N_3323,N_571,N_1091);
or U3324 (N_3324,N_1052,N_1035);
nand U3325 (N_3325,N_126,N_67);
nor U3326 (N_3326,N_548,N_704);
or U3327 (N_3327,N_1543,N_180);
nor U3328 (N_3328,N_436,N_773);
or U3329 (N_3329,N_50,N_1605);
nand U3330 (N_3330,N_293,N_1859);
and U3331 (N_3331,N_1376,N_472);
or U3332 (N_3332,N_1711,N_514);
and U3333 (N_3333,N_1779,N_926);
nor U3334 (N_3334,N_1728,N_242);
nand U3335 (N_3335,N_1571,N_759);
nor U3336 (N_3336,N_587,N_264);
and U3337 (N_3337,N_60,N_416);
or U3338 (N_3338,N_1159,N_1545);
nor U3339 (N_3339,N_675,N_1299);
nand U3340 (N_3340,N_1051,N_185);
nor U3341 (N_3341,N_1184,N_1731);
xor U3342 (N_3342,N_1432,N_1589);
or U3343 (N_3343,N_1919,N_1974);
or U3344 (N_3344,N_147,N_307);
nor U3345 (N_3345,N_551,N_677);
nor U3346 (N_3346,N_460,N_1721);
or U3347 (N_3347,N_1418,N_1748);
nor U3348 (N_3348,N_873,N_1769);
nor U3349 (N_3349,N_1748,N_1570);
or U3350 (N_3350,N_438,N_1472);
and U3351 (N_3351,N_688,N_408);
nor U3352 (N_3352,N_294,N_16);
nand U3353 (N_3353,N_1345,N_588);
and U3354 (N_3354,N_223,N_1847);
or U3355 (N_3355,N_1361,N_1463);
nor U3356 (N_3356,N_1079,N_156);
nand U3357 (N_3357,N_1889,N_1862);
xor U3358 (N_3358,N_958,N_497);
nand U3359 (N_3359,N_757,N_1451);
nand U3360 (N_3360,N_414,N_340);
xnor U3361 (N_3361,N_464,N_280);
nand U3362 (N_3362,N_475,N_462);
nand U3363 (N_3363,N_1063,N_1449);
nor U3364 (N_3364,N_1566,N_763);
nand U3365 (N_3365,N_252,N_1004);
or U3366 (N_3366,N_1962,N_580);
nand U3367 (N_3367,N_1984,N_8);
nor U3368 (N_3368,N_1807,N_1166);
nor U3369 (N_3369,N_1551,N_362);
nand U3370 (N_3370,N_854,N_732);
nor U3371 (N_3371,N_1339,N_1569);
nand U3372 (N_3372,N_254,N_132);
and U3373 (N_3373,N_201,N_554);
nor U3374 (N_3374,N_893,N_1280);
nor U3375 (N_3375,N_904,N_1146);
nor U3376 (N_3376,N_1857,N_455);
nor U3377 (N_3377,N_411,N_1345);
and U3378 (N_3378,N_1476,N_1658);
and U3379 (N_3379,N_503,N_1049);
nand U3380 (N_3380,N_900,N_67);
nor U3381 (N_3381,N_1245,N_946);
or U3382 (N_3382,N_340,N_310);
and U3383 (N_3383,N_5,N_645);
nand U3384 (N_3384,N_1925,N_616);
nor U3385 (N_3385,N_705,N_1189);
and U3386 (N_3386,N_623,N_1646);
nand U3387 (N_3387,N_851,N_750);
or U3388 (N_3388,N_964,N_567);
and U3389 (N_3389,N_1503,N_297);
and U3390 (N_3390,N_1123,N_699);
xor U3391 (N_3391,N_157,N_223);
and U3392 (N_3392,N_1806,N_669);
xnor U3393 (N_3393,N_1171,N_997);
and U3394 (N_3394,N_201,N_1711);
and U3395 (N_3395,N_1877,N_772);
and U3396 (N_3396,N_1083,N_279);
nand U3397 (N_3397,N_536,N_172);
or U3398 (N_3398,N_1533,N_23);
nand U3399 (N_3399,N_1054,N_1841);
and U3400 (N_3400,N_270,N_654);
nor U3401 (N_3401,N_277,N_1079);
or U3402 (N_3402,N_1082,N_1225);
xnor U3403 (N_3403,N_1964,N_1455);
nor U3404 (N_3404,N_1435,N_1251);
nand U3405 (N_3405,N_718,N_143);
and U3406 (N_3406,N_1261,N_1800);
or U3407 (N_3407,N_1678,N_638);
or U3408 (N_3408,N_1922,N_1614);
nand U3409 (N_3409,N_897,N_1894);
nor U3410 (N_3410,N_1725,N_1745);
nor U3411 (N_3411,N_1685,N_109);
xor U3412 (N_3412,N_1543,N_942);
nand U3413 (N_3413,N_1914,N_817);
nor U3414 (N_3414,N_929,N_913);
nor U3415 (N_3415,N_502,N_1178);
xnor U3416 (N_3416,N_1255,N_1998);
nand U3417 (N_3417,N_930,N_1530);
nand U3418 (N_3418,N_710,N_620);
xnor U3419 (N_3419,N_464,N_1398);
xor U3420 (N_3420,N_1795,N_1181);
or U3421 (N_3421,N_1980,N_758);
and U3422 (N_3422,N_131,N_1452);
nand U3423 (N_3423,N_1644,N_551);
nor U3424 (N_3424,N_1235,N_1919);
nor U3425 (N_3425,N_1576,N_768);
nand U3426 (N_3426,N_23,N_525);
or U3427 (N_3427,N_1673,N_63);
or U3428 (N_3428,N_896,N_1977);
xor U3429 (N_3429,N_1205,N_188);
and U3430 (N_3430,N_1060,N_868);
and U3431 (N_3431,N_717,N_1194);
nand U3432 (N_3432,N_1646,N_1701);
nor U3433 (N_3433,N_43,N_967);
xor U3434 (N_3434,N_1684,N_1406);
nand U3435 (N_3435,N_702,N_1496);
nor U3436 (N_3436,N_1977,N_676);
and U3437 (N_3437,N_1337,N_701);
nor U3438 (N_3438,N_1522,N_1085);
nand U3439 (N_3439,N_1692,N_1049);
nand U3440 (N_3440,N_1249,N_471);
and U3441 (N_3441,N_1497,N_1404);
and U3442 (N_3442,N_528,N_502);
nor U3443 (N_3443,N_33,N_1023);
and U3444 (N_3444,N_921,N_1039);
xnor U3445 (N_3445,N_648,N_1545);
nand U3446 (N_3446,N_1121,N_525);
or U3447 (N_3447,N_245,N_1243);
nand U3448 (N_3448,N_1610,N_289);
nand U3449 (N_3449,N_1151,N_1801);
nor U3450 (N_3450,N_443,N_534);
xnor U3451 (N_3451,N_393,N_425);
or U3452 (N_3452,N_1591,N_766);
and U3453 (N_3453,N_1763,N_1132);
nor U3454 (N_3454,N_1989,N_482);
nor U3455 (N_3455,N_1281,N_956);
nand U3456 (N_3456,N_1615,N_1788);
or U3457 (N_3457,N_1336,N_228);
nand U3458 (N_3458,N_1077,N_586);
and U3459 (N_3459,N_268,N_210);
and U3460 (N_3460,N_190,N_505);
or U3461 (N_3461,N_1147,N_1652);
or U3462 (N_3462,N_289,N_421);
or U3463 (N_3463,N_1533,N_710);
nor U3464 (N_3464,N_106,N_1103);
or U3465 (N_3465,N_951,N_1721);
and U3466 (N_3466,N_1824,N_1787);
and U3467 (N_3467,N_841,N_102);
nor U3468 (N_3468,N_1313,N_949);
and U3469 (N_3469,N_1241,N_53);
and U3470 (N_3470,N_1007,N_1608);
nor U3471 (N_3471,N_232,N_1285);
nor U3472 (N_3472,N_247,N_697);
and U3473 (N_3473,N_1629,N_483);
nor U3474 (N_3474,N_412,N_990);
or U3475 (N_3475,N_897,N_290);
and U3476 (N_3476,N_89,N_1017);
xor U3477 (N_3477,N_1907,N_1619);
or U3478 (N_3478,N_276,N_1707);
nand U3479 (N_3479,N_107,N_890);
or U3480 (N_3480,N_1860,N_889);
xor U3481 (N_3481,N_584,N_478);
nor U3482 (N_3482,N_1443,N_304);
xnor U3483 (N_3483,N_1344,N_582);
nor U3484 (N_3484,N_1954,N_405);
nand U3485 (N_3485,N_877,N_29);
or U3486 (N_3486,N_582,N_54);
xor U3487 (N_3487,N_1370,N_1411);
and U3488 (N_3488,N_1998,N_724);
xnor U3489 (N_3489,N_1370,N_796);
and U3490 (N_3490,N_312,N_496);
nand U3491 (N_3491,N_947,N_1578);
xor U3492 (N_3492,N_96,N_241);
and U3493 (N_3493,N_1446,N_868);
nor U3494 (N_3494,N_1258,N_590);
or U3495 (N_3495,N_424,N_1247);
nand U3496 (N_3496,N_674,N_1536);
nor U3497 (N_3497,N_66,N_1047);
nand U3498 (N_3498,N_458,N_1781);
nand U3499 (N_3499,N_1917,N_1041);
nor U3500 (N_3500,N_1813,N_942);
nand U3501 (N_3501,N_1464,N_1495);
or U3502 (N_3502,N_1259,N_1736);
nor U3503 (N_3503,N_1567,N_1283);
or U3504 (N_3504,N_196,N_1308);
or U3505 (N_3505,N_951,N_1416);
or U3506 (N_3506,N_1576,N_1463);
nor U3507 (N_3507,N_113,N_713);
or U3508 (N_3508,N_905,N_1023);
nor U3509 (N_3509,N_1918,N_1912);
and U3510 (N_3510,N_1222,N_1278);
xor U3511 (N_3511,N_161,N_37);
nand U3512 (N_3512,N_417,N_857);
or U3513 (N_3513,N_1114,N_824);
and U3514 (N_3514,N_1324,N_111);
and U3515 (N_3515,N_138,N_1055);
or U3516 (N_3516,N_34,N_54);
or U3517 (N_3517,N_1811,N_1719);
or U3518 (N_3518,N_2,N_1364);
or U3519 (N_3519,N_928,N_1872);
and U3520 (N_3520,N_1586,N_1079);
or U3521 (N_3521,N_1668,N_174);
nand U3522 (N_3522,N_1771,N_1420);
and U3523 (N_3523,N_330,N_731);
and U3524 (N_3524,N_1352,N_1710);
nand U3525 (N_3525,N_340,N_104);
nand U3526 (N_3526,N_797,N_202);
nor U3527 (N_3527,N_1309,N_859);
and U3528 (N_3528,N_1828,N_948);
or U3529 (N_3529,N_1596,N_442);
nor U3530 (N_3530,N_1466,N_979);
nor U3531 (N_3531,N_760,N_1842);
nor U3532 (N_3532,N_1854,N_1251);
nand U3533 (N_3533,N_1739,N_915);
or U3534 (N_3534,N_1153,N_1281);
and U3535 (N_3535,N_1186,N_1518);
and U3536 (N_3536,N_1440,N_731);
and U3537 (N_3537,N_488,N_198);
and U3538 (N_3538,N_118,N_123);
nand U3539 (N_3539,N_1786,N_1525);
or U3540 (N_3540,N_917,N_240);
or U3541 (N_3541,N_1783,N_1450);
or U3542 (N_3542,N_1642,N_595);
or U3543 (N_3543,N_1834,N_831);
nand U3544 (N_3544,N_1884,N_774);
and U3545 (N_3545,N_1206,N_1225);
nor U3546 (N_3546,N_1213,N_293);
or U3547 (N_3547,N_1538,N_1793);
nor U3548 (N_3548,N_1047,N_1800);
or U3549 (N_3549,N_1387,N_1857);
nor U3550 (N_3550,N_1741,N_1538);
nor U3551 (N_3551,N_1017,N_1682);
nand U3552 (N_3552,N_917,N_1683);
xor U3553 (N_3553,N_7,N_273);
xor U3554 (N_3554,N_1082,N_1041);
or U3555 (N_3555,N_1721,N_1740);
nor U3556 (N_3556,N_274,N_354);
and U3557 (N_3557,N_1398,N_291);
or U3558 (N_3558,N_350,N_697);
or U3559 (N_3559,N_1321,N_966);
nor U3560 (N_3560,N_662,N_234);
nor U3561 (N_3561,N_1038,N_1404);
and U3562 (N_3562,N_1926,N_1183);
nand U3563 (N_3563,N_1133,N_1703);
and U3564 (N_3564,N_1121,N_582);
xor U3565 (N_3565,N_948,N_633);
nor U3566 (N_3566,N_1755,N_1604);
nor U3567 (N_3567,N_993,N_237);
nand U3568 (N_3568,N_5,N_446);
nand U3569 (N_3569,N_958,N_724);
nor U3570 (N_3570,N_1412,N_1588);
nor U3571 (N_3571,N_582,N_944);
nor U3572 (N_3572,N_917,N_1902);
xor U3573 (N_3573,N_1368,N_1715);
nor U3574 (N_3574,N_681,N_1788);
and U3575 (N_3575,N_648,N_1810);
nand U3576 (N_3576,N_1632,N_1766);
nand U3577 (N_3577,N_734,N_985);
and U3578 (N_3578,N_1352,N_481);
nand U3579 (N_3579,N_1927,N_377);
or U3580 (N_3580,N_541,N_1357);
nand U3581 (N_3581,N_618,N_1081);
nor U3582 (N_3582,N_1657,N_1495);
nor U3583 (N_3583,N_580,N_604);
nor U3584 (N_3584,N_1816,N_1244);
and U3585 (N_3585,N_451,N_426);
nor U3586 (N_3586,N_1958,N_998);
nor U3587 (N_3587,N_1928,N_1455);
nor U3588 (N_3588,N_1303,N_1190);
and U3589 (N_3589,N_997,N_537);
or U3590 (N_3590,N_1636,N_234);
nand U3591 (N_3591,N_1791,N_850);
or U3592 (N_3592,N_597,N_112);
and U3593 (N_3593,N_738,N_1329);
xnor U3594 (N_3594,N_1677,N_1406);
or U3595 (N_3595,N_1277,N_482);
nor U3596 (N_3596,N_95,N_1306);
or U3597 (N_3597,N_970,N_630);
nor U3598 (N_3598,N_1024,N_992);
or U3599 (N_3599,N_1038,N_200);
nand U3600 (N_3600,N_112,N_1921);
and U3601 (N_3601,N_380,N_858);
nand U3602 (N_3602,N_1025,N_1128);
nand U3603 (N_3603,N_1826,N_1305);
nand U3604 (N_3604,N_80,N_641);
nor U3605 (N_3605,N_643,N_593);
nand U3606 (N_3606,N_299,N_1504);
nand U3607 (N_3607,N_1091,N_6);
or U3608 (N_3608,N_1540,N_1979);
nor U3609 (N_3609,N_877,N_1707);
and U3610 (N_3610,N_16,N_1157);
nor U3611 (N_3611,N_1982,N_685);
or U3612 (N_3612,N_233,N_1113);
nand U3613 (N_3613,N_293,N_1920);
nor U3614 (N_3614,N_1804,N_15);
and U3615 (N_3615,N_1232,N_1955);
nand U3616 (N_3616,N_1127,N_1185);
and U3617 (N_3617,N_1692,N_607);
and U3618 (N_3618,N_963,N_495);
nand U3619 (N_3619,N_1151,N_412);
and U3620 (N_3620,N_756,N_1891);
nor U3621 (N_3621,N_1864,N_1737);
xor U3622 (N_3622,N_158,N_1812);
nor U3623 (N_3623,N_1705,N_1973);
nor U3624 (N_3624,N_747,N_1975);
xnor U3625 (N_3625,N_1993,N_22);
nand U3626 (N_3626,N_1141,N_1285);
xnor U3627 (N_3627,N_1800,N_1711);
nor U3628 (N_3628,N_146,N_1615);
nor U3629 (N_3629,N_52,N_1533);
nand U3630 (N_3630,N_27,N_356);
nor U3631 (N_3631,N_653,N_1366);
xnor U3632 (N_3632,N_1907,N_500);
nand U3633 (N_3633,N_1738,N_421);
and U3634 (N_3634,N_1098,N_440);
nand U3635 (N_3635,N_1026,N_181);
or U3636 (N_3636,N_1946,N_324);
xor U3637 (N_3637,N_730,N_1687);
and U3638 (N_3638,N_1514,N_212);
xnor U3639 (N_3639,N_1202,N_1527);
or U3640 (N_3640,N_465,N_1173);
nor U3641 (N_3641,N_1441,N_643);
or U3642 (N_3642,N_1272,N_264);
nand U3643 (N_3643,N_169,N_526);
nand U3644 (N_3644,N_1748,N_675);
nor U3645 (N_3645,N_1961,N_1514);
xor U3646 (N_3646,N_1068,N_235);
xor U3647 (N_3647,N_1801,N_977);
and U3648 (N_3648,N_78,N_1870);
and U3649 (N_3649,N_817,N_710);
nand U3650 (N_3650,N_1203,N_289);
or U3651 (N_3651,N_1897,N_1169);
and U3652 (N_3652,N_1347,N_1751);
nor U3653 (N_3653,N_1188,N_515);
nor U3654 (N_3654,N_21,N_364);
or U3655 (N_3655,N_1050,N_1743);
and U3656 (N_3656,N_925,N_1591);
and U3657 (N_3657,N_1610,N_986);
and U3658 (N_3658,N_285,N_1942);
xnor U3659 (N_3659,N_668,N_1975);
or U3660 (N_3660,N_961,N_65);
nor U3661 (N_3661,N_1244,N_1990);
or U3662 (N_3662,N_1607,N_1437);
and U3663 (N_3663,N_601,N_686);
or U3664 (N_3664,N_1737,N_1227);
and U3665 (N_3665,N_1767,N_1000);
and U3666 (N_3666,N_1940,N_866);
or U3667 (N_3667,N_1402,N_167);
and U3668 (N_3668,N_909,N_1947);
nor U3669 (N_3669,N_1366,N_1296);
nand U3670 (N_3670,N_763,N_850);
xnor U3671 (N_3671,N_1792,N_576);
nand U3672 (N_3672,N_689,N_315);
and U3673 (N_3673,N_1541,N_288);
xor U3674 (N_3674,N_1861,N_626);
nor U3675 (N_3675,N_969,N_146);
nand U3676 (N_3676,N_1945,N_1221);
xnor U3677 (N_3677,N_1315,N_529);
or U3678 (N_3678,N_188,N_443);
xor U3679 (N_3679,N_1874,N_1575);
nand U3680 (N_3680,N_1939,N_371);
nor U3681 (N_3681,N_1584,N_678);
and U3682 (N_3682,N_1098,N_412);
or U3683 (N_3683,N_13,N_93);
and U3684 (N_3684,N_314,N_1129);
or U3685 (N_3685,N_230,N_1701);
or U3686 (N_3686,N_1088,N_73);
and U3687 (N_3687,N_1348,N_130);
xnor U3688 (N_3688,N_114,N_269);
nand U3689 (N_3689,N_1242,N_177);
xnor U3690 (N_3690,N_1425,N_1586);
nor U3691 (N_3691,N_1746,N_31);
nor U3692 (N_3692,N_1873,N_345);
nor U3693 (N_3693,N_1959,N_352);
nor U3694 (N_3694,N_854,N_1735);
nor U3695 (N_3695,N_238,N_528);
nor U3696 (N_3696,N_1899,N_1944);
nor U3697 (N_3697,N_1745,N_1529);
nand U3698 (N_3698,N_938,N_1268);
or U3699 (N_3699,N_662,N_1254);
nor U3700 (N_3700,N_1397,N_1592);
and U3701 (N_3701,N_1667,N_1577);
xor U3702 (N_3702,N_1604,N_549);
nand U3703 (N_3703,N_1509,N_696);
nor U3704 (N_3704,N_1828,N_80);
nor U3705 (N_3705,N_1965,N_151);
xor U3706 (N_3706,N_156,N_1559);
nor U3707 (N_3707,N_1483,N_1595);
or U3708 (N_3708,N_1023,N_676);
or U3709 (N_3709,N_126,N_264);
xor U3710 (N_3710,N_1335,N_1244);
and U3711 (N_3711,N_1644,N_1601);
nand U3712 (N_3712,N_424,N_1041);
nand U3713 (N_3713,N_227,N_541);
nor U3714 (N_3714,N_1275,N_373);
nand U3715 (N_3715,N_866,N_885);
nor U3716 (N_3716,N_881,N_216);
or U3717 (N_3717,N_183,N_1849);
xor U3718 (N_3718,N_1880,N_520);
and U3719 (N_3719,N_1087,N_276);
or U3720 (N_3720,N_170,N_1364);
or U3721 (N_3721,N_1180,N_1642);
or U3722 (N_3722,N_804,N_679);
nor U3723 (N_3723,N_379,N_670);
and U3724 (N_3724,N_478,N_792);
and U3725 (N_3725,N_584,N_146);
nor U3726 (N_3726,N_130,N_155);
nand U3727 (N_3727,N_1239,N_584);
nand U3728 (N_3728,N_1782,N_1792);
xor U3729 (N_3729,N_1927,N_741);
nor U3730 (N_3730,N_1552,N_1228);
or U3731 (N_3731,N_1622,N_753);
or U3732 (N_3732,N_688,N_957);
and U3733 (N_3733,N_640,N_1162);
or U3734 (N_3734,N_453,N_1027);
and U3735 (N_3735,N_1811,N_1625);
nand U3736 (N_3736,N_1255,N_1764);
or U3737 (N_3737,N_862,N_974);
nand U3738 (N_3738,N_884,N_1657);
nand U3739 (N_3739,N_1878,N_1464);
nor U3740 (N_3740,N_1191,N_1991);
nor U3741 (N_3741,N_1087,N_1115);
nand U3742 (N_3742,N_1276,N_1167);
and U3743 (N_3743,N_1834,N_718);
and U3744 (N_3744,N_469,N_291);
and U3745 (N_3745,N_1986,N_426);
or U3746 (N_3746,N_1829,N_877);
nand U3747 (N_3747,N_4,N_1122);
and U3748 (N_3748,N_659,N_1262);
nand U3749 (N_3749,N_1995,N_1303);
or U3750 (N_3750,N_1405,N_649);
nand U3751 (N_3751,N_887,N_136);
xnor U3752 (N_3752,N_1998,N_116);
nand U3753 (N_3753,N_1650,N_1459);
nand U3754 (N_3754,N_1664,N_301);
nor U3755 (N_3755,N_1586,N_796);
and U3756 (N_3756,N_1054,N_1064);
or U3757 (N_3757,N_1608,N_1414);
and U3758 (N_3758,N_1772,N_1442);
nor U3759 (N_3759,N_958,N_233);
or U3760 (N_3760,N_979,N_681);
nor U3761 (N_3761,N_708,N_1451);
nor U3762 (N_3762,N_1125,N_1839);
or U3763 (N_3763,N_538,N_62);
or U3764 (N_3764,N_1477,N_1602);
or U3765 (N_3765,N_97,N_1636);
nor U3766 (N_3766,N_322,N_1196);
nand U3767 (N_3767,N_1593,N_473);
nand U3768 (N_3768,N_65,N_1813);
nor U3769 (N_3769,N_1421,N_278);
xnor U3770 (N_3770,N_1444,N_530);
and U3771 (N_3771,N_905,N_1981);
nand U3772 (N_3772,N_1680,N_1041);
or U3773 (N_3773,N_1057,N_444);
or U3774 (N_3774,N_785,N_1976);
and U3775 (N_3775,N_986,N_1580);
nand U3776 (N_3776,N_957,N_348);
nor U3777 (N_3777,N_1058,N_599);
and U3778 (N_3778,N_703,N_230);
nor U3779 (N_3779,N_1028,N_692);
or U3780 (N_3780,N_1184,N_330);
and U3781 (N_3781,N_292,N_1166);
or U3782 (N_3782,N_1514,N_613);
nor U3783 (N_3783,N_1898,N_1598);
nor U3784 (N_3784,N_791,N_1931);
nor U3785 (N_3785,N_660,N_969);
or U3786 (N_3786,N_1966,N_591);
or U3787 (N_3787,N_695,N_1394);
or U3788 (N_3788,N_912,N_1344);
or U3789 (N_3789,N_608,N_1837);
and U3790 (N_3790,N_1722,N_581);
nor U3791 (N_3791,N_820,N_1496);
nor U3792 (N_3792,N_562,N_493);
xor U3793 (N_3793,N_29,N_980);
or U3794 (N_3794,N_1560,N_1781);
nand U3795 (N_3795,N_732,N_202);
or U3796 (N_3796,N_1007,N_903);
nand U3797 (N_3797,N_1072,N_220);
nor U3798 (N_3798,N_1044,N_1732);
and U3799 (N_3799,N_625,N_216);
nand U3800 (N_3800,N_1190,N_545);
and U3801 (N_3801,N_1696,N_1318);
or U3802 (N_3802,N_211,N_993);
and U3803 (N_3803,N_763,N_1959);
nor U3804 (N_3804,N_1949,N_71);
nand U3805 (N_3805,N_1292,N_1726);
or U3806 (N_3806,N_336,N_52);
and U3807 (N_3807,N_1602,N_1044);
nand U3808 (N_3808,N_291,N_981);
xor U3809 (N_3809,N_3,N_1128);
nand U3810 (N_3810,N_1533,N_75);
xor U3811 (N_3811,N_904,N_447);
or U3812 (N_3812,N_737,N_1853);
nand U3813 (N_3813,N_1499,N_1284);
or U3814 (N_3814,N_832,N_378);
or U3815 (N_3815,N_520,N_1291);
nand U3816 (N_3816,N_1602,N_831);
nand U3817 (N_3817,N_444,N_1365);
nand U3818 (N_3818,N_1960,N_143);
nand U3819 (N_3819,N_71,N_337);
nor U3820 (N_3820,N_992,N_1925);
nor U3821 (N_3821,N_959,N_1285);
nand U3822 (N_3822,N_1587,N_1183);
nor U3823 (N_3823,N_814,N_1213);
nor U3824 (N_3824,N_1448,N_616);
nand U3825 (N_3825,N_1626,N_1755);
nor U3826 (N_3826,N_902,N_193);
and U3827 (N_3827,N_114,N_233);
or U3828 (N_3828,N_1447,N_490);
xor U3829 (N_3829,N_1011,N_1047);
xor U3830 (N_3830,N_1080,N_919);
xor U3831 (N_3831,N_35,N_406);
nand U3832 (N_3832,N_727,N_1857);
and U3833 (N_3833,N_602,N_961);
or U3834 (N_3834,N_1214,N_1586);
nand U3835 (N_3835,N_982,N_283);
nand U3836 (N_3836,N_15,N_215);
nor U3837 (N_3837,N_487,N_342);
and U3838 (N_3838,N_176,N_268);
nor U3839 (N_3839,N_72,N_1269);
or U3840 (N_3840,N_30,N_43);
or U3841 (N_3841,N_172,N_821);
and U3842 (N_3842,N_884,N_831);
or U3843 (N_3843,N_1590,N_1053);
nor U3844 (N_3844,N_1324,N_1632);
nor U3845 (N_3845,N_1060,N_216);
nand U3846 (N_3846,N_732,N_1366);
and U3847 (N_3847,N_139,N_574);
nand U3848 (N_3848,N_1327,N_1019);
xnor U3849 (N_3849,N_1798,N_214);
xnor U3850 (N_3850,N_1186,N_1594);
nand U3851 (N_3851,N_1611,N_1178);
nand U3852 (N_3852,N_1021,N_464);
nor U3853 (N_3853,N_1110,N_631);
nor U3854 (N_3854,N_80,N_1460);
or U3855 (N_3855,N_1879,N_152);
xnor U3856 (N_3856,N_1512,N_189);
nor U3857 (N_3857,N_295,N_1259);
nor U3858 (N_3858,N_191,N_216);
nand U3859 (N_3859,N_776,N_297);
nand U3860 (N_3860,N_21,N_425);
nor U3861 (N_3861,N_578,N_1543);
nand U3862 (N_3862,N_449,N_161);
nor U3863 (N_3863,N_23,N_1500);
nand U3864 (N_3864,N_37,N_1989);
and U3865 (N_3865,N_442,N_84);
or U3866 (N_3866,N_1155,N_706);
nand U3867 (N_3867,N_1363,N_1751);
and U3868 (N_3868,N_1703,N_344);
and U3869 (N_3869,N_735,N_980);
nor U3870 (N_3870,N_1279,N_612);
nor U3871 (N_3871,N_845,N_758);
nor U3872 (N_3872,N_1254,N_1017);
nor U3873 (N_3873,N_742,N_1130);
nand U3874 (N_3874,N_1333,N_1321);
or U3875 (N_3875,N_1771,N_1472);
and U3876 (N_3876,N_1418,N_1415);
or U3877 (N_3877,N_726,N_1971);
and U3878 (N_3878,N_201,N_116);
and U3879 (N_3879,N_1340,N_864);
and U3880 (N_3880,N_861,N_28);
and U3881 (N_3881,N_1829,N_881);
nand U3882 (N_3882,N_489,N_946);
and U3883 (N_3883,N_962,N_441);
nor U3884 (N_3884,N_1542,N_1332);
xnor U3885 (N_3885,N_534,N_1898);
nor U3886 (N_3886,N_974,N_1050);
nand U3887 (N_3887,N_1562,N_1724);
or U3888 (N_3888,N_431,N_1205);
or U3889 (N_3889,N_266,N_570);
or U3890 (N_3890,N_645,N_1262);
and U3891 (N_3891,N_269,N_1124);
and U3892 (N_3892,N_857,N_914);
nand U3893 (N_3893,N_1853,N_1973);
or U3894 (N_3894,N_1512,N_1743);
or U3895 (N_3895,N_1583,N_791);
nor U3896 (N_3896,N_1055,N_501);
xnor U3897 (N_3897,N_1227,N_1282);
or U3898 (N_3898,N_1918,N_917);
xnor U3899 (N_3899,N_1301,N_333);
nor U3900 (N_3900,N_1701,N_1878);
or U3901 (N_3901,N_96,N_704);
nand U3902 (N_3902,N_386,N_1802);
nand U3903 (N_3903,N_454,N_1307);
nand U3904 (N_3904,N_1760,N_167);
and U3905 (N_3905,N_797,N_698);
nand U3906 (N_3906,N_467,N_742);
nand U3907 (N_3907,N_232,N_915);
and U3908 (N_3908,N_974,N_50);
nand U3909 (N_3909,N_313,N_1064);
nand U3910 (N_3910,N_295,N_959);
nand U3911 (N_3911,N_261,N_1270);
nor U3912 (N_3912,N_1427,N_1587);
xnor U3913 (N_3913,N_1119,N_517);
nor U3914 (N_3914,N_446,N_1416);
nand U3915 (N_3915,N_1110,N_1983);
xor U3916 (N_3916,N_1575,N_1377);
and U3917 (N_3917,N_1920,N_211);
or U3918 (N_3918,N_330,N_982);
and U3919 (N_3919,N_1072,N_1950);
or U3920 (N_3920,N_1315,N_968);
and U3921 (N_3921,N_279,N_499);
nor U3922 (N_3922,N_360,N_136);
nor U3923 (N_3923,N_1851,N_357);
xor U3924 (N_3924,N_1187,N_1734);
or U3925 (N_3925,N_1021,N_1133);
or U3926 (N_3926,N_849,N_80);
nand U3927 (N_3927,N_120,N_815);
or U3928 (N_3928,N_1279,N_1231);
or U3929 (N_3929,N_385,N_1503);
nand U3930 (N_3930,N_1587,N_1314);
xnor U3931 (N_3931,N_457,N_1589);
and U3932 (N_3932,N_1974,N_575);
nor U3933 (N_3933,N_334,N_1583);
or U3934 (N_3934,N_793,N_981);
or U3935 (N_3935,N_850,N_1927);
or U3936 (N_3936,N_84,N_268);
nor U3937 (N_3937,N_1100,N_376);
nand U3938 (N_3938,N_1887,N_353);
and U3939 (N_3939,N_67,N_673);
nand U3940 (N_3940,N_10,N_358);
nand U3941 (N_3941,N_116,N_1786);
nand U3942 (N_3942,N_1220,N_301);
and U3943 (N_3943,N_568,N_943);
nand U3944 (N_3944,N_1257,N_789);
or U3945 (N_3945,N_1299,N_1662);
nor U3946 (N_3946,N_107,N_202);
nor U3947 (N_3947,N_902,N_1757);
and U3948 (N_3948,N_968,N_639);
nor U3949 (N_3949,N_466,N_1146);
nand U3950 (N_3950,N_1836,N_1272);
or U3951 (N_3951,N_308,N_881);
and U3952 (N_3952,N_280,N_1714);
nor U3953 (N_3953,N_85,N_163);
nor U3954 (N_3954,N_288,N_1231);
nor U3955 (N_3955,N_138,N_1344);
nor U3956 (N_3956,N_1175,N_162);
and U3957 (N_3957,N_852,N_1477);
and U3958 (N_3958,N_1862,N_1001);
nand U3959 (N_3959,N_1403,N_1523);
nand U3960 (N_3960,N_1811,N_540);
nand U3961 (N_3961,N_907,N_653);
nand U3962 (N_3962,N_439,N_635);
nor U3963 (N_3963,N_1444,N_487);
nor U3964 (N_3964,N_673,N_737);
or U3965 (N_3965,N_1307,N_91);
and U3966 (N_3966,N_342,N_589);
or U3967 (N_3967,N_1781,N_1518);
nor U3968 (N_3968,N_32,N_201);
or U3969 (N_3969,N_1187,N_534);
or U3970 (N_3970,N_1345,N_709);
or U3971 (N_3971,N_635,N_627);
or U3972 (N_3972,N_1240,N_192);
and U3973 (N_3973,N_1992,N_1323);
nor U3974 (N_3974,N_1167,N_1175);
nor U3975 (N_3975,N_542,N_538);
nor U3976 (N_3976,N_1931,N_1698);
nor U3977 (N_3977,N_1971,N_1035);
nor U3978 (N_3978,N_1909,N_126);
or U3979 (N_3979,N_1219,N_982);
and U3980 (N_3980,N_1497,N_85);
and U3981 (N_3981,N_686,N_520);
nand U3982 (N_3982,N_1087,N_939);
xor U3983 (N_3983,N_1279,N_1919);
or U3984 (N_3984,N_1780,N_1562);
nand U3985 (N_3985,N_287,N_817);
nor U3986 (N_3986,N_403,N_1773);
nor U3987 (N_3987,N_780,N_1178);
nand U3988 (N_3988,N_326,N_906);
and U3989 (N_3989,N_164,N_1030);
nor U3990 (N_3990,N_1750,N_1460);
nand U3991 (N_3991,N_1150,N_1199);
and U3992 (N_3992,N_1358,N_78);
nand U3993 (N_3993,N_1713,N_455);
xnor U3994 (N_3994,N_1567,N_1526);
nand U3995 (N_3995,N_1232,N_1367);
nand U3996 (N_3996,N_346,N_896);
nor U3997 (N_3997,N_500,N_616);
nand U3998 (N_3998,N_373,N_947);
xor U3999 (N_3999,N_111,N_295);
nand U4000 (N_4000,N_3469,N_2848);
and U4001 (N_4001,N_2429,N_2136);
or U4002 (N_4002,N_2526,N_3333);
and U4003 (N_4003,N_2660,N_3755);
and U4004 (N_4004,N_3199,N_3956);
and U4005 (N_4005,N_2251,N_2466);
and U4006 (N_4006,N_2989,N_2804);
nor U4007 (N_4007,N_3726,N_2884);
xor U4008 (N_4008,N_2836,N_3890);
nor U4009 (N_4009,N_2758,N_2109);
and U4010 (N_4010,N_3182,N_3514);
nand U4011 (N_4011,N_3319,N_3688);
and U4012 (N_4012,N_2365,N_3098);
xnor U4013 (N_4013,N_2847,N_3952);
and U4014 (N_4014,N_2636,N_2972);
nand U4015 (N_4015,N_2936,N_2003);
or U4016 (N_4016,N_3522,N_2368);
nor U4017 (N_4017,N_2385,N_3998);
xnor U4018 (N_4018,N_2265,N_2846);
nand U4019 (N_4019,N_3864,N_3450);
nand U4020 (N_4020,N_3009,N_2226);
or U4021 (N_4021,N_3055,N_3154);
xor U4022 (N_4022,N_3627,N_3288);
and U4023 (N_4023,N_2014,N_3428);
nor U4024 (N_4024,N_3230,N_2092);
nand U4025 (N_4025,N_2702,N_2039);
nand U4026 (N_4026,N_3844,N_2337);
nand U4027 (N_4027,N_2865,N_3003);
xor U4028 (N_4028,N_3853,N_2218);
nor U4029 (N_4029,N_2731,N_3895);
or U4030 (N_4030,N_2872,N_2220);
nor U4031 (N_4031,N_3074,N_3015);
and U4032 (N_4032,N_3252,N_2939);
or U4033 (N_4033,N_2011,N_2481);
nor U4034 (N_4034,N_3723,N_3856);
or U4035 (N_4035,N_2344,N_2871);
nor U4036 (N_4036,N_3986,N_2719);
nand U4037 (N_4037,N_2963,N_2695);
xor U4038 (N_4038,N_2837,N_2934);
and U4039 (N_4039,N_3056,N_3134);
or U4040 (N_4040,N_3122,N_3232);
xnor U4041 (N_4041,N_3085,N_2807);
nor U4042 (N_4042,N_3259,N_3115);
nor U4043 (N_4043,N_3955,N_3209);
or U4044 (N_4044,N_3073,N_2384);
or U4045 (N_4045,N_3740,N_3017);
or U4046 (N_4046,N_3948,N_2511);
nor U4047 (N_4047,N_2703,N_2883);
and U4048 (N_4048,N_3316,N_2819);
and U4049 (N_4049,N_3198,N_3538);
nand U4050 (N_4050,N_3808,N_3769);
or U4051 (N_4051,N_3692,N_3082);
or U4052 (N_4052,N_2557,N_2652);
nor U4053 (N_4053,N_3240,N_2735);
and U4054 (N_4054,N_3599,N_3881);
or U4055 (N_4055,N_2315,N_2093);
nor U4056 (N_4056,N_2122,N_3594);
and U4057 (N_4057,N_2459,N_3529);
nand U4058 (N_4058,N_3180,N_3010);
nor U4059 (N_4059,N_2887,N_2005);
and U4060 (N_4060,N_3771,N_3159);
nor U4061 (N_4061,N_3058,N_2911);
and U4062 (N_4062,N_2516,N_2546);
and U4063 (N_4063,N_3924,N_2988);
or U4064 (N_4064,N_2886,N_2442);
and U4065 (N_4065,N_3087,N_3343);
nand U4066 (N_4066,N_2103,N_2177);
or U4067 (N_4067,N_2155,N_2034);
nor U4068 (N_4068,N_2256,N_2644);
and U4069 (N_4069,N_2188,N_3476);
nand U4070 (N_4070,N_2351,N_3752);
and U4071 (N_4071,N_2302,N_3565);
or U4072 (N_4072,N_2680,N_2739);
and U4073 (N_4073,N_3291,N_3426);
nor U4074 (N_4074,N_2941,N_3094);
or U4075 (N_4075,N_2568,N_2498);
xnor U4076 (N_4076,N_3527,N_3984);
or U4077 (N_4077,N_2669,N_2392);
and U4078 (N_4078,N_2990,N_3466);
or U4079 (N_4079,N_2182,N_2086);
or U4080 (N_4080,N_3361,N_2767);
nand U4081 (N_4081,N_3045,N_3649);
or U4082 (N_4082,N_2785,N_2019);
or U4083 (N_4083,N_3967,N_2041);
xor U4084 (N_4084,N_3489,N_3312);
and U4085 (N_4085,N_2390,N_3208);
nor U4086 (N_4086,N_2806,N_2107);
nand U4087 (N_4087,N_3616,N_3324);
and U4088 (N_4088,N_3852,N_3753);
nor U4089 (N_4089,N_3261,N_2559);
or U4090 (N_4090,N_2399,N_2065);
xor U4091 (N_4091,N_3893,N_3326);
and U4092 (N_4092,N_3443,N_3422);
nand U4093 (N_4093,N_3185,N_3170);
and U4094 (N_4094,N_2831,N_2185);
or U4095 (N_4095,N_2482,N_3663);
nand U4096 (N_4096,N_2986,N_2937);
and U4097 (N_4097,N_3862,N_2604);
nand U4098 (N_4098,N_2212,N_3169);
and U4099 (N_4099,N_3378,N_2576);
nand U4100 (N_4100,N_3979,N_2905);
nor U4101 (N_4101,N_2771,N_2876);
and U4102 (N_4102,N_2582,N_3581);
or U4103 (N_4103,N_3069,N_2920);
xor U4104 (N_4104,N_3144,N_3281);
or U4105 (N_4105,N_2575,N_2391);
nor U4106 (N_4106,N_2691,N_3381);
and U4107 (N_4107,N_2762,N_2594);
or U4108 (N_4108,N_3247,N_2353);
and U4109 (N_4109,N_3721,N_3517);
and U4110 (N_4110,N_2563,N_3146);
nor U4111 (N_4111,N_2634,N_3732);
or U4112 (N_4112,N_3496,N_3941);
nor U4113 (N_4113,N_2722,N_2628);
nand U4114 (N_4114,N_3137,N_2115);
nor U4115 (N_4115,N_3654,N_3111);
nand U4116 (N_4116,N_3099,N_3520);
or U4117 (N_4117,N_3646,N_3976);
and U4118 (N_4118,N_3917,N_3664);
or U4119 (N_4119,N_2009,N_2613);
nand U4120 (N_4120,N_2469,N_2446);
nand U4121 (N_4121,N_2348,N_2268);
and U4122 (N_4122,N_3491,N_2027);
or U4123 (N_4123,N_2418,N_3392);
and U4124 (N_4124,N_2354,N_3382);
and U4125 (N_4125,N_3127,N_3791);
xnor U4126 (N_4126,N_3101,N_3005);
nor U4127 (N_4127,N_2023,N_2487);
or U4128 (N_4128,N_3191,N_3996);
nand U4129 (N_4129,N_3898,N_2436);
nor U4130 (N_4130,N_3104,N_2232);
and U4131 (N_4131,N_3222,N_2873);
or U4132 (N_4132,N_3606,N_2471);
xnor U4133 (N_4133,N_2055,N_3540);
nor U4134 (N_4134,N_2321,N_3077);
or U4135 (N_4135,N_2761,N_2879);
and U4136 (N_4136,N_3710,N_3637);
and U4137 (N_4137,N_3783,N_3286);
nor U4138 (N_4138,N_2732,N_3341);
nor U4139 (N_4139,N_2640,N_2741);
nand U4140 (N_4140,N_2250,N_3197);
nand U4141 (N_4141,N_3810,N_3748);
and U4142 (N_4142,N_2227,N_2547);
or U4143 (N_4143,N_3901,N_2172);
and U4144 (N_4144,N_3190,N_3455);
nand U4145 (N_4145,N_3597,N_2889);
and U4146 (N_4146,N_2089,N_2455);
nand U4147 (N_4147,N_2169,N_3394);
or U4148 (N_4148,N_2603,N_3814);
or U4149 (N_4149,N_3595,N_2470);
nor U4150 (N_4150,N_2533,N_3705);
or U4151 (N_4151,N_2813,N_2726);
xor U4152 (N_4152,N_2914,N_3619);
xnor U4153 (N_4153,N_3966,N_2906);
nand U4154 (N_4154,N_3798,N_2863);
xnor U4155 (N_4155,N_3910,N_3231);
or U4156 (N_4156,N_3393,N_2283);
and U4157 (N_4157,N_3766,N_2991);
nand U4158 (N_4158,N_3415,N_3062);
nor U4159 (N_4159,N_2209,N_2102);
and U4160 (N_4160,N_3537,N_3915);
nand U4161 (N_4161,N_3989,N_3310);
and U4162 (N_4162,N_3084,N_2156);
and U4163 (N_4163,N_2295,N_2564);
or U4164 (N_4164,N_2791,N_3429);
nand U4165 (N_4165,N_2852,N_2608);
and U4166 (N_4166,N_2468,N_3579);
or U4167 (N_4167,N_3757,N_3696);
and U4168 (N_4168,N_2549,N_3117);
or U4169 (N_4169,N_2021,N_3916);
nand U4170 (N_4170,N_2062,N_2921);
and U4171 (N_4171,N_2671,N_2662);
nor U4172 (N_4172,N_3867,N_2870);
nand U4173 (N_4173,N_3060,N_2318);
nor U4174 (N_4174,N_2975,N_2207);
or U4175 (N_4175,N_3161,N_2326);
and U4176 (N_4176,N_3969,N_2168);
nand U4177 (N_4177,N_3059,N_2782);
and U4178 (N_4178,N_3874,N_2462);
nor U4179 (N_4179,N_3079,N_3824);
or U4180 (N_4180,N_2350,N_2580);
or U4181 (N_4181,N_3615,N_2061);
nor U4182 (N_4182,N_3631,N_3013);
nand U4183 (N_4183,N_2666,N_2796);
nor U4184 (N_4184,N_3703,N_3997);
and U4185 (N_4185,N_2451,N_2631);
nor U4186 (N_4186,N_2002,N_2298);
nand U4187 (N_4187,N_2304,N_3386);
or U4188 (N_4188,N_3092,N_3136);
and U4189 (N_4189,N_3020,N_3212);
nand U4190 (N_4190,N_3465,N_2605);
nand U4191 (N_4191,N_3822,N_3061);
or U4192 (N_4192,N_2668,N_2052);
nor U4193 (N_4193,N_3293,N_3733);
nand U4194 (N_4194,N_2131,N_2678);
or U4195 (N_4195,N_3065,N_3746);
or U4196 (N_4196,N_2581,N_2823);
xnor U4197 (N_4197,N_2210,N_3744);
nor U4198 (N_4198,N_2742,N_2656);
and U4199 (N_4199,N_2948,N_3528);
nor U4200 (N_4200,N_2561,N_3600);
nor U4201 (N_4201,N_3628,N_2534);
nor U4202 (N_4202,N_2503,N_3456);
or U4203 (N_4203,N_3156,N_2046);
or U4204 (N_4204,N_3891,N_3759);
nand U4205 (N_4205,N_2917,N_2331);
nand U4206 (N_4206,N_3018,N_2569);
or U4207 (N_4207,N_3926,N_2877);
or U4208 (N_4208,N_3183,N_2781);
or U4209 (N_4209,N_2790,N_2382);
xor U4210 (N_4210,N_2084,N_2913);
and U4211 (N_4211,N_2137,N_2943);
nand U4212 (N_4212,N_3970,N_3749);
nand U4213 (N_4213,N_3411,N_2515);
nor U4214 (N_4214,N_3963,N_2674);
xnor U4215 (N_4215,N_2060,N_2809);
or U4216 (N_4216,N_3719,N_3131);
nor U4217 (N_4217,N_2165,N_3019);
and U4218 (N_4218,N_3214,N_2282);
or U4219 (N_4219,N_3307,N_2982);
and U4220 (N_4220,N_2372,N_3427);
and U4221 (N_4221,N_2783,N_3314);
or U4222 (N_4222,N_3743,N_2708);
nand U4223 (N_4223,N_2454,N_2006);
nand U4224 (N_4224,N_3667,N_3632);
nor U4225 (N_4225,N_3380,N_3306);
and U4226 (N_4226,N_3225,N_2772);
nor U4227 (N_4227,N_3143,N_2415);
and U4228 (N_4228,N_2689,N_2746);
xor U4229 (N_4229,N_3118,N_2743);
nor U4230 (N_4230,N_3888,N_3196);
nand U4231 (N_4231,N_2157,N_3138);
nand U4232 (N_4232,N_3585,N_2439);
or U4233 (N_4233,N_3506,N_3035);
nor U4234 (N_4234,N_3267,N_3897);
and U4235 (N_4235,N_2775,N_3408);
or U4236 (N_4236,N_2773,N_2186);
or U4237 (N_4237,N_2252,N_2312);
and U4238 (N_4238,N_2658,N_3571);
nor U4239 (N_4239,N_3793,N_2694);
nor U4240 (N_4240,N_2303,N_3256);
nor U4241 (N_4241,N_2189,N_2076);
and U4242 (N_4242,N_3516,N_3462);
or U4243 (N_4243,N_2035,N_3959);
or U4244 (N_4244,N_2343,N_3772);
or U4245 (N_4245,N_3534,N_2119);
nand U4246 (N_4246,N_2619,N_3471);
nand U4247 (N_4247,N_2297,N_2273);
nor U4248 (N_4248,N_3570,N_2422);
or U4249 (N_4249,N_3054,N_2330);
nand U4250 (N_4250,N_3295,N_3368);
nor U4251 (N_4251,N_3367,N_2647);
nand U4252 (N_4252,N_2681,N_2589);
or U4253 (N_4253,N_3438,N_2334);
and U4254 (N_4254,N_2067,N_2940);
nand U4255 (N_4255,N_2254,N_2536);
xnor U4256 (N_4256,N_3044,N_2373);
or U4257 (N_4257,N_3270,N_2274);
and U4258 (N_4258,N_2340,N_2457);
nor U4259 (N_4259,N_2489,N_3109);
or U4260 (N_4260,N_3181,N_2463);
or U4261 (N_4261,N_3266,N_3350);
nor U4262 (N_4262,N_2585,N_2435);
xnor U4263 (N_4263,N_2241,N_3975);
or U4264 (N_4264,N_3102,N_2045);
or U4265 (N_4265,N_3021,N_3357);
nand U4266 (N_4266,N_3671,N_2788);
nand U4267 (N_4267,N_3362,N_2090);
or U4268 (N_4268,N_3276,N_3106);
nand U4269 (N_4269,N_3336,N_2787);
and U4270 (N_4270,N_2964,N_3882);
or U4271 (N_4271,N_2145,N_3611);
and U4272 (N_4272,N_3727,N_2474);
and U4273 (N_4273,N_3912,N_2031);
nand U4274 (N_4274,N_2335,N_3608);
nand U4275 (N_4275,N_2627,N_2506);
nor U4276 (N_4276,N_2441,N_2854);
or U4277 (N_4277,N_3364,N_3464);
and U4278 (N_4278,N_2857,N_2665);
or U4279 (N_4279,N_2057,N_3813);
and U4280 (N_4280,N_3334,N_3700);
xor U4281 (N_4281,N_2311,N_2687);
and U4282 (N_4282,N_2352,N_3435);
nor U4283 (N_4283,N_3470,N_3909);
nand U4284 (N_4284,N_2545,N_3690);
nand U4285 (N_4285,N_2322,N_3346);
nor U4286 (N_4286,N_2355,N_3968);
xor U4287 (N_4287,N_2024,N_3556);
nand U4288 (N_4288,N_3586,N_3848);
nor U4289 (N_4289,N_3189,N_3487);
nand U4290 (N_4290,N_2779,N_3301);
nor U4291 (N_4291,N_3397,N_3830);
or U4292 (N_4292,N_3873,N_3327);
nor U4293 (N_4293,N_3254,N_3174);
and U4294 (N_4294,N_2626,N_2793);
nand U4295 (N_4295,N_2153,N_3737);
and U4296 (N_4296,N_3679,N_3513);
and U4297 (N_4297,N_3175,N_3220);
or U4298 (N_4298,N_2510,N_3861);
and U4299 (N_4299,N_2505,N_3318);
nand U4300 (N_4300,N_2542,N_2231);
or U4301 (N_4301,N_2234,N_2987);
and U4302 (N_4302,N_3072,N_3578);
and U4303 (N_4303,N_2737,N_3081);
or U4304 (N_4304,N_2633,N_3883);
or U4305 (N_4305,N_3779,N_2161);
nor U4306 (N_4306,N_2705,N_2010);
or U4307 (N_4307,N_3770,N_3447);
nor U4308 (N_4308,N_3217,N_3503);
xor U4309 (N_4309,N_2638,N_3943);
or U4310 (N_4310,N_2308,N_2993);
nor U4311 (N_4311,N_2673,N_3905);
nor U4312 (N_4312,N_2257,N_2359);
or U4313 (N_4313,N_3778,N_2263);
or U4314 (N_4314,N_3030,N_2162);
nor U4315 (N_4315,N_3258,N_3289);
and U4316 (N_4316,N_3510,N_3954);
and U4317 (N_4317,N_2931,N_3931);
or U4318 (N_4318,N_3562,N_3285);
or U4319 (N_4319,N_2799,N_3929);
or U4320 (N_4320,N_3625,N_2339);
or U4321 (N_4321,N_3287,N_3133);
xor U4322 (N_4322,N_2117,N_2213);
or U4323 (N_4323,N_3933,N_2140);
nand U4324 (N_4324,N_3945,N_3173);
nor U4325 (N_4325,N_2692,N_3730);
or U4326 (N_4326,N_2197,N_2635);
nand U4327 (N_4327,N_2786,N_3339);
nand U4328 (N_4328,N_2728,N_2930);
nor U4329 (N_4329,N_3396,N_3234);
or U4330 (N_4330,N_3985,N_2704);
nand U4331 (N_4331,N_3053,N_2126);
and U4332 (N_4332,N_3728,N_3780);
nor U4333 (N_4333,N_3972,N_2393);
nand U4334 (N_4334,N_2805,N_3995);
xnor U4335 (N_4335,N_3602,N_2037);
or U4336 (N_4336,N_2507,N_2670);
nand U4337 (N_4337,N_3229,N_3794);
nor U4338 (N_4338,N_3100,N_2950);
or U4339 (N_4339,N_3572,N_2479);
nor U4340 (N_4340,N_2313,N_2574);
nor U4341 (N_4341,N_3454,N_2379);
nand U4342 (N_4342,N_2878,N_2424);
nor U4343 (N_4343,N_2944,N_3715);
nand U4344 (N_4344,N_2043,N_3063);
xnor U4345 (N_4345,N_3832,N_3661);
and U4346 (N_4346,N_2414,N_2166);
or U4347 (N_4347,N_2133,N_3297);
nor U4348 (N_4348,N_2198,N_2983);
nand U4349 (N_4349,N_3981,N_3802);
nor U4350 (N_4350,N_3908,N_2272);
or U4351 (N_4351,N_3541,N_2036);
or U4352 (N_4352,N_2998,N_2228);
nand U4353 (N_4353,N_3338,N_3919);
nor U4354 (N_4354,N_3598,N_3720);
nand U4355 (N_4355,N_3090,N_2148);
and U4356 (N_4356,N_2332,N_3763);
and U4357 (N_4357,N_3036,N_3803);
nand U4358 (N_4358,N_3472,N_3950);
and U4359 (N_4359,N_2492,N_3290);
or U4360 (N_4360,N_3839,N_2999);
and U4361 (N_4361,N_2306,N_3512);
xor U4362 (N_4362,N_2286,N_2551);
nor U4363 (N_4363,N_3634,N_3651);
or U4364 (N_4364,N_3702,N_2992);
nand U4365 (N_4365,N_3374,N_3605);
nor U4366 (N_4366,N_3292,N_3795);
nor U4367 (N_4367,N_3195,N_2817);
nor U4368 (N_4368,N_3303,N_3155);
or U4369 (N_4369,N_3041,N_2087);
or U4370 (N_4370,N_3383,N_2048);
nand U4371 (N_4371,N_3250,N_3255);
nand U4372 (N_4372,N_3167,N_3329);
nor U4373 (N_4373,N_2425,N_3675);
and U4374 (N_4374,N_2108,N_3211);
or U4375 (N_4375,N_3242,N_3006);
nor U4376 (N_4376,N_3947,N_3275);
or U4377 (N_4377,N_3958,N_2646);
xor U4378 (N_4378,N_3992,N_3886);
xnor U4379 (N_4379,N_3530,N_3937);
nand U4380 (N_4380,N_2612,N_2349);
or U4381 (N_4381,N_2152,N_3463);
nor U4382 (N_4382,N_2450,N_2610);
nor U4383 (N_4383,N_3701,N_2537);
or U4384 (N_4384,N_3603,N_2706);
and U4385 (N_4385,N_3023,N_3553);
and U4386 (N_4386,N_3828,N_3680);
or U4387 (N_4387,N_2181,N_2413);
and U4388 (N_4388,N_3268,N_3563);
xnor U4389 (N_4389,N_2955,N_3166);
and U4390 (N_4390,N_2432,N_2094);
nand U4391 (N_4391,N_2229,N_2573);
nand U4392 (N_4392,N_3097,N_2649);
nand U4393 (N_4393,N_2622,N_3235);
nand U4394 (N_4394,N_3369,N_3677);
nand U4395 (N_4395,N_2291,N_2849);
and U4396 (N_4396,N_2552,N_2756);
and U4397 (N_4397,N_3228,N_2467);
or U4398 (N_4398,N_3200,N_2683);
nor U4399 (N_4399,N_3308,N_3495);
xor U4400 (N_4400,N_3508,N_3940);
and U4401 (N_4401,N_2584,N_3441);
and U4402 (N_4402,N_3193,N_2721);
nor U4403 (N_4403,N_2480,N_2236);
nor U4404 (N_4404,N_3300,N_3402);
nand U4405 (N_4405,N_3849,N_2240);
or U4406 (N_4406,N_3206,N_2243);
and U4407 (N_4407,N_3332,N_2832);
and U4408 (N_4408,N_2058,N_3096);
and U4409 (N_4409,N_2738,N_3294);
or U4410 (N_4410,N_3405,N_2609);
nand U4411 (N_4411,N_3918,N_3284);
or U4412 (N_4412,N_3168,N_2176);
and U4413 (N_4413,N_3492,N_2184);
nor U4414 (N_4414,N_3150,N_2759);
and U4415 (N_4415,N_3384,N_3774);
or U4416 (N_4416,N_3792,N_2111);
xor U4417 (N_4417,N_2219,N_2460);
nor U4418 (N_4418,N_2066,N_2850);
nand U4419 (N_4419,N_3302,N_3375);
and U4420 (N_4420,N_2615,N_2278);
and U4421 (N_4421,N_3507,N_2158);
nor U4422 (N_4422,N_3145,N_2802);
nand U4423 (N_4423,N_2553,N_3140);
xor U4424 (N_4424,N_3549,N_2765);
nand U4425 (N_4425,N_2770,N_2833);
or U4426 (N_4426,N_2866,N_2639);
or U4427 (N_4427,N_3999,N_2118);
and U4428 (N_4428,N_3542,N_2645);
nor U4429 (N_4429,N_2897,N_3736);
nand U4430 (N_4430,N_3414,N_2134);
nand U4431 (N_4431,N_3827,N_3580);
nand U4432 (N_4432,N_2709,N_2453);
or U4433 (N_4433,N_3171,N_3245);
nand U4434 (N_4434,N_2433,N_3983);
nand U4435 (N_4435,N_3444,N_3739);
nor U4436 (N_4436,N_3934,N_3475);
nand U4437 (N_4437,N_2927,N_2591);
and U4438 (N_4438,N_2287,N_2376);
nand U4439 (N_4439,N_3551,N_3391);
and U4440 (N_4440,N_3582,N_2881);
or U4441 (N_4441,N_2042,N_2016);
nor U4442 (N_4442,N_3876,N_2859);
nand U4443 (N_4443,N_3365,N_2517);
and U4444 (N_4444,N_2053,N_2113);
and U4445 (N_4445,N_2485,N_2280);
nor U4446 (N_4446,N_3067,N_3555);
xnor U4447 (N_4447,N_2715,N_3113);
nand U4448 (N_4448,N_3760,N_2730);
and U4449 (N_4449,N_3676,N_3296);
nand U4450 (N_4450,N_3371,N_2030);
nor U4451 (N_4451,N_3773,N_3921);
xnor U4452 (N_4452,N_2797,N_3674);
nor U4453 (N_4453,N_2123,N_2578);
and U4454 (N_4454,N_2821,N_3358);
nand U4455 (N_4455,N_3105,N_3359);
nand U4456 (N_4456,N_3709,N_2292);
nand U4457 (N_4457,N_3788,N_2980);
or U4458 (N_4458,N_3811,N_2729);
nand U4459 (N_4459,N_2438,N_3153);
and U4460 (N_4460,N_3467,N_2171);
or U4461 (N_4461,N_2079,N_3348);
and U4462 (N_4462,N_2932,N_2617);
or U4463 (N_4463,N_3707,N_2394);
nand U4464 (N_4464,N_2532,N_3939);
nand U4465 (N_4465,N_2899,N_2789);
or U4466 (N_4466,N_2653,N_2997);
nand U4467 (N_4467,N_3001,N_3165);
nand U4468 (N_4468,N_2333,N_2745);
xnor U4469 (N_4469,N_3532,N_3000);
nand U4470 (N_4470,N_3207,N_3500);
xnor U4471 (N_4471,N_3659,N_3340);
nand U4472 (N_4472,N_2149,N_2183);
nand U4473 (N_4473,N_3626,N_3622);
nand U4474 (N_4474,N_3088,N_2882);
or U4475 (N_4475,N_2869,N_2180);
xnor U4476 (N_4476,N_3223,N_2701);
nand U4477 (N_4477,N_2146,N_3139);
or U4478 (N_4478,N_2903,N_2497);
and U4479 (N_4479,N_2902,N_2203);
or U4480 (N_4480,N_2143,N_3640);
nand U4481 (N_4481,N_3103,N_2004);
nor U4482 (N_4482,N_2923,N_3277);
nor U4483 (N_4483,N_3961,N_3902);
or U4484 (N_4484,N_3716,N_2417);
nor U4485 (N_4485,N_2714,N_2405);
or U4486 (N_4486,N_2179,N_3596);
or U4487 (N_4487,N_2924,N_2363);
or U4488 (N_4488,N_3840,N_3545);
xnor U4489 (N_4489,N_3880,N_2527);
and U4490 (N_4490,N_2411,N_2851);
xnor U4491 (N_4491,N_3025,N_3401);
nand U4492 (N_4492,N_3558,N_3552);
or U4493 (N_4493,N_3835,N_2301);
and U4494 (N_4494,N_2248,N_3875);
and U4495 (N_4495,N_3870,N_2211);
nand U4496 (N_4496,N_2679,N_3907);
or U4497 (N_4497,N_2395,N_2476);
or U4498 (N_4498,N_3434,N_2688);
nand U4499 (N_4499,N_2216,N_2530);
nor U4500 (N_4500,N_3666,N_2400);
or U4501 (N_4501,N_2676,N_2598);
nor U4502 (N_4502,N_3914,N_2947);
nor U4503 (N_4503,N_3768,N_2565);
and U4504 (N_4504,N_3896,N_3978);
and U4505 (N_4505,N_3468,N_2524);
nand U4506 (N_4506,N_3638,N_2106);
nand U4507 (N_4507,N_3913,N_2520);
nor U4508 (N_4508,N_3283,N_2538);
or U4509 (N_4509,N_3282,N_3847);
nor U4510 (N_4510,N_2440,N_2096);
nor U4511 (N_4511,N_3860,N_2402);
nand U4512 (N_4512,N_3618,N_2570);
nor U4513 (N_4513,N_2979,N_2925);
or U4514 (N_4514,N_3697,N_3711);
and U4515 (N_4515,N_2910,N_3630);
nor U4516 (N_4516,N_3356,N_3859);
and U4517 (N_4517,N_2431,N_2810);
and U4518 (N_4518,N_2040,N_2675);
nand U4519 (N_4519,N_2543,N_3724);
nand U4520 (N_4520,N_3704,N_3162);
nand U4521 (N_4521,N_2267,N_2361);
nand U4522 (N_4522,N_3057,N_3900);
nor U4523 (N_4523,N_3879,N_3204);
nand U4524 (N_4524,N_3821,N_3936);
nand U4525 (N_4525,N_3385,N_3461);
or U4526 (N_4526,N_2364,N_3107);
nor U4527 (N_4527,N_3331,N_3523);
nand U4528 (N_4528,N_2430,N_3610);
or U4529 (N_4529,N_2560,N_2523);
and U4530 (N_4530,N_2864,N_2822);
xnor U4531 (N_4531,N_2513,N_2867);
and U4532 (N_4532,N_2744,N_2217);
and U4533 (N_4533,N_2461,N_2378);
nor U4534 (N_4534,N_2495,N_3248);
nor U4535 (N_4535,N_2159,N_3123);
and U4536 (N_4536,N_2614,N_2445);
xnor U4537 (N_4537,N_3448,N_2142);
or U4538 (N_4538,N_2261,N_2978);
xor U4539 (N_4539,N_2753,N_3095);
xnor U4540 (N_4540,N_2514,N_2755);
or U4541 (N_4541,N_3387,N_3452);
and U4542 (N_4542,N_2050,N_3273);
nand U4543 (N_4543,N_3642,N_3244);
or U4544 (N_4544,N_2898,N_2063);
nor U4545 (N_4545,N_3758,N_3501);
or U4546 (N_4546,N_3911,N_3635);
or U4547 (N_4547,N_2369,N_2190);
and U4548 (N_4548,N_2178,N_2977);
and U4549 (N_4549,N_2713,N_3388);
nand U4550 (N_4550,N_3866,N_2223);
and U4551 (N_4551,N_2175,N_3928);
nand U4552 (N_4552,N_2724,N_3186);
nor U4553 (N_4553,N_2001,N_2033);
nand U4554 (N_4554,N_2407,N_2077);
xnor U4555 (N_4555,N_3591,N_3560);
nor U4556 (N_4556,N_3718,N_2244);
nor U4557 (N_4557,N_2047,N_3446);
xor U4558 (N_4558,N_2970,N_2531);
and U4559 (N_4559,N_3842,N_3641);
nand U4560 (N_4560,N_2193,N_2483);
nand U4561 (N_4561,N_2071,N_2116);
xor U4562 (N_4562,N_2026,N_3187);
nand U4563 (N_4563,N_2825,N_3342);
or U4564 (N_4564,N_2725,N_2012);
xnor U4565 (N_4565,N_3815,N_2270);
or U4566 (N_4566,N_2808,N_2398);
nand U4567 (N_4567,N_2812,N_3395);
nor U4568 (N_4568,N_2984,N_2623);
or U4569 (N_4569,N_3946,N_3543);
and U4570 (N_4570,N_2025,N_3672);
xnor U4571 (N_4571,N_3052,N_3012);
nor U4572 (N_4572,N_3315,N_3483);
and U4573 (N_4573,N_2056,N_3568);
nand U4574 (N_4574,N_3604,N_3617);
and U4575 (N_4575,N_3845,N_2693);
nor U4576 (N_4576,N_3505,N_2082);
or U4577 (N_4577,N_2685,N_2512);
and U4578 (N_4578,N_2661,N_3877);
and U4579 (N_4579,N_3431,N_3526);
and U4580 (N_4580,N_3389,N_2484);
nand U4581 (N_4581,N_2592,N_3202);
nand U4582 (N_4582,N_2752,N_3257);
xor U4583 (N_4583,N_3042,N_3777);
and U4584 (N_4584,N_2170,N_2754);
nand U4585 (N_4585,N_2651,N_2929);
xnor U4586 (N_4586,N_3784,N_2500);
nand U4587 (N_4587,N_2196,N_3458);
and U4588 (N_4588,N_3493,N_2994);
or U4589 (N_4589,N_3249,N_2766);
or U4590 (N_4590,N_2586,N_3789);
or U4591 (N_4591,N_2206,N_3238);
nor U4592 (N_4592,N_3533,N_2127);
or U4593 (N_4593,N_2579,N_2655);
and U4594 (N_4594,N_2070,N_3993);
nand U4595 (N_4595,N_3762,N_2928);
nor U4596 (N_4596,N_2345,N_3991);
nand U4597 (N_4597,N_2973,N_2624);
nor U4598 (N_4598,N_3872,N_2032);
and U4599 (N_4599,N_3765,N_2734);
nand U4600 (N_4600,N_3083,N_3712);
nand U4601 (N_4601,N_2829,N_3751);
or U4602 (N_4602,N_3673,N_3110);
and U4603 (N_4603,N_2114,N_2587);
nor U4604 (N_4604,N_2967,N_3725);
nand U4605 (N_4605,N_2294,N_2915);
and U4606 (N_4606,N_3002,N_3353);
nor U4607 (N_4607,N_2926,N_3372);
or U4608 (N_4608,N_3750,N_3790);
nor U4609 (N_4609,N_3141,N_2478);
nand U4610 (N_4610,N_2472,N_2894);
nand U4611 (N_4611,N_3227,N_2659);
nand U4612 (N_4612,N_3511,N_3264);
nor U4613 (N_4613,N_3224,N_3246);
xor U4614 (N_4614,N_2933,N_2890);
nor U4615 (N_4615,N_3149,N_3192);
or U4616 (N_4616,N_2375,N_3108);
or U4617 (N_4617,N_3218,N_3412);
nor U4618 (N_4618,N_3609,N_3885);
or U4619 (N_4619,N_3804,N_3004);
nor U4620 (N_4620,N_3480,N_2632);
or U4621 (N_4621,N_3089,N_3574);
and U4622 (N_4622,N_2757,N_3775);
and U4623 (N_4623,N_3116,N_3203);
nand U4624 (N_4624,N_2128,N_2488);
nand U4625 (N_4625,N_3620,N_3960);
nand U4626 (N_4626,N_2784,N_3280);
and U4627 (N_4627,N_3028,N_2360);
nand U4628 (N_4628,N_2015,N_3241);
nand U4629 (N_4629,N_3691,N_2412);
nor U4630 (N_4630,N_3957,N_3655);
nand U4631 (N_4631,N_3320,N_2262);
or U4632 (N_4632,N_3575,N_2828);
or U4633 (N_4633,N_3576,N_3430);
nor U4634 (N_4634,N_3129,N_3416);
nor U4635 (N_4635,N_3829,N_2141);
nor U4636 (N_4636,N_2951,N_3624);
nor U4637 (N_4637,N_3884,N_2602);
nor U4638 (N_4638,N_3253,N_3419);
nand U4639 (N_4639,N_3317,N_3951);
nand U4640 (N_4640,N_2643,N_2528);
nand U4641 (N_4641,N_2763,N_2795);
or U4642 (N_4642,N_2945,N_3722);
or U4643 (N_4643,N_2452,N_2101);
and U4644 (N_4644,N_2853,N_2965);
nand U4645 (N_4645,N_2276,N_3262);
nor U4646 (N_4646,N_2904,N_2173);
nand U4647 (N_4647,N_3120,N_3660);
nand U4648 (N_4648,N_3561,N_2299);
nor U4649 (N_4649,N_2341,N_2868);
and U4650 (N_4650,N_3379,N_2167);
nand U4651 (N_4651,N_3502,N_2253);
or U4652 (N_4652,N_3987,N_3330);
nand U4653 (N_4653,N_3432,N_2447);
nand U4654 (N_4654,N_3298,N_2764);
and U4655 (N_4655,N_3305,N_3816);
and U4656 (N_4656,N_3988,N_2205);
or U4657 (N_4657,N_2293,N_3299);
nor U4658 (N_4658,N_3647,N_3459);
or U4659 (N_4659,N_2464,N_3274);
nand U4660 (N_4660,N_3662,N_2616);
xor U4661 (N_4661,N_2269,N_2522);
nor U4662 (N_4662,N_2242,N_2588);
and U4663 (N_4663,N_2075,N_3440);
nor U4664 (N_4664,N_2717,N_3683);
nor U4665 (N_4665,N_2249,N_2953);
or U4666 (N_4666,N_3188,N_3008);
nand U4667 (N_4667,N_3964,N_3124);
or U4668 (N_4668,N_3990,N_2509);
or U4669 (N_4669,N_2289,N_3007);
or U4670 (N_4670,N_2187,N_2401);
or U4671 (N_4671,N_3226,N_2596);
or U4672 (N_4672,N_2607,N_3243);
and U4673 (N_4673,N_2502,N_3417);
nand U4674 (N_4674,N_2969,N_3474);
or U4675 (N_4675,N_3504,N_3977);
or U4676 (N_4676,N_3418,N_2121);
nor U4677 (N_4677,N_2064,N_3152);
and U4678 (N_4678,N_2072,N_3142);
or U4679 (N_4679,N_2195,N_3557);
nand U4680 (N_4680,N_2907,N_3524);
nand U4681 (N_4681,N_3278,N_3064);
or U4682 (N_4682,N_3490,N_3029);
nand U4683 (N_4683,N_3834,N_2727);
or U4684 (N_4684,N_2410,N_3742);
and U4685 (N_4685,N_2408,N_2700);
and U4686 (N_4686,N_2690,N_2996);
nor U4687 (N_4687,N_3125,N_2132);
or U4688 (N_4688,N_2577,N_2960);
xor U4689 (N_4689,N_3026,N_2535);
nand U4690 (N_4690,N_3652,N_2597);
or U4691 (N_4691,N_2583,N_2160);
nor U4692 (N_4692,N_2409,N_3436);
nor U4693 (N_4693,N_2191,N_2264);
and U4694 (N_4694,N_3695,N_2396);
and U4695 (N_4695,N_2309,N_3347);
and U4696 (N_4696,N_2129,N_2000);
nor U4697 (N_4697,N_2091,N_3785);
or U4698 (N_4698,N_3451,N_2529);
nor U4699 (N_4699,N_3614,N_2374);
or U4700 (N_4700,N_3445,N_2493);
or U4701 (N_4701,N_3130,N_3352);
and U4702 (N_4702,N_3163,N_2305);
nand U4703 (N_4703,N_2861,N_3982);
or U4704 (N_4704,N_2225,N_3799);
or U4705 (N_4705,N_2317,N_3566);
or U4706 (N_4706,N_3215,N_3554);
nor U4707 (N_4707,N_3738,N_2699);
xor U4708 (N_4708,N_3022,N_2711);
or U4709 (N_4709,N_3400,N_2112);
nand U4710 (N_4710,N_2599,N_2957);
nand U4711 (N_4711,N_2120,N_2519);
or U4712 (N_4712,N_2909,N_2540);
nor U4713 (N_4713,N_3922,N_3498);
nor U4714 (N_4714,N_3657,N_3569);
or U4715 (N_4715,N_3114,N_2918);
and U4716 (N_4716,N_3335,N_3974);
and U4717 (N_4717,N_3892,N_3157);
nand U4718 (N_4718,N_2088,N_2377);
or U4719 (N_4719,N_2801,N_2138);
nand U4720 (N_4720,N_2222,N_2814);
and U4721 (N_4721,N_2811,N_2028);
nor U4722 (N_4722,N_2059,N_2642);
nor U4723 (N_4723,N_2388,N_2239);
and U4724 (N_4724,N_2855,N_2329);
and U4725 (N_4725,N_2750,N_2327);
nand U4726 (N_4726,N_2860,N_2038);
or U4727 (N_4727,N_3850,N_2663);
or U4728 (N_4728,N_3826,N_2397);
or U4729 (N_4729,N_2245,N_2406);
nand U4730 (N_4730,N_3764,N_3589);
and U4731 (N_4731,N_3925,N_2266);
or U4732 (N_4732,N_3851,N_3216);
and U4733 (N_4733,N_3040,N_3370);
nor U4734 (N_4734,N_3323,N_3831);
and U4735 (N_4735,N_3584,N_3399);
nand U4736 (N_4736,N_3376,N_3836);
or U4737 (N_4737,N_2749,N_3398);
and U4738 (N_4738,N_2820,N_2566);
and U4739 (N_4739,N_3587,N_2518);
nand U4740 (N_4740,N_2499,N_3349);
and U4741 (N_4741,N_2099,N_2625);
xor U4742 (N_4742,N_3269,N_3546);
and U4743 (N_4743,N_3938,N_3682);
xor U4744 (N_4744,N_2271,N_2935);
nor U4745 (N_4745,N_3547,N_2097);
or U4746 (N_4746,N_3184,N_3894);
and U4747 (N_4747,N_3363,N_2080);
or U4748 (N_4748,N_2641,N_2421);
nor U4749 (N_4749,N_3525,N_2630);
nor U4750 (N_4750,N_3818,N_2818);
nand U4751 (N_4751,N_2800,N_2420);
xnor U4752 (N_4752,N_3694,N_3251);
nand U4753 (N_4753,N_2202,N_2277);
and U4754 (N_4754,N_2285,N_2448);
xnor U4755 (N_4755,N_3237,N_3070);
nor U4756 (N_4756,N_2491,N_3899);
nand U4757 (N_4757,N_2154,N_2104);
nand U4758 (N_4758,N_2716,N_3066);
or U4759 (N_4759,N_2712,N_2667);
nor U4760 (N_4760,N_2650,N_3457);
nand U4761 (N_4761,N_3179,N_3477);
or U4762 (N_4762,N_3033,N_3449);
nand U4763 (N_4763,N_2275,N_2672);
or U4764 (N_4764,N_3590,N_3796);
or U4765 (N_4765,N_3686,N_3735);
xor U4766 (N_4766,N_3903,N_2201);
or U4767 (N_4767,N_2556,N_2985);
nor U4768 (N_4768,N_2826,N_3973);
or U4769 (N_4769,N_3812,N_2139);
and U4770 (N_4770,N_2371,N_2769);
and U4771 (N_4771,N_2606,N_3887);
nand U4772 (N_4772,N_3039,N_3645);
nand U4773 (N_4773,N_2380,N_3573);
nor U4774 (N_4774,N_3309,N_2358);
nor U4775 (N_4775,N_3403,N_3653);
or U4776 (N_4776,N_2387,N_2020);
nor U4777 (N_4777,N_2260,N_3263);
nor U4778 (N_4778,N_3354,N_3693);
or U4779 (N_4779,N_2098,N_3920);
or U4780 (N_4780,N_2281,N_3178);
nor U4781 (N_4781,N_2900,N_2130);
nor U4782 (N_4782,N_2555,N_2314);
or U4783 (N_4783,N_2428,N_2834);
nor U4784 (N_4784,N_3550,N_2475);
nand U4785 (N_4785,N_2238,N_3636);
nor U4786 (N_4786,N_2600,N_3433);
and U4787 (N_4787,N_2383,N_2949);
or U4788 (N_4788,N_2558,N_2443);
or U4789 (N_4789,N_2437,N_2328);
xor U4790 (N_4790,N_2875,N_2959);
nand U4791 (N_4791,N_2427,N_2733);
or U4792 (N_4792,N_2357,N_3858);
nand U4793 (N_4793,N_3854,N_2300);
nor U4794 (N_4794,N_3043,N_2224);
and U4795 (N_4795,N_2230,N_3745);
nor U4796 (N_4796,N_2508,N_3767);
nor U4797 (N_4797,N_2362,N_2288);
nand U4798 (N_4798,N_3478,N_3863);
and U4799 (N_4799,N_2049,N_3668);
nor U4800 (N_4800,N_3485,N_3479);
nand U4801 (N_4801,N_2444,N_3272);
and U4802 (N_4802,N_3051,N_2029);
nand U4803 (N_4803,N_2473,N_2893);
xnor U4804 (N_4804,N_3404,N_3855);
and U4805 (N_4805,N_3151,N_3437);
xor U4806 (N_4806,N_3819,N_2827);
and U4807 (N_4807,N_3927,N_3031);
nor U4808 (N_4808,N_2842,N_2290);
or U4809 (N_4809,N_3685,N_2324);
xnor U4810 (N_4810,N_3825,N_2664);
nor U4811 (N_4811,N_2803,N_2525);
nor U4812 (N_4812,N_2367,N_3037);
xor U4813 (N_4813,N_3971,N_2389);
nor U4814 (N_4814,N_3425,N_2776);
nor U4815 (N_4815,N_3126,N_3078);
and U4816 (N_4816,N_2496,N_2338);
nand U4817 (N_4817,N_2748,N_2740);
nor U4818 (N_4818,N_2885,N_2539);
or U4819 (N_4819,N_3038,N_2710);
nor U4820 (N_4820,N_2880,N_3588);
xor U4821 (N_4821,N_3698,N_2611);
nor U4822 (N_4822,N_2974,N_3509);
xor U4823 (N_4823,N_2572,N_2976);
or U4824 (N_4824,N_3442,N_3176);
xor U4825 (N_4825,N_2595,N_3583);
and U4826 (N_4826,N_2707,N_2590);
or U4827 (N_4827,N_3016,N_2521);
nor U4828 (N_4828,N_3648,N_3699);
nand U4829 (N_4829,N_2541,N_2208);
nand U4830 (N_4830,N_3714,N_3843);
nand U4831 (N_4831,N_3518,N_3439);
nand U4832 (N_4832,N_3410,N_2233);
xnor U4833 (N_4833,N_2874,N_2637);
or U4834 (N_4834,N_3729,N_3213);
or U4835 (N_4835,N_2916,N_2751);
nor U4836 (N_4836,N_3210,N_3741);
or U4837 (N_4837,N_2490,N_3484);
and U4838 (N_4838,N_2798,N_2550);
and U4839 (N_4839,N_3592,N_3544);
and U4840 (N_4840,N_3076,N_2073);
or U4841 (N_4841,N_3613,N_3539);
or U4842 (N_4842,N_3011,N_2494);
nand U4843 (N_4843,N_2629,N_2621);
nor U4844 (N_4844,N_2593,N_2843);
and U4845 (N_4845,N_2919,N_3423);
nand U4846 (N_4846,N_2456,N_2215);
or U4847 (N_4847,N_2054,N_3279);
or U4848 (N_4848,N_2844,N_3049);
or U4849 (N_4849,N_2501,N_2654);
or U4850 (N_4850,N_2247,N_3684);
nor U4851 (N_4851,N_3121,N_2938);
or U4852 (N_4852,N_3413,N_2954);
xor U4853 (N_4853,N_3047,N_2961);
or U4854 (N_4854,N_3820,N_3219);
nand U4855 (N_4855,N_2151,N_3935);
nor U4856 (N_4856,N_3325,N_3754);
or U4857 (N_4857,N_2841,N_3871);
nand U4858 (N_4858,N_3128,N_3311);
nand U4859 (N_4859,N_2320,N_2204);
or U4860 (N_4860,N_3164,N_3665);
or U4861 (N_4861,N_3112,N_3841);
nor U4862 (N_4862,N_3805,N_3787);
nand U4863 (N_4863,N_2682,N_2296);
nor U4864 (N_4864,N_2135,N_2554);
nor U4865 (N_4865,N_2386,N_3846);
xor U4866 (N_4866,N_3421,N_2069);
nor U4867 (N_4867,N_3669,N_2017);
nand U4868 (N_4868,N_2235,N_2200);
or U4869 (N_4869,N_3239,N_3656);
nand U4870 (N_4870,N_2194,N_3782);
and U4871 (N_4871,N_3906,N_3132);
and U4872 (N_4872,N_2458,N_2995);
nand U4873 (N_4873,N_2971,N_3328);
and U4874 (N_4874,N_3865,N_3482);
nand U4875 (N_4875,N_2620,N_2571);
or U4876 (N_4876,N_3048,N_3962);
and U4877 (N_4877,N_3014,N_3409);
nor U4878 (N_4878,N_2423,N_2105);
and U4879 (N_4879,N_2370,N_3024);
or U4880 (N_4880,N_3797,N_3420);
nor U4881 (N_4881,N_3119,N_3878);
or U4882 (N_4882,N_2601,N_3265);
and U4883 (N_4883,N_3406,N_2840);
nor U4884 (N_4884,N_3838,N_3373);
and U4885 (N_4885,N_2403,N_2258);
xor U4886 (N_4886,N_2962,N_2416);
or U4887 (N_4887,N_3027,N_3857);
nor U4888 (N_4888,N_3080,N_3708);
xor U4889 (N_4889,N_3519,N_2150);
or U4890 (N_4890,N_2342,N_3776);
xnor U4891 (N_4891,N_3869,N_3071);
nor U4892 (N_4892,N_2815,N_2085);
nor U4893 (N_4893,N_3086,N_3868);
nor U4894 (N_4894,N_3355,N_3515);
nand U4895 (N_4895,N_2794,N_3786);
or U4896 (N_4896,N_2013,N_2908);
nor U4897 (N_4897,N_2174,N_3271);
nor U4898 (N_4898,N_2648,N_2747);
nor U4899 (N_4899,N_2319,N_3075);
nand U4900 (N_4900,N_2696,N_2237);
or U4901 (N_4901,N_3221,N_2718);
nor U4902 (N_4902,N_3965,N_2465);
nand U4903 (N_4903,N_3678,N_2255);
or U4904 (N_4904,N_2284,N_3473);
and U4905 (N_4905,N_2760,N_3670);
and U4906 (N_4906,N_2768,N_2723);
or U4907 (N_4907,N_2774,N_2862);
and U4908 (N_4908,N_3322,N_2858);
nand U4909 (N_4909,N_3800,N_3407);
xnor U4910 (N_4910,N_3923,N_2845);
or U4911 (N_4911,N_3535,N_2981);
and U4912 (N_4912,N_3260,N_3536);
nor U4913 (N_4913,N_2548,N_2366);
or U4914 (N_4914,N_2824,N_3321);
or U4915 (N_4915,N_2657,N_3930);
nand U4916 (N_4916,N_2922,N_2068);
nor U4917 (N_4917,N_3046,N_3639);
or U4918 (N_4918,N_3658,N_3093);
nor U4919 (N_4919,N_2686,N_2095);
nor U4920 (N_4920,N_2956,N_3481);
or U4921 (N_4921,N_2214,N_3781);
nand U4922 (N_4922,N_2125,N_3453);
and U4923 (N_4923,N_3994,N_2958);
and U4924 (N_4924,N_3531,N_2892);
or U4925 (N_4925,N_2968,N_3904);
or U4926 (N_4926,N_2083,N_2891);
or U4927 (N_4927,N_3837,N_3629);
and U4928 (N_4928,N_2778,N_3366);
nor U4929 (N_4929,N_3345,N_3521);
or U4930 (N_4930,N_3486,N_2147);
and U4931 (N_4931,N_3390,N_2449);
and U4932 (N_4932,N_3621,N_2259);
nand U4933 (N_4933,N_3817,N_2081);
or U4934 (N_4934,N_3889,N_2246);
or U4935 (N_4935,N_2325,N_2356);
or U4936 (N_4936,N_2816,N_2896);
and U4937 (N_4937,N_2434,N_3607);
or U4938 (N_4938,N_2777,N_2544);
nand U4939 (N_4939,N_2839,N_3494);
nor U4940 (N_4940,N_3233,N_2736);
and U4941 (N_4941,N_2684,N_3731);
nor U4942 (N_4942,N_2830,N_3953);
xor U4943 (N_4943,N_3135,N_2618);
nor U4944 (N_4944,N_3980,N_3032);
nand U4945 (N_4945,N_3304,N_2677);
and U4946 (N_4946,N_2912,N_3942);
or U4947 (N_4947,N_3497,N_3689);
and U4948 (N_4948,N_3633,N_2486);
nor U4949 (N_4949,N_3148,N_2562);
or U4950 (N_4950,N_2952,N_3344);
xnor U4951 (N_4951,N_3177,N_2110);
nand U4952 (N_4952,N_3687,N_2780);
nor U4953 (N_4953,N_3499,N_3601);
and U4954 (N_4954,N_2346,N_3949);
and U4955 (N_4955,N_3091,N_2698);
nor U4956 (N_4956,N_2942,N_2966);
nand U4957 (N_4957,N_2279,N_3612);
nand U4958 (N_4958,N_3756,N_3577);
nand U4959 (N_4959,N_2720,N_3337);
or U4960 (N_4960,N_3567,N_3806);
nor U4961 (N_4961,N_3932,N_3801);
xnor U4962 (N_4962,N_2504,N_3623);
and U4963 (N_4963,N_2835,N_2792);
xor U4964 (N_4964,N_3068,N_2946);
xnor U4965 (N_4965,N_3377,N_3747);
nor U4966 (N_4966,N_3194,N_3201);
and U4967 (N_4967,N_2477,N_2100);
and U4968 (N_4968,N_3944,N_3313);
xor U4969 (N_4969,N_2199,N_2078);
nor U4970 (N_4970,N_2163,N_3424);
and U4971 (N_4971,N_2051,N_2007);
or U4972 (N_4972,N_3706,N_3564);
nand U4973 (N_4973,N_2697,N_2124);
nor U4974 (N_4974,N_2426,N_2901);
nor U4975 (N_4975,N_3360,N_2336);
nor U4976 (N_4976,N_3236,N_2381);
xor U4977 (N_4977,N_3548,N_3650);
nor U4978 (N_4978,N_3158,N_2419);
or U4979 (N_4979,N_2144,N_2347);
nor U4980 (N_4980,N_3761,N_3717);
or U4981 (N_4981,N_3050,N_2221);
nand U4982 (N_4982,N_2895,N_2022);
or U4983 (N_4983,N_3833,N_2164);
nor U4984 (N_4984,N_2323,N_3713);
and U4985 (N_4985,N_2856,N_2310);
xor U4986 (N_4986,N_3593,N_3809);
xnor U4987 (N_4987,N_3160,N_2316);
nor U4988 (N_4988,N_2404,N_3644);
nand U4989 (N_4989,N_2044,N_3681);
and U4990 (N_4990,N_2074,N_2888);
or U4991 (N_4991,N_3205,N_2018);
nand U4992 (N_4992,N_3488,N_3351);
or U4993 (N_4993,N_3460,N_3734);
nand U4994 (N_4994,N_3807,N_2567);
and U4995 (N_4995,N_3034,N_3147);
or U4996 (N_4996,N_3559,N_3172);
xnor U4997 (N_4997,N_2192,N_3643);
and U4998 (N_4998,N_2008,N_3823);
or U4999 (N_4999,N_2838,N_2307);
xnor U5000 (N_5000,N_2549,N_3554);
and U5001 (N_5001,N_3389,N_3709);
or U5002 (N_5002,N_3436,N_2114);
nand U5003 (N_5003,N_2637,N_3145);
and U5004 (N_5004,N_2922,N_3246);
xor U5005 (N_5005,N_3830,N_3817);
and U5006 (N_5006,N_3660,N_2162);
and U5007 (N_5007,N_3827,N_2300);
and U5008 (N_5008,N_2605,N_2469);
or U5009 (N_5009,N_3880,N_3457);
and U5010 (N_5010,N_3818,N_3239);
and U5011 (N_5011,N_3483,N_2402);
nand U5012 (N_5012,N_2069,N_2060);
nand U5013 (N_5013,N_2402,N_3969);
nor U5014 (N_5014,N_3781,N_2875);
and U5015 (N_5015,N_3722,N_2411);
nand U5016 (N_5016,N_3556,N_2506);
and U5017 (N_5017,N_3243,N_2520);
and U5018 (N_5018,N_2427,N_3325);
xor U5019 (N_5019,N_3802,N_3885);
and U5020 (N_5020,N_3379,N_3408);
nand U5021 (N_5021,N_3312,N_3590);
nand U5022 (N_5022,N_2075,N_3908);
xnor U5023 (N_5023,N_3522,N_3940);
and U5024 (N_5024,N_2237,N_3951);
and U5025 (N_5025,N_2146,N_2269);
nand U5026 (N_5026,N_2099,N_3002);
nand U5027 (N_5027,N_2826,N_3224);
or U5028 (N_5028,N_3807,N_2202);
and U5029 (N_5029,N_2381,N_3507);
and U5030 (N_5030,N_2660,N_3547);
and U5031 (N_5031,N_3498,N_3678);
nand U5032 (N_5032,N_3877,N_2528);
nand U5033 (N_5033,N_3902,N_2785);
or U5034 (N_5034,N_3576,N_3490);
and U5035 (N_5035,N_2328,N_3635);
and U5036 (N_5036,N_3169,N_2183);
nand U5037 (N_5037,N_3345,N_2811);
nor U5038 (N_5038,N_3612,N_2546);
nand U5039 (N_5039,N_2932,N_2597);
and U5040 (N_5040,N_3543,N_3180);
nand U5041 (N_5041,N_3563,N_3451);
and U5042 (N_5042,N_2557,N_3849);
xnor U5043 (N_5043,N_3746,N_2514);
nand U5044 (N_5044,N_2582,N_2544);
or U5045 (N_5045,N_2393,N_2778);
xnor U5046 (N_5046,N_3545,N_3249);
and U5047 (N_5047,N_2996,N_3440);
nor U5048 (N_5048,N_3315,N_2710);
nand U5049 (N_5049,N_2676,N_3074);
nand U5050 (N_5050,N_3682,N_3713);
and U5051 (N_5051,N_2536,N_3633);
or U5052 (N_5052,N_3543,N_3076);
and U5053 (N_5053,N_2830,N_2045);
xnor U5054 (N_5054,N_2692,N_2053);
nand U5055 (N_5055,N_3141,N_3634);
and U5056 (N_5056,N_2911,N_3390);
nand U5057 (N_5057,N_2646,N_2803);
nor U5058 (N_5058,N_2726,N_3793);
or U5059 (N_5059,N_3504,N_3307);
and U5060 (N_5060,N_3664,N_2316);
nor U5061 (N_5061,N_2639,N_3700);
or U5062 (N_5062,N_2592,N_2297);
or U5063 (N_5063,N_3907,N_2622);
nand U5064 (N_5064,N_2827,N_3989);
xor U5065 (N_5065,N_3129,N_2663);
xnor U5066 (N_5066,N_2244,N_2977);
nor U5067 (N_5067,N_2527,N_2195);
nand U5068 (N_5068,N_2730,N_2258);
nor U5069 (N_5069,N_3201,N_2740);
xor U5070 (N_5070,N_2334,N_2562);
and U5071 (N_5071,N_2237,N_3560);
xor U5072 (N_5072,N_2510,N_3403);
xnor U5073 (N_5073,N_3988,N_2790);
nor U5074 (N_5074,N_3523,N_3965);
and U5075 (N_5075,N_2721,N_3041);
and U5076 (N_5076,N_3502,N_2898);
and U5077 (N_5077,N_2343,N_3907);
nor U5078 (N_5078,N_3052,N_3277);
nand U5079 (N_5079,N_3025,N_3188);
or U5080 (N_5080,N_2713,N_3969);
nand U5081 (N_5081,N_3213,N_2917);
nor U5082 (N_5082,N_3669,N_2428);
nor U5083 (N_5083,N_2031,N_3429);
or U5084 (N_5084,N_2924,N_3955);
or U5085 (N_5085,N_3390,N_2149);
xor U5086 (N_5086,N_2022,N_3313);
and U5087 (N_5087,N_3755,N_2336);
and U5088 (N_5088,N_2081,N_2968);
nand U5089 (N_5089,N_3637,N_3412);
or U5090 (N_5090,N_3521,N_3569);
nor U5091 (N_5091,N_3193,N_3583);
nand U5092 (N_5092,N_3759,N_2709);
xor U5093 (N_5093,N_3644,N_3768);
nor U5094 (N_5094,N_2031,N_2537);
nor U5095 (N_5095,N_3567,N_2300);
xor U5096 (N_5096,N_3747,N_2403);
nor U5097 (N_5097,N_3294,N_2620);
and U5098 (N_5098,N_3326,N_2589);
nand U5099 (N_5099,N_3317,N_2682);
nand U5100 (N_5100,N_2907,N_2852);
nor U5101 (N_5101,N_2657,N_3465);
nand U5102 (N_5102,N_3210,N_2232);
or U5103 (N_5103,N_3659,N_3521);
or U5104 (N_5104,N_2750,N_2660);
nor U5105 (N_5105,N_2957,N_3647);
or U5106 (N_5106,N_2270,N_2076);
or U5107 (N_5107,N_2148,N_2864);
nor U5108 (N_5108,N_2691,N_2106);
and U5109 (N_5109,N_3558,N_3373);
or U5110 (N_5110,N_3917,N_2191);
and U5111 (N_5111,N_3998,N_2703);
or U5112 (N_5112,N_3292,N_2833);
nand U5113 (N_5113,N_3998,N_3729);
and U5114 (N_5114,N_2678,N_2985);
nor U5115 (N_5115,N_3067,N_2564);
and U5116 (N_5116,N_2123,N_2864);
and U5117 (N_5117,N_3941,N_2665);
xnor U5118 (N_5118,N_3067,N_3892);
nand U5119 (N_5119,N_2675,N_2922);
nand U5120 (N_5120,N_2349,N_2900);
nand U5121 (N_5121,N_2692,N_2042);
xor U5122 (N_5122,N_3055,N_3303);
or U5123 (N_5123,N_2536,N_2121);
and U5124 (N_5124,N_3179,N_3232);
nor U5125 (N_5125,N_2737,N_2138);
xnor U5126 (N_5126,N_2847,N_2797);
nor U5127 (N_5127,N_2167,N_3823);
nand U5128 (N_5128,N_3162,N_3077);
nand U5129 (N_5129,N_2665,N_3923);
nand U5130 (N_5130,N_2603,N_3937);
or U5131 (N_5131,N_3580,N_3019);
nand U5132 (N_5132,N_2269,N_2377);
or U5133 (N_5133,N_2628,N_2484);
and U5134 (N_5134,N_2761,N_3917);
and U5135 (N_5135,N_2342,N_2021);
or U5136 (N_5136,N_3583,N_2095);
nor U5137 (N_5137,N_2444,N_2124);
nor U5138 (N_5138,N_3850,N_2185);
nor U5139 (N_5139,N_3516,N_3259);
or U5140 (N_5140,N_3140,N_2873);
and U5141 (N_5141,N_2342,N_3347);
or U5142 (N_5142,N_3021,N_2446);
nand U5143 (N_5143,N_2373,N_2604);
or U5144 (N_5144,N_2086,N_3524);
nor U5145 (N_5145,N_3301,N_2726);
nand U5146 (N_5146,N_3349,N_2934);
nand U5147 (N_5147,N_3726,N_3089);
and U5148 (N_5148,N_2528,N_2458);
xor U5149 (N_5149,N_2060,N_3317);
or U5150 (N_5150,N_2617,N_3318);
nand U5151 (N_5151,N_3901,N_2328);
xnor U5152 (N_5152,N_3009,N_3532);
nand U5153 (N_5153,N_2515,N_2160);
and U5154 (N_5154,N_2083,N_2725);
nor U5155 (N_5155,N_3884,N_3951);
nand U5156 (N_5156,N_2864,N_2853);
nor U5157 (N_5157,N_2139,N_3728);
nor U5158 (N_5158,N_3118,N_3394);
nor U5159 (N_5159,N_3158,N_3206);
nor U5160 (N_5160,N_2230,N_3246);
and U5161 (N_5161,N_3712,N_2790);
nand U5162 (N_5162,N_3288,N_3248);
xor U5163 (N_5163,N_2501,N_2021);
or U5164 (N_5164,N_2625,N_2210);
and U5165 (N_5165,N_2903,N_2071);
or U5166 (N_5166,N_2609,N_2987);
or U5167 (N_5167,N_3975,N_2454);
nor U5168 (N_5168,N_2215,N_2439);
nand U5169 (N_5169,N_3356,N_3729);
and U5170 (N_5170,N_2654,N_3172);
nor U5171 (N_5171,N_2218,N_2654);
nand U5172 (N_5172,N_2310,N_2280);
nand U5173 (N_5173,N_3641,N_3485);
xor U5174 (N_5174,N_3345,N_2327);
nand U5175 (N_5175,N_3001,N_2012);
or U5176 (N_5176,N_2392,N_3589);
nor U5177 (N_5177,N_2148,N_2952);
xor U5178 (N_5178,N_2209,N_3572);
nand U5179 (N_5179,N_3791,N_3022);
nor U5180 (N_5180,N_3884,N_3983);
or U5181 (N_5181,N_2963,N_3978);
nor U5182 (N_5182,N_3733,N_2622);
nor U5183 (N_5183,N_3677,N_3995);
nor U5184 (N_5184,N_3285,N_3650);
or U5185 (N_5185,N_2401,N_2298);
nor U5186 (N_5186,N_3606,N_2387);
nand U5187 (N_5187,N_3801,N_2788);
or U5188 (N_5188,N_3169,N_2901);
nand U5189 (N_5189,N_2634,N_3182);
nand U5190 (N_5190,N_2041,N_2218);
nor U5191 (N_5191,N_3593,N_2216);
nand U5192 (N_5192,N_2466,N_2278);
and U5193 (N_5193,N_2879,N_3275);
nor U5194 (N_5194,N_3192,N_2699);
and U5195 (N_5195,N_2148,N_3109);
and U5196 (N_5196,N_3927,N_3173);
nor U5197 (N_5197,N_3969,N_3326);
and U5198 (N_5198,N_3273,N_3167);
nand U5199 (N_5199,N_3342,N_2611);
xor U5200 (N_5200,N_2554,N_2039);
nor U5201 (N_5201,N_3858,N_2980);
and U5202 (N_5202,N_2581,N_2221);
or U5203 (N_5203,N_2466,N_2106);
nor U5204 (N_5204,N_3982,N_2045);
xnor U5205 (N_5205,N_2067,N_2287);
nand U5206 (N_5206,N_3231,N_2475);
nor U5207 (N_5207,N_3153,N_2688);
and U5208 (N_5208,N_3653,N_3675);
or U5209 (N_5209,N_2797,N_2829);
nor U5210 (N_5210,N_2118,N_2275);
and U5211 (N_5211,N_2534,N_3261);
nor U5212 (N_5212,N_2984,N_3883);
nand U5213 (N_5213,N_2723,N_3118);
nand U5214 (N_5214,N_2436,N_2388);
xnor U5215 (N_5215,N_3109,N_2508);
nand U5216 (N_5216,N_3604,N_3193);
and U5217 (N_5217,N_2280,N_3077);
nand U5218 (N_5218,N_2632,N_2904);
nor U5219 (N_5219,N_3547,N_2995);
or U5220 (N_5220,N_3139,N_3135);
nand U5221 (N_5221,N_2494,N_2825);
and U5222 (N_5222,N_2818,N_2489);
and U5223 (N_5223,N_3969,N_2268);
nor U5224 (N_5224,N_3261,N_3879);
or U5225 (N_5225,N_2299,N_3502);
nor U5226 (N_5226,N_2341,N_2449);
or U5227 (N_5227,N_3393,N_2066);
or U5228 (N_5228,N_2851,N_3212);
nand U5229 (N_5229,N_3152,N_3296);
and U5230 (N_5230,N_3921,N_3956);
or U5231 (N_5231,N_3515,N_2763);
xor U5232 (N_5232,N_2740,N_2850);
nor U5233 (N_5233,N_3272,N_3257);
nor U5234 (N_5234,N_3646,N_2469);
xor U5235 (N_5235,N_3155,N_3788);
and U5236 (N_5236,N_2790,N_3485);
nand U5237 (N_5237,N_3471,N_2075);
or U5238 (N_5238,N_3584,N_3190);
nor U5239 (N_5239,N_3065,N_3849);
and U5240 (N_5240,N_3755,N_2975);
nor U5241 (N_5241,N_3518,N_2270);
nand U5242 (N_5242,N_3325,N_3231);
nand U5243 (N_5243,N_3655,N_3741);
and U5244 (N_5244,N_3857,N_2133);
nand U5245 (N_5245,N_3985,N_2624);
nand U5246 (N_5246,N_3981,N_3168);
and U5247 (N_5247,N_2988,N_3610);
or U5248 (N_5248,N_3126,N_2958);
nor U5249 (N_5249,N_3700,N_2583);
nor U5250 (N_5250,N_2790,N_3658);
nor U5251 (N_5251,N_3455,N_2207);
nor U5252 (N_5252,N_3947,N_3043);
and U5253 (N_5253,N_2070,N_2135);
nand U5254 (N_5254,N_3788,N_3569);
or U5255 (N_5255,N_2718,N_2209);
nor U5256 (N_5256,N_3677,N_3471);
and U5257 (N_5257,N_3130,N_2601);
nor U5258 (N_5258,N_2393,N_3235);
nor U5259 (N_5259,N_2247,N_3374);
and U5260 (N_5260,N_3056,N_3130);
or U5261 (N_5261,N_3168,N_2356);
nand U5262 (N_5262,N_2265,N_2809);
and U5263 (N_5263,N_3968,N_3709);
nor U5264 (N_5264,N_2268,N_3805);
xor U5265 (N_5265,N_2396,N_2862);
nand U5266 (N_5266,N_3723,N_2869);
nand U5267 (N_5267,N_2333,N_2953);
or U5268 (N_5268,N_3981,N_2329);
nand U5269 (N_5269,N_3098,N_2303);
or U5270 (N_5270,N_2039,N_2527);
and U5271 (N_5271,N_3084,N_2594);
nor U5272 (N_5272,N_3946,N_3409);
and U5273 (N_5273,N_3210,N_3620);
and U5274 (N_5274,N_3441,N_2810);
and U5275 (N_5275,N_2202,N_3449);
and U5276 (N_5276,N_2119,N_3200);
nor U5277 (N_5277,N_3262,N_2459);
and U5278 (N_5278,N_2290,N_3887);
nand U5279 (N_5279,N_3338,N_3110);
nand U5280 (N_5280,N_2984,N_2844);
and U5281 (N_5281,N_3924,N_2852);
and U5282 (N_5282,N_3274,N_3316);
or U5283 (N_5283,N_3259,N_2684);
nand U5284 (N_5284,N_3947,N_2783);
nor U5285 (N_5285,N_3498,N_2414);
nor U5286 (N_5286,N_2105,N_3104);
and U5287 (N_5287,N_2161,N_3834);
or U5288 (N_5288,N_2031,N_2247);
or U5289 (N_5289,N_3785,N_2335);
or U5290 (N_5290,N_3846,N_2766);
nand U5291 (N_5291,N_3079,N_2316);
nor U5292 (N_5292,N_2034,N_3249);
or U5293 (N_5293,N_3100,N_2951);
nand U5294 (N_5294,N_3184,N_3222);
and U5295 (N_5295,N_2583,N_2123);
and U5296 (N_5296,N_2348,N_2950);
xor U5297 (N_5297,N_3976,N_3738);
nor U5298 (N_5298,N_2303,N_3060);
nand U5299 (N_5299,N_2126,N_3626);
or U5300 (N_5300,N_2014,N_3134);
or U5301 (N_5301,N_2805,N_3209);
or U5302 (N_5302,N_3895,N_3336);
and U5303 (N_5303,N_2757,N_3652);
xnor U5304 (N_5304,N_2355,N_3214);
or U5305 (N_5305,N_3891,N_3412);
nand U5306 (N_5306,N_2259,N_3786);
nor U5307 (N_5307,N_3123,N_3560);
and U5308 (N_5308,N_2664,N_3726);
nand U5309 (N_5309,N_2605,N_3027);
nor U5310 (N_5310,N_3279,N_2580);
nand U5311 (N_5311,N_2536,N_2476);
and U5312 (N_5312,N_3646,N_3464);
or U5313 (N_5313,N_3135,N_3540);
nor U5314 (N_5314,N_2287,N_3721);
and U5315 (N_5315,N_2109,N_2239);
or U5316 (N_5316,N_3403,N_3645);
or U5317 (N_5317,N_3475,N_3369);
or U5318 (N_5318,N_2752,N_3387);
nor U5319 (N_5319,N_3671,N_2948);
nor U5320 (N_5320,N_2169,N_3666);
nor U5321 (N_5321,N_3912,N_3309);
nor U5322 (N_5322,N_2840,N_3340);
and U5323 (N_5323,N_2226,N_2302);
and U5324 (N_5324,N_3799,N_3010);
or U5325 (N_5325,N_2151,N_3597);
xor U5326 (N_5326,N_2081,N_3645);
xnor U5327 (N_5327,N_2759,N_2329);
nand U5328 (N_5328,N_2880,N_3914);
nand U5329 (N_5329,N_3059,N_2370);
xor U5330 (N_5330,N_2469,N_3697);
nand U5331 (N_5331,N_2470,N_2747);
xnor U5332 (N_5332,N_2268,N_3290);
or U5333 (N_5333,N_2151,N_3538);
nor U5334 (N_5334,N_3949,N_2584);
or U5335 (N_5335,N_3045,N_3886);
nand U5336 (N_5336,N_2103,N_3018);
or U5337 (N_5337,N_2731,N_2944);
nor U5338 (N_5338,N_3950,N_3874);
nor U5339 (N_5339,N_3920,N_3025);
and U5340 (N_5340,N_3197,N_2269);
or U5341 (N_5341,N_3051,N_2060);
and U5342 (N_5342,N_3874,N_2030);
and U5343 (N_5343,N_3083,N_3883);
nor U5344 (N_5344,N_3603,N_3703);
nand U5345 (N_5345,N_3685,N_2662);
or U5346 (N_5346,N_3253,N_3752);
and U5347 (N_5347,N_2061,N_3453);
and U5348 (N_5348,N_3905,N_3470);
nand U5349 (N_5349,N_3838,N_2304);
nor U5350 (N_5350,N_3664,N_3192);
nand U5351 (N_5351,N_2491,N_2578);
nor U5352 (N_5352,N_2880,N_3076);
nand U5353 (N_5353,N_2115,N_3601);
or U5354 (N_5354,N_2792,N_2897);
nand U5355 (N_5355,N_3345,N_2902);
and U5356 (N_5356,N_2801,N_2772);
nor U5357 (N_5357,N_2066,N_2166);
nor U5358 (N_5358,N_2833,N_2197);
and U5359 (N_5359,N_3490,N_2665);
or U5360 (N_5360,N_2109,N_2481);
nand U5361 (N_5361,N_2896,N_2968);
nand U5362 (N_5362,N_2799,N_3437);
nor U5363 (N_5363,N_2262,N_2261);
and U5364 (N_5364,N_3876,N_2716);
nand U5365 (N_5365,N_3666,N_2004);
nand U5366 (N_5366,N_2255,N_3225);
nor U5367 (N_5367,N_3121,N_3057);
nand U5368 (N_5368,N_3280,N_2456);
or U5369 (N_5369,N_3793,N_2028);
or U5370 (N_5370,N_3249,N_2838);
nand U5371 (N_5371,N_3334,N_3482);
nor U5372 (N_5372,N_3939,N_3556);
and U5373 (N_5373,N_2356,N_3566);
nor U5374 (N_5374,N_2985,N_3142);
or U5375 (N_5375,N_2892,N_3145);
or U5376 (N_5376,N_3672,N_2129);
or U5377 (N_5377,N_2203,N_3094);
and U5378 (N_5378,N_2965,N_2167);
or U5379 (N_5379,N_2634,N_2921);
or U5380 (N_5380,N_3957,N_2022);
nand U5381 (N_5381,N_2552,N_2362);
or U5382 (N_5382,N_3580,N_3949);
or U5383 (N_5383,N_2213,N_2037);
nor U5384 (N_5384,N_2062,N_2279);
xnor U5385 (N_5385,N_3033,N_3582);
nor U5386 (N_5386,N_3845,N_2867);
nand U5387 (N_5387,N_3417,N_2034);
or U5388 (N_5388,N_2458,N_3768);
and U5389 (N_5389,N_2346,N_3443);
or U5390 (N_5390,N_3023,N_3156);
xnor U5391 (N_5391,N_3361,N_2559);
nor U5392 (N_5392,N_2858,N_2970);
nor U5393 (N_5393,N_3386,N_3825);
nand U5394 (N_5394,N_2029,N_3202);
nor U5395 (N_5395,N_3126,N_2621);
nand U5396 (N_5396,N_3687,N_2761);
nor U5397 (N_5397,N_2177,N_2688);
or U5398 (N_5398,N_2965,N_3169);
xor U5399 (N_5399,N_3262,N_3264);
nor U5400 (N_5400,N_3548,N_2959);
or U5401 (N_5401,N_2935,N_2493);
nand U5402 (N_5402,N_2518,N_2525);
nor U5403 (N_5403,N_3626,N_3655);
and U5404 (N_5404,N_3512,N_2521);
nor U5405 (N_5405,N_3118,N_3921);
nor U5406 (N_5406,N_2419,N_3693);
and U5407 (N_5407,N_2497,N_3678);
or U5408 (N_5408,N_3001,N_2366);
and U5409 (N_5409,N_3731,N_2408);
xnor U5410 (N_5410,N_3928,N_3104);
and U5411 (N_5411,N_3366,N_3885);
nand U5412 (N_5412,N_3377,N_2795);
nand U5413 (N_5413,N_3676,N_2534);
and U5414 (N_5414,N_2357,N_2934);
nor U5415 (N_5415,N_3368,N_2498);
and U5416 (N_5416,N_2526,N_3709);
nand U5417 (N_5417,N_2840,N_2201);
nor U5418 (N_5418,N_3706,N_2708);
nor U5419 (N_5419,N_3409,N_2654);
nor U5420 (N_5420,N_2559,N_2915);
and U5421 (N_5421,N_3920,N_3060);
nand U5422 (N_5422,N_3592,N_2255);
and U5423 (N_5423,N_3931,N_2907);
or U5424 (N_5424,N_3391,N_3181);
nand U5425 (N_5425,N_3575,N_3849);
and U5426 (N_5426,N_3139,N_3580);
nor U5427 (N_5427,N_2468,N_2285);
or U5428 (N_5428,N_3873,N_3399);
or U5429 (N_5429,N_3108,N_3539);
or U5430 (N_5430,N_2064,N_3896);
and U5431 (N_5431,N_2442,N_2679);
nand U5432 (N_5432,N_3460,N_3150);
and U5433 (N_5433,N_3063,N_3266);
and U5434 (N_5434,N_2243,N_3821);
and U5435 (N_5435,N_2569,N_3668);
nand U5436 (N_5436,N_3342,N_3161);
xor U5437 (N_5437,N_2258,N_2007);
xnor U5438 (N_5438,N_2879,N_2148);
and U5439 (N_5439,N_3639,N_3670);
nand U5440 (N_5440,N_3080,N_3440);
nor U5441 (N_5441,N_2022,N_2052);
and U5442 (N_5442,N_3776,N_3242);
nor U5443 (N_5443,N_2216,N_3125);
or U5444 (N_5444,N_3387,N_3521);
nand U5445 (N_5445,N_2146,N_2143);
or U5446 (N_5446,N_2396,N_3526);
or U5447 (N_5447,N_2539,N_3080);
nor U5448 (N_5448,N_3717,N_2805);
and U5449 (N_5449,N_3689,N_3383);
xor U5450 (N_5450,N_2818,N_2984);
nor U5451 (N_5451,N_2395,N_2955);
and U5452 (N_5452,N_2853,N_2571);
and U5453 (N_5453,N_2497,N_2137);
nand U5454 (N_5454,N_3883,N_2704);
or U5455 (N_5455,N_3336,N_3154);
and U5456 (N_5456,N_2127,N_2671);
nand U5457 (N_5457,N_2724,N_3454);
and U5458 (N_5458,N_2042,N_3574);
or U5459 (N_5459,N_3036,N_2378);
xnor U5460 (N_5460,N_3514,N_3967);
or U5461 (N_5461,N_3431,N_2120);
nor U5462 (N_5462,N_3843,N_2298);
or U5463 (N_5463,N_2948,N_2416);
and U5464 (N_5464,N_3353,N_2060);
or U5465 (N_5465,N_3614,N_3668);
nor U5466 (N_5466,N_2127,N_3355);
nor U5467 (N_5467,N_3116,N_3070);
nor U5468 (N_5468,N_2868,N_3505);
nor U5469 (N_5469,N_2861,N_2742);
nor U5470 (N_5470,N_3444,N_2060);
or U5471 (N_5471,N_2614,N_2896);
and U5472 (N_5472,N_2318,N_3562);
nand U5473 (N_5473,N_3862,N_2522);
or U5474 (N_5474,N_3055,N_2450);
xnor U5475 (N_5475,N_2109,N_2148);
and U5476 (N_5476,N_3494,N_3113);
and U5477 (N_5477,N_2669,N_2698);
and U5478 (N_5478,N_3808,N_3421);
or U5479 (N_5479,N_2261,N_3355);
and U5480 (N_5480,N_3325,N_3042);
nor U5481 (N_5481,N_2323,N_3291);
nor U5482 (N_5482,N_3685,N_2340);
and U5483 (N_5483,N_3304,N_3429);
or U5484 (N_5484,N_2992,N_3872);
nor U5485 (N_5485,N_3529,N_3592);
xor U5486 (N_5486,N_3476,N_2775);
nor U5487 (N_5487,N_3462,N_3750);
or U5488 (N_5488,N_2981,N_3513);
nor U5489 (N_5489,N_2439,N_2198);
nand U5490 (N_5490,N_3976,N_3792);
xor U5491 (N_5491,N_3166,N_3184);
or U5492 (N_5492,N_2539,N_2925);
nand U5493 (N_5493,N_3712,N_3416);
and U5494 (N_5494,N_2598,N_2436);
and U5495 (N_5495,N_2966,N_3180);
nand U5496 (N_5496,N_3647,N_2490);
and U5497 (N_5497,N_2887,N_2738);
and U5498 (N_5498,N_3765,N_2892);
or U5499 (N_5499,N_3961,N_3049);
nand U5500 (N_5500,N_2357,N_3592);
or U5501 (N_5501,N_3871,N_2798);
and U5502 (N_5502,N_3986,N_2452);
nor U5503 (N_5503,N_3596,N_3516);
nor U5504 (N_5504,N_2060,N_3954);
nor U5505 (N_5505,N_3588,N_3261);
nand U5506 (N_5506,N_2299,N_2522);
nor U5507 (N_5507,N_2880,N_3654);
nand U5508 (N_5508,N_3749,N_2167);
or U5509 (N_5509,N_3306,N_2839);
nor U5510 (N_5510,N_2782,N_2605);
or U5511 (N_5511,N_2855,N_2875);
nor U5512 (N_5512,N_2143,N_3195);
nor U5513 (N_5513,N_3333,N_2593);
nand U5514 (N_5514,N_2643,N_3308);
xor U5515 (N_5515,N_3140,N_3276);
or U5516 (N_5516,N_3777,N_2495);
or U5517 (N_5517,N_2289,N_3377);
nand U5518 (N_5518,N_3777,N_2971);
or U5519 (N_5519,N_2447,N_3782);
nor U5520 (N_5520,N_3197,N_3620);
nand U5521 (N_5521,N_2326,N_2944);
and U5522 (N_5522,N_3397,N_2816);
or U5523 (N_5523,N_2058,N_3621);
or U5524 (N_5524,N_2315,N_3701);
or U5525 (N_5525,N_3195,N_2761);
and U5526 (N_5526,N_3951,N_3221);
nor U5527 (N_5527,N_3350,N_3441);
and U5528 (N_5528,N_2738,N_2472);
nand U5529 (N_5529,N_3078,N_2435);
nand U5530 (N_5530,N_2903,N_3681);
nor U5531 (N_5531,N_2827,N_2980);
nor U5532 (N_5532,N_2104,N_3344);
nand U5533 (N_5533,N_2018,N_2837);
nor U5534 (N_5534,N_3845,N_2704);
nand U5535 (N_5535,N_2303,N_3302);
or U5536 (N_5536,N_3265,N_3734);
or U5537 (N_5537,N_3563,N_2961);
nor U5538 (N_5538,N_3986,N_3078);
nand U5539 (N_5539,N_2717,N_2833);
and U5540 (N_5540,N_2078,N_2642);
nor U5541 (N_5541,N_2786,N_2666);
or U5542 (N_5542,N_3666,N_3255);
and U5543 (N_5543,N_2634,N_2547);
nor U5544 (N_5544,N_2184,N_2861);
nand U5545 (N_5545,N_3020,N_2279);
nand U5546 (N_5546,N_2775,N_2180);
nor U5547 (N_5547,N_3036,N_2561);
or U5548 (N_5548,N_2802,N_2576);
or U5549 (N_5549,N_3528,N_3047);
nand U5550 (N_5550,N_2247,N_2616);
nor U5551 (N_5551,N_3032,N_3289);
and U5552 (N_5552,N_3570,N_2404);
nor U5553 (N_5553,N_2913,N_2764);
nor U5554 (N_5554,N_3945,N_2382);
xor U5555 (N_5555,N_2235,N_2780);
xnor U5556 (N_5556,N_3358,N_3165);
nor U5557 (N_5557,N_3194,N_2509);
nand U5558 (N_5558,N_2700,N_2089);
or U5559 (N_5559,N_3267,N_2010);
or U5560 (N_5560,N_3107,N_2859);
and U5561 (N_5561,N_2272,N_2670);
nor U5562 (N_5562,N_2262,N_2184);
nor U5563 (N_5563,N_2646,N_3340);
nor U5564 (N_5564,N_3101,N_3301);
or U5565 (N_5565,N_2235,N_3626);
or U5566 (N_5566,N_3368,N_2308);
or U5567 (N_5567,N_3855,N_2141);
or U5568 (N_5568,N_3735,N_2800);
nand U5569 (N_5569,N_2233,N_3896);
nor U5570 (N_5570,N_2777,N_2964);
and U5571 (N_5571,N_3741,N_2918);
xnor U5572 (N_5572,N_3963,N_3192);
nor U5573 (N_5573,N_3453,N_3320);
nor U5574 (N_5574,N_3260,N_2831);
and U5575 (N_5575,N_3275,N_2721);
and U5576 (N_5576,N_2852,N_3878);
nand U5577 (N_5577,N_3584,N_3349);
nor U5578 (N_5578,N_2502,N_3579);
nand U5579 (N_5579,N_2274,N_3441);
or U5580 (N_5580,N_2464,N_2069);
and U5581 (N_5581,N_2912,N_2987);
xnor U5582 (N_5582,N_3546,N_3817);
and U5583 (N_5583,N_2831,N_2956);
xor U5584 (N_5584,N_2192,N_2502);
or U5585 (N_5585,N_3674,N_2763);
xor U5586 (N_5586,N_2836,N_3384);
or U5587 (N_5587,N_2454,N_2668);
nand U5588 (N_5588,N_2570,N_2767);
or U5589 (N_5589,N_3903,N_2453);
and U5590 (N_5590,N_2184,N_3070);
nand U5591 (N_5591,N_3998,N_3246);
xnor U5592 (N_5592,N_3537,N_3353);
nor U5593 (N_5593,N_2036,N_2088);
and U5594 (N_5594,N_3528,N_2361);
nor U5595 (N_5595,N_3266,N_3122);
nand U5596 (N_5596,N_3227,N_3876);
nor U5597 (N_5597,N_3355,N_2184);
nand U5598 (N_5598,N_3284,N_2299);
nor U5599 (N_5599,N_2950,N_2965);
and U5600 (N_5600,N_2049,N_2902);
and U5601 (N_5601,N_2946,N_3158);
or U5602 (N_5602,N_2972,N_2556);
nand U5603 (N_5603,N_3630,N_2981);
nor U5604 (N_5604,N_3174,N_3297);
xor U5605 (N_5605,N_2108,N_2326);
nor U5606 (N_5606,N_2965,N_3267);
or U5607 (N_5607,N_2123,N_2989);
and U5608 (N_5608,N_2747,N_3092);
nor U5609 (N_5609,N_2148,N_3796);
nor U5610 (N_5610,N_3722,N_2135);
or U5611 (N_5611,N_3828,N_3759);
nor U5612 (N_5612,N_3932,N_3266);
and U5613 (N_5613,N_3262,N_2839);
and U5614 (N_5614,N_3602,N_3486);
or U5615 (N_5615,N_2237,N_3269);
nor U5616 (N_5616,N_2417,N_2121);
or U5617 (N_5617,N_2032,N_2878);
or U5618 (N_5618,N_2625,N_2812);
or U5619 (N_5619,N_2446,N_3033);
or U5620 (N_5620,N_3838,N_2805);
nor U5621 (N_5621,N_2453,N_3346);
xor U5622 (N_5622,N_2481,N_3411);
nor U5623 (N_5623,N_3919,N_3456);
or U5624 (N_5624,N_2996,N_2727);
xor U5625 (N_5625,N_2797,N_2835);
and U5626 (N_5626,N_2747,N_3171);
nand U5627 (N_5627,N_2458,N_2374);
nand U5628 (N_5628,N_3769,N_2815);
or U5629 (N_5629,N_2681,N_2959);
nor U5630 (N_5630,N_2873,N_3321);
nand U5631 (N_5631,N_2719,N_2084);
and U5632 (N_5632,N_2509,N_2912);
nor U5633 (N_5633,N_2522,N_2179);
nor U5634 (N_5634,N_2943,N_3611);
or U5635 (N_5635,N_3466,N_2549);
and U5636 (N_5636,N_2452,N_2906);
nand U5637 (N_5637,N_2360,N_3926);
or U5638 (N_5638,N_3712,N_3008);
nand U5639 (N_5639,N_2959,N_2055);
or U5640 (N_5640,N_3593,N_3959);
nand U5641 (N_5641,N_2092,N_2225);
or U5642 (N_5642,N_3957,N_3977);
and U5643 (N_5643,N_2536,N_3464);
nor U5644 (N_5644,N_2919,N_3557);
nor U5645 (N_5645,N_3884,N_2102);
and U5646 (N_5646,N_2260,N_3006);
and U5647 (N_5647,N_3628,N_2212);
and U5648 (N_5648,N_2563,N_2300);
nor U5649 (N_5649,N_2697,N_2239);
nor U5650 (N_5650,N_2291,N_3673);
nand U5651 (N_5651,N_3428,N_3480);
nor U5652 (N_5652,N_3748,N_3993);
and U5653 (N_5653,N_2432,N_2819);
and U5654 (N_5654,N_3380,N_2923);
nor U5655 (N_5655,N_2971,N_3249);
nor U5656 (N_5656,N_2175,N_2801);
nand U5657 (N_5657,N_3052,N_3576);
and U5658 (N_5658,N_3027,N_3281);
nand U5659 (N_5659,N_3970,N_2172);
nor U5660 (N_5660,N_2182,N_2157);
nor U5661 (N_5661,N_2986,N_3647);
xor U5662 (N_5662,N_2571,N_3193);
and U5663 (N_5663,N_2973,N_2302);
nand U5664 (N_5664,N_2226,N_3219);
and U5665 (N_5665,N_3705,N_3975);
or U5666 (N_5666,N_3770,N_2298);
nor U5667 (N_5667,N_2064,N_3173);
or U5668 (N_5668,N_3716,N_3298);
or U5669 (N_5669,N_2265,N_3866);
nor U5670 (N_5670,N_3415,N_2942);
or U5671 (N_5671,N_3363,N_3908);
and U5672 (N_5672,N_2689,N_3441);
nand U5673 (N_5673,N_3148,N_2191);
and U5674 (N_5674,N_3147,N_2735);
nand U5675 (N_5675,N_2424,N_3799);
or U5676 (N_5676,N_2840,N_3441);
or U5677 (N_5677,N_2549,N_2676);
xnor U5678 (N_5678,N_2521,N_2253);
and U5679 (N_5679,N_2935,N_3300);
nand U5680 (N_5680,N_2191,N_3190);
nor U5681 (N_5681,N_2215,N_2229);
xnor U5682 (N_5682,N_2018,N_3664);
nand U5683 (N_5683,N_3849,N_2833);
nor U5684 (N_5684,N_2630,N_2159);
nor U5685 (N_5685,N_2553,N_2463);
and U5686 (N_5686,N_2091,N_3692);
nor U5687 (N_5687,N_2280,N_2664);
or U5688 (N_5688,N_3860,N_3132);
nor U5689 (N_5689,N_2357,N_3872);
or U5690 (N_5690,N_3679,N_3816);
or U5691 (N_5691,N_2802,N_3509);
nand U5692 (N_5692,N_2368,N_3319);
nand U5693 (N_5693,N_2572,N_2807);
xnor U5694 (N_5694,N_3117,N_2563);
xnor U5695 (N_5695,N_3202,N_3722);
nand U5696 (N_5696,N_2784,N_2114);
nand U5697 (N_5697,N_2607,N_3191);
nor U5698 (N_5698,N_2871,N_3371);
and U5699 (N_5699,N_3517,N_2131);
or U5700 (N_5700,N_3628,N_3224);
and U5701 (N_5701,N_3223,N_2290);
xor U5702 (N_5702,N_3222,N_2509);
and U5703 (N_5703,N_3991,N_2642);
nand U5704 (N_5704,N_3488,N_3910);
or U5705 (N_5705,N_3753,N_2703);
nand U5706 (N_5706,N_3958,N_3101);
and U5707 (N_5707,N_2737,N_2934);
nor U5708 (N_5708,N_2158,N_2048);
nand U5709 (N_5709,N_3034,N_3390);
and U5710 (N_5710,N_2660,N_3999);
xnor U5711 (N_5711,N_3493,N_3944);
nor U5712 (N_5712,N_3113,N_2720);
and U5713 (N_5713,N_2417,N_3444);
and U5714 (N_5714,N_2715,N_3242);
or U5715 (N_5715,N_2163,N_2852);
and U5716 (N_5716,N_3885,N_3739);
nand U5717 (N_5717,N_3960,N_3444);
or U5718 (N_5718,N_2509,N_3601);
xnor U5719 (N_5719,N_3188,N_2188);
nand U5720 (N_5720,N_2964,N_2607);
xor U5721 (N_5721,N_3812,N_2453);
or U5722 (N_5722,N_3014,N_2181);
and U5723 (N_5723,N_3518,N_2959);
xor U5724 (N_5724,N_2217,N_2194);
or U5725 (N_5725,N_3766,N_2569);
nand U5726 (N_5726,N_3361,N_2429);
nand U5727 (N_5727,N_3553,N_3685);
and U5728 (N_5728,N_3278,N_3967);
nand U5729 (N_5729,N_2273,N_2072);
or U5730 (N_5730,N_2791,N_3372);
or U5731 (N_5731,N_2837,N_3829);
and U5732 (N_5732,N_3735,N_3250);
nand U5733 (N_5733,N_2882,N_2048);
xnor U5734 (N_5734,N_2779,N_3651);
xnor U5735 (N_5735,N_2177,N_3982);
nor U5736 (N_5736,N_2973,N_3253);
or U5737 (N_5737,N_2710,N_2459);
nand U5738 (N_5738,N_3751,N_3202);
nor U5739 (N_5739,N_2149,N_2519);
nand U5740 (N_5740,N_3740,N_2298);
and U5741 (N_5741,N_2831,N_3115);
nand U5742 (N_5742,N_3815,N_2902);
nor U5743 (N_5743,N_3649,N_2140);
nor U5744 (N_5744,N_3925,N_3257);
or U5745 (N_5745,N_3131,N_2653);
or U5746 (N_5746,N_2825,N_2858);
or U5747 (N_5747,N_2812,N_2754);
nor U5748 (N_5748,N_2682,N_2117);
and U5749 (N_5749,N_3258,N_2211);
or U5750 (N_5750,N_3099,N_2548);
xnor U5751 (N_5751,N_3236,N_2588);
and U5752 (N_5752,N_3374,N_2074);
xor U5753 (N_5753,N_3384,N_2536);
and U5754 (N_5754,N_3054,N_2145);
and U5755 (N_5755,N_2017,N_3735);
or U5756 (N_5756,N_3294,N_2837);
and U5757 (N_5757,N_3906,N_3772);
nand U5758 (N_5758,N_3003,N_3668);
nor U5759 (N_5759,N_3140,N_3999);
nand U5760 (N_5760,N_2888,N_2059);
xor U5761 (N_5761,N_3428,N_2138);
nor U5762 (N_5762,N_2945,N_2934);
nor U5763 (N_5763,N_3026,N_3072);
nand U5764 (N_5764,N_3696,N_3443);
and U5765 (N_5765,N_2217,N_2252);
nor U5766 (N_5766,N_3281,N_2439);
nor U5767 (N_5767,N_3322,N_2222);
or U5768 (N_5768,N_2563,N_3549);
or U5769 (N_5769,N_3813,N_3746);
nand U5770 (N_5770,N_2778,N_3740);
and U5771 (N_5771,N_3212,N_2926);
xor U5772 (N_5772,N_2082,N_3261);
nand U5773 (N_5773,N_3651,N_3696);
nand U5774 (N_5774,N_3434,N_2083);
nand U5775 (N_5775,N_2854,N_3627);
nand U5776 (N_5776,N_2776,N_3506);
nand U5777 (N_5777,N_3882,N_2522);
xor U5778 (N_5778,N_2388,N_3567);
nor U5779 (N_5779,N_3593,N_2478);
xor U5780 (N_5780,N_3660,N_2340);
nand U5781 (N_5781,N_3689,N_3941);
nand U5782 (N_5782,N_2499,N_2341);
nand U5783 (N_5783,N_3063,N_2512);
and U5784 (N_5784,N_3769,N_3838);
and U5785 (N_5785,N_2234,N_2952);
and U5786 (N_5786,N_3693,N_2906);
nor U5787 (N_5787,N_2419,N_2194);
nor U5788 (N_5788,N_2883,N_2662);
and U5789 (N_5789,N_2600,N_2252);
and U5790 (N_5790,N_3126,N_2932);
nand U5791 (N_5791,N_2121,N_3077);
and U5792 (N_5792,N_2772,N_3865);
or U5793 (N_5793,N_3791,N_3861);
nor U5794 (N_5794,N_3337,N_2752);
or U5795 (N_5795,N_3433,N_2228);
nor U5796 (N_5796,N_3640,N_3625);
and U5797 (N_5797,N_2046,N_2611);
or U5798 (N_5798,N_3176,N_2001);
nand U5799 (N_5799,N_2641,N_2986);
nor U5800 (N_5800,N_2238,N_3042);
and U5801 (N_5801,N_2814,N_2893);
or U5802 (N_5802,N_2946,N_3169);
nand U5803 (N_5803,N_3242,N_2728);
nand U5804 (N_5804,N_3898,N_3502);
and U5805 (N_5805,N_2609,N_3070);
nand U5806 (N_5806,N_3437,N_3572);
nand U5807 (N_5807,N_2536,N_3923);
nand U5808 (N_5808,N_3997,N_2260);
or U5809 (N_5809,N_3517,N_2687);
nor U5810 (N_5810,N_2205,N_3403);
nand U5811 (N_5811,N_3352,N_2297);
nor U5812 (N_5812,N_3503,N_2552);
nor U5813 (N_5813,N_2947,N_2130);
nor U5814 (N_5814,N_3237,N_3357);
and U5815 (N_5815,N_3282,N_3187);
xnor U5816 (N_5816,N_2738,N_3217);
and U5817 (N_5817,N_2571,N_3937);
nand U5818 (N_5818,N_2550,N_3481);
xor U5819 (N_5819,N_3577,N_3523);
nand U5820 (N_5820,N_3219,N_2040);
or U5821 (N_5821,N_2138,N_2547);
nand U5822 (N_5822,N_3749,N_3945);
nand U5823 (N_5823,N_2051,N_2412);
and U5824 (N_5824,N_2324,N_3376);
nand U5825 (N_5825,N_2268,N_3165);
nor U5826 (N_5826,N_2114,N_3306);
nor U5827 (N_5827,N_3738,N_2490);
or U5828 (N_5828,N_3343,N_2416);
or U5829 (N_5829,N_2675,N_2254);
and U5830 (N_5830,N_3907,N_2005);
nor U5831 (N_5831,N_3755,N_3398);
or U5832 (N_5832,N_3568,N_2045);
and U5833 (N_5833,N_2889,N_3121);
and U5834 (N_5834,N_2834,N_2687);
nand U5835 (N_5835,N_2680,N_3789);
and U5836 (N_5836,N_2013,N_2185);
or U5837 (N_5837,N_3164,N_3951);
nor U5838 (N_5838,N_2548,N_2507);
and U5839 (N_5839,N_3584,N_2761);
nor U5840 (N_5840,N_3569,N_2597);
and U5841 (N_5841,N_3866,N_3588);
nand U5842 (N_5842,N_2205,N_2963);
nor U5843 (N_5843,N_3481,N_3414);
or U5844 (N_5844,N_3550,N_2146);
nand U5845 (N_5845,N_2943,N_3851);
or U5846 (N_5846,N_2114,N_2475);
and U5847 (N_5847,N_2570,N_3718);
xor U5848 (N_5848,N_2462,N_3105);
xnor U5849 (N_5849,N_2253,N_2379);
or U5850 (N_5850,N_3685,N_2217);
or U5851 (N_5851,N_2763,N_2762);
and U5852 (N_5852,N_2288,N_2637);
and U5853 (N_5853,N_2179,N_2418);
xnor U5854 (N_5854,N_3410,N_2778);
and U5855 (N_5855,N_2763,N_2993);
and U5856 (N_5856,N_3540,N_2116);
nand U5857 (N_5857,N_2476,N_2190);
and U5858 (N_5858,N_3003,N_3782);
nor U5859 (N_5859,N_2594,N_3345);
or U5860 (N_5860,N_2312,N_3763);
nor U5861 (N_5861,N_3964,N_3046);
nor U5862 (N_5862,N_2281,N_3244);
nand U5863 (N_5863,N_3400,N_2899);
nand U5864 (N_5864,N_3798,N_3369);
nand U5865 (N_5865,N_2318,N_2755);
nand U5866 (N_5866,N_3733,N_2307);
and U5867 (N_5867,N_2378,N_2590);
nor U5868 (N_5868,N_2865,N_2920);
nor U5869 (N_5869,N_2390,N_2094);
nor U5870 (N_5870,N_2053,N_3572);
nand U5871 (N_5871,N_2765,N_2333);
nand U5872 (N_5872,N_3290,N_2052);
nand U5873 (N_5873,N_3303,N_3611);
or U5874 (N_5874,N_3587,N_3488);
and U5875 (N_5875,N_2349,N_2302);
nand U5876 (N_5876,N_2064,N_3876);
nor U5877 (N_5877,N_3997,N_2436);
xor U5878 (N_5878,N_2764,N_2575);
or U5879 (N_5879,N_2304,N_2635);
and U5880 (N_5880,N_2001,N_2822);
nor U5881 (N_5881,N_3653,N_2018);
or U5882 (N_5882,N_3903,N_3218);
nand U5883 (N_5883,N_3424,N_2234);
or U5884 (N_5884,N_2834,N_3129);
xor U5885 (N_5885,N_2387,N_3347);
nor U5886 (N_5886,N_3432,N_2557);
or U5887 (N_5887,N_3157,N_3720);
and U5888 (N_5888,N_3628,N_2423);
nand U5889 (N_5889,N_3564,N_2614);
and U5890 (N_5890,N_2993,N_3164);
nor U5891 (N_5891,N_2035,N_3457);
and U5892 (N_5892,N_2773,N_3350);
nand U5893 (N_5893,N_2506,N_2134);
and U5894 (N_5894,N_3005,N_2119);
nand U5895 (N_5895,N_3398,N_2245);
nand U5896 (N_5896,N_2246,N_3011);
or U5897 (N_5897,N_2095,N_3630);
nand U5898 (N_5898,N_2405,N_2289);
nor U5899 (N_5899,N_2578,N_3933);
and U5900 (N_5900,N_3133,N_2331);
xnor U5901 (N_5901,N_2889,N_2156);
nor U5902 (N_5902,N_3893,N_2456);
nand U5903 (N_5903,N_3532,N_2641);
or U5904 (N_5904,N_3972,N_2189);
or U5905 (N_5905,N_3275,N_2234);
nor U5906 (N_5906,N_2396,N_2528);
and U5907 (N_5907,N_3916,N_3497);
and U5908 (N_5908,N_3808,N_3728);
nand U5909 (N_5909,N_3789,N_3317);
nand U5910 (N_5910,N_2694,N_2169);
nor U5911 (N_5911,N_3879,N_3581);
nand U5912 (N_5912,N_2450,N_2900);
or U5913 (N_5913,N_3889,N_2121);
or U5914 (N_5914,N_3008,N_3055);
nor U5915 (N_5915,N_2449,N_3051);
xor U5916 (N_5916,N_2604,N_2842);
and U5917 (N_5917,N_2586,N_3378);
and U5918 (N_5918,N_2564,N_3044);
and U5919 (N_5919,N_3635,N_2959);
or U5920 (N_5920,N_3587,N_2039);
xnor U5921 (N_5921,N_3909,N_3389);
xnor U5922 (N_5922,N_3699,N_3955);
nand U5923 (N_5923,N_2929,N_2370);
nand U5924 (N_5924,N_2810,N_2184);
and U5925 (N_5925,N_3679,N_2044);
or U5926 (N_5926,N_2166,N_2147);
or U5927 (N_5927,N_3282,N_3121);
or U5928 (N_5928,N_3640,N_2788);
or U5929 (N_5929,N_3109,N_2743);
or U5930 (N_5930,N_3294,N_2612);
nand U5931 (N_5931,N_2069,N_2676);
nand U5932 (N_5932,N_2674,N_2954);
and U5933 (N_5933,N_3193,N_3332);
and U5934 (N_5934,N_2115,N_2018);
and U5935 (N_5935,N_3070,N_2320);
and U5936 (N_5936,N_3970,N_2239);
xnor U5937 (N_5937,N_2017,N_2006);
and U5938 (N_5938,N_2577,N_3087);
and U5939 (N_5939,N_2759,N_3598);
or U5940 (N_5940,N_3546,N_2915);
xnor U5941 (N_5941,N_3775,N_3192);
nor U5942 (N_5942,N_2850,N_2361);
nor U5943 (N_5943,N_3484,N_3553);
or U5944 (N_5944,N_2361,N_2825);
and U5945 (N_5945,N_2979,N_3397);
nand U5946 (N_5946,N_3175,N_3369);
nand U5947 (N_5947,N_2554,N_3968);
nor U5948 (N_5948,N_2018,N_3103);
xor U5949 (N_5949,N_3128,N_3913);
or U5950 (N_5950,N_2314,N_2173);
or U5951 (N_5951,N_3944,N_2310);
xor U5952 (N_5952,N_2621,N_2494);
xnor U5953 (N_5953,N_2593,N_3018);
nor U5954 (N_5954,N_3321,N_3890);
xor U5955 (N_5955,N_3456,N_2039);
or U5956 (N_5956,N_2470,N_3283);
or U5957 (N_5957,N_3892,N_2290);
and U5958 (N_5958,N_2351,N_3693);
nand U5959 (N_5959,N_3998,N_2500);
nor U5960 (N_5960,N_2773,N_2314);
and U5961 (N_5961,N_2308,N_2930);
or U5962 (N_5962,N_2488,N_2081);
and U5963 (N_5963,N_2940,N_2472);
and U5964 (N_5964,N_3211,N_3990);
xnor U5965 (N_5965,N_3814,N_2909);
or U5966 (N_5966,N_3619,N_3130);
nor U5967 (N_5967,N_2272,N_2050);
and U5968 (N_5968,N_2259,N_2266);
nand U5969 (N_5969,N_2823,N_2226);
nor U5970 (N_5970,N_3854,N_2584);
or U5971 (N_5971,N_3653,N_3769);
nand U5972 (N_5972,N_3294,N_2713);
nor U5973 (N_5973,N_2657,N_2413);
nand U5974 (N_5974,N_3641,N_2609);
nand U5975 (N_5975,N_2543,N_2605);
nand U5976 (N_5976,N_2014,N_2674);
nand U5977 (N_5977,N_3862,N_3936);
nor U5978 (N_5978,N_3722,N_2013);
nor U5979 (N_5979,N_2281,N_3254);
nor U5980 (N_5980,N_2514,N_2120);
or U5981 (N_5981,N_3781,N_2220);
nand U5982 (N_5982,N_3717,N_2447);
nand U5983 (N_5983,N_2018,N_3537);
nor U5984 (N_5984,N_2092,N_2619);
and U5985 (N_5985,N_2406,N_3391);
and U5986 (N_5986,N_3911,N_2344);
nand U5987 (N_5987,N_3774,N_2367);
xnor U5988 (N_5988,N_2985,N_2045);
or U5989 (N_5989,N_3956,N_3881);
or U5990 (N_5990,N_2539,N_2650);
nand U5991 (N_5991,N_2947,N_3857);
or U5992 (N_5992,N_2984,N_2432);
nor U5993 (N_5993,N_2884,N_2928);
nand U5994 (N_5994,N_2138,N_3761);
nor U5995 (N_5995,N_2177,N_3851);
nand U5996 (N_5996,N_2917,N_3656);
nand U5997 (N_5997,N_3740,N_3074);
or U5998 (N_5998,N_2582,N_3065);
or U5999 (N_5999,N_3456,N_2306);
nor U6000 (N_6000,N_5338,N_4414);
nand U6001 (N_6001,N_5875,N_4003);
nand U6002 (N_6002,N_5166,N_4220);
nor U6003 (N_6003,N_4671,N_4288);
or U6004 (N_6004,N_5915,N_4664);
nor U6005 (N_6005,N_4468,N_5836);
and U6006 (N_6006,N_5137,N_4890);
nor U6007 (N_6007,N_5202,N_5860);
and U6008 (N_6008,N_4542,N_4294);
nand U6009 (N_6009,N_4802,N_4804);
or U6010 (N_6010,N_4669,N_5061);
and U6011 (N_6011,N_4856,N_4160);
nor U6012 (N_6012,N_4501,N_5211);
or U6013 (N_6013,N_5617,N_5120);
and U6014 (N_6014,N_4008,N_4385);
nor U6015 (N_6015,N_5932,N_4038);
or U6016 (N_6016,N_4833,N_4982);
nor U6017 (N_6017,N_5995,N_5079);
and U6018 (N_6018,N_4720,N_5019);
nor U6019 (N_6019,N_4550,N_4048);
nand U6020 (N_6020,N_5601,N_5741);
nand U6021 (N_6021,N_4739,N_4445);
nand U6022 (N_6022,N_5411,N_4015);
or U6023 (N_6023,N_4123,N_4309);
and U6024 (N_6024,N_5893,N_5378);
and U6025 (N_6025,N_4749,N_5027);
nand U6026 (N_6026,N_5450,N_4692);
and U6027 (N_6027,N_5577,N_4311);
or U6028 (N_6028,N_4539,N_5827);
xnor U6029 (N_6029,N_5650,N_5623);
xor U6030 (N_6030,N_5538,N_4180);
or U6031 (N_6031,N_4226,N_4054);
and U6032 (N_6032,N_4926,N_5606);
nor U6033 (N_6033,N_4987,N_5585);
or U6034 (N_6034,N_5908,N_5635);
nor U6035 (N_6035,N_5221,N_4505);
and U6036 (N_6036,N_5196,N_5907);
nand U6037 (N_6037,N_5543,N_4570);
xor U6038 (N_6038,N_4830,N_5064);
and U6039 (N_6039,N_4456,N_5700);
or U6040 (N_6040,N_4246,N_5541);
and U6041 (N_6041,N_4057,N_5399);
xor U6042 (N_6042,N_4346,N_4829);
and U6043 (N_6043,N_5573,N_5274);
or U6044 (N_6044,N_5036,N_5212);
and U6045 (N_6045,N_4431,N_4460);
nand U6046 (N_6046,N_5158,N_4217);
nor U6047 (N_6047,N_4243,N_5840);
or U6048 (N_6048,N_5763,N_4238);
xnor U6049 (N_6049,N_4183,N_5754);
nand U6050 (N_6050,N_5356,N_5990);
nor U6051 (N_6051,N_4549,N_5613);
nor U6052 (N_6052,N_5765,N_5997);
or U6053 (N_6053,N_5928,N_4757);
xor U6054 (N_6054,N_4489,N_4188);
or U6055 (N_6055,N_5375,N_4134);
nor U6056 (N_6056,N_4167,N_5812);
xnor U6057 (N_6057,N_5420,N_4174);
nand U6058 (N_6058,N_5505,N_4264);
or U6059 (N_6059,N_4016,N_4766);
nand U6060 (N_6060,N_5444,N_4439);
nor U6061 (N_6061,N_4053,N_4083);
nand U6062 (N_6062,N_4703,N_5225);
and U6063 (N_6063,N_5834,N_5746);
or U6064 (N_6064,N_5900,N_4317);
and U6065 (N_6065,N_4098,N_4129);
nand U6066 (N_6066,N_5565,N_4230);
or U6067 (N_6067,N_5764,N_4150);
or U6068 (N_6068,N_4056,N_4882);
and U6069 (N_6069,N_5651,N_5994);
nand U6070 (N_6070,N_4970,N_4981);
nand U6071 (N_6071,N_4168,N_5548);
nor U6072 (N_6072,N_5000,N_4910);
and U6073 (N_6073,N_5798,N_4143);
nand U6074 (N_6074,N_4023,N_5435);
nand U6075 (N_6075,N_5144,N_4801);
or U6076 (N_6076,N_4383,N_5493);
nor U6077 (N_6077,N_4778,N_4303);
or U6078 (N_6078,N_4892,N_5287);
and U6079 (N_6079,N_4117,N_5398);
or U6080 (N_6080,N_4787,N_4300);
and U6081 (N_6081,N_4088,N_4957);
and U6082 (N_6082,N_4058,N_5434);
nor U6083 (N_6083,N_4396,N_4625);
xnor U6084 (N_6084,N_4965,N_5696);
nand U6085 (N_6085,N_5920,N_5269);
or U6086 (N_6086,N_5286,N_4518);
and U6087 (N_6087,N_4603,N_4421);
nor U6088 (N_6088,N_5239,N_5261);
nor U6089 (N_6089,N_5597,N_5030);
nand U6090 (N_6090,N_4667,N_5666);
nand U6091 (N_6091,N_4477,N_4363);
and U6092 (N_6092,N_5627,N_4797);
and U6093 (N_6093,N_4320,N_5664);
nor U6094 (N_6094,N_5360,N_5410);
and U6095 (N_6095,N_4478,N_4194);
nand U6096 (N_6096,N_5561,N_5800);
xnor U6097 (N_6097,N_5340,N_4722);
nor U6098 (N_6098,N_5169,N_5583);
or U6099 (N_6099,N_5751,N_4086);
and U6100 (N_6100,N_4263,N_5742);
or U6101 (N_6101,N_4103,N_5766);
nor U6102 (N_6102,N_4480,N_5039);
and U6103 (N_6103,N_5107,N_4277);
xnor U6104 (N_6104,N_5319,N_5544);
nand U6105 (N_6105,N_5524,N_4213);
or U6106 (N_6106,N_4257,N_5949);
or U6107 (N_6107,N_5222,N_5619);
nand U6108 (N_6108,N_5453,N_4157);
or U6109 (N_6109,N_4869,N_5887);
or U6110 (N_6110,N_4712,N_5787);
xnor U6111 (N_6111,N_5018,N_4607);
and U6112 (N_6112,N_4052,N_5810);
or U6113 (N_6113,N_4163,N_5026);
nor U6114 (N_6114,N_4398,N_5084);
or U6115 (N_6115,N_4716,N_4545);
or U6116 (N_6116,N_5686,N_4350);
or U6117 (N_6117,N_4292,N_5953);
nor U6118 (N_6118,N_5255,N_4784);
nor U6119 (N_6119,N_5251,N_4474);
or U6120 (N_6120,N_4629,N_5587);
nand U6121 (N_6121,N_5526,N_5494);
and U6122 (N_6122,N_4858,N_5406);
or U6123 (N_6123,N_5404,N_5760);
and U6124 (N_6124,N_4064,N_4295);
or U6125 (N_6125,N_5337,N_5795);
xor U6126 (N_6126,N_5189,N_4792);
nand U6127 (N_6127,N_4028,N_4321);
and U6128 (N_6128,N_4921,N_5752);
or U6129 (N_6129,N_4424,N_4281);
and U6130 (N_6130,N_5886,N_5046);
or U6131 (N_6131,N_5841,N_5940);
and U6132 (N_6132,N_5271,N_4777);
nand U6133 (N_6133,N_5258,N_4872);
and U6134 (N_6134,N_4336,N_4914);
nor U6135 (N_6135,N_5514,N_5710);
xor U6136 (N_6136,N_4151,N_5910);
nand U6137 (N_6137,N_4632,N_4630);
or U6138 (N_6138,N_5558,N_5096);
and U6139 (N_6139,N_5067,N_5880);
nand U6140 (N_6140,N_4517,N_5111);
or U6141 (N_6141,N_5888,N_5794);
nand U6142 (N_6142,N_5807,N_4218);
nand U6143 (N_6143,N_4090,N_4837);
and U6144 (N_6144,N_4759,N_4031);
or U6145 (N_6145,N_5648,N_4041);
nor U6146 (N_6146,N_5391,N_5244);
or U6147 (N_6147,N_5102,N_4822);
and U6148 (N_6148,N_4568,N_4106);
nor U6149 (N_6149,N_4108,N_5466);
nor U6150 (N_6150,N_4679,N_5618);
or U6151 (N_6151,N_5223,N_5140);
nand U6152 (N_6152,N_5173,N_4340);
xnor U6153 (N_6153,N_5489,N_5925);
and U6154 (N_6154,N_5599,N_4659);
or U6155 (N_6155,N_4475,N_5233);
nand U6156 (N_6156,N_4237,N_4532);
nor U6157 (N_6157,N_5304,N_5724);
and U6158 (N_6158,N_4100,N_4627);
or U6159 (N_6159,N_5778,N_5121);
nand U6160 (N_6160,N_5495,N_5820);
nor U6161 (N_6161,N_5072,N_4061);
nand U6162 (N_6162,N_4197,N_5693);
nor U6163 (N_6163,N_5793,N_5625);
xnor U6164 (N_6164,N_5151,N_4484);
nand U6165 (N_6165,N_5715,N_5339);
or U6166 (N_6166,N_4933,N_4932);
nand U6167 (N_6167,N_4618,N_5328);
or U6168 (N_6168,N_4771,N_4588);
or U6169 (N_6169,N_4844,N_5732);
xor U6170 (N_6170,N_5503,N_5791);
xnor U6171 (N_6171,N_4206,N_4533);
xnor U6172 (N_6172,N_5642,N_4683);
nand U6173 (N_6173,N_4345,N_4121);
nand U6174 (N_6174,N_5331,N_5591);
and U6175 (N_6175,N_5769,N_5872);
and U6176 (N_6176,N_5197,N_4190);
or U6177 (N_6177,N_4794,N_4668);
nor U6178 (N_6178,N_5245,N_5954);
and U6179 (N_6179,N_5939,N_4595);
nor U6180 (N_6180,N_4462,N_5744);
and U6181 (N_6181,N_4769,N_4556);
nand U6182 (N_6182,N_4620,N_4455);
and U6183 (N_6183,N_4196,N_5262);
nand U6184 (N_6184,N_4762,N_5534);
xnor U6185 (N_6185,N_4327,N_5971);
xor U6186 (N_6186,N_5981,N_5032);
xor U6187 (N_6187,N_4552,N_5329);
nand U6188 (N_6188,N_4063,N_4084);
or U6189 (N_6189,N_5332,N_5057);
nand U6190 (N_6190,N_4405,N_4242);
nand U6191 (N_6191,N_5437,N_5813);
nand U6192 (N_6192,N_4075,N_5240);
or U6193 (N_6193,N_5230,N_4723);
or U6194 (N_6194,N_5458,N_5736);
nor U6195 (N_6195,N_4947,N_4419);
and U6196 (N_6196,N_4099,N_4073);
nor U6197 (N_6197,N_5238,N_5743);
and U6198 (N_6198,N_4389,N_5659);
nor U6199 (N_6199,N_4172,N_4537);
or U6200 (N_6200,N_5870,N_4354);
and U6201 (N_6201,N_5101,N_5403);
nor U6202 (N_6202,N_4258,N_5695);
nor U6203 (N_6203,N_4347,N_5848);
or U6204 (N_6204,N_4262,N_4225);
and U6205 (N_6205,N_5014,N_5816);
nor U6206 (N_6206,N_4840,N_5361);
nor U6207 (N_6207,N_5143,N_5692);
and U6208 (N_6208,N_5883,N_5414);
nor U6209 (N_6209,N_5963,N_4156);
nand U6210 (N_6210,N_5445,N_4516);
and U6211 (N_6211,N_5074,N_5707);
nand U6212 (N_6212,N_4254,N_4753);
nand U6213 (N_6213,N_4409,N_4531);
nor U6214 (N_6214,N_5839,N_5967);
nor U6215 (N_6215,N_5242,N_5578);
or U6216 (N_6216,N_4316,N_4481);
and U6217 (N_6217,N_4875,N_5308);
and U6218 (N_6218,N_5837,N_4373);
nand U6219 (N_6219,N_5347,N_5063);
and U6220 (N_6220,N_5980,N_4381);
or U6221 (N_6221,N_4724,N_5809);
or U6222 (N_6222,N_4265,N_4789);
nor U6223 (N_6223,N_4996,N_5139);
or U6224 (N_6224,N_4181,N_5138);
nor U6225 (N_6225,N_4706,N_4461);
xnor U6226 (N_6226,N_4368,N_4298);
xnor U6227 (N_6227,N_4865,N_5824);
nand U6228 (N_6228,N_5673,N_4575);
or U6229 (N_6229,N_5348,N_5785);
and U6230 (N_6230,N_4096,N_5106);
nand U6231 (N_6231,N_4142,N_4847);
nand U6232 (N_6232,N_4813,N_4644);
or U6233 (N_6233,N_4535,N_5232);
nand U6234 (N_6234,N_4135,N_5250);
xnor U6235 (N_6235,N_4714,N_4170);
xnor U6236 (N_6236,N_5449,N_4102);
or U6237 (N_6237,N_5124,N_4818);
nor U6238 (N_6238,N_4042,N_5297);
nor U6239 (N_6239,N_4912,N_4558);
and U6240 (N_6240,N_5210,N_5964);
and U6241 (N_6241,N_5969,N_5116);
nor U6242 (N_6242,N_5080,N_4171);
and U6243 (N_6243,N_5480,N_4945);
or U6244 (N_6244,N_4110,N_5996);
nand U6245 (N_6245,N_5610,N_5060);
and U6246 (N_6246,N_5048,N_4602);
or U6247 (N_6247,N_5085,N_4325);
or U6248 (N_6248,N_5713,N_4029);
nand U6249 (N_6249,N_5652,N_5934);
nand U6250 (N_6250,N_5772,N_4826);
and U6251 (N_6251,N_5277,N_4189);
nand U6252 (N_6252,N_4105,N_5640);
nand U6253 (N_6253,N_5010,N_5464);
nor U6254 (N_6254,N_5560,N_5002);
nand U6255 (N_6255,N_5914,N_4357);
nor U6256 (N_6256,N_4546,N_5598);
and U6257 (N_6257,N_4293,N_5845);
nor U6258 (N_6258,N_4423,N_4819);
xnor U6259 (N_6259,N_4919,N_4718);
nand U6260 (N_6260,N_5334,N_5336);
or U6261 (N_6261,N_5656,N_5866);
or U6262 (N_6262,N_5525,N_5719);
nor U6263 (N_6263,N_4686,N_4879);
nand U6264 (N_6264,N_5823,N_4403);
or U6265 (N_6265,N_5737,N_5115);
and U6266 (N_6266,N_4344,N_5413);
nor U6267 (N_6267,N_4494,N_4782);
and U6268 (N_6268,N_4069,N_5191);
nand U6269 (N_6269,N_4946,N_4074);
or U6270 (N_6270,N_5424,N_4312);
and U6271 (N_6271,N_5916,N_5472);
xor U6272 (N_6272,N_4287,N_4687);
nand U6273 (N_6273,N_5477,N_5564);
and U6274 (N_6274,N_4375,N_5306);
nor U6275 (N_6275,N_5045,N_4304);
or U6276 (N_6276,N_5469,N_5109);
nand U6277 (N_6277,N_5025,N_5344);
and U6278 (N_6278,N_5327,N_4755);
nor U6279 (N_6279,N_4889,N_5438);
xnor U6280 (N_6280,N_5068,N_4394);
and U6281 (N_6281,N_4473,N_4227);
nor U6282 (N_6282,N_5595,N_4235);
or U6283 (N_6283,N_4615,N_5460);
nand U6284 (N_6284,N_5629,N_4988);
nor U6285 (N_6285,N_5050,N_4781);
and U6286 (N_6286,N_4569,N_4365);
or U6287 (N_6287,N_5099,N_4776);
nand U6288 (N_6288,N_5687,N_5885);
nor U6289 (N_6289,N_5055,N_4682);
or U6290 (N_6290,N_4467,N_5976);
or U6291 (N_6291,N_4796,N_4541);
or U6292 (N_6292,N_4124,N_5804);
nand U6293 (N_6293,N_5185,N_4536);
xnor U6294 (N_6294,N_4018,N_4547);
nand U6295 (N_6295,N_5390,N_4348);
or U6296 (N_6296,N_4502,N_4690);
nand U6297 (N_6297,N_5163,N_4415);
and U6298 (N_6298,N_4594,N_4693);
nor U6299 (N_6299,N_4395,N_5141);
nand U6300 (N_6300,N_4922,N_5362);
xnor U6301 (N_6301,N_4775,N_4178);
nor U6302 (N_6302,N_4512,N_4033);
nor U6303 (N_6303,N_4754,N_5432);
nand U6304 (N_6304,N_4047,N_4845);
nand U6305 (N_6305,N_5042,N_5389);
xnor U6306 (N_6306,N_4223,N_5470);
nor U6307 (N_6307,N_4130,N_4200);
nand U6308 (N_6308,N_4485,N_4913);
or U6309 (N_6309,N_5229,N_5318);
or U6310 (N_6310,N_4606,N_5180);
xnor U6311 (N_6311,N_5098,N_5259);
and U6312 (N_6312,N_5755,N_5672);
nor U6313 (N_6313,N_4245,N_5759);
nor U6314 (N_6314,N_5694,N_4049);
nand U6315 (N_6315,N_5966,N_4283);
nand U6316 (N_6316,N_5802,N_4613);
nor U6317 (N_6317,N_5132,N_4772);
or U6318 (N_6318,N_5621,N_5037);
xnor U6319 (N_6319,N_5468,N_4880);
and U6320 (N_6320,N_4930,N_5822);
nand U6321 (N_6321,N_4624,N_5983);
nor U6322 (N_6322,N_5236,N_4068);
or U6323 (N_6323,N_4694,N_5709);
nand U6324 (N_6324,N_4447,N_5545);
or U6325 (N_6325,N_5609,N_4670);
nand U6326 (N_6326,N_4799,N_4944);
nor U6327 (N_6327,N_4622,N_4446);
or U6328 (N_6328,N_5162,N_5868);
nand U6329 (N_6329,N_4162,N_4916);
nor U6330 (N_6330,N_5624,N_5911);
nor U6331 (N_6331,N_4269,N_5083);
and U6332 (N_6332,N_5582,N_5753);
or U6333 (N_6333,N_4806,N_4326);
nand U6334 (N_6334,N_5007,N_5559);
nor U6335 (N_6335,N_4623,N_5706);
and U6336 (N_6336,N_4700,N_5448);
nor U6337 (N_6337,N_4506,N_4486);
nand U6338 (N_6338,N_4175,N_5022);
and U6339 (N_6339,N_5333,N_5090);
nor U6340 (N_6340,N_4356,N_5001);
nand U6341 (N_6341,N_4253,N_4616);
nor U6342 (N_6342,N_4666,N_5523);
nand U6343 (N_6343,N_4490,N_4949);
nand U6344 (N_6344,N_5214,N_4719);
and U6345 (N_6345,N_4885,N_5190);
nand U6346 (N_6346,N_5292,N_5487);
nand U6347 (N_6347,N_5576,N_4995);
nor U6348 (N_6348,N_5838,N_4508);
or U6349 (N_6349,N_4697,N_4332);
nand U6350 (N_6350,N_4585,N_4626);
and U6351 (N_6351,N_4962,N_4593);
nand U6352 (N_6352,N_4990,N_4499);
nor U6353 (N_6353,N_5227,N_5248);
nand U6354 (N_6354,N_4855,N_4852);
or U6355 (N_6355,N_4001,N_5669);
nand U6356 (N_6356,N_5850,N_4884);
and U6357 (N_6357,N_4557,N_5011);
nand U6358 (N_6358,N_5295,N_5588);
xnor U6359 (N_6359,N_4109,N_5462);
nand U6360 (N_6360,N_4634,N_4843);
or U6361 (N_6361,N_4026,N_4521);
nor U6362 (N_6362,N_4094,N_5792);
xor U6363 (N_6363,N_4729,N_4997);
nand U6364 (N_6364,N_4379,N_4425);
nand U6365 (N_6365,N_5913,N_5113);
nand U6366 (N_6366,N_5276,N_4907);
nand U6367 (N_6367,N_5853,N_5518);
and U6368 (N_6368,N_4070,N_5443);
and U6369 (N_6369,N_5433,N_5828);
nand U6370 (N_6370,N_5415,N_5316);
or U6371 (N_6371,N_5796,N_5296);
nor U6372 (N_6372,N_4648,N_4176);
nor U6373 (N_6373,N_5024,N_5641);
nand U6374 (N_6374,N_4768,N_5546);
and U6375 (N_6375,N_4195,N_5510);
nor U6376 (N_6376,N_4184,N_4491);
nand U6377 (N_6377,N_4993,N_5833);
nand U6378 (N_6378,N_4240,N_5569);
and U6379 (N_6379,N_5421,N_4812);
and U6380 (N_6380,N_4544,N_4428);
and U6381 (N_6381,N_5683,N_4451);
nor U6382 (N_6382,N_4915,N_5921);
or U6383 (N_6383,N_4250,N_4654);
or U6384 (N_6384,N_4268,N_5412);
nor U6385 (N_6385,N_5504,N_4816);
or U6386 (N_6386,N_5314,N_4551);
nand U6387 (N_6387,N_4761,N_4011);
or U6388 (N_6388,N_4136,N_4572);
nor U6389 (N_6389,N_4330,N_5726);
nand U6390 (N_6390,N_4685,N_5884);
and U6391 (N_6391,N_4637,N_4967);
nor U6392 (N_6392,N_5771,N_5035);
or U6393 (N_6393,N_5580,N_5728);
or U6394 (N_6394,N_5867,N_5958);
or U6395 (N_6395,N_4931,N_5354);
and U6396 (N_6396,N_4021,N_4393);
nand U6397 (N_6397,N_4495,N_4275);
nand U6398 (N_6398,N_5335,N_5571);
or U6399 (N_6399,N_5408,N_4870);
nor U6400 (N_6400,N_4255,N_4377);
or U6401 (N_6401,N_5734,N_5174);
nand U6402 (N_6402,N_5878,N_5987);
nand U6403 (N_6403,N_5017,N_5442);
and U6404 (N_6404,N_5622,N_4386);
xnor U6405 (N_6405,N_4444,N_5986);
or U6406 (N_6406,N_4927,N_5478);
or U6407 (N_6407,N_5550,N_4305);
and U6408 (N_6408,N_5465,N_5991);
nor U6409 (N_6409,N_4566,N_4208);
nand U6410 (N_6410,N_5178,N_5439);
xnor U6411 (N_6411,N_5890,N_4798);
xnor U6412 (N_6412,N_5697,N_5607);
or U6413 (N_6413,N_5662,N_5467);
or U6414 (N_6414,N_5922,N_5454);
and U6415 (N_6415,N_4929,N_5639);
xor U6416 (N_6416,N_5382,N_5486);
and U6417 (N_6417,N_4387,N_5108);
or U6418 (N_6418,N_4333,N_4645);
and U6419 (N_6419,N_5179,N_5829);
xor U6420 (N_6420,N_4441,N_4203);
or U6421 (N_6421,N_5293,N_5234);
xnor U6422 (N_6422,N_4672,N_5198);
or U6423 (N_6423,N_4120,N_5213);
or U6424 (N_6424,N_4341,N_4113);
or U6425 (N_6425,N_4284,N_4006);
or U6426 (N_6426,N_4448,N_4037);
nand U6427 (N_6427,N_4636,N_5253);
nand U6428 (N_6428,N_5877,N_4740);
and U6429 (N_6429,N_4201,N_5950);
xor U6430 (N_6430,N_4743,N_4482);
and U6431 (N_6431,N_4153,N_4905);
nor U6432 (N_6432,N_5311,N_4342);
or U6433 (N_6433,N_4432,N_5291);
and U6434 (N_6434,N_5509,N_4165);
or U6435 (N_6435,N_5654,N_5135);
nor U6436 (N_6436,N_5906,N_5087);
xnor U6437 (N_6437,N_4874,N_5549);
or U6438 (N_6438,N_5006,N_5671);
nor U6439 (N_6439,N_4586,N_4285);
and U6440 (N_6440,N_4289,N_4902);
and U6441 (N_6441,N_4411,N_4525);
nor U6442 (N_6442,N_5767,N_4097);
nor U6443 (N_6443,N_4527,N_5740);
nand U6444 (N_6444,N_4867,N_4334);
nor U6445 (N_6445,N_5757,N_5423);
nand U6446 (N_6446,N_4891,N_5655);
and U6447 (N_6447,N_5555,N_4752);
or U6448 (N_6448,N_4611,N_5711);
nand U6449 (N_6449,N_4973,N_5149);
xnor U6450 (N_6450,N_5902,N_5858);
nand U6451 (N_6451,N_4435,N_5532);
xor U6452 (N_6452,N_5563,N_5873);
and U6453 (N_6453,N_4941,N_5854);
nand U6454 (N_6454,N_5073,N_5517);
or U6455 (N_6455,N_4115,N_4426);
and U6456 (N_6456,N_5371,N_5547);
nand U6457 (N_6457,N_4515,N_5579);
nor U6458 (N_6458,N_4406,N_4961);
nand U6459 (N_6459,N_4811,N_4564);
nand U6460 (N_6460,N_4315,N_4849);
nor U6461 (N_6461,N_5722,N_4943);
nand U6462 (N_6462,N_4853,N_4252);
nor U6463 (N_6463,N_4555,N_5181);
nand U6464 (N_6464,N_4738,N_5831);
and U6465 (N_6465,N_4689,N_5077);
nor U6466 (N_6466,N_5235,N_5876);
and U6467 (N_6467,N_4571,N_4132);
nor U6468 (N_6468,N_5249,N_5894);
or U6469 (N_6469,N_5630,N_5739);
nand U6470 (N_6470,N_5220,N_4991);
and U6471 (N_6471,N_4876,N_5313);
xnor U6472 (N_6472,N_5041,N_5118);
or U6473 (N_6473,N_4338,N_5370);
and U6474 (N_6474,N_4147,N_4166);
and U6475 (N_6475,N_5170,N_5484);
or U6476 (N_6476,N_4139,N_4886);
and U6477 (N_6477,N_4358,N_4846);
or U6478 (N_6478,N_4024,N_5909);
nand U6479 (N_6479,N_4009,N_5431);
xor U6480 (N_6480,N_5136,N_4600);
or U6481 (N_6481,N_4207,N_5015);
nor U6482 (N_6482,N_5633,N_4040);
nand U6483 (N_6483,N_5537,N_5199);
and U6484 (N_6484,N_5730,N_4133);
and U6485 (N_6485,N_5596,N_4998);
or U6486 (N_6486,N_5680,N_5790);
and U6487 (N_6487,N_4036,N_5372);
or U6488 (N_6488,N_4434,N_4903);
xor U6489 (N_6489,N_4464,N_4917);
xor U6490 (N_6490,N_4361,N_5355);
or U6491 (N_6491,N_5552,N_5407);
xor U6492 (N_6492,N_5756,N_4179);
and U6493 (N_6493,N_4976,N_5069);
nand U6494 (N_6494,N_5643,N_5065);
or U6495 (N_6495,N_5009,N_5270);
nor U6496 (N_6496,N_5044,N_4430);
nand U6497 (N_6497,N_5252,N_4820);
nor U6498 (N_6498,N_4610,N_5033);
nor U6499 (N_6499,N_4887,N_4427);
nor U6500 (N_6500,N_5300,N_4836);
nor U6501 (N_6501,N_5961,N_5342);
nand U6502 (N_6502,N_4051,N_5727);
or U6503 (N_6503,N_5278,N_4067);
nand U6504 (N_6504,N_5944,N_5374);
or U6505 (N_6505,N_4860,N_5243);
nor U6506 (N_6506,N_5703,N_5978);
and U6507 (N_6507,N_4249,N_5119);
nor U6508 (N_6508,N_4701,N_5201);
and U6509 (N_6509,N_5784,N_5531);
nor U6510 (N_6510,N_4509,N_5626);
nand U6511 (N_6511,N_5941,N_5979);
or U6512 (N_6512,N_5636,N_5657);
nand U6513 (N_6513,N_4360,N_5317);
or U6514 (N_6514,N_5658,N_4198);
nand U6515 (N_6515,N_5152,N_4522);
and U6516 (N_6516,N_4906,N_4248);
or U6517 (N_6517,N_5315,N_4511);
nor U6518 (N_6518,N_5681,N_4675);
nor U6519 (N_6519,N_5566,N_4212);
nand U6520 (N_6520,N_5895,N_4408);
nand U6521 (N_6521,N_4635,N_5114);
xnor U6522 (N_6522,N_5473,N_4507);
or U6523 (N_6523,N_4436,N_5684);
nor U6524 (N_6524,N_5951,N_5943);
nor U6525 (N_6525,N_4280,N_5075);
xor U6526 (N_6526,N_5016,N_4193);
nor U6527 (N_6527,N_4000,N_4140);
nor U6528 (N_6528,N_4384,N_5776);
nor U6529 (N_6529,N_5945,N_5447);
nand U6530 (N_6530,N_5843,N_4479);
nor U6531 (N_6531,N_5889,N_5206);
or U6532 (N_6532,N_4442,N_4382);
or U6533 (N_6533,N_4077,N_5955);
or U6534 (N_6534,N_5312,N_5898);
nor U6535 (N_6535,N_4050,N_4737);
and U6536 (N_6536,N_4764,N_4896);
xor U6537 (N_6537,N_5422,N_5156);
nand U6538 (N_6538,N_4433,N_4107);
nor U6539 (N_6539,N_5379,N_5584);
or U6540 (N_6540,N_4873,N_4540);
or U6541 (N_6541,N_4402,N_4391);
and U6542 (N_6542,N_4022,N_5175);
or U6543 (N_6543,N_5040,N_5973);
nor U6544 (N_6544,N_5062,N_5209);
xor U6545 (N_6545,N_4319,N_4487);
nor U6546 (N_6546,N_5305,N_5507);
nor U6547 (N_6547,N_4895,N_4370);
nor U6548 (N_6548,N_5218,N_5070);
or U6549 (N_6549,N_4236,N_4969);
nor U6550 (N_6550,N_5380,N_4986);
nand U6551 (N_6551,N_5499,N_5992);
and U6552 (N_6552,N_5852,N_4786);
and U6553 (N_6553,N_4673,N_5901);
nor U6554 (N_6554,N_5047,N_5299);
or U6555 (N_6555,N_4221,N_4082);
xor U6556 (N_6556,N_4727,N_5615);
nor U6557 (N_6557,N_5704,N_5533);
nor U6558 (N_6558,N_5948,N_4825);
nand U6559 (N_6559,N_5008,N_4958);
xor U6560 (N_6560,N_5999,N_5723);
xor U6561 (N_6561,N_4012,N_5129);
or U6562 (N_6562,N_4019,N_5215);
and U6563 (N_6563,N_4817,N_4647);
nand U6564 (N_6564,N_4144,N_5112);
xnor U6565 (N_6565,N_5265,N_4923);
or U6566 (N_6566,N_4702,N_4814);
nor U6567 (N_6567,N_4631,N_4314);
nand U6568 (N_6568,N_5918,N_5699);
or U6569 (N_6569,N_5965,N_4691);
or U6570 (N_6570,N_5377,N_5803);
nor U6571 (N_6571,N_4695,N_4400);
nand U6572 (N_6572,N_5457,N_4968);
nor U6573 (N_6573,N_4125,N_4824);
or U6574 (N_6574,N_5148,N_5257);
nor U6575 (N_6575,N_4034,N_5428);
xor U6576 (N_6576,N_5511,N_4128);
nand U6577 (N_6577,N_5539,N_4060);
and U6578 (N_6578,N_5436,N_4823);
nor U6579 (N_6579,N_5134,N_4938);
nand U6580 (N_6580,N_5384,N_5301);
nand U6581 (N_6581,N_5401,N_5417);
nand U6582 (N_6582,N_5282,N_5021);
and U6583 (N_6583,N_4587,N_4864);
nand U6584 (N_6584,N_5701,N_5677);
nor U6585 (N_6585,N_5161,N_4095);
and U6586 (N_6586,N_5485,N_4530);
and U6587 (N_6587,N_4114,N_5528);
nor U6588 (N_6588,N_4831,N_5556);
nor U6589 (N_6589,N_5364,N_5307);
or U6590 (N_6590,N_5071,N_4746);
and U6591 (N_6591,N_5678,N_4955);
nor U6592 (N_6592,N_5392,N_5104);
or U6593 (N_6593,N_5052,N_5516);
nor U6594 (N_6594,N_4979,N_4582);
nor U6595 (N_6595,N_5092,N_5957);
and U6596 (N_6596,N_4091,N_4039);
xor U6597 (N_6597,N_4756,N_4299);
or U6598 (N_6598,N_5892,N_4633);
xor U6599 (N_6599,N_4104,N_4747);
or U6600 (N_6600,N_5586,N_5177);
nor U6601 (N_6601,N_5645,N_4247);
or U6602 (N_6602,N_4617,N_4399);
and U6603 (N_6603,N_5649,N_5459);
nand U6604 (N_6604,N_4790,N_5266);
nand U6605 (N_6605,N_4560,N_4563);
and U6606 (N_6606,N_5183,N_4177);
nor U6607 (N_6607,N_4827,N_5634);
or U6608 (N_6608,N_5935,N_5463);
nor U6609 (N_6609,N_5602,N_5679);
or U6610 (N_6610,N_4216,N_5690);
or U6611 (N_6611,N_4210,N_5782);
and U6612 (N_6612,N_5100,N_5646);
and U6613 (N_6613,N_4007,N_4619);
nor U6614 (N_6614,N_4122,N_5110);
nor U6615 (N_6615,N_4025,N_4261);
and U6616 (N_6616,N_5089,N_5912);
nand U6617 (N_6617,N_4032,N_4985);
xor U6618 (N_6618,N_5205,N_4861);
nor U6619 (N_6619,N_4851,N_4388);
or U6620 (N_6620,N_4392,N_4888);
nand U6621 (N_6621,N_5388,N_4653);
and U6622 (N_6622,N_5705,N_4883);
nor U6623 (N_6623,N_5324,N_4821);
nand U6624 (N_6624,N_4717,N_4577);
or U6625 (N_6625,N_5998,N_4751);
and U6626 (N_6626,N_4202,N_5394);
nor U6627 (N_6627,N_5688,N_4848);
nand U6628 (N_6628,N_5325,N_5500);
nor U6629 (N_6629,N_5535,N_5988);
nor U6630 (N_6630,N_5562,N_4677);
or U6631 (N_6631,N_5799,N_5284);
nand U6632 (N_6632,N_5975,N_4800);
nand U6633 (N_6633,N_5302,N_4413);
nor U6634 (N_6634,N_4807,N_5133);
or U6635 (N_6635,N_4500,N_5984);
and U6636 (N_6636,N_4404,N_4035);
and U6637 (N_6637,N_5851,N_5702);
nor U6638 (N_6638,N_5195,N_4978);
and U6639 (N_6639,N_4169,N_4989);
or U6640 (N_6640,N_5446,N_4710);
nand U6641 (N_6641,N_4362,N_5353);
xor U6642 (N_6642,N_4278,N_5184);
xor U6643 (N_6643,N_4939,N_4715);
nor U6644 (N_6644,N_5094,N_5806);
xnor U6645 (N_6645,N_5020,N_5130);
or U6646 (N_6646,N_5721,N_5855);
nor U6647 (N_6647,N_4224,N_4279);
or U6648 (N_6648,N_5346,N_4286);
or U6649 (N_6649,N_5387,N_4452);
nor U6650 (N_6650,N_5691,N_4367);
nand U6651 (N_6651,N_5725,N_4963);
and U6652 (N_6652,N_4553,N_5366);
and U6653 (N_6653,N_5208,N_4964);
and U6654 (N_6654,N_4504,N_4649);
nor U6655 (N_6655,N_4146,N_5761);
xor U6656 (N_6656,N_5519,N_4192);
or U6657 (N_6657,N_4164,N_5279);
and U6658 (N_6658,N_5674,N_5028);
nand U6659 (N_6659,N_5275,N_5665);
and U6660 (N_6660,N_5051,N_5200);
xor U6661 (N_6661,N_5647,N_5430);
and U6662 (N_6662,N_5272,N_5874);
nand U6663 (N_6663,N_5698,N_4005);
nor U6664 (N_6664,N_5038,N_4127);
or U6665 (N_6665,N_4657,N_5357);
nand U6666 (N_6666,N_5747,N_4182);
xnor U6667 (N_6667,N_4731,N_5663);
nor U6668 (N_6668,N_5341,N_4470);
and U6669 (N_6669,N_5859,N_5167);
or U6670 (N_6670,N_5849,N_5054);
and U6671 (N_6671,N_4126,N_5219);
nor U6672 (N_6672,N_5351,N_4092);
or U6673 (N_6673,N_5310,N_5881);
nand U6674 (N_6674,N_5977,N_4046);
or U6675 (N_6675,N_5429,N_5117);
nand U6676 (N_6676,N_5383,N_4578);
nor U6677 (N_6677,N_5508,N_4080);
nand U6678 (N_6678,N_5145,N_4937);
nand U6679 (N_6679,N_5846,N_4418);
or U6680 (N_6680,N_5146,N_5871);
nand U6681 (N_6681,N_5402,N_5122);
xor U6682 (N_6682,N_4276,N_5581);
nor U6683 (N_6683,N_4211,N_4609);
nand U6684 (N_6684,N_5982,N_5942);
xnor U6685 (N_6685,N_5594,N_4897);
nor U6686 (N_6686,N_5590,N_5226);
nor U6687 (N_6687,N_5228,N_5929);
nand U6688 (N_6688,N_5369,N_5280);
nand U6689 (N_6689,N_5376,N_4267);
or U6690 (N_6690,N_4308,N_4688);
xor U6691 (N_6691,N_4137,N_4758);
or U6692 (N_6692,N_5187,N_5830);
nand U6693 (N_6693,N_4204,N_5127);
or U6694 (N_6694,N_5154,N_5427);
nand U6695 (N_6695,N_5749,N_4767);
or U6696 (N_6696,N_5923,N_4471);
or U6697 (N_6697,N_5554,N_4651);
or U6698 (N_6698,N_4828,N_5023);
and U6699 (N_6699,N_5005,N_5817);
or U6700 (N_6700,N_4072,N_5825);
or U6701 (N_6701,N_5689,N_5738);
nor U6702 (N_6702,N_5452,N_5862);
and U6703 (N_6703,N_4323,N_4734);
or U6704 (N_6704,N_4601,N_4270);
and U6705 (N_6705,N_5919,N_5103);
or U6706 (N_6706,N_4791,N_4661);
and U6707 (N_6707,N_5536,N_5400);
or U6708 (N_6708,N_4805,N_4735);
and U6709 (N_6709,N_5350,N_4863);
and U6710 (N_6710,N_4584,N_4656);
and U6711 (N_6711,N_5029,N_4498);
xnor U6712 (N_6712,N_4089,N_5775);
and U6713 (N_6713,N_4854,N_4707);
nor U6714 (N_6714,N_5471,N_5865);
nor U6715 (N_6715,N_4523,N_4894);
nor U6716 (N_6716,N_4158,N_5078);
nand U6717 (N_6717,N_5298,N_5363);
or U6718 (N_6718,N_4959,N_4788);
xnor U6719 (N_6719,N_5530,N_4936);
and U6720 (N_6720,N_5086,N_4972);
nand U6721 (N_6721,N_4810,N_4256);
nand U6722 (N_6722,N_4266,N_4878);
xor U6723 (N_6723,N_5081,N_4960);
nand U6724 (N_6724,N_4119,N_5733);
or U6725 (N_6725,N_5381,N_5637);
and U6726 (N_6726,N_4592,N_5482);
or U6727 (N_6727,N_4380,N_5899);
xnor U6728 (N_6728,N_5515,N_5731);
or U6729 (N_6729,N_4760,N_5474);
or U6730 (N_6730,N_5720,N_4974);
or U6731 (N_6731,N_4138,N_5283);
nand U6732 (N_6732,N_5479,N_4928);
and U6733 (N_6733,N_4598,N_4608);
nor U6734 (N_6734,N_4850,N_4559);
nor U6735 (N_6735,N_4359,N_4841);
nand U6736 (N_6736,N_5644,N_5947);
nand U6737 (N_6737,N_5281,N_5066);
and U6738 (N_6738,N_5289,N_4655);
or U6739 (N_6739,N_4372,N_4526);
nand U6740 (N_6740,N_5612,N_5670);
or U6741 (N_6741,N_5811,N_5638);
and U6742 (N_6742,N_4186,N_4838);
nand U6743 (N_6743,N_4520,N_4925);
nor U6744 (N_6744,N_5611,N_5589);
and U6745 (N_6745,N_4369,N_4343);
xor U6746 (N_6746,N_5352,N_4259);
nor U6747 (N_6747,N_4839,N_5542);
and U6748 (N_6748,N_4770,N_4199);
xnor U6749 (N_6749,N_4222,N_5013);
or U6750 (N_6750,N_4412,N_4793);
or U6751 (N_6751,N_5204,N_4519);
or U6752 (N_6752,N_5451,N_4244);
and U6753 (N_6753,N_5031,N_5685);
nand U6754 (N_6754,N_4899,N_4065);
or U6755 (N_6755,N_5193,N_5551);
or U6756 (N_6756,N_4736,N_4780);
or U6757 (N_6757,N_5676,N_5714);
nor U6758 (N_6758,N_5924,N_4465);
or U6759 (N_6759,N_5962,N_5959);
xnor U6760 (N_6760,N_4641,N_5247);
nor U6761 (N_6761,N_4774,N_4328);
xnor U6762 (N_6762,N_4980,N_5631);
nor U6763 (N_6763,N_5735,N_4364);
or U6764 (N_6764,N_4483,N_4231);
and U6765 (N_6765,N_5632,N_5157);
xor U6766 (N_6766,N_4950,N_4696);
or U6767 (N_6767,N_5405,N_4868);
or U6768 (N_6768,N_5273,N_4185);
and U6769 (N_6769,N_4476,N_5522);
and U6770 (N_6770,N_5093,N_4628);
nand U6771 (N_6771,N_4282,N_4658);
or U6772 (N_6772,N_4161,N_4043);
nand U6773 (N_6773,N_4524,N_5182);
nor U6774 (N_6774,N_4463,N_5832);
nor U6775 (N_6775,N_5491,N_4909);
xnor U6776 (N_6776,N_5131,N_4087);
and U6777 (N_6777,N_4085,N_4866);
nor U6778 (N_6778,N_5821,N_4579);
or U6779 (N_6779,N_4322,N_5989);
nand U6780 (N_6780,N_5770,N_5034);
or U6781 (N_6781,N_5418,N_4859);
nand U6782 (N_6782,N_5574,N_5882);
nor U6783 (N_6783,N_5864,N_5529);
and U6784 (N_6784,N_5168,N_4014);
or U6785 (N_6785,N_4251,N_5256);
and U6786 (N_6786,N_4966,N_5572);
nor U6787 (N_6787,N_4698,N_4145);
nand U6788 (N_6788,N_4599,N_4472);
and U6789 (N_6789,N_5425,N_5956);
nand U6790 (N_6790,N_5176,N_4004);
and U6791 (N_6791,N_5904,N_4862);
nand U6792 (N_6792,N_4842,N_4745);
or U6793 (N_6793,N_4785,N_5294);
nor U6794 (N_6794,N_5675,N_4614);
nor U6795 (N_6795,N_4952,N_4904);
and U6796 (N_6796,N_4612,N_4510);
and U6797 (N_6797,N_5368,N_4030);
nand U6798 (N_6798,N_4597,N_5863);
nor U6799 (N_6799,N_5396,N_4901);
or U6800 (N_6800,N_5773,N_4561);
nand U6801 (N_6801,N_4900,N_5567);
nand U6802 (N_6802,N_4313,N_4676);
nor U6803 (N_6803,N_5203,N_5303);
nor U6804 (N_6804,N_5835,N_5492);
xor U6805 (N_6805,N_5777,N_5668);
nor U6806 (N_6806,N_4159,N_5207);
and U6807 (N_6807,N_5708,N_4748);
nand U6808 (N_6808,N_4589,N_5088);
or U6809 (N_6809,N_5153,N_4378);
or U6810 (N_6810,N_4940,N_4815);
or U6811 (N_6811,N_4335,N_5426);
and U6812 (N_6812,N_5216,N_4834);
nor U6813 (N_6813,N_5779,N_5123);
nor U6814 (N_6814,N_4721,N_4209);
nand U6815 (N_6815,N_5488,N_5501);
xor U6816 (N_6816,N_5513,N_5186);
nor U6817 (N_6817,N_5527,N_5896);
or U6818 (N_6818,N_5521,N_5933);
nor U6819 (N_6819,N_4681,N_5603);
nand U6820 (N_6820,N_4548,N_5224);
nor U6821 (N_6821,N_5105,N_4652);
nand U6822 (N_6822,N_5367,N_4574);
nand U6823 (N_6823,N_5322,N_5575);
or U6824 (N_6824,N_5667,N_5593);
or U6825 (N_6825,N_4497,N_4353);
nor U6826 (N_6826,N_5520,N_5783);
xor U6827 (N_6827,N_5780,N_5267);
and U6828 (N_6828,N_4458,N_5797);
or U6829 (N_6829,N_5891,N_4272);
and U6830 (N_6830,N_4055,N_4116);
xnor U6831 (N_6831,N_4076,N_4239);
nor U6832 (N_6832,N_4438,N_5926);
and U6833 (N_6833,N_5600,N_4044);
nor U6834 (N_6834,N_4646,N_4027);
nor U6835 (N_6835,N_5082,N_5164);
and U6836 (N_6836,N_5058,N_4773);
or U6837 (N_6837,N_5416,N_4410);
or U6838 (N_6838,N_4241,N_5004);
and U6839 (N_6839,N_5805,N_5718);
or U6840 (N_6840,N_5952,N_5155);
and U6841 (N_6841,N_4215,N_5540);
and U6842 (N_6842,N_5661,N_4573);
and U6843 (N_6843,N_5897,N_4062);
nand U6844 (N_6844,N_4013,N_5241);
nand U6845 (N_6845,N_4954,N_5917);
or U6846 (N_6846,N_4407,N_5320);
nand U6847 (N_6847,N_5268,N_4449);
and U6848 (N_6848,N_5049,N_4352);
nand U6849 (N_6849,N_5254,N_5604);
and U6850 (N_6850,N_4492,N_5774);
or U6851 (N_6851,N_4148,N_5856);
and U6852 (N_6852,N_4078,N_5490);
xnor U6853 (N_6853,N_5869,N_4741);
and U6854 (N_6854,N_4554,N_4877);
or U6855 (N_6855,N_5616,N_4401);
and U6856 (N_6856,N_4643,N_4081);
or U6857 (N_6857,N_4576,N_5285);
xnor U6858 (N_6858,N_4131,N_4942);
or U6859 (N_6859,N_4271,N_5819);
and U6860 (N_6860,N_4795,N_4296);
and U6861 (N_6861,N_4329,N_4908);
and U6862 (N_6862,N_5349,N_5419);
and U6863 (N_6863,N_4744,N_5970);
or U6864 (N_6864,N_4469,N_5968);
and U6865 (N_6865,N_5801,N_4567);
nor U6866 (N_6866,N_4205,N_5815);
xnor U6867 (N_6867,N_5818,N_4898);
nand U6868 (N_6868,N_5938,N_5395);
or U6869 (N_6869,N_5326,N_4355);
nand U6870 (N_6870,N_5653,N_4711);
or U6871 (N_6871,N_5748,N_5159);
xnor U6872 (N_6872,N_4071,N_5788);
nand U6873 (N_6873,N_4605,N_5762);
and U6874 (N_6874,N_5397,N_4466);
and U6875 (N_6875,N_5192,N_4219);
nand U6876 (N_6876,N_4660,N_5497);
and U6877 (N_6877,N_4538,N_5188);
xor U6878 (N_6878,N_5844,N_4152);
and U6879 (N_6879,N_4935,N_4457);
nand U6880 (N_6880,N_5142,N_4010);
or U6881 (N_6881,N_4528,N_5125);
nand U6882 (N_6882,N_4450,N_5608);
and U6883 (N_6883,N_4066,N_4663);
nor U6884 (N_6884,N_5365,N_4596);
nand U6885 (N_6885,N_4290,N_5717);
or U6886 (N_6886,N_4983,N_4590);
nor U6887 (N_6887,N_5097,N_5053);
xnor U6888 (N_6888,N_5095,N_4459);
nor U6889 (N_6889,N_4543,N_4591);
nand U6890 (N_6890,N_5786,N_5441);
and U6891 (N_6891,N_5931,N_4857);
and U6892 (N_6892,N_4306,N_4453);
nand U6893 (N_6893,N_4763,N_4020);
nand U6894 (N_6894,N_5373,N_5345);
and U6895 (N_6895,N_5246,N_5927);
nand U6896 (N_6896,N_4366,N_4496);
nor U6897 (N_6897,N_5758,N_4488);
nor U6898 (N_6898,N_5359,N_4918);
and U6899 (N_6899,N_4079,N_4999);
xnor U6900 (N_6900,N_4733,N_4260);
nand U6901 (N_6901,N_5150,N_5993);
nand U6902 (N_6902,N_5842,N_4141);
or U6903 (N_6903,N_4101,N_4956);
and U6904 (N_6904,N_4374,N_4893);
nand U6905 (N_6905,N_5343,N_4232);
nor U6906 (N_6906,N_4339,N_5385);
nor U6907 (N_6907,N_5660,N_4920);
nor U6908 (N_6908,N_4665,N_4376);
and U6909 (N_6909,N_4680,N_4274);
or U6910 (N_6910,N_4742,N_4118);
nand U6911 (N_6911,N_5905,N_4971);
nand U6912 (N_6912,N_5974,N_4291);
nor U6913 (N_6913,N_4704,N_4713);
xnor U6914 (N_6914,N_5128,N_5260);
xnor U6915 (N_6915,N_5323,N_5568);
and U6916 (N_6916,N_5960,N_4002);
and U6917 (N_6917,N_5461,N_5985);
xor U6918 (N_6918,N_5570,N_5264);
nand U6919 (N_6919,N_5231,N_4708);
or U6920 (N_6920,N_4604,N_5614);
nand U6921 (N_6921,N_4984,N_4732);
and U6922 (N_6922,N_4709,N_4417);
nor U6923 (N_6923,N_4149,N_4728);
nand U6924 (N_6924,N_5605,N_4565);
nor U6925 (N_6925,N_4422,N_5903);
nand U6926 (N_6926,N_5321,N_4750);
nand U6927 (N_6927,N_5936,N_4765);
nor U6928 (N_6928,N_5750,N_4934);
nor U6929 (N_6929,N_5506,N_4017);
xnor U6930 (N_6930,N_5475,N_5768);
and U6931 (N_6931,N_5172,N_5808);
nand U6932 (N_6932,N_4881,N_4674);
nor U6933 (N_6933,N_5937,N_4351);
or U6934 (N_6934,N_4154,N_4534);
and U6935 (N_6935,N_4725,N_4059);
and U6936 (N_6936,N_4513,N_4581);
nand U6937 (N_6937,N_5076,N_4318);
nand U6938 (N_6938,N_5194,N_4835);
nor U6939 (N_6939,N_4684,N_4173);
or U6940 (N_6940,N_4562,N_5814);
or U6941 (N_6941,N_4234,N_4429);
nor U6942 (N_6942,N_4437,N_4699);
or U6943 (N_6943,N_4297,N_5456);
nand U6944 (N_6944,N_4662,N_5091);
or U6945 (N_6945,N_5729,N_5476);
nand U6946 (N_6946,N_5972,N_4705);
or U6947 (N_6947,N_5288,N_5620);
and U6948 (N_6948,N_5330,N_4994);
nand U6949 (N_6949,N_4924,N_4443);
nor U6950 (N_6950,N_4397,N_4977);
xor U6951 (N_6951,N_5879,N_4093);
xnor U6952 (N_6952,N_5126,N_4678);
nor U6953 (N_6953,N_4440,N_4529);
or U6954 (N_6954,N_5237,N_4809);
xnor U6955 (N_6955,N_4992,N_5409);
nor U6956 (N_6956,N_5043,N_4187);
or U6957 (N_6957,N_5358,N_5481);
and U6958 (N_6958,N_5557,N_4228);
and U6959 (N_6959,N_5217,N_4191);
and U6960 (N_6960,N_4730,N_5857);
nor U6961 (N_6961,N_4302,N_5496);
nor U6962 (N_6962,N_5309,N_5930);
nor U6963 (N_6963,N_4803,N_4640);
nor U6964 (N_6964,N_5502,N_5826);
nand U6965 (N_6965,N_5861,N_5386);
or U6966 (N_6966,N_4371,N_4493);
and U6967 (N_6967,N_5003,N_4808);
and U6968 (N_6968,N_5290,N_5628);
nand U6969 (N_6969,N_5012,N_4583);
nor U6970 (N_6970,N_4503,N_4301);
xor U6971 (N_6971,N_4454,N_5781);
or U6972 (N_6972,N_5059,N_5789);
nor U6973 (N_6973,N_5056,N_4948);
or U6974 (N_6974,N_4214,N_5712);
or U6975 (N_6975,N_4951,N_5498);
nand U6976 (N_6976,N_5483,N_4337);
nand U6977 (N_6977,N_4416,N_4779);
nor U6978 (N_6978,N_4638,N_4871);
or U6979 (N_6979,N_5847,N_5553);
or U6980 (N_6980,N_5147,N_4514);
nand U6981 (N_6981,N_5716,N_4045);
or U6982 (N_6982,N_4580,N_5512);
nor U6983 (N_6983,N_4349,N_5165);
or U6984 (N_6984,N_4832,N_4420);
nand U6985 (N_6985,N_4273,N_4331);
or U6986 (N_6986,N_4310,N_4975);
nand U6987 (N_6987,N_4112,N_5455);
or U6988 (N_6988,N_4621,N_5592);
nand U6989 (N_6989,N_4390,N_4307);
and U6990 (N_6990,N_5171,N_5440);
xnor U6991 (N_6991,N_4229,N_5745);
nor U6992 (N_6992,N_4642,N_4911);
and U6993 (N_6993,N_5393,N_4783);
or U6994 (N_6994,N_4155,N_4650);
or U6995 (N_6995,N_4953,N_4111);
nand U6996 (N_6996,N_4639,N_5160);
and U6997 (N_6997,N_4233,N_5263);
nand U6998 (N_6998,N_4726,N_5946);
nand U6999 (N_6999,N_4324,N_5682);
and U7000 (N_7000,N_4901,N_5993);
and U7001 (N_7001,N_5967,N_5711);
xor U7002 (N_7002,N_4836,N_5378);
and U7003 (N_7003,N_5403,N_4918);
or U7004 (N_7004,N_5318,N_5596);
xor U7005 (N_7005,N_4830,N_4372);
nand U7006 (N_7006,N_4001,N_4417);
nand U7007 (N_7007,N_5989,N_4949);
xnor U7008 (N_7008,N_5163,N_4435);
and U7009 (N_7009,N_5825,N_5100);
nor U7010 (N_7010,N_5233,N_5494);
or U7011 (N_7011,N_5380,N_5612);
nor U7012 (N_7012,N_4691,N_5366);
and U7013 (N_7013,N_4255,N_4408);
xnor U7014 (N_7014,N_4277,N_4758);
or U7015 (N_7015,N_5233,N_4897);
nor U7016 (N_7016,N_5529,N_4805);
nand U7017 (N_7017,N_5525,N_5602);
or U7018 (N_7018,N_4584,N_5257);
or U7019 (N_7019,N_5377,N_5425);
xor U7020 (N_7020,N_5893,N_4984);
and U7021 (N_7021,N_5804,N_5938);
and U7022 (N_7022,N_5487,N_4072);
or U7023 (N_7023,N_4372,N_4596);
nor U7024 (N_7024,N_5904,N_5610);
nor U7025 (N_7025,N_5208,N_5435);
nand U7026 (N_7026,N_4542,N_5460);
nand U7027 (N_7027,N_5395,N_4811);
nor U7028 (N_7028,N_5519,N_5603);
or U7029 (N_7029,N_5767,N_5922);
nand U7030 (N_7030,N_5847,N_5688);
and U7031 (N_7031,N_4638,N_5277);
or U7032 (N_7032,N_4422,N_5028);
xor U7033 (N_7033,N_4957,N_4300);
and U7034 (N_7034,N_5851,N_4879);
and U7035 (N_7035,N_4860,N_4338);
nor U7036 (N_7036,N_4292,N_4778);
nor U7037 (N_7037,N_4093,N_4890);
and U7038 (N_7038,N_4158,N_4006);
or U7039 (N_7039,N_4332,N_5275);
or U7040 (N_7040,N_5249,N_5978);
nor U7041 (N_7041,N_5980,N_4308);
nand U7042 (N_7042,N_4822,N_5270);
nand U7043 (N_7043,N_4867,N_4132);
xnor U7044 (N_7044,N_5828,N_5039);
nand U7045 (N_7045,N_4536,N_4520);
and U7046 (N_7046,N_5098,N_4432);
nand U7047 (N_7047,N_5828,N_5956);
and U7048 (N_7048,N_5361,N_5209);
or U7049 (N_7049,N_5171,N_5202);
or U7050 (N_7050,N_4036,N_5449);
or U7051 (N_7051,N_4908,N_4884);
nor U7052 (N_7052,N_5155,N_5941);
or U7053 (N_7053,N_4239,N_4608);
nor U7054 (N_7054,N_4020,N_4613);
or U7055 (N_7055,N_4320,N_5108);
or U7056 (N_7056,N_4829,N_5180);
xnor U7057 (N_7057,N_5682,N_4296);
or U7058 (N_7058,N_4786,N_4295);
nor U7059 (N_7059,N_5546,N_4796);
nor U7060 (N_7060,N_4747,N_5735);
or U7061 (N_7061,N_4072,N_4146);
nor U7062 (N_7062,N_4939,N_4207);
nand U7063 (N_7063,N_5873,N_4998);
nor U7064 (N_7064,N_4246,N_5491);
nor U7065 (N_7065,N_4992,N_4578);
nor U7066 (N_7066,N_5914,N_4481);
nor U7067 (N_7067,N_4453,N_5001);
nand U7068 (N_7068,N_4869,N_5437);
or U7069 (N_7069,N_4727,N_4756);
and U7070 (N_7070,N_4742,N_4057);
and U7071 (N_7071,N_5371,N_5868);
nand U7072 (N_7072,N_5940,N_5141);
nand U7073 (N_7073,N_5007,N_4256);
or U7074 (N_7074,N_4081,N_4298);
and U7075 (N_7075,N_5139,N_4332);
or U7076 (N_7076,N_5813,N_5561);
nor U7077 (N_7077,N_5922,N_4360);
nand U7078 (N_7078,N_4670,N_5546);
nor U7079 (N_7079,N_4506,N_4162);
and U7080 (N_7080,N_4394,N_4893);
or U7081 (N_7081,N_4479,N_4735);
nand U7082 (N_7082,N_4991,N_5135);
xor U7083 (N_7083,N_5757,N_5868);
or U7084 (N_7084,N_4692,N_4915);
nand U7085 (N_7085,N_5256,N_4555);
or U7086 (N_7086,N_4860,N_5279);
nand U7087 (N_7087,N_5978,N_5712);
nor U7088 (N_7088,N_5910,N_4355);
or U7089 (N_7089,N_4869,N_5636);
nor U7090 (N_7090,N_4836,N_4800);
nor U7091 (N_7091,N_4368,N_4681);
or U7092 (N_7092,N_4864,N_5304);
or U7093 (N_7093,N_5793,N_5949);
nand U7094 (N_7094,N_4280,N_4742);
nand U7095 (N_7095,N_5189,N_5218);
nand U7096 (N_7096,N_5432,N_4519);
nand U7097 (N_7097,N_4830,N_4508);
nand U7098 (N_7098,N_5420,N_4239);
nor U7099 (N_7099,N_4512,N_5359);
nor U7100 (N_7100,N_5829,N_5069);
nand U7101 (N_7101,N_4884,N_4048);
nand U7102 (N_7102,N_4293,N_4091);
and U7103 (N_7103,N_4285,N_4639);
nand U7104 (N_7104,N_4052,N_4364);
and U7105 (N_7105,N_4569,N_4717);
or U7106 (N_7106,N_4416,N_4777);
and U7107 (N_7107,N_5815,N_5879);
and U7108 (N_7108,N_5133,N_5009);
nand U7109 (N_7109,N_4054,N_4395);
and U7110 (N_7110,N_5157,N_5126);
nand U7111 (N_7111,N_4530,N_4814);
and U7112 (N_7112,N_4440,N_4045);
xnor U7113 (N_7113,N_4704,N_4549);
nor U7114 (N_7114,N_5715,N_5643);
nor U7115 (N_7115,N_5700,N_4269);
nand U7116 (N_7116,N_5511,N_5489);
or U7117 (N_7117,N_5631,N_5010);
nand U7118 (N_7118,N_5188,N_5470);
or U7119 (N_7119,N_4475,N_5239);
and U7120 (N_7120,N_4917,N_4149);
xnor U7121 (N_7121,N_4892,N_5419);
and U7122 (N_7122,N_4186,N_4888);
and U7123 (N_7123,N_5337,N_5403);
and U7124 (N_7124,N_4328,N_4418);
nor U7125 (N_7125,N_4418,N_4937);
nand U7126 (N_7126,N_4519,N_4064);
or U7127 (N_7127,N_5655,N_4382);
and U7128 (N_7128,N_4558,N_5164);
and U7129 (N_7129,N_5932,N_5941);
and U7130 (N_7130,N_5892,N_5038);
or U7131 (N_7131,N_4214,N_4775);
or U7132 (N_7132,N_4364,N_4063);
nor U7133 (N_7133,N_4818,N_5899);
xor U7134 (N_7134,N_4235,N_5145);
nand U7135 (N_7135,N_5109,N_4478);
or U7136 (N_7136,N_5052,N_5529);
or U7137 (N_7137,N_5701,N_4126);
nand U7138 (N_7138,N_4464,N_4522);
or U7139 (N_7139,N_4949,N_4186);
or U7140 (N_7140,N_5910,N_4827);
xor U7141 (N_7141,N_5755,N_4798);
nor U7142 (N_7142,N_5885,N_5382);
nand U7143 (N_7143,N_4350,N_5989);
and U7144 (N_7144,N_5058,N_5702);
nand U7145 (N_7145,N_4127,N_5962);
nor U7146 (N_7146,N_4135,N_5277);
nor U7147 (N_7147,N_5571,N_5418);
nor U7148 (N_7148,N_5638,N_4478);
nor U7149 (N_7149,N_5383,N_5784);
nand U7150 (N_7150,N_4866,N_5159);
and U7151 (N_7151,N_4900,N_5377);
or U7152 (N_7152,N_4122,N_4747);
nand U7153 (N_7153,N_5180,N_5010);
nor U7154 (N_7154,N_5473,N_5016);
or U7155 (N_7155,N_5178,N_4408);
or U7156 (N_7156,N_5696,N_4695);
xor U7157 (N_7157,N_5144,N_5263);
and U7158 (N_7158,N_5591,N_4782);
nand U7159 (N_7159,N_4515,N_4936);
xor U7160 (N_7160,N_4885,N_5449);
nor U7161 (N_7161,N_5172,N_4516);
and U7162 (N_7162,N_4489,N_4396);
nor U7163 (N_7163,N_5411,N_4799);
nor U7164 (N_7164,N_4366,N_4028);
nand U7165 (N_7165,N_5618,N_5266);
xor U7166 (N_7166,N_4739,N_5571);
xor U7167 (N_7167,N_5365,N_5456);
xor U7168 (N_7168,N_5341,N_5838);
nand U7169 (N_7169,N_5105,N_5585);
nand U7170 (N_7170,N_4005,N_4147);
nor U7171 (N_7171,N_5836,N_4338);
nand U7172 (N_7172,N_5977,N_4131);
nor U7173 (N_7173,N_5601,N_5865);
nor U7174 (N_7174,N_4085,N_4665);
nor U7175 (N_7175,N_4238,N_4991);
or U7176 (N_7176,N_4399,N_5237);
nor U7177 (N_7177,N_4595,N_4625);
xnor U7178 (N_7178,N_5754,N_5157);
or U7179 (N_7179,N_5588,N_5322);
or U7180 (N_7180,N_4846,N_4120);
or U7181 (N_7181,N_4031,N_5294);
and U7182 (N_7182,N_5760,N_4950);
nand U7183 (N_7183,N_5671,N_4665);
nor U7184 (N_7184,N_4571,N_4666);
nand U7185 (N_7185,N_4450,N_5664);
nand U7186 (N_7186,N_5347,N_5686);
nor U7187 (N_7187,N_5736,N_4485);
xnor U7188 (N_7188,N_5361,N_5756);
and U7189 (N_7189,N_5006,N_4014);
nor U7190 (N_7190,N_4567,N_5379);
and U7191 (N_7191,N_4729,N_4993);
and U7192 (N_7192,N_4097,N_4349);
xor U7193 (N_7193,N_5478,N_4784);
nor U7194 (N_7194,N_4245,N_4154);
nor U7195 (N_7195,N_5584,N_4988);
nand U7196 (N_7196,N_4925,N_4422);
nor U7197 (N_7197,N_5886,N_4503);
nor U7198 (N_7198,N_4006,N_4226);
and U7199 (N_7199,N_4563,N_4852);
and U7200 (N_7200,N_5522,N_5596);
nand U7201 (N_7201,N_5001,N_5866);
nand U7202 (N_7202,N_5496,N_5332);
or U7203 (N_7203,N_5304,N_4501);
xor U7204 (N_7204,N_5965,N_5273);
or U7205 (N_7205,N_5781,N_4068);
nor U7206 (N_7206,N_5808,N_5747);
or U7207 (N_7207,N_5294,N_4887);
nand U7208 (N_7208,N_4111,N_5676);
xor U7209 (N_7209,N_5410,N_5978);
xnor U7210 (N_7210,N_5541,N_4401);
nand U7211 (N_7211,N_5602,N_4097);
or U7212 (N_7212,N_5622,N_4935);
nor U7213 (N_7213,N_5098,N_4580);
nor U7214 (N_7214,N_5887,N_4366);
nor U7215 (N_7215,N_5096,N_5485);
or U7216 (N_7216,N_4031,N_4140);
and U7217 (N_7217,N_5125,N_4828);
nor U7218 (N_7218,N_4631,N_5075);
nor U7219 (N_7219,N_5234,N_4072);
or U7220 (N_7220,N_5710,N_4164);
and U7221 (N_7221,N_4791,N_5975);
or U7222 (N_7222,N_5574,N_4771);
or U7223 (N_7223,N_5193,N_4634);
and U7224 (N_7224,N_4719,N_4792);
nand U7225 (N_7225,N_5120,N_5040);
nor U7226 (N_7226,N_5710,N_5197);
and U7227 (N_7227,N_5531,N_4518);
and U7228 (N_7228,N_4583,N_4235);
nand U7229 (N_7229,N_5562,N_4352);
nor U7230 (N_7230,N_4542,N_5361);
and U7231 (N_7231,N_5179,N_5700);
xor U7232 (N_7232,N_4760,N_5872);
or U7233 (N_7233,N_4883,N_5147);
nor U7234 (N_7234,N_4776,N_5359);
nor U7235 (N_7235,N_5764,N_5601);
and U7236 (N_7236,N_5024,N_5972);
or U7237 (N_7237,N_4715,N_5935);
or U7238 (N_7238,N_5159,N_4365);
nor U7239 (N_7239,N_4481,N_4963);
nand U7240 (N_7240,N_4700,N_5785);
and U7241 (N_7241,N_4030,N_5873);
nand U7242 (N_7242,N_5600,N_5471);
or U7243 (N_7243,N_4745,N_4766);
or U7244 (N_7244,N_4636,N_4739);
and U7245 (N_7245,N_4238,N_5814);
or U7246 (N_7246,N_4852,N_5571);
or U7247 (N_7247,N_4434,N_5273);
nand U7248 (N_7248,N_5326,N_5565);
and U7249 (N_7249,N_4860,N_4893);
nor U7250 (N_7250,N_4355,N_5366);
nand U7251 (N_7251,N_5038,N_5549);
and U7252 (N_7252,N_4954,N_5207);
or U7253 (N_7253,N_5067,N_4511);
nor U7254 (N_7254,N_5740,N_5715);
nand U7255 (N_7255,N_4962,N_5774);
or U7256 (N_7256,N_4378,N_4858);
nand U7257 (N_7257,N_5746,N_5994);
or U7258 (N_7258,N_4414,N_4374);
or U7259 (N_7259,N_4925,N_4300);
nor U7260 (N_7260,N_4082,N_4411);
nor U7261 (N_7261,N_5751,N_4316);
nand U7262 (N_7262,N_4652,N_4479);
xnor U7263 (N_7263,N_4395,N_5361);
and U7264 (N_7264,N_4215,N_4060);
or U7265 (N_7265,N_5922,N_4379);
or U7266 (N_7266,N_4427,N_5333);
and U7267 (N_7267,N_4727,N_4497);
nand U7268 (N_7268,N_5015,N_5752);
nor U7269 (N_7269,N_4418,N_4267);
nor U7270 (N_7270,N_5645,N_5164);
nand U7271 (N_7271,N_4052,N_4241);
xnor U7272 (N_7272,N_5438,N_5377);
nor U7273 (N_7273,N_5645,N_4283);
nor U7274 (N_7274,N_5107,N_5916);
or U7275 (N_7275,N_5639,N_5628);
nand U7276 (N_7276,N_5026,N_4784);
nor U7277 (N_7277,N_5263,N_5064);
nor U7278 (N_7278,N_5891,N_4949);
or U7279 (N_7279,N_4579,N_5212);
xor U7280 (N_7280,N_4353,N_5386);
nor U7281 (N_7281,N_5999,N_4888);
nand U7282 (N_7282,N_5938,N_4886);
nor U7283 (N_7283,N_5671,N_5864);
nor U7284 (N_7284,N_4733,N_4116);
nor U7285 (N_7285,N_5432,N_5261);
or U7286 (N_7286,N_5722,N_5626);
and U7287 (N_7287,N_5358,N_4659);
nand U7288 (N_7288,N_4068,N_5665);
xnor U7289 (N_7289,N_5838,N_5910);
nor U7290 (N_7290,N_5841,N_5028);
nor U7291 (N_7291,N_5468,N_5614);
and U7292 (N_7292,N_4512,N_4305);
and U7293 (N_7293,N_5664,N_5154);
nor U7294 (N_7294,N_5268,N_5817);
xor U7295 (N_7295,N_4854,N_4775);
nor U7296 (N_7296,N_5038,N_4310);
and U7297 (N_7297,N_4365,N_4918);
or U7298 (N_7298,N_5822,N_5572);
and U7299 (N_7299,N_5310,N_5671);
nor U7300 (N_7300,N_5253,N_4702);
nor U7301 (N_7301,N_4896,N_5740);
and U7302 (N_7302,N_5324,N_4132);
or U7303 (N_7303,N_4839,N_4676);
nor U7304 (N_7304,N_4128,N_5561);
and U7305 (N_7305,N_5483,N_4084);
or U7306 (N_7306,N_4221,N_5138);
nor U7307 (N_7307,N_5400,N_5291);
nor U7308 (N_7308,N_5102,N_5687);
nor U7309 (N_7309,N_4693,N_4673);
and U7310 (N_7310,N_5076,N_4706);
nand U7311 (N_7311,N_4847,N_5638);
xor U7312 (N_7312,N_4982,N_4813);
nor U7313 (N_7313,N_4799,N_5244);
nor U7314 (N_7314,N_5004,N_5099);
or U7315 (N_7315,N_5721,N_4985);
nand U7316 (N_7316,N_5717,N_4070);
nor U7317 (N_7317,N_5627,N_4338);
nand U7318 (N_7318,N_4993,N_4890);
nand U7319 (N_7319,N_4779,N_5596);
and U7320 (N_7320,N_4885,N_5081);
or U7321 (N_7321,N_4614,N_5627);
or U7322 (N_7322,N_5437,N_4398);
nand U7323 (N_7323,N_5187,N_5172);
and U7324 (N_7324,N_4651,N_5896);
nor U7325 (N_7325,N_5016,N_4829);
nand U7326 (N_7326,N_5358,N_4200);
and U7327 (N_7327,N_4681,N_5048);
nand U7328 (N_7328,N_5837,N_4569);
nor U7329 (N_7329,N_4991,N_5700);
or U7330 (N_7330,N_4259,N_4230);
nand U7331 (N_7331,N_4903,N_5411);
nand U7332 (N_7332,N_4447,N_4448);
nand U7333 (N_7333,N_5883,N_5140);
nor U7334 (N_7334,N_5621,N_5394);
xor U7335 (N_7335,N_5481,N_5642);
nand U7336 (N_7336,N_4951,N_4936);
nor U7337 (N_7337,N_5612,N_4977);
and U7338 (N_7338,N_4576,N_4282);
and U7339 (N_7339,N_5118,N_4529);
and U7340 (N_7340,N_4785,N_5575);
or U7341 (N_7341,N_5229,N_4893);
and U7342 (N_7342,N_4644,N_4591);
nor U7343 (N_7343,N_5801,N_5855);
nand U7344 (N_7344,N_5308,N_5707);
nor U7345 (N_7345,N_5402,N_5882);
or U7346 (N_7346,N_4043,N_4073);
nand U7347 (N_7347,N_5368,N_4110);
nor U7348 (N_7348,N_5966,N_4917);
nor U7349 (N_7349,N_4159,N_4294);
nand U7350 (N_7350,N_4989,N_4506);
and U7351 (N_7351,N_5538,N_4579);
or U7352 (N_7352,N_5640,N_4653);
nand U7353 (N_7353,N_5091,N_4575);
and U7354 (N_7354,N_4850,N_5429);
or U7355 (N_7355,N_5150,N_4133);
nand U7356 (N_7356,N_4118,N_5492);
or U7357 (N_7357,N_4764,N_4091);
or U7358 (N_7358,N_4166,N_5961);
nand U7359 (N_7359,N_5009,N_5912);
xor U7360 (N_7360,N_4585,N_4839);
or U7361 (N_7361,N_5413,N_4844);
nand U7362 (N_7362,N_5361,N_4617);
nand U7363 (N_7363,N_4492,N_4575);
nor U7364 (N_7364,N_4489,N_5889);
or U7365 (N_7365,N_5461,N_4295);
and U7366 (N_7366,N_4576,N_5752);
and U7367 (N_7367,N_4234,N_4277);
nand U7368 (N_7368,N_4682,N_5382);
xnor U7369 (N_7369,N_5129,N_4801);
nand U7370 (N_7370,N_4604,N_5124);
nand U7371 (N_7371,N_5476,N_5726);
nor U7372 (N_7372,N_4861,N_5822);
xnor U7373 (N_7373,N_4793,N_5110);
and U7374 (N_7374,N_4602,N_5930);
xor U7375 (N_7375,N_5891,N_5982);
or U7376 (N_7376,N_5025,N_4188);
and U7377 (N_7377,N_4305,N_5407);
or U7378 (N_7378,N_5518,N_4754);
nor U7379 (N_7379,N_5905,N_5201);
nor U7380 (N_7380,N_5523,N_4391);
or U7381 (N_7381,N_5419,N_5782);
nand U7382 (N_7382,N_5842,N_5295);
or U7383 (N_7383,N_5160,N_4615);
or U7384 (N_7384,N_5479,N_5413);
nand U7385 (N_7385,N_4008,N_4372);
nand U7386 (N_7386,N_4833,N_4831);
nor U7387 (N_7387,N_4540,N_5376);
nand U7388 (N_7388,N_5213,N_5146);
xnor U7389 (N_7389,N_5752,N_5184);
and U7390 (N_7390,N_5134,N_4092);
or U7391 (N_7391,N_4682,N_4093);
nand U7392 (N_7392,N_5947,N_5910);
nor U7393 (N_7393,N_5596,N_4823);
or U7394 (N_7394,N_5391,N_5821);
nor U7395 (N_7395,N_4130,N_4522);
and U7396 (N_7396,N_5081,N_4449);
or U7397 (N_7397,N_4639,N_5353);
nand U7398 (N_7398,N_5211,N_5787);
nand U7399 (N_7399,N_4776,N_5463);
and U7400 (N_7400,N_4413,N_4200);
or U7401 (N_7401,N_4110,N_4581);
and U7402 (N_7402,N_5497,N_5965);
and U7403 (N_7403,N_4088,N_4069);
or U7404 (N_7404,N_5362,N_4295);
or U7405 (N_7405,N_5332,N_5221);
and U7406 (N_7406,N_5127,N_5842);
and U7407 (N_7407,N_4541,N_4074);
nand U7408 (N_7408,N_5054,N_5794);
nor U7409 (N_7409,N_5010,N_4007);
nand U7410 (N_7410,N_5708,N_4387);
and U7411 (N_7411,N_4666,N_5089);
or U7412 (N_7412,N_4780,N_5179);
nand U7413 (N_7413,N_4301,N_4405);
nand U7414 (N_7414,N_5773,N_4443);
or U7415 (N_7415,N_5694,N_5486);
and U7416 (N_7416,N_5959,N_4940);
nand U7417 (N_7417,N_4381,N_5629);
nand U7418 (N_7418,N_5432,N_5894);
nand U7419 (N_7419,N_5353,N_4888);
and U7420 (N_7420,N_4979,N_4556);
nand U7421 (N_7421,N_4731,N_4643);
nor U7422 (N_7422,N_4980,N_4589);
xor U7423 (N_7423,N_4344,N_5728);
and U7424 (N_7424,N_4441,N_5122);
or U7425 (N_7425,N_4368,N_4444);
and U7426 (N_7426,N_5247,N_4827);
and U7427 (N_7427,N_4619,N_4053);
nor U7428 (N_7428,N_4971,N_4441);
nor U7429 (N_7429,N_5319,N_4374);
or U7430 (N_7430,N_4077,N_5205);
xnor U7431 (N_7431,N_5426,N_5956);
xor U7432 (N_7432,N_4496,N_4049);
or U7433 (N_7433,N_5134,N_5586);
and U7434 (N_7434,N_5632,N_5532);
nand U7435 (N_7435,N_5766,N_4673);
nand U7436 (N_7436,N_5617,N_4570);
or U7437 (N_7437,N_5803,N_4404);
or U7438 (N_7438,N_4835,N_5953);
nor U7439 (N_7439,N_5873,N_4202);
and U7440 (N_7440,N_5103,N_5636);
xnor U7441 (N_7441,N_5158,N_4647);
and U7442 (N_7442,N_4131,N_5911);
and U7443 (N_7443,N_5830,N_4335);
nand U7444 (N_7444,N_5673,N_4153);
and U7445 (N_7445,N_4288,N_4889);
nand U7446 (N_7446,N_5589,N_5179);
nor U7447 (N_7447,N_5758,N_4514);
nor U7448 (N_7448,N_4898,N_4219);
or U7449 (N_7449,N_4983,N_4366);
nand U7450 (N_7450,N_4621,N_4054);
xor U7451 (N_7451,N_5473,N_4646);
nor U7452 (N_7452,N_5197,N_5191);
nor U7453 (N_7453,N_5427,N_5663);
nor U7454 (N_7454,N_4160,N_4026);
nor U7455 (N_7455,N_4465,N_4942);
or U7456 (N_7456,N_5037,N_4683);
or U7457 (N_7457,N_5408,N_4389);
or U7458 (N_7458,N_5194,N_4647);
or U7459 (N_7459,N_5230,N_5153);
nand U7460 (N_7460,N_4567,N_5629);
and U7461 (N_7461,N_5028,N_5165);
or U7462 (N_7462,N_5767,N_4143);
nand U7463 (N_7463,N_5519,N_5799);
or U7464 (N_7464,N_4716,N_5473);
nand U7465 (N_7465,N_5711,N_5832);
or U7466 (N_7466,N_4465,N_4542);
nand U7467 (N_7467,N_5161,N_5419);
and U7468 (N_7468,N_5486,N_5221);
nand U7469 (N_7469,N_4240,N_4516);
nor U7470 (N_7470,N_4331,N_5312);
nor U7471 (N_7471,N_4085,N_5626);
and U7472 (N_7472,N_5110,N_4653);
or U7473 (N_7473,N_5039,N_4275);
xnor U7474 (N_7474,N_4791,N_5722);
nor U7475 (N_7475,N_5118,N_5159);
xnor U7476 (N_7476,N_5326,N_5622);
nor U7477 (N_7477,N_4654,N_5443);
xor U7478 (N_7478,N_4887,N_4366);
or U7479 (N_7479,N_5386,N_4536);
nor U7480 (N_7480,N_4071,N_5631);
nor U7481 (N_7481,N_4513,N_4228);
and U7482 (N_7482,N_4020,N_5033);
nand U7483 (N_7483,N_4882,N_4000);
or U7484 (N_7484,N_4981,N_4896);
or U7485 (N_7485,N_5425,N_4829);
and U7486 (N_7486,N_4768,N_5586);
nor U7487 (N_7487,N_5293,N_4395);
nand U7488 (N_7488,N_4885,N_5090);
or U7489 (N_7489,N_4812,N_4363);
nor U7490 (N_7490,N_5958,N_4402);
or U7491 (N_7491,N_5009,N_4660);
and U7492 (N_7492,N_5231,N_4123);
or U7493 (N_7493,N_4207,N_4598);
nor U7494 (N_7494,N_5294,N_5366);
or U7495 (N_7495,N_5823,N_5000);
nor U7496 (N_7496,N_4305,N_5554);
nor U7497 (N_7497,N_4363,N_5230);
nand U7498 (N_7498,N_4095,N_5334);
nand U7499 (N_7499,N_5263,N_5886);
nand U7500 (N_7500,N_4360,N_5219);
nor U7501 (N_7501,N_4913,N_4760);
and U7502 (N_7502,N_4367,N_4218);
and U7503 (N_7503,N_5223,N_4007);
nor U7504 (N_7504,N_4333,N_5684);
or U7505 (N_7505,N_4886,N_5073);
nor U7506 (N_7506,N_4487,N_4746);
and U7507 (N_7507,N_4655,N_4620);
or U7508 (N_7508,N_5397,N_5894);
or U7509 (N_7509,N_4496,N_5750);
or U7510 (N_7510,N_4198,N_4738);
or U7511 (N_7511,N_4375,N_4327);
nand U7512 (N_7512,N_5478,N_5727);
and U7513 (N_7513,N_5948,N_5412);
or U7514 (N_7514,N_4973,N_5805);
or U7515 (N_7515,N_4771,N_5735);
nand U7516 (N_7516,N_5284,N_5441);
nor U7517 (N_7517,N_5212,N_5994);
and U7518 (N_7518,N_4452,N_4793);
nand U7519 (N_7519,N_4308,N_5999);
and U7520 (N_7520,N_4449,N_4166);
nor U7521 (N_7521,N_5620,N_4614);
and U7522 (N_7522,N_5399,N_4434);
nand U7523 (N_7523,N_4360,N_5491);
nand U7524 (N_7524,N_4887,N_5714);
nor U7525 (N_7525,N_5900,N_4378);
or U7526 (N_7526,N_4223,N_4905);
or U7527 (N_7527,N_5711,N_5942);
nand U7528 (N_7528,N_4966,N_4180);
nand U7529 (N_7529,N_5926,N_5678);
nor U7530 (N_7530,N_4883,N_5237);
nor U7531 (N_7531,N_4078,N_4369);
or U7532 (N_7532,N_4490,N_4954);
xnor U7533 (N_7533,N_5224,N_4029);
or U7534 (N_7534,N_4257,N_5712);
nand U7535 (N_7535,N_4809,N_4892);
and U7536 (N_7536,N_4198,N_4617);
nand U7537 (N_7537,N_5718,N_5287);
nor U7538 (N_7538,N_4551,N_5218);
and U7539 (N_7539,N_5306,N_4365);
nor U7540 (N_7540,N_4444,N_4950);
or U7541 (N_7541,N_5099,N_4105);
nor U7542 (N_7542,N_5348,N_5795);
nor U7543 (N_7543,N_4446,N_5270);
and U7544 (N_7544,N_5583,N_4336);
nor U7545 (N_7545,N_4154,N_4617);
nand U7546 (N_7546,N_4233,N_4213);
or U7547 (N_7547,N_4736,N_4140);
and U7548 (N_7548,N_5551,N_4336);
nand U7549 (N_7549,N_5740,N_5601);
and U7550 (N_7550,N_5632,N_4734);
nor U7551 (N_7551,N_5415,N_5767);
xnor U7552 (N_7552,N_5142,N_5533);
xor U7553 (N_7553,N_5306,N_5998);
xor U7554 (N_7554,N_5808,N_5730);
and U7555 (N_7555,N_4193,N_4400);
and U7556 (N_7556,N_4709,N_5470);
nor U7557 (N_7557,N_5774,N_4435);
and U7558 (N_7558,N_4885,N_5091);
nand U7559 (N_7559,N_5872,N_5948);
or U7560 (N_7560,N_4077,N_5781);
nor U7561 (N_7561,N_4671,N_4167);
nand U7562 (N_7562,N_5750,N_4830);
or U7563 (N_7563,N_5684,N_5303);
nor U7564 (N_7564,N_5557,N_5690);
or U7565 (N_7565,N_4626,N_5364);
nand U7566 (N_7566,N_5601,N_5610);
or U7567 (N_7567,N_5065,N_5957);
nand U7568 (N_7568,N_4207,N_5293);
nand U7569 (N_7569,N_4499,N_4265);
and U7570 (N_7570,N_5187,N_4121);
xor U7571 (N_7571,N_4275,N_5572);
nand U7572 (N_7572,N_4436,N_5981);
or U7573 (N_7573,N_4907,N_5790);
or U7574 (N_7574,N_4198,N_5218);
and U7575 (N_7575,N_4789,N_5480);
nand U7576 (N_7576,N_5347,N_5301);
nand U7577 (N_7577,N_5868,N_5608);
nand U7578 (N_7578,N_4023,N_5335);
or U7579 (N_7579,N_4952,N_5367);
nand U7580 (N_7580,N_5511,N_4166);
nor U7581 (N_7581,N_5765,N_4100);
nor U7582 (N_7582,N_4745,N_5038);
nor U7583 (N_7583,N_4064,N_4803);
or U7584 (N_7584,N_5786,N_4253);
or U7585 (N_7585,N_4957,N_5086);
nor U7586 (N_7586,N_5829,N_4525);
nand U7587 (N_7587,N_4954,N_5661);
nor U7588 (N_7588,N_4541,N_4960);
and U7589 (N_7589,N_5330,N_5703);
nor U7590 (N_7590,N_4094,N_5112);
and U7591 (N_7591,N_4815,N_4737);
nor U7592 (N_7592,N_4119,N_4508);
nor U7593 (N_7593,N_5586,N_5608);
xor U7594 (N_7594,N_4837,N_5572);
or U7595 (N_7595,N_4606,N_5274);
nor U7596 (N_7596,N_4815,N_4357);
nand U7597 (N_7597,N_4684,N_4796);
nor U7598 (N_7598,N_4390,N_5258);
nand U7599 (N_7599,N_5018,N_5486);
nand U7600 (N_7600,N_5999,N_4780);
nand U7601 (N_7601,N_5195,N_5510);
nor U7602 (N_7602,N_4799,N_5634);
nor U7603 (N_7603,N_4366,N_5021);
nand U7604 (N_7604,N_5337,N_5023);
nand U7605 (N_7605,N_4280,N_5691);
nor U7606 (N_7606,N_4538,N_4836);
nand U7607 (N_7607,N_5479,N_4454);
or U7608 (N_7608,N_4109,N_5198);
nor U7609 (N_7609,N_5888,N_4505);
xnor U7610 (N_7610,N_4533,N_4415);
nor U7611 (N_7611,N_4508,N_5294);
nand U7612 (N_7612,N_4737,N_5448);
nor U7613 (N_7613,N_4212,N_4582);
and U7614 (N_7614,N_4142,N_4994);
nand U7615 (N_7615,N_4521,N_5459);
or U7616 (N_7616,N_4900,N_4313);
or U7617 (N_7617,N_4934,N_4214);
nor U7618 (N_7618,N_4835,N_4296);
nor U7619 (N_7619,N_5702,N_5383);
or U7620 (N_7620,N_5443,N_5791);
nor U7621 (N_7621,N_4640,N_4556);
and U7622 (N_7622,N_5790,N_4199);
nor U7623 (N_7623,N_4100,N_4663);
and U7624 (N_7624,N_4189,N_5799);
nor U7625 (N_7625,N_5210,N_5572);
nor U7626 (N_7626,N_5809,N_5641);
nand U7627 (N_7627,N_4340,N_5933);
nand U7628 (N_7628,N_4421,N_5877);
and U7629 (N_7629,N_4648,N_5150);
and U7630 (N_7630,N_5598,N_5531);
xor U7631 (N_7631,N_4049,N_4846);
or U7632 (N_7632,N_5361,N_5088);
or U7633 (N_7633,N_4446,N_5178);
or U7634 (N_7634,N_4809,N_5758);
nand U7635 (N_7635,N_5062,N_5107);
nor U7636 (N_7636,N_5409,N_4798);
nand U7637 (N_7637,N_4506,N_4414);
nand U7638 (N_7638,N_4236,N_4434);
nor U7639 (N_7639,N_4610,N_5787);
nand U7640 (N_7640,N_4548,N_4198);
nand U7641 (N_7641,N_5256,N_4667);
nand U7642 (N_7642,N_4545,N_4996);
and U7643 (N_7643,N_4307,N_4306);
xnor U7644 (N_7644,N_4772,N_5264);
or U7645 (N_7645,N_5961,N_5974);
nor U7646 (N_7646,N_5610,N_5367);
or U7647 (N_7647,N_4977,N_4439);
nand U7648 (N_7648,N_4973,N_4449);
nor U7649 (N_7649,N_4903,N_4021);
nand U7650 (N_7650,N_4266,N_5712);
and U7651 (N_7651,N_4520,N_4310);
nand U7652 (N_7652,N_4910,N_5322);
nor U7653 (N_7653,N_4253,N_4924);
and U7654 (N_7654,N_5230,N_4234);
nor U7655 (N_7655,N_4715,N_5448);
and U7656 (N_7656,N_5869,N_5569);
xor U7657 (N_7657,N_4880,N_5428);
nand U7658 (N_7658,N_5425,N_4106);
or U7659 (N_7659,N_5147,N_5803);
and U7660 (N_7660,N_5493,N_5621);
nand U7661 (N_7661,N_5562,N_4488);
nand U7662 (N_7662,N_4477,N_5849);
and U7663 (N_7663,N_4376,N_5436);
or U7664 (N_7664,N_5370,N_4192);
or U7665 (N_7665,N_4385,N_5437);
nor U7666 (N_7666,N_4238,N_5347);
and U7667 (N_7667,N_4182,N_4264);
and U7668 (N_7668,N_4099,N_5028);
or U7669 (N_7669,N_5111,N_5793);
nor U7670 (N_7670,N_4746,N_5001);
nand U7671 (N_7671,N_5928,N_4741);
nor U7672 (N_7672,N_4467,N_5107);
and U7673 (N_7673,N_5457,N_5663);
nand U7674 (N_7674,N_4252,N_4599);
nor U7675 (N_7675,N_5572,N_5330);
or U7676 (N_7676,N_4444,N_5253);
or U7677 (N_7677,N_5200,N_4000);
nand U7678 (N_7678,N_5129,N_5906);
and U7679 (N_7679,N_5093,N_5283);
nor U7680 (N_7680,N_4307,N_4581);
or U7681 (N_7681,N_5419,N_5008);
or U7682 (N_7682,N_5096,N_5981);
and U7683 (N_7683,N_5819,N_4487);
xor U7684 (N_7684,N_5846,N_5016);
and U7685 (N_7685,N_5228,N_5193);
and U7686 (N_7686,N_5518,N_4620);
and U7687 (N_7687,N_4850,N_5401);
or U7688 (N_7688,N_4731,N_5395);
and U7689 (N_7689,N_5202,N_5144);
nand U7690 (N_7690,N_4429,N_4036);
and U7691 (N_7691,N_4352,N_5999);
or U7692 (N_7692,N_4102,N_4654);
nand U7693 (N_7693,N_4579,N_5421);
xor U7694 (N_7694,N_5158,N_4421);
or U7695 (N_7695,N_5548,N_4859);
or U7696 (N_7696,N_4817,N_4315);
and U7697 (N_7697,N_5072,N_4800);
or U7698 (N_7698,N_4239,N_5708);
or U7699 (N_7699,N_5455,N_5050);
and U7700 (N_7700,N_5543,N_4218);
or U7701 (N_7701,N_5845,N_4732);
and U7702 (N_7702,N_5990,N_5243);
nand U7703 (N_7703,N_4174,N_5390);
nor U7704 (N_7704,N_5561,N_4274);
xor U7705 (N_7705,N_4731,N_5669);
or U7706 (N_7706,N_5873,N_4846);
nor U7707 (N_7707,N_4206,N_5287);
nor U7708 (N_7708,N_5987,N_4963);
nor U7709 (N_7709,N_5176,N_4380);
or U7710 (N_7710,N_4264,N_5204);
xor U7711 (N_7711,N_5888,N_5452);
xor U7712 (N_7712,N_4851,N_5293);
and U7713 (N_7713,N_5263,N_4832);
nor U7714 (N_7714,N_4128,N_4248);
nand U7715 (N_7715,N_5593,N_5316);
nor U7716 (N_7716,N_5060,N_5048);
and U7717 (N_7717,N_5760,N_4785);
or U7718 (N_7718,N_4804,N_4208);
nor U7719 (N_7719,N_5185,N_5021);
or U7720 (N_7720,N_4585,N_5756);
xor U7721 (N_7721,N_5749,N_4802);
nand U7722 (N_7722,N_5027,N_4123);
nand U7723 (N_7723,N_4892,N_4044);
nor U7724 (N_7724,N_4656,N_5416);
nand U7725 (N_7725,N_4601,N_4792);
nand U7726 (N_7726,N_5007,N_5552);
nor U7727 (N_7727,N_4159,N_4362);
nand U7728 (N_7728,N_4437,N_4776);
or U7729 (N_7729,N_4862,N_4800);
nor U7730 (N_7730,N_4538,N_4989);
nand U7731 (N_7731,N_5288,N_4735);
nand U7732 (N_7732,N_4629,N_4861);
and U7733 (N_7733,N_4266,N_4719);
nor U7734 (N_7734,N_4044,N_4159);
or U7735 (N_7735,N_4125,N_5720);
xnor U7736 (N_7736,N_5421,N_5216);
nor U7737 (N_7737,N_5018,N_5825);
and U7738 (N_7738,N_4786,N_4085);
and U7739 (N_7739,N_5009,N_4627);
nand U7740 (N_7740,N_4778,N_5159);
nor U7741 (N_7741,N_4112,N_4901);
or U7742 (N_7742,N_5336,N_5495);
or U7743 (N_7743,N_4061,N_5315);
and U7744 (N_7744,N_5385,N_4515);
and U7745 (N_7745,N_4853,N_5655);
nor U7746 (N_7746,N_5174,N_5766);
and U7747 (N_7747,N_4290,N_4928);
xor U7748 (N_7748,N_4240,N_5000);
xor U7749 (N_7749,N_5671,N_5687);
nand U7750 (N_7750,N_4819,N_4451);
nand U7751 (N_7751,N_5091,N_4543);
or U7752 (N_7752,N_4933,N_5324);
or U7753 (N_7753,N_5693,N_4535);
or U7754 (N_7754,N_5464,N_4339);
nor U7755 (N_7755,N_5656,N_4383);
xnor U7756 (N_7756,N_5164,N_5139);
and U7757 (N_7757,N_4775,N_5027);
and U7758 (N_7758,N_4487,N_4669);
nor U7759 (N_7759,N_5422,N_4034);
xor U7760 (N_7760,N_4873,N_4178);
or U7761 (N_7761,N_5242,N_4728);
and U7762 (N_7762,N_4748,N_5086);
or U7763 (N_7763,N_4700,N_4722);
nand U7764 (N_7764,N_5979,N_4901);
nand U7765 (N_7765,N_5883,N_5078);
nor U7766 (N_7766,N_5748,N_5415);
nor U7767 (N_7767,N_5629,N_4866);
and U7768 (N_7768,N_5964,N_5795);
or U7769 (N_7769,N_4655,N_4596);
nand U7770 (N_7770,N_4424,N_4078);
nand U7771 (N_7771,N_4282,N_5241);
nor U7772 (N_7772,N_4409,N_5556);
nand U7773 (N_7773,N_5922,N_5707);
xnor U7774 (N_7774,N_4210,N_5361);
nand U7775 (N_7775,N_5999,N_5088);
nor U7776 (N_7776,N_5047,N_5081);
or U7777 (N_7777,N_5915,N_4644);
and U7778 (N_7778,N_5768,N_5307);
and U7779 (N_7779,N_5764,N_5615);
xnor U7780 (N_7780,N_4269,N_5471);
nor U7781 (N_7781,N_5102,N_4686);
and U7782 (N_7782,N_4475,N_4073);
nand U7783 (N_7783,N_4613,N_4152);
or U7784 (N_7784,N_4404,N_5150);
and U7785 (N_7785,N_5606,N_5854);
nand U7786 (N_7786,N_4674,N_4299);
nor U7787 (N_7787,N_4188,N_4416);
or U7788 (N_7788,N_5585,N_5717);
and U7789 (N_7789,N_5114,N_4627);
nand U7790 (N_7790,N_4271,N_5570);
xor U7791 (N_7791,N_4086,N_4964);
nand U7792 (N_7792,N_5651,N_4697);
nand U7793 (N_7793,N_4764,N_5349);
nor U7794 (N_7794,N_5734,N_5789);
nor U7795 (N_7795,N_5339,N_5874);
or U7796 (N_7796,N_4956,N_4915);
or U7797 (N_7797,N_5004,N_4932);
or U7798 (N_7798,N_4524,N_5018);
nor U7799 (N_7799,N_4276,N_5456);
and U7800 (N_7800,N_4111,N_5025);
and U7801 (N_7801,N_5853,N_5597);
or U7802 (N_7802,N_4437,N_4375);
or U7803 (N_7803,N_5893,N_4105);
nor U7804 (N_7804,N_5559,N_5939);
or U7805 (N_7805,N_4248,N_4018);
or U7806 (N_7806,N_4858,N_4744);
nand U7807 (N_7807,N_4736,N_4666);
nor U7808 (N_7808,N_5008,N_4596);
and U7809 (N_7809,N_4448,N_4533);
nand U7810 (N_7810,N_4955,N_5211);
and U7811 (N_7811,N_4909,N_5722);
nor U7812 (N_7812,N_5133,N_4730);
or U7813 (N_7813,N_5794,N_4309);
and U7814 (N_7814,N_5042,N_5175);
and U7815 (N_7815,N_5059,N_5495);
and U7816 (N_7816,N_5927,N_5333);
nand U7817 (N_7817,N_4765,N_5889);
and U7818 (N_7818,N_5602,N_5083);
or U7819 (N_7819,N_4658,N_5823);
nor U7820 (N_7820,N_5020,N_5056);
nand U7821 (N_7821,N_4181,N_4165);
and U7822 (N_7822,N_5907,N_4544);
and U7823 (N_7823,N_5296,N_4098);
and U7824 (N_7824,N_5013,N_5198);
or U7825 (N_7825,N_4148,N_5040);
or U7826 (N_7826,N_4940,N_5527);
and U7827 (N_7827,N_4102,N_5368);
nand U7828 (N_7828,N_4079,N_4703);
nand U7829 (N_7829,N_5873,N_4391);
and U7830 (N_7830,N_4891,N_5976);
nand U7831 (N_7831,N_5278,N_5693);
xor U7832 (N_7832,N_5843,N_4719);
and U7833 (N_7833,N_5750,N_5203);
nor U7834 (N_7834,N_5127,N_5625);
and U7835 (N_7835,N_4074,N_5260);
nand U7836 (N_7836,N_5379,N_4443);
nand U7837 (N_7837,N_4089,N_4684);
xnor U7838 (N_7838,N_4063,N_5875);
nand U7839 (N_7839,N_4622,N_4920);
nand U7840 (N_7840,N_5005,N_4445);
nor U7841 (N_7841,N_4847,N_5998);
nor U7842 (N_7842,N_5101,N_4409);
and U7843 (N_7843,N_5749,N_5153);
nand U7844 (N_7844,N_4960,N_4804);
or U7845 (N_7845,N_4400,N_5240);
and U7846 (N_7846,N_5503,N_5088);
or U7847 (N_7847,N_4844,N_4738);
and U7848 (N_7848,N_4068,N_4951);
nand U7849 (N_7849,N_4899,N_4539);
nand U7850 (N_7850,N_5733,N_5894);
nor U7851 (N_7851,N_4582,N_5495);
nor U7852 (N_7852,N_5565,N_4073);
and U7853 (N_7853,N_5497,N_5479);
or U7854 (N_7854,N_4582,N_5764);
or U7855 (N_7855,N_4612,N_4945);
and U7856 (N_7856,N_5730,N_4083);
or U7857 (N_7857,N_5864,N_5255);
or U7858 (N_7858,N_4709,N_5683);
nor U7859 (N_7859,N_5209,N_5227);
nor U7860 (N_7860,N_5272,N_4259);
nand U7861 (N_7861,N_5696,N_5876);
nand U7862 (N_7862,N_4783,N_5726);
and U7863 (N_7863,N_4596,N_4832);
and U7864 (N_7864,N_5928,N_4963);
and U7865 (N_7865,N_5531,N_5932);
and U7866 (N_7866,N_4455,N_5924);
and U7867 (N_7867,N_4803,N_5862);
nand U7868 (N_7868,N_4519,N_5548);
nor U7869 (N_7869,N_4470,N_4808);
nor U7870 (N_7870,N_4099,N_4598);
xor U7871 (N_7871,N_4079,N_5257);
nor U7872 (N_7872,N_5171,N_5242);
nor U7873 (N_7873,N_5529,N_5275);
or U7874 (N_7874,N_5514,N_5072);
xnor U7875 (N_7875,N_5068,N_4074);
nor U7876 (N_7876,N_4925,N_4032);
and U7877 (N_7877,N_4190,N_4660);
or U7878 (N_7878,N_5199,N_4263);
nor U7879 (N_7879,N_4842,N_4835);
nor U7880 (N_7880,N_4158,N_4760);
and U7881 (N_7881,N_5255,N_4812);
nand U7882 (N_7882,N_4044,N_5603);
and U7883 (N_7883,N_5023,N_5145);
nand U7884 (N_7884,N_4399,N_4029);
nand U7885 (N_7885,N_5640,N_4085);
or U7886 (N_7886,N_5024,N_5887);
nand U7887 (N_7887,N_5455,N_5988);
nand U7888 (N_7888,N_4929,N_4154);
or U7889 (N_7889,N_5263,N_5468);
nor U7890 (N_7890,N_5688,N_4307);
or U7891 (N_7891,N_5997,N_5722);
nand U7892 (N_7892,N_4082,N_4862);
xor U7893 (N_7893,N_5444,N_4848);
nand U7894 (N_7894,N_4621,N_5411);
nor U7895 (N_7895,N_5618,N_5151);
or U7896 (N_7896,N_4915,N_5606);
or U7897 (N_7897,N_4133,N_4063);
and U7898 (N_7898,N_5951,N_4900);
and U7899 (N_7899,N_4052,N_4377);
xor U7900 (N_7900,N_4572,N_4611);
nand U7901 (N_7901,N_4377,N_4963);
or U7902 (N_7902,N_4636,N_4344);
or U7903 (N_7903,N_4221,N_5024);
and U7904 (N_7904,N_5285,N_5133);
and U7905 (N_7905,N_4101,N_5106);
or U7906 (N_7906,N_5508,N_5397);
nand U7907 (N_7907,N_5564,N_5126);
and U7908 (N_7908,N_5767,N_5230);
xor U7909 (N_7909,N_5937,N_5578);
and U7910 (N_7910,N_4812,N_5878);
or U7911 (N_7911,N_5021,N_5031);
or U7912 (N_7912,N_4562,N_4032);
nand U7913 (N_7913,N_5342,N_4469);
or U7914 (N_7914,N_4104,N_4694);
nand U7915 (N_7915,N_5286,N_5356);
nor U7916 (N_7916,N_4011,N_5991);
and U7917 (N_7917,N_4098,N_5394);
and U7918 (N_7918,N_5743,N_5923);
nor U7919 (N_7919,N_5288,N_5964);
and U7920 (N_7920,N_4445,N_4201);
or U7921 (N_7921,N_5178,N_5402);
and U7922 (N_7922,N_5795,N_4809);
and U7923 (N_7923,N_5491,N_4870);
and U7924 (N_7924,N_4943,N_4085);
nand U7925 (N_7925,N_5206,N_5463);
nor U7926 (N_7926,N_5599,N_4030);
nor U7927 (N_7927,N_5398,N_4802);
or U7928 (N_7928,N_4820,N_4378);
and U7929 (N_7929,N_5001,N_4065);
nor U7930 (N_7930,N_4075,N_4001);
or U7931 (N_7931,N_5911,N_5421);
or U7932 (N_7932,N_4795,N_5986);
nand U7933 (N_7933,N_4228,N_4250);
nor U7934 (N_7934,N_4740,N_5056);
nand U7935 (N_7935,N_4939,N_4032);
or U7936 (N_7936,N_4676,N_5556);
nand U7937 (N_7937,N_4229,N_4266);
nand U7938 (N_7938,N_5226,N_5957);
and U7939 (N_7939,N_4052,N_5819);
and U7940 (N_7940,N_5753,N_5447);
nand U7941 (N_7941,N_5361,N_5422);
and U7942 (N_7942,N_4010,N_4409);
or U7943 (N_7943,N_5932,N_4525);
nand U7944 (N_7944,N_4555,N_5044);
nand U7945 (N_7945,N_5980,N_5261);
and U7946 (N_7946,N_5652,N_4665);
nor U7947 (N_7947,N_4951,N_5469);
nand U7948 (N_7948,N_4696,N_5588);
nand U7949 (N_7949,N_5516,N_5846);
nor U7950 (N_7950,N_4747,N_4380);
or U7951 (N_7951,N_4892,N_5146);
nand U7952 (N_7952,N_4732,N_5273);
and U7953 (N_7953,N_4193,N_5315);
nor U7954 (N_7954,N_4388,N_4547);
nand U7955 (N_7955,N_5412,N_5913);
or U7956 (N_7956,N_5614,N_4358);
or U7957 (N_7957,N_4421,N_4495);
and U7958 (N_7958,N_4797,N_5815);
nand U7959 (N_7959,N_4462,N_4762);
and U7960 (N_7960,N_4785,N_4704);
or U7961 (N_7961,N_4983,N_5868);
nor U7962 (N_7962,N_5099,N_4676);
nor U7963 (N_7963,N_4467,N_4428);
nand U7964 (N_7964,N_5782,N_5379);
nand U7965 (N_7965,N_4766,N_5405);
and U7966 (N_7966,N_4687,N_4762);
or U7967 (N_7967,N_4326,N_5716);
or U7968 (N_7968,N_4166,N_5999);
and U7969 (N_7969,N_4561,N_5571);
or U7970 (N_7970,N_5903,N_5605);
nor U7971 (N_7971,N_4265,N_4310);
or U7972 (N_7972,N_5402,N_5488);
nor U7973 (N_7973,N_5164,N_4271);
nor U7974 (N_7974,N_5097,N_4958);
and U7975 (N_7975,N_4913,N_5084);
nand U7976 (N_7976,N_5937,N_4692);
and U7977 (N_7977,N_4356,N_5528);
or U7978 (N_7978,N_5751,N_4415);
nor U7979 (N_7979,N_4448,N_4002);
and U7980 (N_7980,N_4214,N_4479);
or U7981 (N_7981,N_5949,N_5098);
nand U7982 (N_7982,N_4184,N_4794);
or U7983 (N_7983,N_4686,N_4739);
xor U7984 (N_7984,N_5538,N_5940);
nor U7985 (N_7985,N_4682,N_5806);
nand U7986 (N_7986,N_4537,N_4808);
or U7987 (N_7987,N_5778,N_4951);
or U7988 (N_7988,N_4868,N_4845);
or U7989 (N_7989,N_5573,N_4921);
and U7990 (N_7990,N_4974,N_4355);
or U7991 (N_7991,N_4886,N_4615);
or U7992 (N_7992,N_4091,N_5794);
and U7993 (N_7993,N_4257,N_4901);
nand U7994 (N_7994,N_5572,N_4015);
and U7995 (N_7995,N_4032,N_5253);
nor U7996 (N_7996,N_5235,N_4210);
or U7997 (N_7997,N_5230,N_5335);
nand U7998 (N_7998,N_5585,N_4940);
nand U7999 (N_7999,N_5280,N_4280);
nor U8000 (N_8000,N_7746,N_7611);
nand U8001 (N_8001,N_7044,N_7473);
xor U8002 (N_8002,N_6089,N_7916);
or U8003 (N_8003,N_6648,N_6001);
or U8004 (N_8004,N_6238,N_7087);
xnor U8005 (N_8005,N_7743,N_7265);
nand U8006 (N_8006,N_7450,N_7342);
nor U8007 (N_8007,N_6680,N_6787);
nor U8008 (N_8008,N_6927,N_7992);
xnor U8009 (N_8009,N_6370,N_6615);
nor U8010 (N_8010,N_7229,N_7672);
nand U8011 (N_8011,N_6990,N_6818);
or U8012 (N_8012,N_7481,N_6695);
nand U8013 (N_8013,N_6933,N_6505);
nor U8014 (N_8014,N_7008,N_7736);
and U8015 (N_8015,N_7370,N_7027);
or U8016 (N_8016,N_6525,N_6811);
or U8017 (N_8017,N_6110,N_7272);
nand U8018 (N_8018,N_6778,N_7814);
nor U8019 (N_8019,N_7789,N_6214);
or U8020 (N_8020,N_7693,N_7129);
or U8021 (N_8021,N_6373,N_6616);
nor U8022 (N_8022,N_7492,N_7117);
xor U8023 (N_8023,N_6286,N_6762);
and U8024 (N_8024,N_7251,N_7768);
nor U8025 (N_8025,N_7505,N_6497);
xnor U8026 (N_8026,N_6984,N_6488);
nor U8027 (N_8027,N_6071,N_6064);
or U8028 (N_8028,N_7862,N_6069);
or U8029 (N_8029,N_6922,N_7994);
or U8030 (N_8030,N_7310,N_6183);
xor U8031 (N_8031,N_7841,N_7617);
and U8032 (N_8032,N_6063,N_6607);
nand U8033 (N_8033,N_6813,N_6008);
xnor U8034 (N_8034,N_6605,N_7828);
nor U8035 (N_8035,N_6639,N_6832);
nor U8036 (N_8036,N_7501,N_7023);
xor U8037 (N_8037,N_7578,N_6205);
nand U8038 (N_8038,N_7856,N_7902);
or U8039 (N_8039,N_6002,N_6260);
or U8040 (N_8040,N_6215,N_6926);
nand U8041 (N_8041,N_6796,N_7248);
nand U8042 (N_8042,N_7514,N_7622);
nor U8043 (N_8043,N_6599,N_6576);
nand U8044 (N_8044,N_7852,N_7685);
nand U8045 (N_8045,N_6500,N_7052);
nor U8046 (N_8046,N_7085,N_6170);
or U8047 (N_8047,N_6073,N_7754);
nor U8048 (N_8048,N_6782,N_7966);
or U8049 (N_8049,N_7084,N_6232);
and U8050 (N_8050,N_7016,N_6257);
and U8051 (N_8051,N_7772,N_7075);
xor U8052 (N_8052,N_6406,N_7451);
and U8053 (N_8053,N_7638,N_6708);
and U8054 (N_8054,N_7267,N_6612);
xnor U8055 (N_8055,N_6660,N_7006);
or U8056 (N_8056,N_7946,N_6719);
or U8057 (N_8057,N_7998,N_6472);
and U8058 (N_8058,N_7329,N_7669);
or U8059 (N_8059,N_7896,N_7215);
nor U8060 (N_8060,N_6822,N_7857);
nor U8061 (N_8061,N_7463,N_7159);
nor U8062 (N_8062,N_6724,N_6770);
xnor U8063 (N_8063,N_6530,N_6654);
or U8064 (N_8064,N_7634,N_7065);
nand U8065 (N_8065,N_7025,N_6960);
nor U8066 (N_8066,N_6919,N_7456);
or U8067 (N_8067,N_6746,N_7604);
nor U8068 (N_8068,N_6491,N_7162);
nand U8069 (N_8069,N_6803,N_6819);
and U8070 (N_8070,N_7756,N_7525);
xnor U8071 (N_8071,N_7537,N_6240);
or U8072 (N_8072,N_6457,N_7679);
and U8073 (N_8073,N_6084,N_7869);
xor U8074 (N_8074,N_6835,N_7437);
nor U8075 (N_8075,N_6634,N_7628);
nor U8076 (N_8076,N_6829,N_6333);
and U8077 (N_8077,N_7017,N_6589);
xor U8078 (N_8078,N_6833,N_7769);
and U8079 (N_8079,N_6184,N_6595);
and U8080 (N_8080,N_6230,N_7396);
nor U8081 (N_8081,N_6976,N_6425);
nor U8082 (N_8082,N_7262,N_7566);
or U8083 (N_8083,N_7898,N_7987);
or U8084 (N_8084,N_7901,N_6156);
nor U8085 (N_8085,N_7795,N_7101);
nor U8086 (N_8086,N_6195,N_7784);
nand U8087 (N_8087,N_6206,N_6011);
xnor U8088 (N_8088,N_7985,N_7963);
xnor U8089 (N_8089,N_7427,N_6414);
and U8090 (N_8090,N_7173,N_6097);
nand U8091 (N_8091,N_6498,N_7429);
nand U8092 (N_8092,N_6278,N_6553);
or U8093 (N_8093,N_6752,N_7011);
nand U8094 (N_8094,N_7300,N_6596);
nor U8095 (N_8095,N_7298,N_6867);
xnor U8096 (N_8096,N_7171,N_7867);
nor U8097 (N_8097,N_6999,N_7078);
and U8098 (N_8098,N_7252,N_7938);
and U8099 (N_8099,N_7706,N_7147);
nor U8100 (N_8100,N_7840,N_7647);
or U8101 (N_8101,N_7472,N_6633);
or U8102 (N_8102,N_6885,N_7707);
nand U8103 (N_8103,N_6606,N_7741);
nor U8104 (N_8104,N_7076,N_6928);
nor U8105 (N_8105,N_7573,N_6027);
nor U8106 (N_8106,N_6443,N_7710);
and U8107 (N_8107,N_7656,N_6854);
or U8108 (N_8108,N_6776,N_6858);
nand U8109 (N_8109,N_7822,N_6336);
nand U8110 (N_8110,N_6964,N_6555);
xor U8111 (N_8111,N_6850,N_7311);
and U8112 (N_8112,N_6880,N_7060);
and U8113 (N_8113,N_7221,N_6690);
nor U8114 (N_8114,N_7616,N_7132);
and U8115 (N_8115,N_6954,N_7353);
and U8116 (N_8116,N_7696,N_6729);
nand U8117 (N_8117,N_7546,N_7895);
nand U8118 (N_8118,N_7335,N_7127);
and U8119 (N_8119,N_6010,N_6989);
and U8120 (N_8120,N_6619,N_6845);
and U8121 (N_8121,N_6407,N_6542);
nor U8122 (N_8122,N_7281,N_6468);
xnor U8123 (N_8123,N_7760,N_6944);
and U8124 (N_8124,N_7137,N_6973);
or U8125 (N_8125,N_6900,N_7439);
nor U8126 (N_8126,N_6334,N_7788);
nor U8127 (N_8127,N_7392,N_6072);
nor U8128 (N_8128,N_7844,N_6611);
nand U8129 (N_8129,N_7391,N_6985);
nand U8130 (N_8130,N_6123,N_7453);
and U8131 (N_8131,N_6098,N_6853);
xor U8132 (N_8132,N_6795,N_7909);
xnor U8133 (N_8133,N_6480,N_7028);
and U8134 (N_8134,N_7749,N_7661);
nor U8135 (N_8135,N_6843,N_7791);
xor U8136 (N_8136,N_6039,N_7911);
nor U8137 (N_8137,N_7369,N_6251);
nor U8138 (N_8138,N_6149,N_7351);
nor U8139 (N_8139,N_6629,N_7116);
nand U8140 (N_8140,N_6440,N_7759);
and U8141 (N_8141,N_6115,N_6034);
nor U8142 (N_8142,N_7476,N_7061);
or U8143 (N_8143,N_6473,N_7900);
nor U8144 (N_8144,N_6631,N_7196);
or U8145 (N_8145,N_7846,N_6899);
nor U8146 (N_8146,N_7545,N_7811);
or U8147 (N_8147,N_6499,N_6306);
xnor U8148 (N_8148,N_6826,N_6134);
nand U8149 (N_8149,N_6552,N_7907);
and U8150 (N_8150,N_7771,N_6712);
xnor U8151 (N_8151,N_6735,N_7740);
or U8152 (N_8152,N_6534,N_6083);
nor U8153 (N_8153,N_7599,N_7889);
nor U8154 (N_8154,N_7242,N_6288);
and U8155 (N_8155,N_7090,N_7146);
nor U8156 (N_8156,N_6907,N_6846);
nor U8157 (N_8157,N_7705,N_7040);
and U8158 (N_8158,N_6798,N_7515);
or U8159 (N_8159,N_6330,N_6416);
xor U8160 (N_8160,N_6091,N_6020);
or U8161 (N_8161,N_6549,N_7260);
nor U8162 (N_8162,N_6038,N_6598);
nand U8163 (N_8163,N_6346,N_7411);
or U8164 (N_8164,N_6748,N_6879);
and U8165 (N_8165,N_7534,N_7340);
or U8166 (N_8166,N_6824,N_7465);
and U8167 (N_8167,N_7640,N_7919);
or U8168 (N_8168,N_6754,N_7475);
nand U8169 (N_8169,N_6159,N_6541);
and U8170 (N_8170,N_6424,N_6802);
nand U8171 (N_8171,N_7562,N_6276);
xnor U8172 (N_8172,N_6462,N_6231);
nor U8173 (N_8173,N_6358,N_6940);
and U8174 (N_8174,N_7538,N_7539);
xor U8175 (N_8175,N_6906,N_6731);
nand U8176 (N_8176,N_6095,N_6081);
nor U8177 (N_8177,N_6717,N_6766);
and U8178 (N_8178,N_6299,N_7149);
and U8179 (N_8179,N_6108,N_7013);
or U8180 (N_8180,N_7003,N_6378);
xnor U8181 (N_8181,N_6431,N_6613);
or U8182 (N_8182,N_6580,N_7498);
nand U8183 (N_8183,N_7469,N_7285);
and U8184 (N_8184,N_7842,N_7275);
nor U8185 (N_8185,N_7848,N_6959);
or U8186 (N_8186,N_7099,N_6583);
or U8187 (N_8187,N_7321,N_7245);
and U8188 (N_8188,N_6124,N_7209);
or U8189 (N_8189,N_7041,N_6935);
nor U8190 (N_8190,N_7894,N_6895);
or U8191 (N_8191,N_6982,N_7048);
nand U8192 (N_8192,N_6320,N_7767);
nand U8193 (N_8193,N_7373,N_7261);
and U8194 (N_8194,N_6154,N_6799);
and U8195 (N_8195,N_6079,N_6921);
or U8196 (N_8196,N_7205,N_6908);
nor U8197 (N_8197,N_7214,N_6956);
nor U8198 (N_8198,N_7010,N_6855);
and U8199 (N_8199,N_7884,N_6394);
nand U8200 (N_8200,N_6841,N_7558);
nor U8201 (N_8201,N_6451,N_7400);
and U8202 (N_8202,N_6768,N_6780);
nor U8203 (N_8203,N_7021,N_6318);
or U8204 (N_8204,N_7280,N_6666);
nor U8205 (N_8205,N_6936,N_6788);
and U8206 (N_8206,N_7591,N_6475);
nor U8207 (N_8207,N_7928,N_6347);
nor U8208 (N_8208,N_6705,N_6963);
and U8209 (N_8209,N_7477,N_7226);
xor U8210 (N_8210,N_7720,N_7602);
nand U8211 (N_8211,N_6442,N_7605);
or U8212 (N_8212,N_7951,N_6161);
or U8213 (N_8213,N_6916,N_6630);
nand U8214 (N_8214,N_6942,N_6801);
and U8215 (N_8215,N_7999,N_6859);
nor U8216 (N_8216,N_6688,N_7692);
nor U8217 (N_8217,N_7082,N_7303);
nor U8218 (N_8218,N_6622,N_7153);
xnor U8219 (N_8219,N_6465,N_7703);
nor U8220 (N_8220,N_7601,N_6172);
and U8221 (N_8221,N_6847,N_6151);
or U8222 (N_8222,N_6955,N_7623);
xnor U8223 (N_8223,N_6838,N_6592);
or U8224 (N_8224,N_7495,N_6920);
nor U8225 (N_8225,N_7333,N_7444);
or U8226 (N_8226,N_7947,N_6901);
and U8227 (N_8227,N_6308,N_7181);
nand U8228 (N_8228,N_6777,N_6374);
or U8229 (N_8229,N_6896,N_6434);
and U8230 (N_8230,N_7500,N_7920);
and U8231 (N_8231,N_7056,N_6567);
nand U8232 (N_8232,N_7635,N_7751);
xnor U8233 (N_8233,N_7865,N_7677);
or U8234 (N_8234,N_6352,N_7287);
nor U8235 (N_8235,N_6980,N_7511);
nor U8236 (N_8236,N_7151,N_6139);
nor U8237 (N_8237,N_6842,N_7341);
or U8238 (N_8238,N_6540,N_6645);
xor U8239 (N_8239,N_7940,N_7356);
nor U8240 (N_8240,N_7953,N_7521);
nand U8241 (N_8241,N_6699,N_7432);
nand U8242 (N_8242,N_6016,N_6714);
or U8243 (N_8243,N_6902,N_6272);
nor U8244 (N_8244,N_6495,N_6546);
and U8245 (N_8245,N_7874,N_6253);
and U8246 (N_8246,N_6790,N_6691);
and U8247 (N_8247,N_6486,N_7462);
or U8248 (N_8248,N_7454,N_6628);
nor U8249 (N_8249,N_7140,N_7654);
and U8250 (N_8250,N_7405,N_7175);
nor U8251 (N_8251,N_7383,N_7070);
or U8252 (N_8252,N_7580,N_6166);
xor U8253 (N_8253,N_7847,N_6287);
nor U8254 (N_8254,N_6344,N_7544);
nor U8255 (N_8255,N_6222,N_6225);
nor U8256 (N_8256,N_6506,N_6078);
nand U8257 (N_8257,N_6261,N_7490);
or U8258 (N_8258,N_7727,N_7109);
xor U8259 (N_8259,N_6173,N_7125);
and U8260 (N_8260,N_7496,N_6636);
or U8261 (N_8261,N_7160,N_7589);
or U8262 (N_8262,N_6313,N_7086);
nand U8263 (N_8263,N_6529,N_7694);
or U8264 (N_8264,N_6827,N_6673);
and U8265 (N_8265,N_7952,N_6204);
and U8266 (N_8266,N_6825,N_6958);
xor U8267 (N_8267,N_6521,N_6326);
nor U8268 (N_8268,N_7858,N_7503);
or U8269 (N_8269,N_7404,N_6273);
or U8270 (N_8270,N_6861,N_6925);
nand U8271 (N_8271,N_7408,N_6007);
xnor U8272 (N_8272,N_6175,N_6271);
or U8273 (N_8273,N_6792,N_6755);
or U8274 (N_8274,N_6055,N_7831);
and U8275 (N_8275,N_6548,N_7910);
and U8276 (N_8276,N_6446,N_7830);
nor U8277 (N_8277,N_7633,N_6283);
nor U8278 (N_8278,N_7643,N_6201);
or U8279 (N_8279,N_7547,N_6371);
or U8280 (N_8280,N_7022,N_7112);
nand U8281 (N_8281,N_7887,N_7725);
nor U8282 (N_8282,N_7328,N_7415);
nand U8283 (N_8283,N_6651,N_7827);
nand U8284 (N_8284,N_6456,N_7393);
nand U8285 (N_8285,N_6032,N_7349);
nand U8286 (N_8286,N_7988,N_6972);
nand U8287 (N_8287,N_7197,N_6015);
nor U8288 (N_8288,N_6311,N_6076);
nand U8289 (N_8289,N_7177,N_7785);
and U8290 (N_8290,N_7045,N_7266);
nor U8291 (N_8291,N_7676,N_6126);
and U8292 (N_8292,N_6983,N_6602);
xor U8293 (N_8293,N_7435,N_7564);
nand U8294 (N_8294,N_6181,N_7426);
xnor U8295 (N_8295,N_7375,N_6059);
nand U8296 (N_8296,N_7626,N_7877);
and U8297 (N_8297,N_7712,N_6753);
nand U8298 (N_8298,N_7879,N_7773);
nor U8299 (N_8299,N_7796,N_7046);
xnor U8300 (N_8300,N_7761,N_7838);
and U8301 (N_8301,N_7362,N_6804);
nand U8302 (N_8302,N_7674,N_7449);
nand U8303 (N_8303,N_6676,N_6739);
and U8304 (N_8304,N_7230,N_6898);
nor U8305 (N_8305,N_7113,N_6131);
nand U8306 (N_8306,N_6510,N_6444);
or U8307 (N_8307,N_7105,N_6180);
and U8308 (N_8308,N_7908,N_7397);
and U8309 (N_8309,N_6148,N_7993);
or U8310 (N_8310,N_7050,N_7441);
nor U8311 (N_8311,N_6282,N_7627);
nand U8312 (N_8312,N_7675,N_6128);
xor U8313 (N_8313,N_6279,N_7930);
nor U8314 (N_8314,N_6526,N_7357);
nor U8315 (N_8315,N_7452,N_6242);
xnor U8316 (N_8316,N_6736,N_6939);
nand U8317 (N_8317,N_6913,N_6775);
nand U8318 (N_8318,N_7631,N_7419);
or U8319 (N_8319,N_7430,N_7715);
and U8320 (N_8320,N_7567,N_6952);
or U8321 (N_8321,N_7428,N_6709);
xnor U8322 (N_8322,N_6663,N_6036);
nand U8323 (N_8323,N_6177,N_6684);
and U8324 (N_8324,N_7236,N_6568);
and U8325 (N_8325,N_7990,N_6285);
nand U8326 (N_8326,N_7246,N_7192);
nand U8327 (N_8327,N_7620,N_7783);
or U8328 (N_8328,N_6058,N_7648);
and U8329 (N_8329,N_7359,N_7967);
and U8330 (N_8330,N_6934,N_7782);
and U8331 (N_8331,N_6730,N_6946);
or U8332 (N_8332,N_6828,N_7378);
or U8333 (N_8333,N_7584,N_6514);
nor U8334 (N_8334,N_7174,N_6870);
or U8335 (N_8335,N_7774,N_6535);
and U8336 (N_8336,N_7057,N_6050);
nor U8337 (N_8337,N_6369,N_6127);
nor U8338 (N_8338,N_6507,N_6924);
and U8339 (N_8339,N_7063,N_7199);
or U8340 (N_8340,N_6194,N_7290);
nand U8341 (N_8341,N_7120,N_7517);
nand U8342 (N_8342,N_7543,N_7030);
nand U8343 (N_8343,N_7961,N_6138);
nor U8344 (N_8344,N_7243,N_6044);
or U8345 (N_8345,N_7939,N_6259);
and U8346 (N_8346,N_6863,N_7182);
xor U8347 (N_8347,N_6042,N_7960);
nor U8348 (N_8348,N_6192,N_6196);
nand U8349 (N_8349,N_6150,N_6721);
nor U8350 (N_8350,N_6538,N_6678);
or U8351 (N_8351,N_6547,N_7807);
and U8352 (N_8352,N_6996,N_6626);
and U8353 (N_8353,N_6831,N_6948);
nand U8354 (N_8354,N_6670,N_6893);
or U8355 (N_8355,N_7148,N_6119);
nand U8356 (N_8356,N_6968,N_7365);
and U8357 (N_8357,N_6767,N_7766);
xnor U8358 (N_8358,N_7163,N_6087);
and U8359 (N_8359,N_6275,N_7970);
nor U8360 (N_8360,N_6018,N_7211);
or U8361 (N_8361,N_7519,N_6386);
nor U8362 (N_8362,N_7817,N_6104);
nand U8363 (N_8363,N_6435,N_7222);
xnor U8364 (N_8364,N_6569,N_7824);
nand U8365 (N_8365,N_7289,N_6365);
nand U8366 (N_8366,N_6875,N_6429);
and U8367 (N_8367,N_6280,N_7556);
and U8368 (N_8368,N_7312,N_6823);
nor U8369 (N_8369,N_7716,N_6307);
nand U8370 (N_8370,N_7414,N_6614);
and U8371 (N_8371,N_7377,N_6773);
and U8372 (N_8372,N_7409,N_7664);
xnor U8373 (N_8373,N_6566,N_7541);
xor U8374 (N_8374,N_6448,N_7145);
or U8375 (N_8375,N_6049,N_6881);
or U8376 (N_8376,N_6317,N_7352);
or U8377 (N_8377,N_7363,N_6957);
xor U8378 (N_8378,N_6092,N_6892);
xnor U8379 (N_8379,N_7135,N_7776);
or U8380 (N_8380,N_7187,N_6387);
nand U8381 (N_8381,N_6323,N_7283);
nand U8382 (N_8382,N_7941,N_6783);
and U8383 (N_8383,N_7931,N_7058);
or U8384 (N_8384,N_7739,N_7809);
xor U8385 (N_8385,N_6453,N_7121);
and U8386 (N_8386,N_6364,N_7691);
nor U8387 (N_8387,N_6236,N_6303);
xor U8388 (N_8388,N_6395,N_7093);
nor U8389 (N_8389,N_7512,N_6536);
nor U8390 (N_8390,N_7781,N_6353);
nand U8391 (N_8391,N_6551,N_6508);
nand U8392 (N_8392,N_7755,N_7681);
nor U8393 (N_8393,N_7855,N_7508);
or U8394 (N_8394,N_7374,N_6384);
or U8395 (N_8395,N_6786,N_6143);
nand U8396 (N_8396,N_6221,N_6603);
nor U8397 (N_8397,N_6993,N_6910);
or U8398 (N_8398,N_6579,N_6400);
nand U8399 (N_8399,N_7358,N_7954);
nor U8400 (N_8400,N_6683,N_6393);
or U8401 (N_8401,N_6812,N_6176);
nand U8402 (N_8402,N_6597,N_7819);
or U8403 (N_8403,N_6668,N_6707);
nand U8404 (N_8404,N_7032,N_6375);
xnor U8405 (N_8405,N_6997,N_7764);
nor U8406 (N_8406,N_6856,N_6153);
nor U8407 (N_8407,N_6341,N_7779);
nand U8408 (N_8408,N_7594,N_7216);
and U8409 (N_8409,N_7976,N_6322);
or U8410 (N_8410,N_6392,N_7395);
and U8411 (N_8411,N_7059,N_6327);
nor U8412 (N_8412,N_7188,N_7007);
nor U8413 (N_8413,N_7313,N_7925);
nor U8414 (N_8414,N_7241,N_7097);
nor U8415 (N_8415,N_6970,N_7870);
nor U8416 (N_8416,N_7719,N_6168);
and U8417 (N_8417,N_6677,N_7015);
and U8418 (N_8418,N_7263,N_6671);
nor U8419 (N_8419,N_6995,N_6800);
xnor U8420 (N_8420,N_6740,N_6367);
or U8421 (N_8421,N_7823,N_7816);
xnor U8422 (N_8422,N_7237,N_7786);
nand U8423 (N_8423,N_6931,N_6621);
and U8424 (N_8424,N_6361,N_7055);
and U8425 (N_8425,N_7651,N_6485);
nor U8426 (N_8426,N_7297,N_7001);
nand U8427 (N_8427,N_6966,N_6969);
nand U8428 (N_8428,N_7168,N_7520);
nor U8429 (N_8429,N_7406,N_6235);
nand U8430 (N_8430,N_7098,N_6243);
nor U8431 (N_8431,N_7014,N_6132);
xnor U8432 (N_8432,N_7903,N_7401);
or U8433 (N_8433,N_6099,N_6487);
nor U8434 (N_8434,N_6332,N_7753);
or U8435 (N_8435,N_7973,N_6586);
or U8436 (N_8436,N_7073,N_7306);
or U8437 (N_8437,N_6284,N_7258);
nor U8438 (N_8438,N_7942,N_6074);
or U8439 (N_8439,N_6065,N_6821);
nor U8440 (N_8440,N_6292,N_6624);
and U8441 (N_8441,N_7047,N_7569);
nor U8442 (N_8442,N_6028,N_7202);
or U8443 (N_8443,N_7757,N_7354);
nor U8444 (N_8444,N_7530,N_6789);
or U8445 (N_8445,N_7367,N_7645);
nand U8446 (N_8446,N_7480,N_6022);
nand U8447 (N_8447,N_7386,N_7253);
nor U8448 (N_8448,N_7913,N_7080);
or U8449 (N_8449,N_7882,N_7642);
and U8450 (N_8450,N_7293,N_6986);
nor U8451 (N_8451,N_7667,N_6390);
nor U8452 (N_8452,N_6295,N_7886);
xnor U8453 (N_8453,N_7379,N_7004);
xnor U8454 (N_8454,N_6531,N_7264);
nand U8455 (N_8455,N_6815,N_7979);
nor U8456 (N_8456,N_6264,N_7169);
nor U8457 (N_8457,N_7650,N_6449);
nand U8458 (N_8458,N_6447,N_7596);
and U8459 (N_8459,N_6190,N_7348);
and U8460 (N_8460,N_6522,N_7270);
xnor U8461 (N_8461,N_6075,N_7536);
xor U8462 (N_8462,N_7744,N_7799);
and U8463 (N_8463,N_7583,N_6187);
nor U8464 (N_8464,N_6391,N_6136);
or U8465 (N_8465,N_7726,N_6116);
and U8466 (N_8466,N_7190,N_7559);
and U8467 (N_8467,N_7704,N_6158);
nand U8468 (N_8468,N_7598,N_6558);
nor U8469 (N_8469,N_7522,N_7304);
xnor U8470 (N_8470,N_7549,N_7587);
nor U8471 (N_8471,N_7557,N_6355);
and U8472 (N_8472,N_6247,N_7800);
or U8473 (N_8473,N_6309,N_7944);
nor U8474 (N_8474,N_7005,N_7470);
and U8475 (N_8475,N_6025,N_7618);
xnor U8476 (N_8476,N_6067,N_7975);
nor U8477 (N_8477,N_6869,N_7096);
nand U8478 (N_8478,N_7295,N_7144);
or U8479 (N_8479,N_6426,N_6246);
and U8480 (N_8480,N_6410,N_7042);
and U8481 (N_8481,N_6545,N_6217);
and U8482 (N_8482,N_6665,N_7459);
or U8483 (N_8483,N_6223,N_7069);
nand U8484 (N_8484,N_7191,N_6419);
and U8485 (N_8485,N_6797,N_7875);
nand U8486 (N_8486,N_6675,N_6492);
or U8487 (N_8487,N_6561,N_7416);
nor U8488 (N_8488,N_7964,N_6991);
nand U8489 (N_8489,N_6047,N_7487);
or U8490 (N_8490,N_7899,N_7049);
or U8491 (N_8491,N_6618,N_6021);
nor U8492 (N_8492,N_6100,N_7036);
nor U8493 (N_8493,N_6737,N_6713);
or U8494 (N_8494,N_7418,N_7336);
nand U8495 (N_8495,N_7762,N_6300);
and U8496 (N_8496,N_7550,N_7658);
and U8497 (N_8497,N_6694,N_6031);
xor U8498 (N_8498,N_6733,N_7804);
or U8499 (N_8499,N_6682,N_6040);
or U8500 (N_8500,N_7154,N_6662);
nand U8501 (N_8501,N_6584,N_6112);
nand U8502 (N_8502,N_7257,N_7655);
and U8503 (N_8503,N_7936,N_7102);
or U8504 (N_8504,N_7836,N_7170);
nand U8505 (N_8505,N_6200,N_6887);
nand U8506 (N_8506,N_6199,N_7053);
nor U8507 (N_8507,N_6241,N_7614);
or U8508 (N_8508,N_7646,N_6360);
or U8509 (N_8509,N_7748,N_7315);
nand U8510 (N_8510,N_6174,N_7832);
nand U8511 (N_8511,N_6653,N_6617);
or U8512 (N_8512,N_6565,N_7424);
nand U8513 (N_8513,N_7542,N_7815);
nand U8514 (N_8514,N_7288,N_6994);
nor U8515 (N_8515,N_7853,N_7371);
xor U8516 (N_8516,N_7305,N_6741);
and U8517 (N_8517,N_6297,N_6747);
nor U8518 (N_8518,N_6588,N_6930);
or U8519 (N_8519,N_7972,N_6848);
and U8520 (N_8520,N_6005,N_7206);
nor U8521 (N_8521,N_6179,N_7234);
or U8522 (N_8522,N_7457,N_7745);
nor U8523 (N_8523,N_7235,N_7625);
nor U8524 (N_8524,N_6359,N_7600);
nor U8525 (N_8525,N_7533,N_6321);
or U8526 (N_8526,N_7122,N_6345);
nand U8527 (N_8527,N_7568,N_7504);
and U8528 (N_8528,N_6474,N_6904);
nand U8529 (N_8529,N_6886,N_6593);
and U8530 (N_8530,N_6340,N_6537);
nand U8531 (N_8531,N_7644,N_6220);
or U8532 (N_8532,N_6455,N_7662);
nor U8533 (N_8533,N_6757,N_6977);
nand U8534 (N_8534,N_6239,N_7820);
and U8535 (N_8535,N_6503,N_6820);
nor U8536 (N_8536,N_6539,N_7141);
nand U8537 (N_8537,N_6467,N_7384);
or U8538 (N_8538,N_6572,N_7731);
and U8539 (N_8539,N_7278,N_7714);
nand U8540 (N_8540,N_7043,N_6974);
and U8541 (N_8541,N_7361,N_7621);
nand U8542 (N_8542,N_6274,N_6701);
xnor U8543 (N_8543,N_6923,N_6209);
nor U8544 (N_8544,N_7808,N_6398);
nor U8545 (N_8545,N_7851,N_6248);
nor U8546 (N_8546,N_6610,N_7455);
and U8547 (N_8547,N_7958,N_6113);
nand U8548 (N_8548,N_6105,N_6411);
nand U8549 (N_8549,N_6494,N_6484);
xnor U8550 (N_8550,N_6329,N_7565);
or U8551 (N_8551,N_6385,N_6082);
and U8552 (N_8552,N_7797,N_7179);
nor U8553 (N_8553,N_6490,N_7156);
nand U8554 (N_8554,N_7484,N_7969);
and U8555 (N_8555,N_7029,N_7872);
nand U8556 (N_8556,N_7943,N_6937);
or U8557 (N_8557,N_7031,N_7632);
or U8558 (N_8558,N_6661,N_7826);
nor U8559 (N_8559,N_7284,N_7142);
nand U8560 (N_8560,N_6849,N_6866);
or U8561 (N_8561,N_7552,N_6328);
nor U8562 (N_8562,N_6256,N_6316);
nand U8563 (N_8563,N_7037,N_7423);
nand U8564 (N_8564,N_7167,N_6738);
or U8565 (N_8565,N_7033,N_7307);
nand U8566 (N_8566,N_7124,N_6716);
nor U8567 (N_8567,N_6669,N_6101);
xnor U8568 (N_8568,N_6987,N_6335);
nor U8569 (N_8569,N_7332,N_6878);
nor U8570 (N_8570,N_7986,N_7100);
nor U8571 (N_8571,N_6476,N_6430);
xor U8572 (N_8572,N_6354,N_6758);
and U8573 (N_8573,N_6532,N_7866);
or U8574 (N_8574,N_7347,N_7527);
nor U8575 (N_8575,N_6319,N_7528);
xnor U8576 (N_8576,N_6765,N_6277);
and U8577 (N_8577,N_7213,N_6533);
and U8578 (N_8578,N_7184,N_7666);
or U8579 (N_8579,N_7071,N_7734);
and U8580 (N_8580,N_7548,N_6118);
and U8581 (N_8581,N_7834,N_6702);
and U8582 (N_8582,N_6992,N_6441);
and U8583 (N_8583,N_7412,N_7850);
and U8584 (N_8584,N_7709,N_6404);
or U8585 (N_8585,N_7343,N_7268);
or U8586 (N_8586,N_6627,N_6646);
or U8587 (N_8587,N_7054,N_6160);
or U8588 (N_8588,N_6761,N_6657);
nor U8589 (N_8589,N_6145,N_6315);
nand U8590 (N_8590,N_6213,N_6338);
nand U8591 (N_8591,N_7366,N_6388);
nor U8592 (N_8592,N_7161,N_7372);
or U8593 (N_8593,N_6851,N_6023);
or U8594 (N_8594,N_6269,N_6681);
or U8595 (N_8595,N_7603,N_7535);
nand U8596 (N_8596,N_6844,N_6728);
or U8597 (N_8597,N_7152,N_7700);
nor U8598 (N_8598,N_6650,N_6403);
and U8599 (N_8599,N_7183,N_6590);
and U8600 (N_8600,N_6524,N_7860);
nor U8601 (N_8601,N_6897,N_6637);
nand U8602 (N_8602,N_6122,N_6718);
nand U8603 (N_8603,N_7518,N_7180);
nor U8604 (N_8604,N_6706,N_7684);
or U8605 (N_8605,N_7394,N_6109);
and U8606 (N_8606,N_6003,N_7561);
and U8607 (N_8607,N_7506,N_6017);
or U8608 (N_8608,N_6281,N_6581);
nor U8609 (N_8609,N_6268,N_6967);
or U8610 (N_8610,N_7592,N_6342);
xnor U8611 (N_8611,N_7641,N_6399);
and U8612 (N_8612,N_7721,N_7697);
and U8613 (N_8613,N_6562,N_6903);
or U8614 (N_8614,N_7585,N_6750);
and U8615 (N_8615,N_6950,N_6601);
nor U8616 (N_8616,N_6884,N_7659);
nor U8617 (N_8617,N_6012,N_7493);
nand U8618 (N_8618,N_7034,N_7688);
or U8619 (N_8619,N_6270,N_6077);
nand U8620 (N_8620,N_6703,N_7904);
nand U8621 (N_8621,N_7921,N_6254);
nand U8622 (N_8622,N_7540,N_7572);
nand U8623 (N_8623,N_6185,N_6427);
nor U8624 (N_8624,N_7956,N_7238);
or U8625 (N_8625,N_7730,N_6046);
xnor U8626 (N_8626,N_7989,N_7433);
nor U8627 (N_8627,N_6520,N_7590);
nor U8628 (N_8628,N_7934,N_7271);
and U8629 (N_8629,N_7380,N_6219);
and U8630 (N_8630,N_7917,N_7794);
nand U8631 (N_8631,N_7195,N_6961);
or U8632 (N_8632,N_6401,N_7955);
or U8633 (N_8633,N_6481,N_6417);
nand U8634 (N_8634,N_6685,N_6026);
or U8635 (N_8635,N_7554,N_7223);
and U8636 (N_8636,N_6756,N_6865);
or U8637 (N_8637,N_7448,N_7711);
xor U8638 (N_8638,N_7702,N_6909);
nor U8639 (N_8639,N_7765,N_6111);
nand U8640 (N_8640,N_6193,N_7198);
nand U8641 (N_8641,N_6035,N_7276);
nand U8642 (N_8642,N_7337,N_7000);
nand U8643 (N_8643,N_6226,N_7225);
xor U8644 (N_8644,N_6437,N_7968);
and U8645 (N_8645,N_7957,N_7582);
or U8646 (N_8646,N_7532,N_6054);
or U8647 (N_8647,N_6512,N_7445);
nor U8648 (N_8648,N_6422,N_6428);
nand U8649 (N_8649,N_7713,N_6571);
and U8650 (N_8650,N_6211,N_6772);
nor U8651 (N_8651,N_6785,N_7577);
nand U8652 (N_8652,N_7837,N_7020);
nor U8653 (N_8653,N_7322,N_6656);
nand U8654 (N_8654,N_6343,N_6006);
nand U8655 (N_8655,N_7232,N_6517);
or U8656 (N_8656,N_7106,N_6304);
and U8657 (N_8657,N_7758,N_7612);
nand U8658 (N_8658,N_7325,N_7918);
or U8659 (N_8659,N_6951,N_7239);
or U8660 (N_8660,N_7932,N_7255);
nor U8661 (N_8661,N_6658,N_7510);
nand U8662 (N_8662,N_6249,N_6839);
or U8663 (N_8663,N_6372,N_6258);
nand U8664 (N_8664,N_7608,N_7780);
or U8665 (N_8665,N_6912,N_7402);
nand U8666 (N_8666,N_7868,N_6502);
nand U8667 (N_8667,N_7474,N_7863);
and U8668 (N_8668,N_6037,N_7588);
and U8669 (N_8669,N_7763,N_6623);
nor U8670 (N_8670,N_6169,N_6045);
nor U8671 (N_8671,N_7131,N_6218);
nor U8672 (N_8672,N_7443,N_7890);
and U8673 (N_8673,N_6339,N_7790);
and U8674 (N_8674,N_7390,N_7576);
nor U8675 (N_8675,N_7479,N_7296);
nor U8676 (N_8676,N_6088,N_7478);
and U8677 (N_8677,N_7324,N_7224);
and U8678 (N_8678,N_6167,N_6759);
xor U8679 (N_8679,N_6632,N_6519);
xnor U8680 (N_8680,N_7653,N_6471);
or U8681 (N_8681,N_6771,N_7350);
nor U8682 (N_8682,N_6697,N_6988);
nor U8683 (N_8683,N_6405,N_6182);
and U8684 (N_8684,N_7286,N_6250);
and U8685 (N_8685,N_7081,N_6806);
or U8686 (N_8686,N_7133,N_6096);
nand U8687 (N_8687,N_7555,N_7805);
and U8688 (N_8688,N_6917,N_7812);
nand U8689 (N_8689,N_7802,N_6245);
xnor U8690 (N_8690,N_6080,N_6945);
and U8691 (N_8691,N_6265,N_6725);
nand U8692 (N_8692,N_6482,N_7308);
nor U8693 (N_8693,N_6379,N_7615);
nor U8694 (N_8694,N_7323,N_7927);
nor U8695 (N_8695,N_6860,N_7861);
nand U8696 (N_8696,N_6751,N_7360);
nand U8697 (N_8697,N_7250,N_6979);
and U8698 (N_8698,N_7491,N_6975);
nand U8699 (N_8699,N_6291,N_6817);
or U8700 (N_8700,N_7845,N_6876);
nor U8701 (N_8701,N_6436,N_6030);
nor U8702 (N_8702,N_7813,N_7164);
and U8703 (N_8703,N_7165,N_6560);
nor U8704 (N_8704,N_6723,N_6188);
or U8705 (N_8705,N_6396,N_7438);
or U8706 (N_8706,N_6383,N_6402);
or U8707 (N_8707,N_6478,N_6483);
and U8708 (N_8708,N_6978,N_6382);
or U8709 (N_8709,N_7607,N_7193);
xnor U8710 (N_8710,N_7933,N_6808);
nand U8711 (N_8711,N_6198,N_6672);
or U8712 (N_8712,N_6423,N_7186);
nor U8713 (N_8713,N_6679,N_7442);
xor U8714 (N_8714,N_7126,N_7787);
nor U8715 (N_8715,N_6041,N_7381);
or U8716 (N_8716,N_6152,N_7247);
nand U8717 (N_8717,N_6652,N_7345);
nand U8718 (N_8718,N_7309,N_6504);
and U8719 (N_8719,N_7327,N_6696);
nand U8720 (N_8720,N_6397,N_7778);
or U8721 (N_8721,N_6516,N_6090);
and U8722 (N_8722,N_6244,N_7108);
nor U8723 (N_8723,N_6362,N_7344);
and U8724 (N_8724,N_7570,N_7485);
nor U8725 (N_8725,N_7652,N_6464);
and U8726 (N_8726,N_6809,N_7294);
nor U8727 (N_8727,N_7273,N_6852);
and U8728 (N_8728,N_7368,N_6459);
nand U8729 (N_8729,N_6013,N_6466);
nand U8730 (N_8730,N_7104,N_7138);
xnor U8731 (N_8731,N_6769,N_6877);
nand U8732 (N_8732,N_6556,N_7531);
and U8733 (N_8733,N_6155,N_6544);
xor U8734 (N_8734,N_7924,N_7038);
nand U8735 (N_8735,N_7079,N_6608);
or U8736 (N_8736,N_6454,N_7597);
or U8737 (N_8737,N_7747,N_7434);
or U8738 (N_8738,N_7077,N_6237);
or U8739 (N_8739,N_6147,N_6894);
or U8740 (N_8740,N_7801,N_7945);
nor U8741 (N_8741,N_6094,N_7421);
nor U8742 (N_8742,N_7128,N_7810);
and U8743 (N_8743,N_6998,N_6057);
nand U8744 (N_8744,N_6171,N_7088);
nand U8745 (N_8745,N_7166,N_6644);
nor U8746 (N_8746,N_7482,N_6133);
xor U8747 (N_8747,N_7207,N_7637);
xnor U8748 (N_8748,N_6189,N_6742);
nor U8749 (N_8749,N_7089,N_6178);
and U8750 (N_8750,N_7299,N_7218);
or U8751 (N_8751,N_6061,N_6102);
and U8752 (N_8752,N_6710,N_6162);
or U8753 (N_8753,N_7984,N_7563);
nor U8754 (N_8754,N_6577,N_6068);
nor U8755 (N_8755,N_6791,N_7657);
and U8756 (N_8756,N_6452,N_7732);
nor U8757 (N_8757,N_6513,N_7636);
and U8758 (N_8758,N_6625,N_7876);
and U8759 (N_8759,N_7254,N_7355);
and U8760 (N_8760,N_6301,N_7339);
xor U8761 (N_8761,N_7039,N_6186);
nand U8762 (N_8762,N_6368,N_7157);
nand U8763 (N_8763,N_7948,N_7905);
nor U8764 (N_8764,N_7729,N_6953);
or U8765 (N_8765,N_6381,N_6043);
nand U8766 (N_8766,N_7798,N_6445);
nand U8767 (N_8767,N_6210,N_6229);
nor U8768 (N_8768,N_7581,N_6647);
nor U8769 (N_8769,N_7407,N_6203);
nor U8770 (N_8770,N_6350,N_7971);
xnor U8771 (N_8771,N_7833,N_6489);
nand U8772 (N_8772,N_7864,N_6366);
nand U8773 (N_8773,N_6458,N_6888);
or U8774 (N_8774,N_7064,N_7978);
nand U8775 (N_8775,N_7103,N_7770);
xor U8776 (N_8776,N_6418,N_6305);
or U8777 (N_8777,N_7217,N_6834);
or U8778 (N_8778,N_7935,N_7035);
nor U8779 (N_8779,N_7489,N_6807);
and U8780 (N_8780,N_6029,N_6620);
nand U8781 (N_8781,N_7668,N_6348);
nor U8782 (N_8782,N_7708,N_6915);
or U8783 (N_8783,N_6543,N_6337);
or U8784 (N_8784,N_6052,N_7673);
and U8785 (N_8785,N_7292,N_7571);
xor U8786 (N_8786,N_6314,N_7468);
xor U8787 (N_8787,N_7018,N_6962);
xnor U8788 (N_8788,N_7072,N_7291);
nor U8789 (N_8789,N_6689,N_6294);
or U8790 (N_8790,N_6949,N_7240);
xor U8791 (N_8791,N_7639,N_7923);
nor U8792 (N_8792,N_6570,N_6107);
nor U8793 (N_8793,N_6743,N_6862);
nor U8794 (N_8794,N_6609,N_7891);
nand U8795 (N_8795,N_6635,N_6574);
nand U8796 (N_8796,N_6377,N_6698);
or U8797 (N_8797,N_7095,N_7914);
or U8798 (N_8798,N_6053,N_7486);
nor U8799 (N_8799,N_6763,N_6056);
and U8800 (N_8800,N_7200,N_7977);
and U8801 (N_8801,N_7663,N_7389);
or U8802 (N_8802,N_7466,N_7735);
and U8803 (N_8803,N_6325,N_6700);
nor U8804 (N_8804,N_6130,N_6883);
nor U8805 (N_8805,N_7609,N_6501);
and U8806 (N_8806,N_7203,N_6420);
or U8807 (N_8807,N_7208,N_7051);
and U8808 (N_8808,N_7301,N_7425);
nand U8809 (N_8809,N_7422,N_6929);
nor U8810 (N_8810,N_6106,N_7883);
and U8811 (N_8811,N_7873,N_6137);
nand U8812 (N_8812,N_6421,N_6911);
or U8813 (N_8813,N_6814,N_7915);
nand U8814 (N_8814,N_6310,N_6642);
nor U8815 (N_8815,N_6585,N_7436);
nor U8816 (N_8816,N_6760,N_6349);
and U8817 (N_8817,N_6479,N_6575);
or U8818 (N_8818,N_6024,N_6550);
and U8819 (N_8819,N_7682,N_6296);
or U8820 (N_8820,N_6331,N_7619);
or U8821 (N_8821,N_6600,N_7665);
and U8822 (N_8822,N_6266,N_6591);
and U8823 (N_8823,N_7446,N_7269);
and U8824 (N_8824,N_7733,N_7210);
or U8825 (N_8825,N_7680,N_6009);
nand U8826 (N_8826,N_6263,N_7256);
or U8827 (N_8827,N_6947,N_7410);
nor U8828 (N_8828,N_7630,N_7026);
nor U8829 (N_8829,N_7885,N_7690);
nand U8830 (N_8830,N_7074,N_6062);
xor U8831 (N_8831,N_6874,N_6120);
nand U8832 (N_8832,N_7143,N_7461);
nor U8833 (N_8833,N_6351,N_6103);
and U8834 (N_8834,N_6564,N_7274);
and U8835 (N_8835,N_7024,N_7922);
or U8836 (N_8836,N_7686,N_6060);
nor U8837 (N_8837,N_7185,N_6509);
nand U8838 (N_8838,N_6918,N_6412);
and U8839 (N_8839,N_7382,N_6460);
nand U8840 (N_8840,N_7871,N_7678);
and U8841 (N_8841,N_6692,N_7529);
nand U8842 (N_8842,N_7687,N_7139);
xnor U8843 (N_8843,N_7722,N_7888);
nor U8844 (N_8844,N_7346,N_7440);
or U8845 (N_8845,N_7134,N_7792);
and U8846 (N_8846,N_6704,N_6004);
xnor U8847 (N_8847,N_7399,N_7660);
or U8848 (N_8848,N_6114,N_7067);
nand U8849 (N_8849,N_6674,N_7803);
and U8850 (N_8850,N_7906,N_7115);
nor U8851 (N_8851,N_7695,N_6659);
and U8852 (N_8852,N_6376,N_6890);
nor U8853 (N_8853,N_6212,N_6450);
nor U8854 (N_8854,N_6216,N_7219);
nor U8855 (N_8855,N_6191,N_7793);
nand U8856 (N_8856,N_7912,N_6836);
nor U8857 (N_8857,N_6649,N_6142);
nand U8858 (N_8858,N_6496,N_7937);
nor U8859 (N_8859,N_6722,N_7818);
and U8860 (N_8860,N_7509,N_7233);
nand U8861 (N_8861,N_7316,N_6085);
xnor U8862 (N_8862,N_6805,N_6655);
xor U8863 (N_8863,N_7551,N_6745);
or U8864 (N_8864,N_6965,N_6981);
and U8865 (N_8865,N_7277,N_7728);
and U8866 (N_8866,N_7398,N_6873);
nor U8867 (N_8867,N_6518,N_6781);
nor U8868 (N_8868,N_6882,N_6527);
or U8869 (N_8869,N_7995,N_6228);
and U8870 (N_8870,N_6943,N_6559);
nand U8871 (N_8871,N_6687,N_7494);
nand U8872 (N_8872,N_6711,N_7320);
and U8873 (N_8873,N_7110,N_6554);
nor U8874 (N_8874,N_6582,N_6493);
or U8875 (N_8875,N_7775,N_7483);
nand U8876 (N_8876,N_7388,N_6227);
and U8877 (N_8877,N_7523,N_6816);
nand U8878 (N_8878,N_6938,N_7497);
xnor U8879 (N_8879,N_6312,N_6726);
nand U8880 (N_8880,N_6774,N_7649);
or U8881 (N_8881,N_7777,N_6298);
or U8882 (N_8882,N_6511,N_7574);
and U8883 (N_8883,N_6293,N_7227);
xnor U8884 (N_8884,N_6640,N_6389);
and U8885 (N_8885,N_6267,N_6557);
nand U8886 (N_8886,N_7458,N_7835);
xor U8887 (N_8887,N_7897,N_7318);
nand U8888 (N_8888,N_7279,N_7338);
nor U8889 (N_8889,N_6000,N_6324);
or U8890 (N_8890,N_6732,N_6905);
and U8891 (N_8891,N_7201,N_7991);
or U8892 (N_8892,N_6667,N_6749);
nand U8893 (N_8893,N_7189,N_6197);
nand U8894 (N_8894,N_7194,N_7331);
nand U8895 (N_8895,N_7892,N_7178);
nand U8896 (N_8896,N_7606,N_7507);
and U8897 (N_8897,N_7959,N_7854);
nand U8898 (N_8898,N_7893,N_6380);
or U8899 (N_8899,N_6048,N_6019);
or U8900 (N_8900,N_6727,N_6563);
and U8901 (N_8901,N_7417,N_6871);
nor U8902 (N_8902,N_7431,N_6477);
and U8903 (N_8903,N_7737,N_7949);
nand U8904 (N_8904,N_6810,N_7698);
nand U8905 (N_8905,N_6086,N_7464);
and U8906 (N_8906,N_7881,N_6093);
nor U8907 (N_8907,N_6515,N_7176);
and U8908 (N_8908,N_6840,N_6734);
and U8909 (N_8909,N_7387,N_7624);
and U8910 (N_8910,N_7155,N_7460);
and U8911 (N_8911,N_6914,N_7136);
nor U8912 (N_8912,N_6686,N_6140);
or U8913 (N_8913,N_7843,N_6864);
xnor U8914 (N_8914,N_7249,N_7839);
nor U8915 (N_8915,N_7499,N_7997);
nor U8916 (N_8916,N_7403,N_6357);
and U8917 (N_8917,N_7717,N_7965);
and U8918 (N_8918,N_7880,N_6784);
nand U8919 (N_8919,N_7513,N_6255);
or U8920 (N_8920,N_7066,N_7319);
xnor U8921 (N_8921,N_7119,N_6157);
and U8922 (N_8922,N_6872,N_6409);
or U8923 (N_8923,N_7962,N_6363);
nand U8924 (N_8924,N_7282,N_7750);
nor U8925 (N_8925,N_6432,N_6433);
nand U8926 (N_8926,N_7302,N_6573);
and U8927 (N_8927,N_6971,N_7012);
nand U8928 (N_8928,N_7091,N_7575);
nand U8929 (N_8929,N_7502,N_7228);
nor U8930 (N_8930,N_7524,N_6837);
nand U8931 (N_8931,N_7118,N_7172);
or U8932 (N_8932,N_6070,N_6715);
nand U8933 (N_8933,N_7204,N_6066);
and U8934 (N_8934,N_6469,N_7974);
nand U8935 (N_8935,N_7689,N_7107);
or U8936 (N_8936,N_7718,N_7670);
nor U8937 (N_8937,N_6604,N_7593);
nand U8938 (N_8938,N_7996,N_7560);
xor U8939 (N_8939,N_7114,N_6207);
and U8940 (N_8940,N_7231,N_6463);
nand U8941 (N_8941,N_6356,N_6121);
nor U8942 (N_8942,N_7326,N_6470);
or U8943 (N_8943,N_7244,N_7629);
and U8944 (N_8944,N_7447,N_6302);
nand U8945 (N_8945,N_6932,N_6523);
and U8946 (N_8946,N_6408,N_6830);
nand U8947 (N_8947,N_7586,N_7420);
nand U8948 (N_8948,N_7829,N_7083);
and U8949 (N_8949,N_6587,N_7983);
nand U8950 (N_8950,N_7314,N_6125);
nand U8951 (N_8951,N_6779,N_7130);
nor U8952 (N_8952,N_6594,N_6224);
and U8953 (N_8953,N_6638,N_7738);
nor U8954 (N_8954,N_7926,N_6693);
nor U8955 (N_8955,N_6129,N_6234);
nand U8956 (N_8956,N_7259,N_6438);
nor U8957 (N_8957,N_7683,N_6165);
nand U8958 (N_8958,N_6720,N_7526);
nand U8959 (N_8959,N_6262,N_6033);
nor U8960 (N_8960,N_7981,N_6578);
nand U8961 (N_8961,N_6208,N_6941);
or U8962 (N_8962,N_7825,N_6643);
nor U8963 (N_8963,N_6889,N_6793);
or U8964 (N_8964,N_7123,N_7158);
nor U8965 (N_8965,N_6146,N_7150);
nor U8966 (N_8966,N_7330,N_7471);
or U8967 (N_8967,N_6461,N_6794);
nand U8968 (N_8968,N_7334,N_6289);
and U8969 (N_8969,N_7111,N_7859);
xnor U8970 (N_8970,N_6202,N_7009);
or U8971 (N_8971,N_7752,N_7980);
and U8972 (N_8972,N_6051,N_7821);
and U8973 (N_8973,N_6252,N_6641);
and U8974 (N_8974,N_7488,N_6415);
and U8975 (N_8975,N_7068,N_7376);
or U8976 (N_8976,N_7019,N_6868);
xnor U8977 (N_8977,N_7385,N_7701);
nor U8978 (N_8978,N_6290,N_7929);
and U8979 (N_8979,N_7092,N_7699);
or U8980 (N_8980,N_7317,N_7724);
or U8981 (N_8981,N_6014,N_7364);
nand U8982 (N_8982,N_6664,N_7002);
xor U8983 (N_8983,N_7062,N_7553);
nand U8984 (N_8984,N_6764,N_7613);
or U8985 (N_8985,N_7806,N_6891);
nand U8986 (N_8986,N_7579,N_6413);
or U8987 (N_8987,N_7671,N_6439);
nand U8988 (N_8988,N_7595,N_6144);
nand U8989 (N_8989,N_7516,N_6233);
nor U8990 (N_8990,N_7413,N_6857);
and U8991 (N_8991,N_7742,N_7212);
nor U8992 (N_8992,N_6141,N_7878);
or U8993 (N_8993,N_6163,N_6744);
nand U8994 (N_8994,N_7950,N_7220);
and U8995 (N_8995,N_6117,N_7849);
nor U8996 (N_8996,N_6528,N_6164);
and U8997 (N_8997,N_7610,N_7094);
nor U8998 (N_8998,N_7723,N_6135);
and U8999 (N_8999,N_7467,N_7982);
or U9000 (N_9000,N_6091,N_6093);
and U9001 (N_9001,N_7771,N_7137);
nor U9002 (N_9002,N_6892,N_7126);
nand U9003 (N_9003,N_6137,N_6261);
nor U9004 (N_9004,N_7190,N_6233);
nand U9005 (N_9005,N_7943,N_7524);
xor U9006 (N_9006,N_6677,N_7406);
nor U9007 (N_9007,N_6598,N_7397);
nand U9008 (N_9008,N_6474,N_6949);
nor U9009 (N_9009,N_7586,N_7706);
and U9010 (N_9010,N_7009,N_7432);
nor U9011 (N_9011,N_7866,N_7803);
or U9012 (N_9012,N_7227,N_6207);
nand U9013 (N_9013,N_6570,N_7432);
nand U9014 (N_9014,N_7537,N_7467);
and U9015 (N_9015,N_7312,N_6765);
nand U9016 (N_9016,N_7619,N_7529);
or U9017 (N_9017,N_7893,N_7480);
nor U9018 (N_9018,N_6524,N_6286);
nand U9019 (N_9019,N_6765,N_7642);
xor U9020 (N_9020,N_7207,N_6526);
nand U9021 (N_9021,N_7753,N_7555);
nor U9022 (N_9022,N_7397,N_7863);
or U9023 (N_9023,N_6180,N_7918);
or U9024 (N_9024,N_7685,N_6707);
or U9025 (N_9025,N_6408,N_6522);
or U9026 (N_9026,N_6139,N_6144);
nand U9027 (N_9027,N_7126,N_6032);
nor U9028 (N_9028,N_6788,N_6652);
or U9029 (N_9029,N_6513,N_6680);
xor U9030 (N_9030,N_6493,N_7993);
or U9031 (N_9031,N_6653,N_6984);
nand U9032 (N_9032,N_6692,N_7333);
nand U9033 (N_9033,N_7187,N_7305);
nand U9034 (N_9034,N_7234,N_7944);
or U9035 (N_9035,N_6635,N_6106);
and U9036 (N_9036,N_7965,N_6489);
nor U9037 (N_9037,N_6522,N_7179);
xnor U9038 (N_9038,N_7718,N_6195);
xor U9039 (N_9039,N_6276,N_6891);
or U9040 (N_9040,N_7196,N_6621);
nor U9041 (N_9041,N_7705,N_7867);
or U9042 (N_9042,N_6631,N_6525);
or U9043 (N_9043,N_6867,N_7031);
nand U9044 (N_9044,N_6308,N_6651);
nor U9045 (N_9045,N_7104,N_7721);
and U9046 (N_9046,N_6139,N_6113);
xnor U9047 (N_9047,N_7327,N_6251);
and U9048 (N_9048,N_7936,N_6637);
or U9049 (N_9049,N_6195,N_6048);
or U9050 (N_9050,N_6478,N_6066);
nand U9051 (N_9051,N_6160,N_6768);
and U9052 (N_9052,N_7978,N_7979);
nor U9053 (N_9053,N_6464,N_6209);
or U9054 (N_9054,N_7537,N_6797);
xnor U9055 (N_9055,N_6801,N_6982);
xor U9056 (N_9056,N_7930,N_6644);
and U9057 (N_9057,N_7541,N_6895);
and U9058 (N_9058,N_6813,N_7922);
nand U9059 (N_9059,N_6586,N_7317);
or U9060 (N_9060,N_7162,N_7838);
nor U9061 (N_9061,N_7451,N_7675);
and U9062 (N_9062,N_7104,N_7510);
nand U9063 (N_9063,N_7821,N_6129);
nor U9064 (N_9064,N_7312,N_7753);
xnor U9065 (N_9065,N_7978,N_6182);
nand U9066 (N_9066,N_6223,N_6410);
and U9067 (N_9067,N_6408,N_7134);
or U9068 (N_9068,N_7716,N_7984);
and U9069 (N_9069,N_6083,N_7586);
nand U9070 (N_9070,N_6989,N_6764);
and U9071 (N_9071,N_6569,N_6612);
nand U9072 (N_9072,N_7119,N_7287);
or U9073 (N_9073,N_7341,N_7241);
nand U9074 (N_9074,N_6118,N_7207);
xnor U9075 (N_9075,N_7861,N_7639);
nor U9076 (N_9076,N_7049,N_6753);
xnor U9077 (N_9077,N_6170,N_6254);
and U9078 (N_9078,N_6595,N_7606);
xor U9079 (N_9079,N_6529,N_6731);
nor U9080 (N_9080,N_7157,N_7827);
nor U9081 (N_9081,N_6439,N_6524);
nor U9082 (N_9082,N_6762,N_6118);
or U9083 (N_9083,N_7956,N_6075);
nor U9084 (N_9084,N_7120,N_6026);
nor U9085 (N_9085,N_6319,N_6064);
nor U9086 (N_9086,N_7046,N_6754);
xnor U9087 (N_9087,N_7195,N_6544);
nor U9088 (N_9088,N_6089,N_7401);
nor U9089 (N_9089,N_6358,N_7846);
nor U9090 (N_9090,N_6700,N_7343);
or U9091 (N_9091,N_7820,N_7489);
nor U9092 (N_9092,N_6262,N_6744);
nor U9093 (N_9093,N_6465,N_6878);
or U9094 (N_9094,N_6784,N_6357);
or U9095 (N_9095,N_6967,N_6526);
nor U9096 (N_9096,N_6727,N_6392);
or U9097 (N_9097,N_7067,N_7440);
nor U9098 (N_9098,N_7169,N_6626);
or U9099 (N_9099,N_7325,N_7465);
xnor U9100 (N_9100,N_6596,N_6419);
and U9101 (N_9101,N_7659,N_6456);
nand U9102 (N_9102,N_7025,N_7944);
nor U9103 (N_9103,N_6143,N_7672);
xor U9104 (N_9104,N_7141,N_7003);
and U9105 (N_9105,N_7084,N_6942);
nand U9106 (N_9106,N_7148,N_7448);
and U9107 (N_9107,N_7700,N_7500);
xnor U9108 (N_9108,N_6918,N_6739);
and U9109 (N_9109,N_6423,N_7881);
nand U9110 (N_9110,N_6952,N_6846);
nand U9111 (N_9111,N_6382,N_7550);
nor U9112 (N_9112,N_7124,N_7505);
nand U9113 (N_9113,N_6092,N_7801);
nor U9114 (N_9114,N_7051,N_6018);
xnor U9115 (N_9115,N_6060,N_7007);
or U9116 (N_9116,N_7632,N_6983);
nor U9117 (N_9117,N_7123,N_6522);
nor U9118 (N_9118,N_6419,N_6523);
or U9119 (N_9119,N_6572,N_6362);
or U9120 (N_9120,N_7260,N_6296);
nor U9121 (N_9121,N_6754,N_7958);
or U9122 (N_9122,N_6881,N_6560);
and U9123 (N_9123,N_6010,N_6005);
or U9124 (N_9124,N_7591,N_7794);
nand U9125 (N_9125,N_6190,N_6009);
nand U9126 (N_9126,N_6906,N_7136);
nor U9127 (N_9127,N_6891,N_6550);
nor U9128 (N_9128,N_6696,N_6200);
or U9129 (N_9129,N_6172,N_7567);
nor U9130 (N_9130,N_7652,N_7823);
and U9131 (N_9131,N_7554,N_7701);
xnor U9132 (N_9132,N_7644,N_7373);
nor U9133 (N_9133,N_6129,N_7930);
and U9134 (N_9134,N_7678,N_7941);
and U9135 (N_9135,N_7927,N_6241);
and U9136 (N_9136,N_6211,N_6907);
and U9137 (N_9137,N_7785,N_6069);
and U9138 (N_9138,N_7225,N_7934);
nor U9139 (N_9139,N_7315,N_6977);
xnor U9140 (N_9140,N_6182,N_6565);
nor U9141 (N_9141,N_6504,N_6985);
xor U9142 (N_9142,N_7878,N_7422);
nand U9143 (N_9143,N_7365,N_7693);
nor U9144 (N_9144,N_6344,N_7534);
or U9145 (N_9145,N_6869,N_6194);
xor U9146 (N_9146,N_7613,N_7247);
nor U9147 (N_9147,N_7249,N_7478);
or U9148 (N_9148,N_6389,N_7000);
nand U9149 (N_9149,N_7684,N_6445);
nand U9150 (N_9150,N_7742,N_7090);
nor U9151 (N_9151,N_7122,N_6515);
and U9152 (N_9152,N_7662,N_6194);
or U9153 (N_9153,N_7960,N_7343);
or U9154 (N_9154,N_6473,N_7391);
and U9155 (N_9155,N_7791,N_6263);
and U9156 (N_9156,N_6923,N_7006);
and U9157 (N_9157,N_6839,N_6668);
nand U9158 (N_9158,N_6046,N_6118);
nor U9159 (N_9159,N_7399,N_6293);
nor U9160 (N_9160,N_7432,N_6959);
nor U9161 (N_9161,N_6049,N_6466);
xnor U9162 (N_9162,N_6694,N_7603);
and U9163 (N_9163,N_7256,N_6303);
and U9164 (N_9164,N_7695,N_7542);
xor U9165 (N_9165,N_6134,N_6423);
xor U9166 (N_9166,N_7445,N_6380);
nand U9167 (N_9167,N_7026,N_7771);
nand U9168 (N_9168,N_6848,N_6674);
nand U9169 (N_9169,N_6618,N_6217);
xor U9170 (N_9170,N_6994,N_7716);
and U9171 (N_9171,N_7851,N_6059);
nor U9172 (N_9172,N_7211,N_7600);
and U9173 (N_9173,N_7130,N_7769);
or U9174 (N_9174,N_7660,N_6201);
nand U9175 (N_9175,N_6126,N_7652);
nand U9176 (N_9176,N_6178,N_6763);
nor U9177 (N_9177,N_6787,N_6864);
and U9178 (N_9178,N_7375,N_7126);
nand U9179 (N_9179,N_7538,N_6394);
nand U9180 (N_9180,N_6047,N_6349);
or U9181 (N_9181,N_7857,N_6859);
or U9182 (N_9182,N_6131,N_6146);
nor U9183 (N_9183,N_6276,N_6703);
or U9184 (N_9184,N_7478,N_7587);
or U9185 (N_9185,N_6451,N_7894);
and U9186 (N_9186,N_6523,N_7335);
nor U9187 (N_9187,N_6978,N_6089);
nor U9188 (N_9188,N_7994,N_7601);
nand U9189 (N_9189,N_7375,N_6097);
or U9190 (N_9190,N_7001,N_7088);
and U9191 (N_9191,N_7420,N_6480);
xor U9192 (N_9192,N_7222,N_6066);
nor U9193 (N_9193,N_7581,N_7351);
and U9194 (N_9194,N_7459,N_7223);
or U9195 (N_9195,N_6481,N_6488);
nor U9196 (N_9196,N_7460,N_7950);
nor U9197 (N_9197,N_6296,N_7366);
or U9198 (N_9198,N_6512,N_6975);
nor U9199 (N_9199,N_6256,N_7017);
or U9200 (N_9200,N_7080,N_6394);
and U9201 (N_9201,N_7904,N_7412);
and U9202 (N_9202,N_7838,N_7333);
or U9203 (N_9203,N_7764,N_6863);
and U9204 (N_9204,N_6381,N_6743);
or U9205 (N_9205,N_7299,N_6324);
nand U9206 (N_9206,N_6857,N_6089);
and U9207 (N_9207,N_6916,N_7787);
and U9208 (N_9208,N_7168,N_6253);
xnor U9209 (N_9209,N_6544,N_6255);
and U9210 (N_9210,N_6964,N_6428);
and U9211 (N_9211,N_7364,N_6659);
or U9212 (N_9212,N_6445,N_6363);
and U9213 (N_9213,N_6286,N_6225);
nand U9214 (N_9214,N_6363,N_6138);
and U9215 (N_9215,N_7344,N_7703);
or U9216 (N_9216,N_7107,N_6043);
xor U9217 (N_9217,N_7234,N_6793);
xor U9218 (N_9218,N_6101,N_7574);
xor U9219 (N_9219,N_6101,N_7596);
nor U9220 (N_9220,N_6541,N_7969);
or U9221 (N_9221,N_7847,N_7350);
or U9222 (N_9222,N_6148,N_6431);
and U9223 (N_9223,N_6185,N_7164);
xnor U9224 (N_9224,N_7106,N_7457);
and U9225 (N_9225,N_6183,N_7656);
nor U9226 (N_9226,N_6472,N_6265);
nor U9227 (N_9227,N_7702,N_7159);
nor U9228 (N_9228,N_7735,N_7846);
or U9229 (N_9229,N_6963,N_6278);
nor U9230 (N_9230,N_7443,N_7355);
xnor U9231 (N_9231,N_6877,N_7402);
or U9232 (N_9232,N_7939,N_6240);
nor U9233 (N_9233,N_7119,N_6345);
nand U9234 (N_9234,N_6605,N_7875);
or U9235 (N_9235,N_6751,N_6133);
or U9236 (N_9236,N_7694,N_7869);
and U9237 (N_9237,N_6209,N_6084);
nand U9238 (N_9238,N_6979,N_6977);
nand U9239 (N_9239,N_6568,N_7831);
nand U9240 (N_9240,N_7297,N_6552);
nand U9241 (N_9241,N_7965,N_7483);
or U9242 (N_9242,N_6841,N_6238);
and U9243 (N_9243,N_7305,N_7174);
and U9244 (N_9244,N_7010,N_6037);
or U9245 (N_9245,N_6791,N_7473);
and U9246 (N_9246,N_7186,N_7361);
nor U9247 (N_9247,N_7858,N_7055);
xor U9248 (N_9248,N_6259,N_7911);
nor U9249 (N_9249,N_6409,N_6627);
nand U9250 (N_9250,N_7674,N_7952);
nor U9251 (N_9251,N_7024,N_7450);
nand U9252 (N_9252,N_6272,N_7811);
nand U9253 (N_9253,N_7669,N_7499);
or U9254 (N_9254,N_7475,N_6988);
xor U9255 (N_9255,N_7507,N_7880);
or U9256 (N_9256,N_6323,N_6615);
nand U9257 (N_9257,N_6303,N_6365);
and U9258 (N_9258,N_6363,N_7218);
and U9259 (N_9259,N_7069,N_6174);
and U9260 (N_9260,N_6150,N_7947);
nand U9261 (N_9261,N_7914,N_7776);
nand U9262 (N_9262,N_7361,N_6987);
and U9263 (N_9263,N_6463,N_7774);
and U9264 (N_9264,N_7182,N_6734);
or U9265 (N_9265,N_7470,N_6174);
and U9266 (N_9266,N_6341,N_7499);
nor U9267 (N_9267,N_7934,N_7436);
nand U9268 (N_9268,N_7129,N_6671);
and U9269 (N_9269,N_6141,N_7747);
nand U9270 (N_9270,N_7269,N_6223);
and U9271 (N_9271,N_6400,N_6136);
nand U9272 (N_9272,N_7410,N_7723);
or U9273 (N_9273,N_7636,N_7580);
and U9274 (N_9274,N_6035,N_6864);
or U9275 (N_9275,N_6671,N_6233);
nand U9276 (N_9276,N_6878,N_6891);
or U9277 (N_9277,N_7928,N_6471);
xor U9278 (N_9278,N_7761,N_7471);
or U9279 (N_9279,N_7924,N_6673);
or U9280 (N_9280,N_6835,N_7892);
nor U9281 (N_9281,N_7506,N_6445);
nand U9282 (N_9282,N_7331,N_7446);
or U9283 (N_9283,N_7953,N_7897);
or U9284 (N_9284,N_6236,N_6482);
and U9285 (N_9285,N_7419,N_6133);
or U9286 (N_9286,N_7741,N_7274);
and U9287 (N_9287,N_7110,N_7685);
and U9288 (N_9288,N_6894,N_6789);
nor U9289 (N_9289,N_7017,N_6448);
nor U9290 (N_9290,N_6647,N_6891);
nor U9291 (N_9291,N_7558,N_7374);
and U9292 (N_9292,N_6777,N_7779);
nor U9293 (N_9293,N_7972,N_7347);
nor U9294 (N_9294,N_7957,N_6352);
or U9295 (N_9295,N_6045,N_7119);
or U9296 (N_9296,N_6415,N_6939);
nand U9297 (N_9297,N_7298,N_7570);
or U9298 (N_9298,N_7811,N_6406);
and U9299 (N_9299,N_7022,N_7734);
nor U9300 (N_9300,N_6282,N_6131);
or U9301 (N_9301,N_7156,N_6472);
nor U9302 (N_9302,N_6072,N_7425);
xnor U9303 (N_9303,N_6150,N_7408);
nand U9304 (N_9304,N_6417,N_6086);
and U9305 (N_9305,N_6211,N_6536);
nand U9306 (N_9306,N_6677,N_6760);
nand U9307 (N_9307,N_7147,N_7383);
or U9308 (N_9308,N_6300,N_7670);
and U9309 (N_9309,N_6865,N_6863);
and U9310 (N_9310,N_6405,N_6685);
nand U9311 (N_9311,N_7712,N_7881);
nor U9312 (N_9312,N_7977,N_6700);
or U9313 (N_9313,N_7073,N_7110);
and U9314 (N_9314,N_6803,N_6731);
or U9315 (N_9315,N_6674,N_7176);
or U9316 (N_9316,N_6168,N_6085);
and U9317 (N_9317,N_6393,N_6693);
nand U9318 (N_9318,N_6528,N_7705);
nand U9319 (N_9319,N_6670,N_7871);
or U9320 (N_9320,N_6933,N_7897);
xnor U9321 (N_9321,N_7739,N_7559);
or U9322 (N_9322,N_7911,N_7133);
nand U9323 (N_9323,N_7560,N_6080);
nand U9324 (N_9324,N_7335,N_7919);
and U9325 (N_9325,N_6636,N_7414);
nor U9326 (N_9326,N_7614,N_6363);
or U9327 (N_9327,N_6582,N_6631);
nor U9328 (N_9328,N_7500,N_6177);
or U9329 (N_9329,N_6960,N_7741);
nor U9330 (N_9330,N_6093,N_6146);
or U9331 (N_9331,N_6604,N_7408);
nor U9332 (N_9332,N_7027,N_7080);
xor U9333 (N_9333,N_6188,N_6977);
nor U9334 (N_9334,N_6850,N_7389);
or U9335 (N_9335,N_7741,N_6454);
or U9336 (N_9336,N_7009,N_6634);
nor U9337 (N_9337,N_7517,N_7145);
or U9338 (N_9338,N_7217,N_7515);
nor U9339 (N_9339,N_6829,N_6232);
nand U9340 (N_9340,N_6541,N_7445);
nor U9341 (N_9341,N_7018,N_6450);
nand U9342 (N_9342,N_7063,N_6996);
and U9343 (N_9343,N_7613,N_7992);
nor U9344 (N_9344,N_6139,N_7980);
nand U9345 (N_9345,N_7364,N_6987);
or U9346 (N_9346,N_6561,N_6623);
nand U9347 (N_9347,N_6254,N_7389);
or U9348 (N_9348,N_7725,N_7495);
nor U9349 (N_9349,N_7627,N_7472);
xnor U9350 (N_9350,N_7598,N_6140);
xnor U9351 (N_9351,N_6502,N_7384);
nand U9352 (N_9352,N_7432,N_7188);
and U9353 (N_9353,N_6972,N_7567);
nor U9354 (N_9354,N_6807,N_7000);
nand U9355 (N_9355,N_7275,N_7947);
and U9356 (N_9356,N_7913,N_6470);
nand U9357 (N_9357,N_7631,N_6201);
nand U9358 (N_9358,N_7578,N_7163);
nand U9359 (N_9359,N_7684,N_7178);
nor U9360 (N_9360,N_6031,N_7210);
nor U9361 (N_9361,N_6687,N_7033);
and U9362 (N_9362,N_7910,N_6726);
nand U9363 (N_9363,N_6588,N_7249);
and U9364 (N_9364,N_6486,N_7367);
or U9365 (N_9365,N_6117,N_6551);
or U9366 (N_9366,N_7212,N_6199);
nor U9367 (N_9367,N_6410,N_7054);
and U9368 (N_9368,N_6028,N_7681);
nand U9369 (N_9369,N_6642,N_6073);
and U9370 (N_9370,N_6808,N_7141);
nor U9371 (N_9371,N_6537,N_6090);
and U9372 (N_9372,N_6830,N_7010);
or U9373 (N_9373,N_7554,N_6487);
and U9374 (N_9374,N_6191,N_7666);
and U9375 (N_9375,N_7158,N_7392);
nand U9376 (N_9376,N_6860,N_7795);
and U9377 (N_9377,N_6305,N_7862);
or U9378 (N_9378,N_7773,N_6839);
nor U9379 (N_9379,N_7160,N_7197);
xnor U9380 (N_9380,N_6192,N_7446);
and U9381 (N_9381,N_7632,N_7866);
nor U9382 (N_9382,N_6047,N_6616);
nand U9383 (N_9383,N_7363,N_6875);
nor U9384 (N_9384,N_6168,N_6012);
nand U9385 (N_9385,N_7502,N_7672);
nor U9386 (N_9386,N_6705,N_6878);
and U9387 (N_9387,N_7528,N_7519);
nand U9388 (N_9388,N_6383,N_7008);
nand U9389 (N_9389,N_7605,N_6873);
nor U9390 (N_9390,N_7676,N_7820);
nand U9391 (N_9391,N_6532,N_6701);
nor U9392 (N_9392,N_6625,N_6766);
nor U9393 (N_9393,N_6316,N_7877);
nor U9394 (N_9394,N_6254,N_7543);
or U9395 (N_9395,N_6462,N_7684);
and U9396 (N_9396,N_7819,N_6897);
nor U9397 (N_9397,N_6197,N_7724);
and U9398 (N_9398,N_6637,N_6126);
and U9399 (N_9399,N_6109,N_7128);
and U9400 (N_9400,N_7860,N_7760);
and U9401 (N_9401,N_6574,N_6107);
nor U9402 (N_9402,N_7179,N_6298);
or U9403 (N_9403,N_7967,N_7558);
and U9404 (N_9404,N_7879,N_6671);
nand U9405 (N_9405,N_6089,N_6164);
xnor U9406 (N_9406,N_7366,N_6261);
nand U9407 (N_9407,N_7190,N_6185);
or U9408 (N_9408,N_6771,N_7812);
nand U9409 (N_9409,N_6185,N_7332);
nand U9410 (N_9410,N_6155,N_6829);
xnor U9411 (N_9411,N_6824,N_7651);
and U9412 (N_9412,N_6441,N_7310);
or U9413 (N_9413,N_7493,N_7103);
nor U9414 (N_9414,N_7014,N_7810);
or U9415 (N_9415,N_7636,N_7567);
and U9416 (N_9416,N_7103,N_7879);
nand U9417 (N_9417,N_7965,N_7655);
or U9418 (N_9418,N_7936,N_7035);
nand U9419 (N_9419,N_6822,N_7648);
nand U9420 (N_9420,N_7964,N_6193);
xnor U9421 (N_9421,N_7996,N_6240);
nor U9422 (N_9422,N_6734,N_6020);
xor U9423 (N_9423,N_7251,N_7825);
nand U9424 (N_9424,N_6187,N_6857);
and U9425 (N_9425,N_7943,N_7511);
and U9426 (N_9426,N_6878,N_7877);
nand U9427 (N_9427,N_6594,N_7208);
or U9428 (N_9428,N_6037,N_6179);
nand U9429 (N_9429,N_7265,N_7944);
and U9430 (N_9430,N_7312,N_6883);
nor U9431 (N_9431,N_6940,N_7023);
or U9432 (N_9432,N_7353,N_6615);
nand U9433 (N_9433,N_7763,N_6807);
nor U9434 (N_9434,N_7165,N_7878);
or U9435 (N_9435,N_7994,N_7048);
nor U9436 (N_9436,N_6591,N_6658);
nor U9437 (N_9437,N_6894,N_6980);
xor U9438 (N_9438,N_7761,N_7667);
and U9439 (N_9439,N_6761,N_6786);
nand U9440 (N_9440,N_6380,N_6506);
nor U9441 (N_9441,N_6899,N_7409);
nand U9442 (N_9442,N_6240,N_6660);
and U9443 (N_9443,N_7563,N_6567);
nand U9444 (N_9444,N_7815,N_6445);
nand U9445 (N_9445,N_6315,N_7620);
and U9446 (N_9446,N_7050,N_7523);
nor U9447 (N_9447,N_7408,N_6233);
nand U9448 (N_9448,N_6625,N_6006);
or U9449 (N_9449,N_6625,N_7342);
nor U9450 (N_9450,N_7622,N_7687);
and U9451 (N_9451,N_7856,N_6020);
or U9452 (N_9452,N_7880,N_6388);
xnor U9453 (N_9453,N_6951,N_6790);
nor U9454 (N_9454,N_6129,N_6385);
xor U9455 (N_9455,N_7834,N_6240);
and U9456 (N_9456,N_7673,N_6504);
or U9457 (N_9457,N_6725,N_7363);
or U9458 (N_9458,N_7560,N_6863);
xnor U9459 (N_9459,N_7866,N_7880);
nand U9460 (N_9460,N_7352,N_7223);
or U9461 (N_9461,N_7007,N_7040);
or U9462 (N_9462,N_7603,N_7520);
or U9463 (N_9463,N_7336,N_7230);
nor U9464 (N_9464,N_7101,N_7312);
nor U9465 (N_9465,N_7830,N_6349);
or U9466 (N_9466,N_6880,N_7326);
nand U9467 (N_9467,N_6340,N_7276);
nand U9468 (N_9468,N_7934,N_7524);
nor U9469 (N_9469,N_6390,N_6717);
xnor U9470 (N_9470,N_6551,N_6836);
nor U9471 (N_9471,N_6232,N_7207);
nand U9472 (N_9472,N_7753,N_7185);
nand U9473 (N_9473,N_6340,N_6841);
nor U9474 (N_9474,N_6158,N_7747);
and U9475 (N_9475,N_7755,N_7311);
or U9476 (N_9476,N_7284,N_7880);
nand U9477 (N_9477,N_7229,N_7099);
and U9478 (N_9478,N_6312,N_7345);
nor U9479 (N_9479,N_6073,N_7844);
and U9480 (N_9480,N_6252,N_7593);
nor U9481 (N_9481,N_7167,N_6317);
or U9482 (N_9482,N_6610,N_7177);
nor U9483 (N_9483,N_6352,N_6789);
nand U9484 (N_9484,N_7299,N_6568);
or U9485 (N_9485,N_6055,N_7028);
and U9486 (N_9486,N_6417,N_7130);
xnor U9487 (N_9487,N_7371,N_7040);
nand U9488 (N_9488,N_6795,N_6083);
nor U9489 (N_9489,N_6341,N_6554);
nand U9490 (N_9490,N_6225,N_7462);
or U9491 (N_9491,N_7717,N_7958);
nand U9492 (N_9492,N_7693,N_6292);
or U9493 (N_9493,N_7919,N_6868);
or U9494 (N_9494,N_7692,N_7953);
nor U9495 (N_9495,N_7454,N_7356);
nand U9496 (N_9496,N_7476,N_6130);
nand U9497 (N_9497,N_7012,N_6182);
xor U9498 (N_9498,N_6112,N_7711);
or U9499 (N_9499,N_6777,N_7430);
nand U9500 (N_9500,N_7537,N_7219);
or U9501 (N_9501,N_7513,N_7470);
nand U9502 (N_9502,N_7797,N_6391);
nor U9503 (N_9503,N_6729,N_7752);
and U9504 (N_9504,N_6048,N_6895);
nand U9505 (N_9505,N_7626,N_7285);
nor U9506 (N_9506,N_7996,N_7143);
and U9507 (N_9507,N_6486,N_6448);
or U9508 (N_9508,N_7781,N_6020);
and U9509 (N_9509,N_7372,N_6557);
and U9510 (N_9510,N_6469,N_7576);
and U9511 (N_9511,N_6301,N_6660);
or U9512 (N_9512,N_7342,N_6176);
or U9513 (N_9513,N_7634,N_7129);
and U9514 (N_9514,N_6595,N_6418);
nor U9515 (N_9515,N_7154,N_7996);
nor U9516 (N_9516,N_6776,N_6091);
or U9517 (N_9517,N_7195,N_6365);
or U9518 (N_9518,N_6944,N_6332);
or U9519 (N_9519,N_6023,N_6809);
nand U9520 (N_9520,N_6010,N_7535);
or U9521 (N_9521,N_6313,N_6463);
nand U9522 (N_9522,N_7431,N_7928);
and U9523 (N_9523,N_7269,N_7748);
or U9524 (N_9524,N_6866,N_7740);
and U9525 (N_9525,N_6775,N_6257);
xor U9526 (N_9526,N_7408,N_6479);
xnor U9527 (N_9527,N_7266,N_7937);
and U9528 (N_9528,N_7391,N_7264);
xnor U9529 (N_9529,N_7833,N_6190);
and U9530 (N_9530,N_7447,N_7616);
and U9531 (N_9531,N_7013,N_6721);
nor U9532 (N_9532,N_6242,N_6676);
nand U9533 (N_9533,N_7586,N_6795);
or U9534 (N_9534,N_6244,N_7956);
xor U9535 (N_9535,N_6509,N_7470);
or U9536 (N_9536,N_7793,N_7468);
nor U9537 (N_9537,N_7111,N_6378);
nor U9538 (N_9538,N_6604,N_6530);
or U9539 (N_9539,N_7627,N_6834);
nor U9540 (N_9540,N_7267,N_6434);
or U9541 (N_9541,N_7788,N_6668);
and U9542 (N_9542,N_7174,N_7916);
or U9543 (N_9543,N_6430,N_7920);
nor U9544 (N_9544,N_6483,N_7311);
or U9545 (N_9545,N_6208,N_6953);
nand U9546 (N_9546,N_6613,N_7217);
nand U9547 (N_9547,N_6920,N_6974);
or U9548 (N_9548,N_7891,N_6120);
or U9549 (N_9549,N_7751,N_6794);
or U9550 (N_9550,N_7266,N_7963);
nand U9551 (N_9551,N_6738,N_6944);
nor U9552 (N_9552,N_6001,N_7022);
nand U9553 (N_9553,N_6083,N_6335);
and U9554 (N_9554,N_6514,N_6877);
and U9555 (N_9555,N_7069,N_7103);
or U9556 (N_9556,N_6394,N_7595);
nor U9557 (N_9557,N_7953,N_7315);
and U9558 (N_9558,N_7182,N_6235);
or U9559 (N_9559,N_6168,N_7033);
nor U9560 (N_9560,N_6288,N_6525);
and U9561 (N_9561,N_6655,N_7476);
or U9562 (N_9562,N_7858,N_6312);
and U9563 (N_9563,N_7305,N_6559);
and U9564 (N_9564,N_6335,N_6791);
nor U9565 (N_9565,N_7929,N_7578);
and U9566 (N_9566,N_6953,N_6559);
xor U9567 (N_9567,N_6972,N_6433);
nand U9568 (N_9568,N_7159,N_6015);
xor U9569 (N_9569,N_6584,N_7608);
or U9570 (N_9570,N_7073,N_6819);
and U9571 (N_9571,N_7146,N_6727);
nand U9572 (N_9572,N_7555,N_6962);
nand U9573 (N_9573,N_6094,N_6488);
or U9574 (N_9574,N_6626,N_6672);
nor U9575 (N_9575,N_6399,N_6326);
and U9576 (N_9576,N_6322,N_6771);
and U9577 (N_9577,N_7624,N_7961);
and U9578 (N_9578,N_6358,N_6075);
nor U9579 (N_9579,N_6719,N_6692);
nor U9580 (N_9580,N_6519,N_7205);
nand U9581 (N_9581,N_7968,N_7681);
xor U9582 (N_9582,N_7054,N_7058);
and U9583 (N_9583,N_6411,N_7532);
nor U9584 (N_9584,N_6112,N_7434);
nor U9585 (N_9585,N_6280,N_7853);
nor U9586 (N_9586,N_7388,N_7805);
nor U9587 (N_9587,N_6678,N_6890);
nor U9588 (N_9588,N_7366,N_7211);
nor U9589 (N_9589,N_6440,N_6188);
and U9590 (N_9590,N_7702,N_6910);
xnor U9591 (N_9591,N_7367,N_6574);
nand U9592 (N_9592,N_6735,N_6163);
and U9593 (N_9593,N_7513,N_6219);
or U9594 (N_9594,N_7038,N_6243);
or U9595 (N_9595,N_6801,N_6278);
and U9596 (N_9596,N_7045,N_7507);
nor U9597 (N_9597,N_6268,N_7542);
and U9598 (N_9598,N_7928,N_7821);
xnor U9599 (N_9599,N_6833,N_6227);
or U9600 (N_9600,N_7983,N_6539);
nand U9601 (N_9601,N_7397,N_6596);
nor U9602 (N_9602,N_6974,N_6321);
nor U9603 (N_9603,N_7304,N_6605);
nand U9604 (N_9604,N_7191,N_7285);
nor U9605 (N_9605,N_7293,N_6807);
nor U9606 (N_9606,N_6142,N_7225);
and U9607 (N_9607,N_6317,N_7304);
or U9608 (N_9608,N_7848,N_7536);
nand U9609 (N_9609,N_6895,N_7017);
nor U9610 (N_9610,N_6631,N_6550);
and U9611 (N_9611,N_6311,N_7062);
or U9612 (N_9612,N_7626,N_6102);
and U9613 (N_9613,N_7711,N_7144);
nand U9614 (N_9614,N_7085,N_7793);
or U9615 (N_9615,N_7380,N_6525);
or U9616 (N_9616,N_7436,N_7875);
or U9617 (N_9617,N_7001,N_6201);
nand U9618 (N_9618,N_6244,N_7027);
and U9619 (N_9619,N_7975,N_6096);
or U9620 (N_9620,N_7158,N_6788);
or U9621 (N_9621,N_7254,N_7998);
and U9622 (N_9622,N_6063,N_6325);
nor U9623 (N_9623,N_7791,N_7920);
or U9624 (N_9624,N_7249,N_7668);
nor U9625 (N_9625,N_6570,N_6716);
nor U9626 (N_9626,N_6775,N_7883);
and U9627 (N_9627,N_6046,N_7721);
nor U9628 (N_9628,N_6731,N_6091);
and U9629 (N_9629,N_6473,N_6416);
and U9630 (N_9630,N_6595,N_7107);
and U9631 (N_9631,N_6530,N_7717);
nor U9632 (N_9632,N_6791,N_6660);
nor U9633 (N_9633,N_7529,N_6820);
nor U9634 (N_9634,N_7449,N_7928);
nand U9635 (N_9635,N_6939,N_6468);
or U9636 (N_9636,N_7481,N_6773);
or U9637 (N_9637,N_7080,N_7975);
xor U9638 (N_9638,N_6929,N_6473);
nor U9639 (N_9639,N_6642,N_7395);
or U9640 (N_9640,N_7997,N_6625);
nand U9641 (N_9641,N_6486,N_7662);
nor U9642 (N_9642,N_6581,N_7606);
nand U9643 (N_9643,N_7473,N_7225);
or U9644 (N_9644,N_6067,N_6478);
or U9645 (N_9645,N_7576,N_6617);
or U9646 (N_9646,N_6241,N_6735);
or U9647 (N_9647,N_6365,N_7761);
and U9648 (N_9648,N_7228,N_7355);
xnor U9649 (N_9649,N_7232,N_6461);
or U9650 (N_9650,N_6171,N_6663);
xor U9651 (N_9651,N_7795,N_6618);
or U9652 (N_9652,N_6956,N_7708);
nand U9653 (N_9653,N_7843,N_6265);
nand U9654 (N_9654,N_6021,N_7958);
nor U9655 (N_9655,N_7875,N_6813);
or U9656 (N_9656,N_6476,N_6926);
nor U9657 (N_9657,N_6077,N_7936);
nand U9658 (N_9658,N_7220,N_7816);
nand U9659 (N_9659,N_7757,N_7854);
xnor U9660 (N_9660,N_6414,N_6929);
nand U9661 (N_9661,N_7324,N_7839);
or U9662 (N_9662,N_7303,N_6174);
xnor U9663 (N_9663,N_7179,N_7322);
nor U9664 (N_9664,N_7955,N_6641);
nor U9665 (N_9665,N_6276,N_7907);
and U9666 (N_9666,N_7210,N_6617);
nor U9667 (N_9667,N_7087,N_7237);
and U9668 (N_9668,N_6905,N_7882);
and U9669 (N_9669,N_7206,N_6426);
nand U9670 (N_9670,N_7091,N_7083);
or U9671 (N_9671,N_6226,N_7146);
and U9672 (N_9672,N_6556,N_6794);
or U9673 (N_9673,N_6263,N_6790);
and U9674 (N_9674,N_7188,N_6002);
nand U9675 (N_9675,N_7652,N_7495);
or U9676 (N_9676,N_6906,N_6968);
and U9677 (N_9677,N_6744,N_6748);
and U9678 (N_9678,N_7224,N_6522);
and U9679 (N_9679,N_6788,N_6590);
or U9680 (N_9680,N_7837,N_7204);
and U9681 (N_9681,N_6346,N_6134);
or U9682 (N_9682,N_7837,N_7783);
nand U9683 (N_9683,N_6135,N_7054);
and U9684 (N_9684,N_6935,N_6073);
nor U9685 (N_9685,N_7340,N_6943);
or U9686 (N_9686,N_6397,N_7349);
nor U9687 (N_9687,N_6523,N_6469);
nand U9688 (N_9688,N_6954,N_6950);
nor U9689 (N_9689,N_6196,N_6789);
and U9690 (N_9690,N_7922,N_7929);
and U9691 (N_9691,N_7346,N_6351);
or U9692 (N_9692,N_7707,N_7582);
nand U9693 (N_9693,N_7617,N_6786);
nand U9694 (N_9694,N_6162,N_6182);
nand U9695 (N_9695,N_7250,N_6079);
nand U9696 (N_9696,N_6379,N_6356);
nor U9697 (N_9697,N_7040,N_6366);
nand U9698 (N_9698,N_6202,N_6028);
nor U9699 (N_9699,N_7883,N_7733);
nand U9700 (N_9700,N_6997,N_7471);
and U9701 (N_9701,N_6270,N_7851);
or U9702 (N_9702,N_6871,N_7499);
nand U9703 (N_9703,N_7567,N_7791);
nand U9704 (N_9704,N_6728,N_7640);
and U9705 (N_9705,N_6431,N_6668);
or U9706 (N_9706,N_6919,N_7957);
nand U9707 (N_9707,N_6178,N_6412);
xor U9708 (N_9708,N_6294,N_7598);
nand U9709 (N_9709,N_6403,N_7708);
nand U9710 (N_9710,N_7613,N_7357);
or U9711 (N_9711,N_6134,N_7259);
nor U9712 (N_9712,N_7736,N_6554);
or U9713 (N_9713,N_6013,N_7833);
nor U9714 (N_9714,N_7005,N_6569);
nor U9715 (N_9715,N_6522,N_6699);
nand U9716 (N_9716,N_7716,N_7558);
nor U9717 (N_9717,N_6438,N_7591);
and U9718 (N_9718,N_7190,N_6560);
or U9719 (N_9719,N_6012,N_7336);
nand U9720 (N_9720,N_6617,N_7443);
nand U9721 (N_9721,N_6977,N_6410);
or U9722 (N_9722,N_6073,N_7891);
nor U9723 (N_9723,N_7360,N_7105);
and U9724 (N_9724,N_7009,N_7041);
nand U9725 (N_9725,N_7147,N_7668);
nor U9726 (N_9726,N_7607,N_7388);
nor U9727 (N_9727,N_7296,N_7631);
nor U9728 (N_9728,N_7507,N_6455);
and U9729 (N_9729,N_7547,N_7554);
and U9730 (N_9730,N_6869,N_6523);
or U9731 (N_9731,N_7295,N_7856);
xor U9732 (N_9732,N_6813,N_6574);
or U9733 (N_9733,N_6532,N_6156);
nand U9734 (N_9734,N_7305,N_6401);
nor U9735 (N_9735,N_6562,N_7845);
xor U9736 (N_9736,N_7284,N_6254);
nand U9737 (N_9737,N_7957,N_7286);
nand U9738 (N_9738,N_7421,N_7168);
or U9739 (N_9739,N_7573,N_6196);
nor U9740 (N_9740,N_7158,N_6698);
nor U9741 (N_9741,N_7391,N_6106);
nand U9742 (N_9742,N_6475,N_7159);
nand U9743 (N_9743,N_6824,N_6604);
or U9744 (N_9744,N_7872,N_7685);
nor U9745 (N_9745,N_7996,N_6258);
or U9746 (N_9746,N_7163,N_7434);
and U9747 (N_9747,N_6809,N_7184);
or U9748 (N_9748,N_7970,N_6203);
nand U9749 (N_9749,N_6840,N_7702);
and U9750 (N_9750,N_7824,N_6070);
nor U9751 (N_9751,N_7911,N_7976);
nor U9752 (N_9752,N_7528,N_7379);
nand U9753 (N_9753,N_6042,N_7760);
or U9754 (N_9754,N_7615,N_7616);
or U9755 (N_9755,N_7342,N_7971);
or U9756 (N_9756,N_6486,N_7359);
nor U9757 (N_9757,N_6137,N_7779);
nand U9758 (N_9758,N_6821,N_6928);
xnor U9759 (N_9759,N_7952,N_6977);
nor U9760 (N_9760,N_7221,N_7298);
and U9761 (N_9761,N_6725,N_6396);
nand U9762 (N_9762,N_6004,N_7284);
nand U9763 (N_9763,N_6445,N_6849);
and U9764 (N_9764,N_6921,N_7687);
and U9765 (N_9765,N_7601,N_6576);
nand U9766 (N_9766,N_6318,N_7332);
nand U9767 (N_9767,N_7869,N_7383);
and U9768 (N_9768,N_6668,N_6503);
nor U9769 (N_9769,N_7803,N_7371);
or U9770 (N_9770,N_7194,N_7255);
or U9771 (N_9771,N_6460,N_7669);
nor U9772 (N_9772,N_7136,N_6712);
nor U9773 (N_9773,N_7036,N_6924);
xnor U9774 (N_9774,N_6291,N_6372);
nor U9775 (N_9775,N_7630,N_7914);
nor U9776 (N_9776,N_6938,N_7283);
and U9777 (N_9777,N_7790,N_7835);
and U9778 (N_9778,N_7707,N_7528);
and U9779 (N_9779,N_6410,N_6979);
and U9780 (N_9780,N_7732,N_7210);
nand U9781 (N_9781,N_6669,N_7980);
or U9782 (N_9782,N_6490,N_7565);
and U9783 (N_9783,N_6917,N_6083);
nor U9784 (N_9784,N_6790,N_7269);
and U9785 (N_9785,N_7885,N_7927);
and U9786 (N_9786,N_7043,N_6567);
nor U9787 (N_9787,N_7711,N_6959);
nand U9788 (N_9788,N_6387,N_7999);
and U9789 (N_9789,N_7343,N_7783);
or U9790 (N_9790,N_6777,N_6621);
and U9791 (N_9791,N_6767,N_7214);
nor U9792 (N_9792,N_7816,N_7360);
and U9793 (N_9793,N_6073,N_6400);
nor U9794 (N_9794,N_6505,N_7964);
nor U9795 (N_9795,N_7058,N_6504);
or U9796 (N_9796,N_7187,N_7728);
or U9797 (N_9797,N_7781,N_7152);
or U9798 (N_9798,N_7512,N_7074);
xor U9799 (N_9799,N_7122,N_6866);
xor U9800 (N_9800,N_7795,N_6990);
xnor U9801 (N_9801,N_7670,N_7945);
xor U9802 (N_9802,N_7281,N_7868);
xnor U9803 (N_9803,N_7939,N_7841);
and U9804 (N_9804,N_6975,N_6467);
nor U9805 (N_9805,N_6071,N_6728);
or U9806 (N_9806,N_7449,N_6121);
and U9807 (N_9807,N_6483,N_6169);
xnor U9808 (N_9808,N_7081,N_7239);
or U9809 (N_9809,N_7077,N_6492);
nand U9810 (N_9810,N_7779,N_6865);
nand U9811 (N_9811,N_6233,N_7701);
xor U9812 (N_9812,N_7550,N_7676);
and U9813 (N_9813,N_6904,N_7968);
xnor U9814 (N_9814,N_7656,N_7890);
nor U9815 (N_9815,N_7887,N_6075);
xor U9816 (N_9816,N_7011,N_7941);
nand U9817 (N_9817,N_6884,N_7416);
or U9818 (N_9818,N_6204,N_6833);
xor U9819 (N_9819,N_7195,N_6703);
nand U9820 (N_9820,N_6044,N_6964);
nor U9821 (N_9821,N_7473,N_7682);
and U9822 (N_9822,N_7990,N_7167);
and U9823 (N_9823,N_6689,N_6203);
nor U9824 (N_9824,N_7676,N_6087);
nor U9825 (N_9825,N_7956,N_7448);
or U9826 (N_9826,N_6032,N_6850);
or U9827 (N_9827,N_7096,N_7580);
and U9828 (N_9828,N_6105,N_6571);
nor U9829 (N_9829,N_7742,N_7661);
nand U9830 (N_9830,N_7439,N_6159);
nand U9831 (N_9831,N_6317,N_6588);
and U9832 (N_9832,N_6823,N_7045);
and U9833 (N_9833,N_7267,N_6406);
nand U9834 (N_9834,N_7185,N_6351);
or U9835 (N_9835,N_6087,N_6286);
nand U9836 (N_9836,N_6823,N_7452);
nand U9837 (N_9837,N_7955,N_6847);
and U9838 (N_9838,N_6012,N_6717);
and U9839 (N_9839,N_7102,N_6545);
nand U9840 (N_9840,N_6304,N_6399);
nand U9841 (N_9841,N_7905,N_7669);
and U9842 (N_9842,N_6303,N_6761);
nand U9843 (N_9843,N_7489,N_7948);
and U9844 (N_9844,N_7615,N_6328);
xor U9845 (N_9845,N_6763,N_6275);
nor U9846 (N_9846,N_6226,N_6126);
nor U9847 (N_9847,N_6372,N_6547);
nand U9848 (N_9848,N_7007,N_6709);
nor U9849 (N_9849,N_7465,N_7330);
nor U9850 (N_9850,N_6474,N_6937);
nor U9851 (N_9851,N_7880,N_7941);
or U9852 (N_9852,N_7725,N_6349);
nor U9853 (N_9853,N_6747,N_7494);
or U9854 (N_9854,N_7178,N_7185);
nand U9855 (N_9855,N_7405,N_6707);
or U9856 (N_9856,N_7360,N_7162);
nor U9857 (N_9857,N_7884,N_7353);
or U9858 (N_9858,N_7675,N_6122);
and U9859 (N_9859,N_7111,N_6138);
nand U9860 (N_9860,N_7405,N_6629);
and U9861 (N_9861,N_6434,N_7824);
or U9862 (N_9862,N_7295,N_7814);
and U9863 (N_9863,N_7776,N_6302);
nor U9864 (N_9864,N_7631,N_7871);
or U9865 (N_9865,N_7331,N_7945);
nor U9866 (N_9866,N_6154,N_7996);
nor U9867 (N_9867,N_6836,N_7711);
xnor U9868 (N_9868,N_7161,N_7693);
nor U9869 (N_9869,N_6682,N_7909);
xnor U9870 (N_9870,N_6937,N_7271);
nand U9871 (N_9871,N_6386,N_6743);
and U9872 (N_9872,N_7425,N_7804);
nand U9873 (N_9873,N_7840,N_6756);
nor U9874 (N_9874,N_6547,N_6570);
xnor U9875 (N_9875,N_7758,N_6758);
nand U9876 (N_9876,N_7821,N_7280);
or U9877 (N_9877,N_6231,N_7035);
and U9878 (N_9878,N_6612,N_7122);
or U9879 (N_9879,N_6197,N_7013);
and U9880 (N_9880,N_7248,N_6331);
nor U9881 (N_9881,N_6719,N_7075);
nand U9882 (N_9882,N_7052,N_6183);
or U9883 (N_9883,N_7602,N_6159);
and U9884 (N_9884,N_7888,N_6338);
and U9885 (N_9885,N_6180,N_7591);
and U9886 (N_9886,N_7371,N_6045);
nand U9887 (N_9887,N_6839,N_7877);
nand U9888 (N_9888,N_6406,N_7581);
nor U9889 (N_9889,N_6238,N_7989);
nand U9890 (N_9890,N_7902,N_7288);
or U9891 (N_9891,N_6927,N_7491);
nor U9892 (N_9892,N_7528,N_7608);
xnor U9893 (N_9893,N_6270,N_7959);
nand U9894 (N_9894,N_6944,N_7641);
nor U9895 (N_9895,N_6032,N_7434);
and U9896 (N_9896,N_6109,N_6565);
nor U9897 (N_9897,N_7175,N_7119);
xor U9898 (N_9898,N_7767,N_6888);
or U9899 (N_9899,N_6896,N_7618);
and U9900 (N_9900,N_7545,N_6529);
nand U9901 (N_9901,N_7030,N_7848);
and U9902 (N_9902,N_6363,N_6303);
or U9903 (N_9903,N_7266,N_7073);
nor U9904 (N_9904,N_7147,N_7409);
or U9905 (N_9905,N_6844,N_7073);
nand U9906 (N_9906,N_7732,N_6915);
nand U9907 (N_9907,N_6963,N_7232);
nand U9908 (N_9908,N_6582,N_6976);
and U9909 (N_9909,N_6831,N_6451);
nor U9910 (N_9910,N_7929,N_6734);
or U9911 (N_9911,N_7156,N_6505);
nor U9912 (N_9912,N_6315,N_6697);
or U9913 (N_9913,N_7036,N_7662);
and U9914 (N_9914,N_6801,N_7697);
and U9915 (N_9915,N_6360,N_7084);
or U9916 (N_9916,N_6798,N_7710);
nor U9917 (N_9917,N_6175,N_6135);
and U9918 (N_9918,N_6019,N_7982);
nor U9919 (N_9919,N_7958,N_6795);
or U9920 (N_9920,N_7295,N_6494);
nand U9921 (N_9921,N_6882,N_6288);
nand U9922 (N_9922,N_7723,N_7264);
and U9923 (N_9923,N_7892,N_6514);
xor U9924 (N_9924,N_7062,N_7984);
or U9925 (N_9925,N_7610,N_6484);
or U9926 (N_9926,N_7829,N_7728);
and U9927 (N_9927,N_6613,N_6807);
xor U9928 (N_9928,N_6590,N_7716);
xor U9929 (N_9929,N_6197,N_7831);
or U9930 (N_9930,N_7025,N_6294);
nor U9931 (N_9931,N_7532,N_6146);
nor U9932 (N_9932,N_7903,N_6718);
or U9933 (N_9933,N_7880,N_6834);
or U9934 (N_9934,N_7498,N_7515);
and U9935 (N_9935,N_7277,N_6106);
nor U9936 (N_9936,N_6952,N_7764);
xnor U9937 (N_9937,N_7044,N_6062);
nand U9938 (N_9938,N_6386,N_7919);
nand U9939 (N_9939,N_7066,N_6192);
or U9940 (N_9940,N_6388,N_6516);
or U9941 (N_9941,N_6331,N_6904);
nand U9942 (N_9942,N_7783,N_6576);
nand U9943 (N_9943,N_7258,N_6797);
and U9944 (N_9944,N_7635,N_7859);
nor U9945 (N_9945,N_6100,N_7282);
nand U9946 (N_9946,N_7260,N_7637);
nor U9947 (N_9947,N_7251,N_6497);
nor U9948 (N_9948,N_6332,N_6353);
xnor U9949 (N_9949,N_6912,N_6002);
nand U9950 (N_9950,N_6003,N_6932);
and U9951 (N_9951,N_7897,N_6465);
or U9952 (N_9952,N_6606,N_6096);
or U9953 (N_9953,N_7599,N_7961);
and U9954 (N_9954,N_7021,N_7809);
and U9955 (N_9955,N_6651,N_7455);
nand U9956 (N_9956,N_6124,N_6064);
xnor U9957 (N_9957,N_7854,N_6375);
and U9958 (N_9958,N_7520,N_6105);
xnor U9959 (N_9959,N_7847,N_6382);
nor U9960 (N_9960,N_6747,N_6703);
nor U9961 (N_9961,N_6693,N_6564);
and U9962 (N_9962,N_6122,N_6697);
nor U9963 (N_9963,N_7179,N_7355);
nor U9964 (N_9964,N_7194,N_7382);
nand U9965 (N_9965,N_6645,N_7561);
or U9966 (N_9966,N_6282,N_6341);
nor U9967 (N_9967,N_6039,N_7452);
or U9968 (N_9968,N_7136,N_7818);
nor U9969 (N_9969,N_6925,N_6521);
and U9970 (N_9970,N_7985,N_6242);
and U9971 (N_9971,N_6414,N_6469);
nand U9972 (N_9972,N_7262,N_6113);
and U9973 (N_9973,N_6595,N_7045);
nor U9974 (N_9974,N_6366,N_6363);
nor U9975 (N_9975,N_6687,N_7228);
and U9976 (N_9976,N_7837,N_7189);
nor U9977 (N_9977,N_7154,N_6671);
or U9978 (N_9978,N_6090,N_7066);
and U9979 (N_9979,N_7425,N_7432);
or U9980 (N_9980,N_7553,N_7277);
nand U9981 (N_9981,N_6925,N_6353);
and U9982 (N_9982,N_7676,N_7995);
nand U9983 (N_9983,N_7686,N_6021);
nor U9984 (N_9984,N_6250,N_7037);
nand U9985 (N_9985,N_6876,N_6009);
and U9986 (N_9986,N_7934,N_6179);
or U9987 (N_9987,N_6815,N_7302);
nand U9988 (N_9988,N_6346,N_6276);
xor U9989 (N_9989,N_6861,N_7153);
nor U9990 (N_9990,N_7997,N_7250);
nor U9991 (N_9991,N_7021,N_6981);
nor U9992 (N_9992,N_7448,N_6153);
xor U9993 (N_9993,N_6258,N_7079);
nor U9994 (N_9994,N_6798,N_6590);
nand U9995 (N_9995,N_6586,N_6663);
nand U9996 (N_9996,N_7754,N_7808);
nand U9997 (N_9997,N_7493,N_7407);
and U9998 (N_9998,N_6888,N_7393);
nor U9999 (N_9999,N_6082,N_6242);
nand UO_0 (O_0,N_9660,N_8610);
or UO_1 (O_1,N_8978,N_8233);
nand UO_2 (O_2,N_8885,N_8814);
nor UO_3 (O_3,N_8264,N_8111);
and UO_4 (O_4,N_9415,N_9589);
nor UO_5 (O_5,N_8927,N_9853);
nor UO_6 (O_6,N_9259,N_8381);
nand UO_7 (O_7,N_9898,N_9904);
nor UO_8 (O_8,N_9127,N_8991);
nand UO_9 (O_9,N_8118,N_9646);
or UO_10 (O_10,N_8598,N_9843);
nor UO_11 (O_11,N_9522,N_8386);
or UO_12 (O_12,N_9205,N_9171);
or UO_13 (O_13,N_9573,N_9854);
xnor UO_14 (O_14,N_9796,N_8435);
nand UO_15 (O_15,N_9349,N_9738);
nand UO_16 (O_16,N_9971,N_8252);
or UO_17 (O_17,N_8887,N_8599);
or UO_18 (O_18,N_9094,N_9727);
nand UO_19 (O_19,N_8045,N_9679);
nand UO_20 (O_20,N_9298,N_9504);
or UO_21 (O_21,N_9980,N_9383);
nand UO_22 (O_22,N_9154,N_8857);
or UO_23 (O_23,N_8635,N_8519);
nand UO_24 (O_24,N_8745,N_9882);
or UO_25 (O_25,N_9635,N_9661);
nor UO_26 (O_26,N_9215,N_9655);
nor UO_27 (O_27,N_9217,N_9461);
nand UO_28 (O_28,N_9150,N_9799);
nand UO_29 (O_29,N_9224,N_8260);
and UO_30 (O_30,N_9236,N_8654);
or UO_31 (O_31,N_9385,N_9793);
nand UO_32 (O_32,N_8698,N_8685);
nand UO_33 (O_33,N_9990,N_8113);
xnor UO_34 (O_34,N_9359,N_8426);
nor UO_35 (O_35,N_9707,N_8601);
and UO_36 (O_36,N_8957,N_8695);
and UO_37 (O_37,N_8505,N_8646);
nand UO_38 (O_38,N_9396,N_8358);
and UO_39 (O_39,N_9252,N_8979);
or UO_40 (O_40,N_9828,N_8712);
nor UO_41 (O_41,N_9703,N_8275);
and UO_42 (O_42,N_8158,N_9795);
or UO_43 (O_43,N_8127,N_9879);
xnor UO_44 (O_44,N_9204,N_9960);
and UO_45 (O_45,N_8869,N_9474);
and UO_46 (O_46,N_9031,N_9947);
nor UO_47 (O_47,N_9388,N_8813);
or UO_48 (O_48,N_9005,N_8382);
and UO_49 (O_49,N_8987,N_8247);
or UO_50 (O_50,N_8152,N_9603);
nor UO_51 (O_51,N_8457,N_9791);
and UO_52 (O_52,N_9077,N_8861);
and UO_53 (O_53,N_8076,N_8427);
nor UO_54 (O_54,N_8681,N_9059);
and UO_55 (O_55,N_8863,N_9979);
nand UO_56 (O_56,N_8733,N_8054);
or UO_57 (O_57,N_8725,N_9626);
or UO_58 (O_58,N_8672,N_8121);
and UO_59 (O_59,N_8996,N_9440);
nand UO_60 (O_60,N_8257,N_9051);
or UO_61 (O_61,N_8784,N_8575);
or UO_62 (O_62,N_9157,N_9138);
nor UO_63 (O_63,N_8557,N_8272);
nand UO_64 (O_64,N_8824,N_9426);
nor UO_65 (O_65,N_9446,N_9423);
nand UO_66 (O_66,N_8067,N_9472);
nand UO_67 (O_67,N_9621,N_9049);
and UO_68 (O_68,N_9118,N_8682);
and UO_69 (O_69,N_9546,N_9739);
and UO_70 (O_70,N_9060,N_8029);
and UO_71 (O_71,N_8298,N_9299);
or UO_72 (O_72,N_9038,N_8715);
and UO_73 (O_73,N_8096,N_9903);
xnor UO_74 (O_74,N_8550,N_9514);
nand UO_75 (O_75,N_9111,N_8460);
nor UO_76 (O_76,N_9945,N_9834);
xor UO_77 (O_77,N_9257,N_8352);
nand UO_78 (O_78,N_9761,N_8514);
nand UO_79 (O_79,N_9940,N_9024);
nand UO_80 (O_80,N_9705,N_8923);
nor UO_81 (O_81,N_8953,N_9641);
nand UO_82 (O_82,N_9774,N_8888);
or UO_83 (O_83,N_9428,N_9827);
and UO_84 (O_84,N_9235,N_8277);
or UO_85 (O_85,N_9061,N_9722);
and UO_86 (O_86,N_9422,N_8830);
or UO_87 (O_87,N_9872,N_9473);
nand UO_88 (O_88,N_9672,N_8976);
and UO_89 (O_89,N_8584,N_9728);
or UO_90 (O_90,N_9680,N_9069);
nor UO_91 (O_91,N_9441,N_8545);
xnor UO_92 (O_92,N_8244,N_8699);
and UO_93 (O_93,N_9921,N_8818);
xnor UO_94 (O_94,N_8801,N_8994);
nand UO_95 (O_95,N_8150,N_8255);
nand UO_96 (O_96,N_9911,N_9460);
nor UO_97 (O_97,N_8693,N_9377);
nand UO_98 (O_98,N_8135,N_8259);
and UO_99 (O_99,N_8479,N_8161);
and UO_100 (O_100,N_8778,N_8491);
nand UO_101 (O_101,N_8049,N_9895);
and UO_102 (O_102,N_8729,N_8042);
nor UO_103 (O_103,N_8637,N_8517);
nor UO_104 (O_104,N_8821,N_9730);
nor UO_105 (O_105,N_9407,N_8612);
xnor UO_106 (O_106,N_9449,N_8536);
xnor UO_107 (O_107,N_9245,N_8562);
or UO_108 (O_108,N_9699,N_9319);
and UO_109 (O_109,N_9518,N_9390);
nor UO_110 (O_110,N_9307,N_9140);
and UO_111 (O_111,N_8163,N_8677);
and UO_112 (O_112,N_8675,N_8325);
nor UO_113 (O_113,N_8942,N_8773);
xnor UO_114 (O_114,N_9066,N_9109);
or UO_115 (O_115,N_9794,N_9134);
and UO_116 (O_116,N_8347,N_8825);
nor UO_117 (O_117,N_8577,N_8844);
or UO_118 (O_118,N_9719,N_8159);
and UO_119 (O_119,N_8608,N_9885);
nor UO_120 (O_120,N_8555,N_8753);
or UO_121 (O_121,N_8180,N_8828);
nand UO_122 (O_122,N_8965,N_9075);
nor UO_123 (O_123,N_8787,N_9177);
or UO_124 (O_124,N_8003,N_9628);
or UO_125 (O_125,N_9825,N_9226);
or UO_126 (O_126,N_8777,N_8452);
nand UO_127 (O_127,N_8518,N_8756);
nand UO_128 (O_128,N_8134,N_8687);
nand UO_129 (O_129,N_8549,N_9468);
and UO_130 (O_130,N_8649,N_9042);
and UO_131 (O_131,N_8768,N_9478);
or UO_132 (O_132,N_9491,N_8438);
xor UO_133 (O_133,N_8890,N_8930);
nand UO_134 (O_134,N_8807,N_8786);
and UO_135 (O_135,N_9139,N_9720);
and UO_136 (O_136,N_9992,N_8061);
nor UO_137 (O_137,N_9330,N_9922);
and UO_138 (O_138,N_9736,N_8702);
or UO_139 (O_139,N_8270,N_9327);
and UO_140 (O_140,N_9925,N_8251);
nand UO_141 (O_141,N_9512,N_8243);
nand UO_142 (O_142,N_8176,N_9718);
nor UO_143 (O_143,N_8077,N_8609);
nor UO_144 (O_144,N_8546,N_9143);
nand UO_145 (O_145,N_9897,N_8789);
nand UO_146 (O_146,N_9408,N_8868);
and UO_147 (O_147,N_8525,N_8164);
nor UO_148 (O_148,N_9497,N_8040);
or UO_149 (O_149,N_8922,N_9588);
nand UO_150 (O_150,N_8443,N_8908);
and UO_151 (O_151,N_8153,N_8975);
nor UO_152 (O_152,N_9309,N_9191);
or UO_153 (O_153,N_9886,N_8969);
nand UO_154 (O_154,N_8719,N_8862);
and UO_155 (O_155,N_8019,N_8220);
nand UO_156 (O_156,N_9822,N_9312);
nand UO_157 (O_157,N_9684,N_9759);
and UO_158 (O_158,N_9433,N_9037);
or UO_159 (O_159,N_9905,N_8538);
or UO_160 (O_160,N_9866,N_8423);
or UO_161 (O_161,N_8980,N_8574);
xnor UO_162 (O_162,N_9490,N_8737);
and UO_163 (O_163,N_9214,N_8785);
nor UO_164 (O_164,N_8075,N_9450);
nand UO_165 (O_165,N_9097,N_9760);
or UO_166 (O_166,N_9344,N_9938);
nand UO_167 (O_167,N_8805,N_9606);
and UO_168 (O_168,N_8871,N_9733);
and UO_169 (O_169,N_9342,N_9618);
xnor UO_170 (O_170,N_8916,N_8847);
or UO_171 (O_171,N_9486,N_8812);
nor UO_172 (O_172,N_9852,N_9405);
or UO_173 (O_173,N_8177,N_9009);
and UO_174 (O_174,N_8642,N_9179);
and UO_175 (O_175,N_8455,N_8703);
nor UO_176 (O_176,N_9923,N_9465);
nor UO_177 (O_177,N_9090,N_9984);
or UO_178 (O_178,N_9740,N_9447);
nand UO_179 (O_179,N_9308,N_8328);
and UO_180 (O_180,N_9250,N_9570);
nor UO_181 (O_181,N_8816,N_8605);
xor UO_182 (O_182,N_9837,N_9642);
nand UO_183 (O_183,N_8676,N_9275);
and UO_184 (O_184,N_9329,N_8900);
nand UO_185 (O_185,N_8216,N_8659);
nor UO_186 (O_186,N_9393,N_8701);
nor UO_187 (O_187,N_9244,N_8242);
nand UO_188 (O_188,N_8214,N_9994);
or UO_189 (O_189,N_9578,N_9741);
or UO_190 (O_190,N_8302,N_9597);
xnor UO_191 (O_191,N_8665,N_9399);
and UO_192 (O_192,N_9434,N_9001);
and UO_193 (O_193,N_8779,N_8143);
and UO_194 (O_194,N_8442,N_9869);
and UO_195 (O_195,N_8454,N_8615);
and UO_196 (O_196,N_8149,N_8776);
and UO_197 (O_197,N_8235,N_8772);
and UO_198 (O_198,N_9961,N_9747);
or UO_199 (O_199,N_8058,N_9333);
nand UO_200 (O_200,N_8578,N_8507);
nand UO_201 (O_201,N_9510,N_8241);
nand UO_202 (O_202,N_9262,N_9239);
nand UO_203 (O_203,N_8833,N_9829);
or UO_204 (O_204,N_8450,N_9850);
nor UO_205 (O_205,N_9056,N_9046);
nor UO_206 (O_206,N_9786,N_9779);
xnor UO_207 (O_207,N_9632,N_8846);
and UO_208 (O_208,N_9706,N_8469);
xor UO_209 (O_209,N_8395,N_9755);
and UO_210 (O_210,N_8799,N_9208);
nand UO_211 (O_211,N_8832,N_8686);
and UO_212 (O_212,N_8393,N_8281);
and UO_213 (O_213,N_9062,N_9035);
nor UO_214 (O_214,N_8553,N_9567);
nand UO_215 (O_215,N_8449,N_9146);
or UO_216 (O_216,N_8389,N_9430);
nand UO_217 (O_217,N_8213,N_9800);
or UO_218 (O_218,N_8100,N_8198);
nor UO_219 (O_219,N_8032,N_9225);
and UO_220 (O_220,N_9715,N_9300);
nand UO_221 (O_221,N_8407,N_9653);
nor UO_222 (O_222,N_9219,N_8318);
xor UO_223 (O_223,N_9731,N_9867);
or UO_224 (O_224,N_9640,N_9677);
xnor UO_225 (O_225,N_8591,N_8836);
or UO_226 (O_226,N_8917,N_8629);
nand UO_227 (O_227,N_8261,N_9395);
nand UO_228 (O_228,N_9859,N_8820);
and UO_229 (O_229,N_8937,N_8295);
nor UO_230 (O_230,N_8129,N_9246);
nor UO_231 (O_231,N_8854,N_9935);
nand UO_232 (O_232,N_8633,N_8480);
xor UO_233 (O_233,N_8935,N_9636);
nor UO_234 (O_234,N_9162,N_8477);
or UO_235 (O_235,N_9268,N_8311);
nor UO_236 (O_236,N_8462,N_8005);
or UO_237 (O_237,N_9125,N_8764);
nor UO_238 (O_238,N_9418,N_9571);
nor UO_239 (O_239,N_8586,N_8631);
xor UO_240 (O_240,N_8664,N_8413);
nor UO_241 (O_241,N_8417,N_8502);
or UO_242 (O_242,N_8110,N_8895);
nor UO_243 (O_243,N_9930,N_9172);
or UO_244 (O_244,N_9656,N_9222);
nand UO_245 (O_245,N_9382,N_8950);
or UO_246 (O_246,N_9714,N_9900);
and UO_247 (O_247,N_8012,N_9493);
and UO_248 (O_248,N_9926,N_9917);
or UO_249 (O_249,N_8899,N_9662);
nand UO_250 (O_250,N_8365,N_8466);
or UO_251 (O_251,N_8834,N_8564);
nor UO_252 (O_252,N_9698,N_9713);
and UO_253 (O_253,N_9149,N_9067);
nand UO_254 (O_254,N_8043,N_9193);
nand UO_255 (O_255,N_9682,N_8406);
and UO_256 (O_256,N_8332,N_9856);
nand UO_257 (O_257,N_8498,N_8087);
and UO_258 (O_258,N_9881,N_9598);
nor UO_259 (O_259,N_8094,N_9025);
and UO_260 (O_260,N_8652,N_8835);
xor UO_261 (O_261,N_9517,N_9887);
nand UO_262 (O_262,N_8440,N_8377);
or UO_263 (O_263,N_9784,N_8131);
and UO_264 (O_264,N_9362,N_8998);
xor UO_265 (O_265,N_9509,N_9999);
nand UO_266 (O_266,N_8234,N_8028);
and UO_267 (O_267,N_9894,N_9499);
and UO_268 (O_268,N_8616,N_9564);
nor UO_269 (O_269,N_8170,N_9939);
or UO_270 (O_270,N_8156,N_8112);
or UO_271 (O_271,N_8848,N_8411);
xor UO_272 (O_272,N_8383,N_9110);
nand UO_273 (O_273,N_8752,N_8196);
nor UO_274 (O_274,N_9950,N_9673);
and UO_275 (O_275,N_8239,N_9724);
nor UO_276 (O_276,N_9890,N_9586);
nand UO_277 (O_277,N_8944,N_8582);
or UO_278 (O_278,N_8142,N_9360);
nor UO_279 (O_279,N_8039,N_8203);
and UO_280 (O_280,N_8185,N_8827);
or UO_281 (O_281,N_9845,N_9645);
nand UO_282 (O_282,N_9108,N_8085);
and UO_283 (O_283,N_8169,N_9182);
or UO_284 (O_284,N_8547,N_8762);
nor UO_285 (O_285,N_8329,N_8212);
nand UO_286 (O_286,N_9838,N_9593);
nor UO_287 (O_287,N_8853,N_9243);
nand UO_288 (O_288,N_9379,N_9710);
and UO_289 (O_289,N_8499,N_9954);
nor UO_290 (O_290,N_8750,N_8589);
nand UO_291 (O_291,N_8369,N_9986);
and UO_292 (O_292,N_9376,N_8696);
and UO_293 (O_293,N_8648,N_9700);
and UO_294 (O_294,N_8249,N_9864);
nand UO_295 (O_295,N_9106,N_8181);
nor UO_296 (O_296,N_8690,N_9135);
nand UO_297 (O_297,N_9575,N_8966);
nor UO_298 (O_298,N_9502,N_9389);
and UO_299 (O_299,N_8376,N_9238);
or UO_300 (O_300,N_9516,N_8138);
and UO_301 (O_301,N_9267,N_8179);
or UO_302 (O_302,N_8837,N_8441);
and UO_303 (O_303,N_8183,N_8657);
nor UO_304 (O_304,N_8808,N_8815);
and UO_305 (O_305,N_9664,N_9340);
nor UO_306 (O_306,N_9581,N_9403);
nand UO_307 (O_307,N_9644,N_8911);
and UO_308 (O_308,N_8350,N_9676);
and UO_309 (O_309,N_8428,N_9633);
nor UO_310 (O_310,N_8496,N_8651);
or UO_311 (O_311,N_9220,N_8843);
nor UO_312 (O_312,N_9983,N_9419);
and UO_313 (O_313,N_9432,N_9652);
nand UO_314 (O_314,N_8913,N_9997);
nand UO_315 (O_315,N_9409,N_9544);
and UO_316 (O_316,N_8534,N_8162);
and UO_317 (O_317,N_9666,N_8988);
and UO_318 (O_318,N_8708,N_9233);
or UO_319 (O_319,N_9273,N_9888);
nand UO_320 (O_320,N_9627,N_9539);
nor UO_321 (O_321,N_9937,N_8078);
nor UO_322 (O_322,N_9931,N_9202);
nor UO_323 (O_323,N_9271,N_9506);
nand UO_324 (O_324,N_9792,N_9425);
and UO_325 (O_325,N_8420,N_8803);
xor UO_326 (O_326,N_8684,N_9197);
xnor UO_327 (O_327,N_9093,N_8905);
nor UO_328 (O_328,N_8232,N_8528);
nand UO_329 (O_329,N_8530,N_9967);
and UO_330 (O_330,N_8375,N_9151);
nor UO_331 (O_331,N_9821,N_8458);
nand UO_332 (O_332,N_9557,N_9416);
and UO_333 (O_333,N_8990,N_9036);
and UO_334 (O_334,N_9016,N_9985);
and UO_335 (O_335,N_9975,N_8579);
or UO_336 (O_336,N_8274,N_9401);
xor UO_337 (O_337,N_9012,N_9265);
nor UO_338 (O_338,N_9352,N_9634);
nor UO_339 (O_339,N_8770,N_8007);
and UO_340 (O_340,N_8630,N_8956);
xnor UO_341 (O_341,N_9543,N_9380);
nor UO_342 (O_342,N_8025,N_9290);
xor UO_343 (O_343,N_9186,N_8439);
nand UO_344 (O_344,N_9442,N_9007);
xnor UO_345 (O_345,N_8720,N_9263);
and UO_346 (O_346,N_8120,N_8718);
nand UO_347 (O_347,N_8038,N_8307);
and UO_348 (O_348,N_8157,N_8892);
nand UO_349 (O_349,N_8444,N_8312);
nor UO_350 (O_350,N_9228,N_8873);
and UO_351 (O_351,N_9554,N_9752);
xor UO_352 (O_352,N_8567,N_8650);
and UO_353 (O_353,N_8981,N_8297);
or UO_354 (O_354,N_8875,N_9667);
or UO_355 (O_355,N_9778,N_9915);
xnor UO_356 (O_356,N_9311,N_9577);
and UO_357 (O_357,N_8544,N_9155);
and UO_358 (O_358,N_9443,N_9160);
xor UO_359 (O_359,N_9891,N_9015);
nor UO_360 (O_360,N_9631,N_9797);
nand UO_361 (O_361,N_8709,N_9875);
or UO_362 (O_362,N_8155,N_9648);
xor UO_363 (O_363,N_9584,N_9331);
or UO_364 (O_364,N_8673,N_8585);
and UO_365 (O_365,N_8503,N_8004);
nand UO_366 (O_366,N_9768,N_8408);
nand UO_367 (O_367,N_8540,N_8985);
nand UO_368 (O_368,N_9691,N_9369);
nand UO_369 (O_369,N_9045,N_8119);
and UO_370 (O_370,N_8516,N_9229);
or UO_371 (O_371,N_9034,N_8474);
and UO_372 (O_372,N_8997,N_9384);
xor UO_373 (O_373,N_8740,N_9200);
or UO_374 (O_374,N_9189,N_8174);
xnor UO_375 (O_375,N_9538,N_8581);
or UO_376 (O_376,N_9716,N_9944);
and UO_377 (O_377,N_9972,N_8791);
nor UO_378 (O_378,N_8026,N_8015);
and UO_379 (O_379,N_8678,N_8790);
nor UO_380 (O_380,N_9959,N_8044);
nor UO_381 (O_381,N_9316,N_8064);
nand UO_382 (O_382,N_8509,N_9173);
nor UO_383 (O_383,N_9892,N_8486);
nand UO_384 (O_384,N_9966,N_9366);
and UO_385 (O_385,N_8947,N_8374);
nor UO_386 (O_386,N_8062,N_8201);
xor UO_387 (O_387,N_9167,N_9470);
nand UO_388 (O_388,N_8071,N_8108);
xnor UO_389 (O_389,N_9301,N_9014);
xnor UO_390 (O_390,N_8838,N_8842);
or UO_391 (O_391,N_9746,N_8731);
nand UO_392 (O_392,N_9809,N_8103);
nor UO_393 (O_393,N_8902,N_8995);
nand UO_394 (O_394,N_8563,N_8101);
and UO_395 (O_395,N_8932,N_8253);
nand UO_396 (O_396,N_9453,N_9976);
nor UO_397 (O_397,N_9174,N_8308);
and UO_398 (O_398,N_9701,N_9932);
nor UO_399 (O_399,N_9574,N_9130);
and UO_400 (O_400,N_8128,N_9255);
nor UO_401 (O_401,N_9022,N_9413);
xor UO_402 (O_402,N_8858,N_8596);
or UO_403 (O_403,N_9021,N_9374);
and UO_404 (O_404,N_8034,N_9817);
or UO_405 (O_405,N_8602,N_9524);
xnor UO_406 (O_406,N_9317,N_8219);
or UO_407 (O_407,N_8734,N_9771);
and UO_408 (O_408,N_8983,N_9027);
nand UO_409 (O_409,N_8571,N_9721);
nand UO_410 (O_410,N_9102,N_9084);
nand UO_411 (O_411,N_9375,N_9558);
nor UO_412 (O_412,N_8618,N_9010);
xor UO_413 (O_413,N_8520,N_9696);
nand UO_414 (O_414,N_8016,N_8125);
nor UO_415 (O_415,N_9579,N_8430);
nor UO_416 (O_416,N_9582,N_8471);
nor UO_417 (O_417,N_8668,N_9277);
nand UO_418 (O_418,N_9269,N_8218);
and UO_419 (O_419,N_9241,N_9406);
and UO_420 (O_420,N_9306,N_9734);
nor UO_421 (O_421,N_8327,N_8346);
nand UO_422 (O_422,N_9073,N_9534);
nor UO_423 (O_423,N_9726,N_8556);
nand UO_424 (O_424,N_8324,N_8315);
nand UO_425 (O_425,N_9694,N_9880);
or UO_426 (O_426,N_9671,N_9129);
nor UO_427 (O_427,N_9378,N_9141);
or UO_428 (O_428,N_8529,N_9833);
nand UO_429 (O_429,N_9079,N_8378);
nand UO_430 (O_430,N_9595,N_8191);
nand UO_431 (O_431,N_8590,N_9861);
nand UO_432 (O_432,N_9594,N_8759);
xor UO_433 (O_433,N_8484,N_8224);
nor UO_434 (O_434,N_9583,N_8425);
or UO_435 (O_435,N_9485,N_8860);
and UO_436 (O_436,N_9185,N_8945);
or UO_437 (O_437,N_9013,N_8009);
nor UO_438 (O_438,N_9258,N_9445);
nand UO_439 (O_439,N_8184,N_8344);
xnor UO_440 (O_440,N_8010,N_9487);
nand UO_441 (O_441,N_9203,N_8066);
nor UO_442 (O_442,N_9943,N_9466);
nor UO_443 (O_443,N_9744,N_9924);
or UO_444 (O_444,N_8626,N_9688);
or UO_445 (O_445,N_8645,N_9783);
or UO_446 (O_446,N_8221,N_8380);
nand UO_447 (O_447,N_8931,N_8878);
and UO_448 (O_448,N_8583,N_9424);
and UO_449 (O_449,N_9836,N_9192);
nand UO_450 (O_450,N_9610,N_8788);
and UO_451 (O_451,N_8141,N_8091);
nand UO_452 (O_452,N_9876,N_8929);
nand UO_453 (O_453,N_9417,N_8829);
or UO_454 (O_454,N_9019,N_9743);
or UO_455 (O_455,N_8104,N_9874);
and UO_456 (O_456,N_9540,N_9240);
and UO_457 (O_457,N_9279,N_8876);
nand UO_458 (O_458,N_8114,N_9585);
or UO_459 (O_459,N_8736,N_9758);
nor UO_460 (O_460,N_9089,N_9121);
or UO_461 (O_461,N_8704,N_9974);
nor UO_462 (O_462,N_8299,N_9029);
or UO_463 (O_463,N_9198,N_9043);
nand UO_464 (O_464,N_8939,N_9624);
or UO_465 (O_465,N_9622,N_9293);
nor UO_466 (O_466,N_8122,N_9285);
nor UO_467 (O_467,N_9532,N_8614);
or UO_468 (O_468,N_9372,N_8211);
nor UO_469 (O_469,N_9103,N_8946);
nor UO_470 (O_470,N_9521,N_8802);
and UO_471 (O_471,N_9690,N_9294);
and UO_472 (O_472,N_8504,N_9968);
and UO_473 (O_473,N_8237,N_9429);
nand UO_474 (O_474,N_9776,N_9651);
nand UO_475 (O_475,N_8952,N_8711);
nand UO_476 (O_476,N_9469,N_9865);
or UO_477 (O_477,N_8419,N_8671);
and UO_478 (O_478,N_8065,N_9196);
xor UO_479 (O_479,N_9216,N_9353);
or UO_480 (O_480,N_8187,N_8436);
xor UO_481 (O_481,N_9550,N_9088);
or UO_482 (O_482,N_8949,N_8992);
nor UO_483 (O_483,N_8200,N_8123);
or UO_484 (O_484,N_9658,N_9003);
and UO_485 (O_485,N_9816,N_9617);
nand UO_486 (O_486,N_8881,N_8267);
and UO_487 (O_487,N_9934,N_9625);
nand UO_488 (O_488,N_8296,N_9561);
nor UO_489 (O_489,N_8751,N_8060);
nor UO_490 (O_490,N_9412,N_8470);
nand UO_491 (O_491,N_9823,N_9350);
nor UO_492 (O_492,N_9414,N_9068);
and UO_493 (O_493,N_9076,N_8151);
nand UO_494 (O_494,N_8634,N_9471);
nand UO_495 (O_495,N_8463,N_9846);
and UO_496 (O_496,N_8914,N_8568);
nand UO_497 (O_497,N_9500,N_8048);
nand UO_498 (O_498,N_8051,N_9420);
nor UO_499 (O_499,N_9946,N_8973);
nand UO_500 (O_500,N_8595,N_9970);
nand UO_501 (O_501,N_9452,N_8160);
and UO_502 (O_502,N_9451,N_8293);
or UO_503 (O_503,N_9787,N_8467);
or UO_504 (O_504,N_8742,N_8228);
nand UO_505 (O_505,N_8258,N_8314);
nand UO_506 (O_506,N_9608,N_9187);
nor UO_507 (O_507,N_9234,N_8072);
nor UO_508 (O_508,N_8388,N_9689);
or UO_509 (O_509,N_9087,N_9587);
nand UO_510 (O_510,N_9248,N_8084);
xor UO_511 (O_511,N_8850,N_8001);
xnor UO_512 (O_512,N_9619,N_8081);
nor UO_513 (O_513,N_8559,N_9889);
xor UO_514 (O_514,N_8304,N_9287);
xnor UO_515 (O_515,N_9391,N_9247);
or UO_516 (O_516,N_9123,N_8020);
and UO_517 (O_517,N_9560,N_9064);
and UO_518 (O_518,N_8974,N_9824);
xnor UO_519 (O_519,N_9511,N_8774);
and UO_520 (O_520,N_9848,N_8934);
and UO_521 (O_521,N_9562,N_8222);
or UO_522 (O_522,N_9695,N_9762);
or UO_523 (O_523,N_8628,N_9082);
and UO_524 (O_524,N_8606,N_9981);
nor UO_525 (O_525,N_9789,N_8810);
nor UO_526 (O_526,N_8317,N_8746);
and UO_527 (O_527,N_9548,N_9498);
nand UO_528 (O_528,N_8276,N_9785);
xnor UO_529 (O_529,N_8912,N_9764);
or UO_530 (O_530,N_9569,N_9251);
nor UO_531 (O_531,N_9295,N_8506);
nor UO_532 (O_532,N_9537,N_8250);
nor UO_533 (O_533,N_8494,N_8551);
xnor UO_534 (O_534,N_9116,N_8269);
xnor UO_535 (O_535,N_9844,N_8002);
and UO_536 (O_536,N_8938,N_8489);
nor UO_537 (O_537,N_9769,N_9392);
xnor UO_538 (O_538,N_8399,N_8984);
and UO_539 (O_539,N_8661,N_8760);
nor UO_540 (O_540,N_9335,N_9675);
nand UO_541 (O_541,N_8741,N_8524);
xor UO_542 (O_542,N_9339,N_8368);
nor UO_543 (O_543,N_9284,N_8573);
or UO_544 (O_544,N_9495,N_9920);
and UO_545 (O_545,N_9404,N_9211);
nor UO_546 (O_546,N_8732,N_8620);
or UO_547 (O_547,N_8493,N_9363);
nor UO_548 (O_548,N_8137,N_9811);
nand UO_549 (O_549,N_9368,N_8351);
nor UO_550 (O_550,N_9615,N_8132);
or UO_551 (O_551,N_8468,N_8537);
nor UO_552 (O_552,N_8570,N_8018);
nand UO_553 (O_553,N_8941,N_9386);
nand UO_554 (O_554,N_8891,N_9572);
nand UO_555 (O_555,N_9334,N_8285);
and UO_556 (O_556,N_9810,N_8593);
or UO_557 (O_557,N_9840,N_9508);
or UO_558 (O_558,N_9788,N_8809);
nor UO_559 (O_559,N_9773,N_8739);
or UO_560 (O_560,N_8278,N_9657);
nand UO_561 (O_561,N_8117,N_8670);
nor UO_562 (O_562,N_8330,N_8728);
and UO_563 (O_563,N_8793,N_8880);
nor UO_564 (O_564,N_8580,N_9018);
nor UO_565 (O_565,N_8483,N_9685);
xor UO_566 (O_566,N_9884,N_8268);
nor UO_567 (O_567,N_9777,N_8679);
nand UO_568 (O_568,N_9488,N_9324);
and UO_569 (O_569,N_9126,N_9505);
and UO_570 (O_570,N_8921,N_9052);
nor UO_571 (O_571,N_9351,N_8738);
and UO_572 (O_572,N_9649,N_9080);
or UO_573 (O_573,N_9600,N_9354);
nor UO_574 (O_574,N_9462,N_8190);
or UO_575 (O_575,N_9431,N_9855);
nand UO_576 (O_576,N_9458,N_9563);
and UO_577 (O_577,N_8933,N_8572);
and UO_578 (O_578,N_8033,N_9479);
or UO_579 (O_579,N_9276,N_9100);
nand UO_580 (O_580,N_9529,N_8403);
or UO_581 (O_581,N_9020,N_8986);
or UO_582 (O_582,N_9754,N_8710);
xor UO_583 (O_583,N_9017,N_9832);
and UO_584 (O_584,N_8639,N_9858);
nand UO_585 (O_585,N_9347,N_8961);
nand UO_586 (O_586,N_8387,N_8955);
and UO_587 (O_587,N_8475,N_8204);
and UO_588 (O_588,N_9987,N_9742);
nor UO_589 (O_589,N_9839,N_8429);
xnor UO_590 (O_590,N_8624,N_9048);
nor UO_591 (O_591,N_8031,N_8126);
or UO_592 (O_592,N_8139,N_9242);
nand UO_593 (O_593,N_8341,N_8817);
and UO_594 (O_594,N_9078,N_8333);
and UO_595 (O_595,N_9613,N_9394);
nand UO_596 (O_596,N_8447,N_9614);
and UO_597 (O_597,N_9936,N_9184);
or UO_598 (O_598,N_8806,N_9835);
nor UO_599 (O_599,N_9323,N_8870);
nor UO_600 (O_600,N_9901,N_9847);
nand UO_601 (O_601,N_8412,N_9099);
nor UO_602 (O_602,N_8175,N_9270);
nand UO_603 (O_603,N_8340,N_8240);
nor UO_604 (O_604,N_9604,N_9283);
or UO_605 (O_605,N_9288,N_8982);
nor UO_606 (O_606,N_9542,N_8360);
and UO_607 (O_607,N_8287,N_8757);
or UO_608 (O_608,N_8433,N_9166);
nand UO_609 (O_609,N_9591,N_8348);
nor UO_610 (O_610,N_9011,N_9909);
and UO_611 (O_611,N_8663,N_9128);
and UO_612 (O_612,N_8445,N_8195);
and UO_613 (O_613,N_8587,N_9978);
nand UO_614 (O_614,N_8831,N_9989);
nand UO_615 (O_615,N_8765,N_8721);
and UO_616 (O_616,N_8623,N_9227);
nor UO_617 (O_617,N_8840,N_9918);
nand UO_618 (O_618,N_9919,N_9732);
nand UO_619 (O_619,N_9612,N_8225);
xnor UO_620 (O_620,N_8656,N_8794);
and UO_621 (O_621,N_8106,N_9398);
and UO_622 (O_622,N_8335,N_9503);
nand UO_623 (O_623,N_8924,N_9181);
nor UO_624 (O_624,N_9122,N_8459);
nand UO_625 (O_625,N_8172,N_9798);
nor UO_626 (O_626,N_8006,N_8473);
or UO_627 (O_627,N_8951,N_8822);
or UO_628 (O_628,N_9912,N_8437);
nand UO_629 (O_629,N_9464,N_9152);
nand UO_630 (O_630,N_9630,N_8017);
nor UO_631 (O_631,N_9531,N_9438);
or UO_632 (O_632,N_8342,N_8316);
nand UO_633 (O_633,N_8658,N_9314);
and UO_634 (O_634,N_8600,N_9028);
nand UO_635 (O_635,N_8392,N_8422);
and UO_636 (O_636,N_9801,N_8336);
or UO_637 (O_637,N_8130,N_8508);
and UO_638 (O_638,N_9528,N_8223);
nor UO_639 (O_639,N_8359,N_8967);
nand UO_640 (O_640,N_9536,N_9962);
xnor UO_641 (O_641,N_9927,N_9551);
or UO_642 (O_642,N_8541,N_8173);
nand UO_643 (O_643,N_9332,N_8970);
nand UO_644 (O_644,N_9877,N_8208);
nand UO_645 (O_645,N_8743,N_8036);
and UO_646 (O_646,N_9348,N_9749);
nand UO_647 (O_647,N_8056,N_9343);
nor UO_648 (O_648,N_9004,N_8322);
nor UO_649 (O_649,N_9654,N_9611);
or UO_650 (O_650,N_9638,N_8919);
and UO_651 (O_651,N_8893,N_8478);
nand UO_652 (O_652,N_8410,N_8434);
nand UO_653 (O_653,N_8894,N_9070);
and UO_654 (O_654,N_9209,N_8280);
nor UO_655 (O_655,N_8560,N_8943);
nor UO_656 (O_656,N_9381,N_9717);
nor UO_657 (O_657,N_8047,N_8884);
nor UO_658 (O_658,N_9230,N_8512);
or UO_659 (O_659,N_8373,N_8855);
and UO_660 (O_660,N_9770,N_8099);
and UO_661 (O_661,N_8936,N_9057);
and UO_662 (O_662,N_9144,N_8744);
nor UO_663 (O_663,N_8140,N_9117);
nand UO_664 (O_664,N_9188,N_9993);
nor UO_665 (O_665,N_8898,N_8227);
nor UO_666 (O_666,N_8727,N_8691);
nand UO_667 (O_667,N_8319,N_8532);
nor UO_668 (O_668,N_9302,N_8644);
xor UO_669 (O_669,N_9180,N_8053);
nand UO_670 (O_670,N_8907,N_8217);
nand UO_671 (O_671,N_9147,N_9054);
nand UO_672 (O_672,N_8819,N_9956);
and UO_673 (O_673,N_8409,N_8405);
nor UO_674 (O_674,N_9373,N_9958);
and UO_675 (O_675,N_8798,N_8231);
nand UO_676 (O_676,N_9254,N_8310);
or UO_677 (O_677,N_8714,N_9813);
and UO_678 (O_678,N_9213,N_8305);
nor UO_679 (O_679,N_8683,N_9668);
nand UO_680 (O_680,N_9357,N_8097);
and UO_681 (O_681,N_9325,N_8186);
nor UO_682 (O_682,N_9933,N_8363);
and UO_683 (O_683,N_8092,N_9868);
nor UO_684 (O_684,N_8424,N_8763);
and UO_685 (O_685,N_8074,N_8896);
xor UO_686 (O_686,N_8723,N_8109);
xnor UO_687 (O_687,N_9361,N_8432);
and UO_688 (O_688,N_9568,N_9580);
nand UO_689 (O_689,N_8958,N_9107);
or UO_690 (O_690,N_9893,N_8290);
nand UO_691 (O_691,N_9552,N_9032);
xnor UO_692 (O_692,N_8124,N_9448);
nor UO_693 (O_693,N_9830,N_9723);
nor UO_694 (O_694,N_8766,N_9765);
nor UO_695 (O_695,N_8030,N_9555);
nor UO_696 (O_696,N_9168,N_8500);
or UO_697 (O_697,N_9998,N_9530);
or UO_698 (O_698,N_9136,N_9914);
nor UO_699 (O_699,N_8229,N_9002);
nor UO_700 (O_700,N_9928,N_9454);
xnor UO_701 (O_701,N_9402,N_8248);
or UO_702 (O_702,N_9281,N_9033);
or UO_703 (O_703,N_9525,N_8390);
nand UO_704 (O_704,N_8617,N_8013);
xor UO_705 (O_705,N_9955,N_8115);
nor UO_706 (O_706,N_8371,N_8133);
xnor UO_707 (O_707,N_9218,N_9305);
and UO_708 (O_708,N_8416,N_9133);
or UO_709 (O_709,N_9482,N_8533);
or UO_710 (O_710,N_9605,N_8667);
and UO_711 (O_711,N_8482,N_8926);
and UO_712 (O_712,N_9977,N_8826);
and UO_713 (O_713,N_8999,N_9896);
nor UO_714 (O_714,N_8613,N_9693);
or UO_715 (O_715,N_9870,N_9818);
nor UO_716 (O_716,N_9687,N_8954);
xnor UO_717 (O_717,N_8095,N_8771);
xnor UO_718 (O_718,N_9260,N_8323);
nand UO_719 (O_719,N_8522,N_8057);
nand UO_720 (O_720,N_8554,N_9421);
and UO_721 (O_721,N_9826,N_9763);
nor UO_722 (O_722,N_8666,N_9669);
and UO_723 (O_723,N_9206,N_9535);
nor UO_724 (O_724,N_8611,N_8356);
xor UO_725 (O_725,N_8401,N_8968);
nor UO_726 (O_726,N_8022,N_9364);
nor UO_727 (O_727,N_9397,N_8856);
nor UO_728 (O_728,N_8485,N_9456);
or UO_729 (O_729,N_8797,N_9463);
nand UO_730 (O_730,N_8543,N_9815);
and UO_731 (O_731,N_8397,N_9274);
xor UO_732 (O_732,N_8852,N_8098);
or UO_733 (O_733,N_9310,N_9592);
or UO_734 (O_734,N_8361,N_8147);
nand UO_735 (O_735,N_8526,N_8282);
nor UO_736 (O_736,N_9988,N_8472);
and UO_737 (O_737,N_9475,N_8849);
or UO_738 (O_738,N_8925,N_8338);
nor UO_739 (O_739,N_8288,N_9729);
and UO_740 (O_740,N_9678,N_8379);
xor UO_741 (O_741,N_9804,N_9878);
nand UO_742 (O_742,N_9047,N_8874);
and UO_743 (O_743,N_8603,N_8511);
nand UO_744 (O_744,N_9674,N_9906);
nand UO_745 (O_745,N_9808,N_8404);
or UO_746 (O_746,N_9566,N_8928);
and UO_747 (O_747,N_9681,N_8724);
or UO_748 (O_748,N_9995,N_8767);
xnor UO_749 (O_749,N_8334,N_8027);
nand UO_750 (O_750,N_9253,N_8189);
nand UO_751 (O_751,N_9261,N_9526);
nand UO_752 (O_752,N_8055,N_8889);
and UO_753 (O_753,N_8080,N_8210);
nor UO_754 (O_754,N_9096,N_9437);
nor UO_755 (O_755,N_9686,N_9902);
and UO_756 (O_756,N_9851,N_8492);
and UO_757 (O_757,N_9692,N_8050);
or UO_758 (O_758,N_9515,N_9455);
nor UO_759 (O_759,N_9541,N_8521);
nor UO_760 (O_760,N_9063,N_8070);
or UO_761 (O_761,N_9559,N_9161);
nor UO_762 (O_762,N_9158,N_8088);
or UO_763 (O_763,N_9553,N_8083);
xnor UO_764 (O_764,N_9820,N_8811);
nand UO_765 (O_765,N_8497,N_9751);
xnor UO_766 (O_766,N_9596,N_9637);
nor UO_767 (O_767,N_9549,N_8689);
or UO_768 (O_768,N_8303,N_8301);
xnor UO_769 (O_769,N_9670,N_8755);
or UO_770 (O_770,N_9336,N_9170);
or UO_771 (O_771,N_8904,N_8294);
and UO_772 (O_772,N_8418,N_9142);
and UO_773 (O_773,N_8398,N_9164);
nand UO_774 (O_774,N_8197,N_8021);
nand UO_775 (O_775,N_9756,N_8309);
nor UO_776 (O_776,N_8215,N_9159);
or UO_777 (O_777,N_8523,N_9702);
or UO_778 (O_778,N_9991,N_9436);
and UO_779 (O_779,N_8510,N_9659);
or UO_780 (O_780,N_8697,N_8046);
nand UO_781 (O_781,N_8845,N_9289);
nand UO_782 (O_782,N_8717,N_8313);
xnor UO_783 (O_783,N_9663,N_9266);
nand UO_784 (O_784,N_9480,N_9907);
and UO_785 (O_785,N_8265,N_9282);
or UO_786 (O_786,N_8068,N_9590);
and UO_787 (O_787,N_8604,N_8041);
nor UO_788 (O_788,N_9780,N_9137);
nand UO_789 (O_789,N_8238,N_8972);
nor UO_790 (O_790,N_8089,N_9910);
and UO_791 (O_791,N_9957,N_8758);
and UO_792 (O_792,N_9665,N_9041);
nand UO_793 (O_793,N_9952,N_8607);
and UO_794 (O_794,N_9842,N_8495);
or UO_795 (O_795,N_8839,N_8014);
and UO_796 (O_796,N_8245,N_8431);
or UO_797 (O_797,N_9602,N_8669);
xor UO_798 (O_798,N_9000,N_9643);
nand UO_799 (O_799,N_8680,N_8353);
or UO_800 (O_800,N_9601,N_8722);
xnor UO_801 (O_801,N_8700,N_9086);
or UO_802 (O_802,N_8906,N_9712);
or UO_803 (O_803,N_9095,N_9223);
nand UO_804 (O_804,N_8063,N_9410);
or UO_805 (O_805,N_9292,N_8107);
and UO_806 (O_806,N_9081,N_8362);
and UO_807 (O_807,N_9477,N_9303);
or UO_808 (O_808,N_9124,N_8402);
nor UO_809 (O_809,N_9163,N_8154);
nand UO_810 (O_810,N_9280,N_8339);
xor UO_811 (O_811,N_8576,N_9030);
xnor UO_812 (O_812,N_9708,N_8754);
and UO_813 (O_813,N_9439,N_9023);
or UO_814 (O_814,N_9156,N_8867);
and UO_815 (O_815,N_9629,N_8349);
nor UO_816 (O_816,N_9737,N_8093);
or UO_817 (O_817,N_9767,N_8989);
nor UO_818 (O_818,N_9507,N_9195);
nand UO_819 (O_819,N_9790,N_8069);
or UO_820 (O_820,N_8481,N_8747);
nor UO_821 (O_821,N_8372,N_8209);
xor UO_822 (O_822,N_9313,N_9996);
or UO_823 (O_823,N_8531,N_8877);
and UO_824 (O_824,N_8882,N_8886);
and UO_825 (O_825,N_9153,N_8256);
or UO_826 (O_826,N_9114,N_8289);
and UO_827 (O_827,N_8145,N_8292);
nor UO_828 (O_828,N_8566,N_9320);
nor UO_829 (O_829,N_8539,N_9711);
nor UO_830 (O_830,N_8962,N_9065);
and UO_831 (O_831,N_9058,N_8795);
xor UO_832 (O_832,N_9883,N_8263);
and UO_833 (O_833,N_9607,N_9328);
and UO_834 (O_834,N_9105,N_9545);
nor UO_835 (O_835,N_8082,N_9951);
nand UO_836 (O_836,N_9819,N_8569);
or UO_837 (O_837,N_9871,N_8193);
nand UO_838 (O_838,N_9318,N_8366);
and UO_839 (O_839,N_8488,N_9481);
nor UO_840 (O_840,N_8660,N_8357);
and UO_841 (O_841,N_8713,N_9132);
and UO_842 (O_842,N_8641,N_8761);
and UO_843 (O_843,N_9210,N_8909);
and UO_844 (O_844,N_9750,N_8851);
and UO_845 (O_845,N_8490,N_8625);
nand UO_846 (O_846,N_9286,N_9484);
or UO_847 (O_847,N_8622,N_8592);
nand UO_848 (O_848,N_9427,N_9371);
or UO_849 (O_849,N_9183,N_9873);
or UO_850 (O_850,N_9120,N_9860);
nor UO_851 (O_851,N_8011,N_8674);
or UO_852 (O_852,N_8000,N_8872);
or UO_853 (O_853,N_9341,N_8167);
nor UO_854 (O_854,N_9278,N_8394);
and UO_855 (O_855,N_8273,N_8621);
or UO_856 (O_856,N_9616,N_8090);
xor UO_857 (O_857,N_8102,N_9527);
or UO_858 (O_858,N_9807,N_8627);
xor UO_859 (O_859,N_9941,N_9444);
and UO_860 (O_860,N_9113,N_9264);
xnor UO_861 (O_861,N_9044,N_9337);
and UO_862 (O_862,N_8706,N_8182);
nand UO_863 (O_863,N_8781,N_9346);
and UO_864 (O_864,N_9212,N_9101);
nor UO_865 (O_865,N_8448,N_8476);
and UO_866 (O_866,N_8171,N_9457);
nand UO_867 (O_867,N_8535,N_8948);
and UO_868 (O_868,N_8897,N_8915);
or UO_869 (O_869,N_9599,N_8864);
or UO_870 (O_870,N_9683,N_8859);
nand UO_871 (O_871,N_9841,N_9315);
and UO_872 (O_872,N_8178,N_8594);
nand UO_873 (O_873,N_8964,N_9039);
and UO_874 (O_874,N_8035,N_8086);
and UO_875 (O_875,N_9916,N_8262);
nor UO_876 (O_876,N_9513,N_9942);
and UO_877 (O_877,N_8396,N_8414);
nor UO_878 (O_878,N_9008,N_8037);
and UO_879 (O_879,N_9766,N_9496);
or UO_880 (O_880,N_9411,N_9831);
nor UO_881 (O_881,N_9483,N_9304);
or UO_882 (O_882,N_8271,N_9387);
nor UO_883 (O_883,N_8321,N_8901);
nor UO_884 (O_884,N_9519,N_9321);
nor UO_885 (O_885,N_9501,N_9735);
and UO_886 (O_886,N_8024,N_8782);
or UO_887 (O_887,N_9050,N_8542);
xnor UO_888 (O_888,N_8783,N_8918);
or UO_889 (O_889,N_8391,N_9953);
or UO_890 (O_890,N_9092,N_9083);
or UO_891 (O_891,N_8558,N_9145);
and UO_892 (O_892,N_8453,N_9297);
or UO_893 (O_893,N_8367,N_8775);
nor UO_894 (O_894,N_8279,N_8971);
and UO_895 (O_895,N_8188,N_9806);
nand UO_896 (O_896,N_8236,N_9547);
nor UO_897 (O_897,N_8841,N_8465);
and UO_898 (O_898,N_8769,N_8146);
and UO_899 (O_899,N_8300,N_9775);
nand UO_900 (O_900,N_8246,N_9857);
xor UO_901 (O_901,N_8653,N_9620);
nand UO_902 (O_902,N_9055,N_9757);
or UO_903 (O_903,N_8008,N_9523);
nor UO_904 (O_904,N_9074,N_8735);
nand UO_905 (O_905,N_9576,N_8384);
xnor UO_906 (O_906,N_9355,N_8707);
nor UO_907 (O_907,N_8306,N_8254);
and UO_908 (O_908,N_8694,N_9207);
or UO_909 (O_909,N_9119,N_8903);
and UO_910 (O_910,N_8345,N_8588);
nor UO_911 (O_911,N_8638,N_8207);
or UO_912 (O_912,N_8792,N_9098);
or UO_913 (O_913,N_8385,N_9326);
or UO_914 (O_914,N_8355,N_9494);
nor UO_915 (O_915,N_9849,N_9969);
nand UO_916 (O_916,N_9112,N_8780);
and UO_917 (O_917,N_8206,N_9908);
or UO_918 (O_918,N_9115,N_9709);
nand UO_919 (O_919,N_9520,N_8283);
nand UO_920 (O_920,N_8291,N_8487);
nand UO_921 (O_921,N_8168,N_9169);
nand UO_922 (O_922,N_8513,N_9175);
and UO_923 (O_923,N_8804,N_8865);
and UO_924 (O_924,N_8662,N_9753);
xnor UO_925 (O_925,N_8415,N_8501);
nand UO_926 (O_926,N_9249,N_8552);
and UO_927 (O_927,N_9040,N_9949);
xor UO_928 (O_928,N_8148,N_8515);
and UO_929 (O_929,N_9338,N_9781);
and UO_930 (O_930,N_8116,N_8230);
and UO_931 (O_931,N_8883,N_9623);
nand UO_932 (O_932,N_9072,N_9199);
and UO_933 (O_933,N_9190,N_8079);
or UO_934 (O_934,N_8105,N_9948);
or UO_935 (O_935,N_8421,N_8910);
nand UO_936 (O_936,N_8866,N_8688);
or UO_937 (O_937,N_8284,N_8823);
and UO_938 (O_938,N_8548,N_8716);
nand UO_939 (O_939,N_8266,N_9367);
nand UO_940 (O_940,N_9725,N_9782);
or UO_941 (O_941,N_9296,N_8940);
or UO_942 (O_942,N_8960,N_8456);
nor UO_943 (O_943,N_8730,N_8705);
nand UO_944 (O_944,N_9345,N_9006);
nor UO_945 (O_945,N_9964,N_9091);
nand UO_946 (O_946,N_8354,N_9803);
nand UO_947 (O_947,N_9232,N_8059);
or UO_948 (O_948,N_9435,N_8632);
and UO_949 (O_949,N_9194,N_9973);
or UO_950 (O_950,N_9467,N_9071);
or UO_951 (O_951,N_8286,N_9358);
nand UO_952 (O_952,N_8226,N_8597);
or UO_953 (O_953,N_9609,N_8692);
and UO_954 (O_954,N_8192,N_8647);
or UO_955 (O_955,N_9085,N_9370);
and UO_956 (O_956,N_9148,N_9492);
xnor UO_957 (O_957,N_8166,N_9748);
and UO_958 (O_958,N_9963,N_9650);
or UO_959 (O_959,N_9812,N_8527);
nor UO_960 (O_960,N_9476,N_9639);
xor UO_961 (O_961,N_9697,N_9322);
nand UO_962 (O_962,N_8144,N_8643);
or UO_963 (O_963,N_8165,N_8326);
nand UO_964 (O_964,N_9176,N_9565);
nor UO_965 (O_965,N_9647,N_8748);
or UO_966 (O_966,N_8400,N_9237);
and UO_967 (O_967,N_9459,N_9913);
nand UO_968 (O_968,N_8023,N_9533);
or UO_969 (O_969,N_9231,N_8977);
xor UO_970 (O_970,N_9862,N_9704);
xor UO_971 (O_971,N_8205,N_8963);
or UO_972 (O_972,N_8464,N_8199);
and UO_973 (O_973,N_8796,N_8331);
and UO_974 (O_974,N_9814,N_9863);
and UO_975 (O_975,N_8655,N_9201);
nand UO_976 (O_976,N_8337,N_9982);
nand UO_977 (O_977,N_9221,N_8343);
and UO_978 (O_978,N_9131,N_8993);
nand UO_979 (O_979,N_8461,N_9805);
or UO_980 (O_980,N_9256,N_9026);
nor UO_981 (O_981,N_8879,N_8194);
nand UO_982 (O_982,N_8640,N_8565);
and UO_983 (O_983,N_9178,N_9899);
nand UO_984 (O_984,N_9165,N_9556);
and UO_985 (O_985,N_8136,N_9104);
and UO_986 (O_986,N_9356,N_9400);
nor UO_987 (O_987,N_8451,N_9489);
nand UO_988 (O_988,N_8364,N_8959);
and UO_989 (O_989,N_8726,N_9053);
or UO_990 (O_990,N_9772,N_9745);
xnor UO_991 (O_991,N_8561,N_8052);
or UO_992 (O_992,N_9802,N_9291);
xor UO_993 (O_993,N_9272,N_8202);
nor UO_994 (O_994,N_8749,N_8800);
nand UO_995 (O_995,N_8636,N_8619);
and UO_996 (O_996,N_8320,N_9965);
or UO_997 (O_997,N_9365,N_8073);
nand UO_998 (O_998,N_8446,N_8920);
and UO_999 (O_999,N_9929,N_8370);
or UO_1000 (O_1000,N_9551,N_9268);
xnor UO_1001 (O_1001,N_8603,N_8114);
nand UO_1002 (O_1002,N_8269,N_8093);
xor UO_1003 (O_1003,N_9623,N_9691);
or UO_1004 (O_1004,N_8838,N_9781);
nor UO_1005 (O_1005,N_9734,N_8178);
nor UO_1006 (O_1006,N_9183,N_9320);
and UO_1007 (O_1007,N_9705,N_9644);
nor UO_1008 (O_1008,N_9645,N_8745);
or UO_1009 (O_1009,N_8725,N_8975);
nand UO_1010 (O_1010,N_8855,N_8366);
or UO_1011 (O_1011,N_8406,N_8344);
nand UO_1012 (O_1012,N_8494,N_9816);
nand UO_1013 (O_1013,N_8080,N_8422);
nor UO_1014 (O_1014,N_9818,N_8138);
nand UO_1015 (O_1015,N_9402,N_8368);
and UO_1016 (O_1016,N_9707,N_8142);
xnor UO_1017 (O_1017,N_8514,N_9633);
or UO_1018 (O_1018,N_8981,N_8928);
nor UO_1019 (O_1019,N_8008,N_9872);
xor UO_1020 (O_1020,N_8381,N_8818);
nand UO_1021 (O_1021,N_9140,N_9507);
nand UO_1022 (O_1022,N_9089,N_9067);
or UO_1023 (O_1023,N_9289,N_8967);
nor UO_1024 (O_1024,N_8722,N_9103);
nor UO_1025 (O_1025,N_8738,N_9338);
xnor UO_1026 (O_1026,N_9234,N_9642);
xnor UO_1027 (O_1027,N_9994,N_9971);
nor UO_1028 (O_1028,N_9095,N_8850);
nand UO_1029 (O_1029,N_8086,N_8727);
nor UO_1030 (O_1030,N_9030,N_8912);
or UO_1031 (O_1031,N_9182,N_8093);
and UO_1032 (O_1032,N_8468,N_9932);
or UO_1033 (O_1033,N_8946,N_9897);
and UO_1034 (O_1034,N_8246,N_9771);
or UO_1035 (O_1035,N_9742,N_9418);
nand UO_1036 (O_1036,N_8576,N_8006);
or UO_1037 (O_1037,N_8356,N_9680);
nor UO_1038 (O_1038,N_8150,N_9764);
and UO_1039 (O_1039,N_9711,N_9551);
or UO_1040 (O_1040,N_9517,N_9071);
or UO_1041 (O_1041,N_8395,N_8056);
xor UO_1042 (O_1042,N_8478,N_9654);
nand UO_1043 (O_1043,N_8590,N_8569);
or UO_1044 (O_1044,N_9511,N_9557);
or UO_1045 (O_1045,N_8050,N_9172);
nor UO_1046 (O_1046,N_9234,N_9054);
nor UO_1047 (O_1047,N_8113,N_8451);
nand UO_1048 (O_1048,N_8418,N_9437);
and UO_1049 (O_1049,N_9580,N_9871);
nand UO_1050 (O_1050,N_9756,N_9416);
xor UO_1051 (O_1051,N_8126,N_9430);
or UO_1052 (O_1052,N_9116,N_9907);
and UO_1053 (O_1053,N_8814,N_8219);
and UO_1054 (O_1054,N_9627,N_8129);
nand UO_1055 (O_1055,N_9783,N_9063);
or UO_1056 (O_1056,N_8837,N_9290);
xor UO_1057 (O_1057,N_8102,N_9054);
or UO_1058 (O_1058,N_9703,N_9372);
nand UO_1059 (O_1059,N_8476,N_8750);
nand UO_1060 (O_1060,N_8229,N_9923);
or UO_1061 (O_1061,N_8753,N_9392);
nand UO_1062 (O_1062,N_8666,N_9222);
or UO_1063 (O_1063,N_9052,N_9769);
nor UO_1064 (O_1064,N_8203,N_9643);
or UO_1065 (O_1065,N_9319,N_9981);
nand UO_1066 (O_1066,N_8987,N_9023);
xor UO_1067 (O_1067,N_9844,N_9397);
and UO_1068 (O_1068,N_9348,N_8372);
nand UO_1069 (O_1069,N_8776,N_9178);
or UO_1070 (O_1070,N_9956,N_9172);
and UO_1071 (O_1071,N_9782,N_9471);
nand UO_1072 (O_1072,N_9344,N_9052);
and UO_1073 (O_1073,N_9144,N_8600);
xor UO_1074 (O_1074,N_8674,N_9303);
nand UO_1075 (O_1075,N_8059,N_9119);
and UO_1076 (O_1076,N_9194,N_8020);
or UO_1077 (O_1077,N_9677,N_8448);
or UO_1078 (O_1078,N_8762,N_9571);
nor UO_1079 (O_1079,N_9760,N_8107);
nand UO_1080 (O_1080,N_8498,N_8677);
xor UO_1081 (O_1081,N_9680,N_9115);
nand UO_1082 (O_1082,N_9112,N_9684);
nand UO_1083 (O_1083,N_9144,N_9015);
or UO_1084 (O_1084,N_9827,N_9762);
nor UO_1085 (O_1085,N_8336,N_8163);
nor UO_1086 (O_1086,N_8909,N_8950);
or UO_1087 (O_1087,N_9729,N_9341);
nand UO_1088 (O_1088,N_9873,N_8021);
nor UO_1089 (O_1089,N_8548,N_8444);
nand UO_1090 (O_1090,N_8546,N_8691);
nor UO_1091 (O_1091,N_9026,N_8917);
xor UO_1092 (O_1092,N_9193,N_8372);
and UO_1093 (O_1093,N_9993,N_8012);
nor UO_1094 (O_1094,N_9197,N_8740);
or UO_1095 (O_1095,N_8662,N_9152);
nor UO_1096 (O_1096,N_8503,N_8769);
xnor UO_1097 (O_1097,N_8851,N_8803);
nor UO_1098 (O_1098,N_9681,N_8456);
and UO_1099 (O_1099,N_8270,N_8047);
xor UO_1100 (O_1100,N_8371,N_9028);
and UO_1101 (O_1101,N_9765,N_8612);
and UO_1102 (O_1102,N_8709,N_8595);
or UO_1103 (O_1103,N_9168,N_9509);
xnor UO_1104 (O_1104,N_9305,N_9221);
and UO_1105 (O_1105,N_9280,N_9866);
and UO_1106 (O_1106,N_8037,N_8029);
nor UO_1107 (O_1107,N_9091,N_9532);
or UO_1108 (O_1108,N_8654,N_8145);
nand UO_1109 (O_1109,N_8720,N_8611);
xor UO_1110 (O_1110,N_8428,N_9683);
nand UO_1111 (O_1111,N_8116,N_8602);
xor UO_1112 (O_1112,N_8265,N_8106);
and UO_1113 (O_1113,N_8937,N_9355);
or UO_1114 (O_1114,N_8172,N_8229);
and UO_1115 (O_1115,N_8611,N_9600);
nand UO_1116 (O_1116,N_8718,N_8402);
nor UO_1117 (O_1117,N_9505,N_9253);
and UO_1118 (O_1118,N_9769,N_9729);
or UO_1119 (O_1119,N_8174,N_9623);
nor UO_1120 (O_1120,N_9155,N_9541);
or UO_1121 (O_1121,N_9879,N_9427);
and UO_1122 (O_1122,N_9604,N_9312);
nor UO_1123 (O_1123,N_9098,N_9832);
nand UO_1124 (O_1124,N_9821,N_9022);
and UO_1125 (O_1125,N_8245,N_9043);
xnor UO_1126 (O_1126,N_9713,N_8158);
xor UO_1127 (O_1127,N_8814,N_9781);
xor UO_1128 (O_1128,N_8956,N_9614);
or UO_1129 (O_1129,N_8348,N_8437);
or UO_1130 (O_1130,N_9744,N_8597);
or UO_1131 (O_1131,N_8729,N_9767);
nor UO_1132 (O_1132,N_9919,N_9802);
or UO_1133 (O_1133,N_8087,N_8341);
nand UO_1134 (O_1134,N_9389,N_8222);
xor UO_1135 (O_1135,N_9591,N_9115);
nand UO_1136 (O_1136,N_8894,N_8004);
and UO_1137 (O_1137,N_9950,N_9237);
nand UO_1138 (O_1138,N_9869,N_9125);
xnor UO_1139 (O_1139,N_8092,N_8281);
and UO_1140 (O_1140,N_8773,N_8427);
and UO_1141 (O_1141,N_8082,N_9293);
and UO_1142 (O_1142,N_8366,N_9037);
nand UO_1143 (O_1143,N_8057,N_8929);
and UO_1144 (O_1144,N_8929,N_9410);
nor UO_1145 (O_1145,N_9321,N_9253);
nand UO_1146 (O_1146,N_9571,N_8489);
or UO_1147 (O_1147,N_8817,N_8082);
nor UO_1148 (O_1148,N_8901,N_8510);
nor UO_1149 (O_1149,N_8559,N_9291);
nor UO_1150 (O_1150,N_9868,N_9622);
and UO_1151 (O_1151,N_9167,N_9675);
or UO_1152 (O_1152,N_8752,N_9845);
nand UO_1153 (O_1153,N_9495,N_9656);
nand UO_1154 (O_1154,N_8718,N_9954);
and UO_1155 (O_1155,N_9530,N_9023);
or UO_1156 (O_1156,N_8273,N_8741);
or UO_1157 (O_1157,N_9405,N_8884);
nand UO_1158 (O_1158,N_8751,N_9665);
nor UO_1159 (O_1159,N_8460,N_8714);
nand UO_1160 (O_1160,N_9555,N_8846);
or UO_1161 (O_1161,N_9451,N_9433);
nor UO_1162 (O_1162,N_8700,N_8836);
and UO_1163 (O_1163,N_9843,N_8306);
nor UO_1164 (O_1164,N_9430,N_9323);
and UO_1165 (O_1165,N_8840,N_9642);
or UO_1166 (O_1166,N_8559,N_8501);
nor UO_1167 (O_1167,N_9960,N_8236);
nor UO_1168 (O_1168,N_9165,N_8534);
nor UO_1169 (O_1169,N_8247,N_9923);
or UO_1170 (O_1170,N_9605,N_9579);
and UO_1171 (O_1171,N_9074,N_8188);
nor UO_1172 (O_1172,N_8503,N_8776);
and UO_1173 (O_1173,N_9136,N_8416);
and UO_1174 (O_1174,N_9779,N_8361);
nor UO_1175 (O_1175,N_8526,N_8817);
xnor UO_1176 (O_1176,N_8954,N_8525);
nor UO_1177 (O_1177,N_9827,N_8552);
nand UO_1178 (O_1178,N_9003,N_9060);
and UO_1179 (O_1179,N_9382,N_8919);
xnor UO_1180 (O_1180,N_9267,N_8494);
or UO_1181 (O_1181,N_8132,N_8509);
xor UO_1182 (O_1182,N_8108,N_9489);
nor UO_1183 (O_1183,N_9702,N_9066);
nand UO_1184 (O_1184,N_9581,N_8254);
xor UO_1185 (O_1185,N_8384,N_8136);
and UO_1186 (O_1186,N_9954,N_8646);
or UO_1187 (O_1187,N_8709,N_9948);
nor UO_1188 (O_1188,N_9472,N_9613);
or UO_1189 (O_1189,N_8923,N_9503);
xor UO_1190 (O_1190,N_9309,N_8430);
nand UO_1191 (O_1191,N_8293,N_8956);
nand UO_1192 (O_1192,N_8893,N_8170);
nor UO_1193 (O_1193,N_9594,N_9524);
nand UO_1194 (O_1194,N_9927,N_8225);
nor UO_1195 (O_1195,N_8493,N_9707);
xor UO_1196 (O_1196,N_9388,N_9462);
nor UO_1197 (O_1197,N_9674,N_9507);
nor UO_1198 (O_1198,N_8961,N_8731);
nor UO_1199 (O_1199,N_8868,N_8001);
nor UO_1200 (O_1200,N_8670,N_8960);
and UO_1201 (O_1201,N_8603,N_8400);
or UO_1202 (O_1202,N_8936,N_8004);
xnor UO_1203 (O_1203,N_8752,N_8991);
nor UO_1204 (O_1204,N_8294,N_8792);
nor UO_1205 (O_1205,N_8304,N_9300);
nor UO_1206 (O_1206,N_8134,N_9872);
and UO_1207 (O_1207,N_9642,N_9989);
nor UO_1208 (O_1208,N_9274,N_8517);
and UO_1209 (O_1209,N_9809,N_9316);
xnor UO_1210 (O_1210,N_8900,N_9513);
xnor UO_1211 (O_1211,N_9833,N_9106);
nor UO_1212 (O_1212,N_9585,N_9122);
or UO_1213 (O_1213,N_9666,N_9013);
and UO_1214 (O_1214,N_8753,N_8378);
nor UO_1215 (O_1215,N_9906,N_8823);
nor UO_1216 (O_1216,N_8221,N_8296);
nand UO_1217 (O_1217,N_9944,N_9221);
or UO_1218 (O_1218,N_8057,N_9189);
xnor UO_1219 (O_1219,N_8304,N_9406);
nand UO_1220 (O_1220,N_9260,N_8253);
nor UO_1221 (O_1221,N_9800,N_9209);
xor UO_1222 (O_1222,N_9530,N_9484);
nor UO_1223 (O_1223,N_8573,N_9570);
nor UO_1224 (O_1224,N_9750,N_8897);
nor UO_1225 (O_1225,N_9984,N_9840);
and UO_1226 (O_1226,N_8952,N_9760);
nor UO_1227 (O_1227,N_8702,N_9189);
nor UO_1228 (O_1228,N_9388,N_9791);
nand UO_1229 (O_1229,N_8374,N_8465);
nor UO_1230 (O_1230,N_9857,N_8581);
and UO_1231 (O_1231,N_9055,N_8512);
nor UO_1232 (O_1232,N_8764,N_8857);
or UO_1233 (O_1233,N_8197,N_9046);
nand UO_1234 (O_1234,N_8102,N_8082);
and UO_1235 (O_1235,N_9928,N_9743);
nand UO_1236 (O_1236,N_8886,N_8139);
nor UO_1237 (O_1237,N_8516,N_8491);
and UO_1238 (O_1238,N_8815,N_8861);
nor UO_1239 (O_1239,N_8689,N_9692);
nor UO_1240 (O_1240,N_8732,N_9089);
nand UO_1241 (O_1241,N_9133,N_9889);
xnor UO_1242 (O_1242,N_9079,N_9945);
or UO_1243 (O_1243,N_8238,N_8485);
and UO_1244 (O_1244,N_8780,N_9897);
nor UO_1245 (O_1245,N_8757,N_9489);
or UO_1246 (O_1246,N_9961,N_8551);
nand UO_1247 (O_1247,N_9777,N_8975);
nor UO_1248 (O_1248,N_9037,N_9837);
and UO_1249 (O_1249,N_8492,N_9568);
nor UO_1250 (O_1250,N_9491,N_9026);
or UO_1251 (O_1251,N_8330,N_8240);
xnor UO_1252 (O_1252,N_8949,N_9940);
nand UO_1253 (O_1253,N_9359,N_8332);
nor UO_1254 (O_1254,N_8595,N_8545);
xor UO_1255 (O_1255,N_8013,N_8317);
nand UO_1256 (O_1256,N_8293,N_8616);
and UO_1257 (O_1257,N_8434,N_8689);
nand UO_1258 (O_1258,N_8748,N_9550);
xnor UO_1259 (O_1259,N_8752,N_9626);
xnor UO_1260 (O_1260,N_8833,N_9899);
xnor UO_1261 (O_1261,N_9763,N_9552);
xor UO_1262 (O_1262,N_9887,N_8247);
and UO_1263 (O_1263,N_8516,N_9841);
or UO_1264 (O_1264,N_8306,N_9276);
or UO_1265 (O_1265,N_9684,N_9136);
and UO_1266 (O_1266,N_8699,N_8749);
nand UO_1267 (O_1267,N_9090,N_9918);
or UO_1268 (O_1268,N_8480,N_8519);
or UO_1269 (O_1269,N_9218,N_9908);
nor UO_1270 (O_1270,N_8646,N_8246);
and UO_1271 (O_1271,N_9097,N_9781);
and UO_1272 (O_1272,N_8874,N_9604);
nand UO_1273 (O_1273,N_9003,N_9567);
or UO_1274 (O_1274,N_9651,N_9659);
nand UO_1275 (O_1275,N_9930,N_8602);
nor UO_1276 (O_1276,N_9021,N_8466);
or UO_1277 (O_1277,N_9098,N_8191);
and UO_1278 (O_1278,N_9791,N_8177);
nand UO_1279 (O_1279,N_8409,N_9910);
and UO_1280 (O_1280,N_9913,N_8544);
and UO_1281 (O_1281,N_9399,N_8594);
or UO_1282 (O_1282,N_9794,N_8924);
or UO_1283 (O_1283,N_8102,N_8353);
nand UO_1284 (O_1284,N_9269,N_9610);
nor UO_1285 (O_1285,N_9374,N_8088);
and UO_1286 (O_1286,N_9557,N_9798);
nor UO_1287 (O_1287,N_8514,N_9850);
nor UO_1288 (O_1288,N_8605,N_8308);
and UO_1289 (O_1289,N_8203,N_8751);
nor UO_1290 (O_1290,N_9677,N_9870);
or UO_1291 (O_1291,N_9516,N_8333);
or UO_1292 (O_1292,N_8916,N_9038);
nand UO_1293 (O_1293,N_8874,N_8518);
nor UO_1294 (O_1294,N_8162,N_8090);
nor UO_1295 (O_1295,N_8980,N_8428);
nand UO_1296 (O_1296,N_8012,N_8348);
nand UO_1297 (O_1297,N_8458,N_9537);
or UO_1298 (O_1298,N_8673,N_9428);
or UO_1299 (O_1299,N_9310,N_8423);
nand UO_1300 (O_1300,N_9504,N_8748);
nor UO_1301 (O_1301,N_9722,N_9730);
nand UO_1302 (O_1302,N_9374,N_8736);
nand UO_1303 (O_1303,N_9087,N_8424);
nor UO_1304 (O_1304,N_8684,N_9985);
and UO_1305 (O_1305,N_8412,N_8346);
or UO_1306 (O_1306,N_8745,N_9912);
nor UO_1307 (O_1307,N_8678,N_8648);
or UO_1308 (O_1308,N_8523,N_9503);
or UO_1309 (O_1309,N_9936,N_9728);
and UO_1310 (O_1310,N_8265,N_9661);
and UO_1311 (O_1311,N_8504,N_9721);
or UO_1312 (O_1312,N_9142,N_8386);
nand UO_1313 (O_1313,N_8166,N_9965);
nor UO_1314 (O_1314,N_9359,N_8527);
and UO_1315 (O_1315,N_9611,N_8032);
nor UO_1316 (O_1316,N_9755,N_8712);
nand UO_1317 (O_1317,N_9020,N_8225);
nand UO_1318 (O_1318,N_8160,N_9110);
nand UO_1319 (O_1319,N_8682,N_9530);
nor UO_1320 (O_1320,N_9013,N_9422);
nand UO_1321 (O_1321,N_9936,N_8329);
or UO_1322 (O_1322,N_8183,N_9357);
nand UO_1323 (O_1323,N_9748,N_8941);
nand UO_1324 (O_1324,N_8527,N_8854);
nand UO_1325 (O_1325,N_9441,N_9332);
nor UO_1326 (O_1326,N_9446,N_9188);
or UO_1327 (O_1327,N_9811,N_8513);
or UO_1328 (O_1328,N_8598,N_9910);
nand UO_1329 (O_1329,N_8364,N_9936);
nor UO_1330 (O_1330,N_9730,N_9941);
nor UO_1331 (O_1331,N_8356,N_9479);
nand UO_1332 (O_1332,N_9256,N_8320);
nor UO_1333 (O_1333,N_9616,N_9841);
xnor UO_1334 (O_1334,N_9183,N_8885);
nand UO_1335 (O_1335,N_9752,N_9393);
nor UO_1336 (O_1336,N_8643,N_8254);
and UO_1337 (O_1337,N_9367,N_8795);
and UO_1338 (O_1338,N_9916,N_8172);
nand UO_1339 (O_1339,N_9167,N_9847);
or UO_1340 (O_1340,N_8750,N_9090);
or UO_1341 (O_1341,N_9884,N_9044);
or UO_1342 (O_1342,N_9388,N_9018);
and UO_1343 (O_1343,N_8117,N_8063);
or UO_1344 (O_1344,N_9742,N_9494);
and UO_1345 (O_1345,N_9086,N_8426);
or UO_1346 (O_1346,N_8176,N_9087);
nand UO_1347 (O_1347,N_8130,N_9691);
nor UO_1348 (O_1348,N_8702,N_8451);
xor UO_1349 (O_1349,N_9177,N_8533);
xor UO_1350 (O_1350,N_9660,N_8339);
and UO_1351 (O_1351,N_8185,N_9984);
xnor UO_1352 (O_1352,N_8366,N_8884);
nor UO_1353 (O_1353,N_8224,N_9187);
or UO_1354 (O_1354,N_9532,N_9138);
and UO_1355 (O_1355,N_8042,N_9099);
nand UO_1356 (O_1356,N_8638,N_9630);
nor UO_1357 (O_1357,N_8205,N_8673);
nor UO_1358 (O_1358,N_9615,N_9845);
nand UO_1359 (O_1359,N_9351,N_8515);
and UO_1360 (O_1360,N_9859,N_8153);
and UO_1361 (O_1361,N_9515,N_9029);
and UO_1362 (O_1362,N_9391,N_8029);
nor UO_1363 (O_1363,N_9084,N_9502);
nand UO_1364 (O_1364,N_9348,N_8709);
nand UO_1365 (O_1365,N_8430,N_8306);
nand UO_1366 (O_1366,N_8058,N_9311);
nor UO_1367 (O_1367,N_9490,N_8360);
nor UO_1368 (O_1368,N_9280,N_9761);
or UO_1369 (O_1369,N_8425,N_8359);
nand UO_1370 (O_1370,N_8100,N_9658);
nor UO_1371 (O_1371,N_8090,N_9847);
or UO_1372 (O_1372,N_8485,N_9021);
or UO_1373 (O_1373,N_8500,N_9959);
nor UO_1374 (O_1374,N_8469,N_9979);
and UO_1375 (O_1375,N_8384,N_8171);
nand UO_1376 (O_1376,N_9559,N_8674);
nand UO_1377 (O_1377,N_9169,N_9845);
nor UO_1378 (O_1378,N_9583,N_9492);
and UO_1379 (O_1379,N_8110,N_9645);
or UO_1380 (O_1380,N_8680,N_8364);
or UO_1381 (O_1381,N_8569,N_9249);
xor UO_1382 (O_1382,N_9632,N_8720);
nand UO_1383 (O_1383,N_9763,N_9803);
and UO_1384 (O_1384,N_9466,N_9946);
nand UO_1385 (O_1385,N_8108,N_8444);
nand UO_1386 (O_1386,N_9433,N_8725);
or UO_1387 (O_1387,N_9371,N_8632);
xor UO_1388 (O_1388,N_9079,N_9788);
and UO_1389 (O_1389,N_9751,N_9156);
and UO_1390 (O_1390,N_8936,N_9269);
and UO_1391 (O_1391,N_9142,N_8610);
and UO_1392 (O_1392,N_9676,N_8102);
nand UO_1393 (O_1393,N_8833,N_8681);
or UO_1394 (O_1394,N_9084,N_8895);
nand UO_1395 (O_1395,N_8135,N_9407);
xnor UO_1396 (O_1396,N_8314,N_9649);
nand UO_1397 (O_1397,N_9090,N_9634);
or UO_1398 (O_1398,N_8565,N_8402);
nand UO_1399 (O_1399,N_9017,N_8276);
nand UO_1400 (O_1400,N_9463,N_8011);
and UO_1401 (O_1401,N_8517,N_9893);
nand UO_1402 (O_1402,N_9575,N_9994);
xnor UO_1403 (O_1403,N_8534,N_9995);
or UO_1404 (O_1404,N_9015,N_8660);
and UO_1405 (O_1405,N_8894,N_9084);
nor UO_1406 (O_1406,N_9859,N_9166);
or UO_1407 (O_1407,N_8866,N_8105);
nand UO_1408 (O_1408,N_9428,N_8061);
and UO_1409 (O_1409,N_8252,N_8491);
nor UO_1410 (O_1410,N_9488,N_8807);
or UO_1411 (O_1411,N_9142,N_8289);
nand UO_1412 (O_1412,N_8337,N_9321);
or UO_1413 (O_1413,N_9236,N_8922);
or UO_1414 (O_1414,N_8068,N_8019);
nor UO_1415 (O_1415,N_8154,N_8534);
or UO_1416 (O_1416,N_8185,N_8465);
nor UO_1417 (O_1417,N_8187,N_8720);
nand UO_1418 (O_1418,N_8738,N_9140);
or UO_1419 (O_1419,N_8049,N_9195);
nor UO_1420 (O_1420,N_9956,N_9288);
xor UO_1421 (O_1421,N_8228,N_8035);
or UO_1422 (O_1422,N_8255,N_9803);
or UO_1423 (O_1423,N_9559,N_9557);
nand UO_1424 (O_1424,N_9256,N_8102);
and UO_1425 (O_1425,N_8405,N_9891);
and UO_1426 (O_1426,N_8947,N_9129);
and UO_1427 (O_1427,N_9455,N_8572);
or UO_1428 (O_1428,N_9678,N_9779);
nor UO_1429 (O_1429,N_8731,N_8968);
and UO_1430 (O_1430,N_8302,N_9713);
and UO_1431 (O_1431,N_9016,N_8925);
or UO_1432 (O_1432,N_9121,N_9289);
and UO_1433 (O_1433,N_9709,N_9962);
nand UO_1434 (O_1434,N_9704,N_8887);
nor UO_1435 (O_1435,N_8059,N_9915);
and UO_1436 (O_1436,N_8190,N_8539);
nor UO_1437 (O_1437,N_9116,N_8531);
or UO_1438 (O_1438,N_9473,N_9959);
and UO_1439 (O_1439,N_9676,N_9490);
and UO_1440 (O_1440,N_9582,N_9942);
or UO_1441 (O_1441,N_8529,N_8477);
or UO_1442 (O_1442,N_8706,N_9073);
and UO_1443 (O_1443,N_9896,N_9169);
or UO_1444 (O_1444,N_8743,N_9668);
nor UO_1445 (O_1445,N_8128,N_9789);
and UO_1446 (O_1446,N_8464,N_8712);
and UO_1447 (O_1447,N_9521,N_9529);
nor UO_1448 (O_1448,N_9341,N_9674);
and UO_1449 (O_1449,N_9518,N_8428);
nand UO_1450 (O_1450,N_8525,N_8145);
xnor UO_1451 (O_1451,N_9684,N_9578);
nor UO_1452 (O_1452,N_9101,N_8111);
nand UO_1453 (O_1453,N_8672,N_8267);
nand UO_1454 (O_1454,N_8031,N_8000);
or UO_1455 (O_1455,N_9404,N_9852);
nor UO_1456 (O_1456,N_8028,N_9505);
nor UO_1457 (O_1457,N_8662,N_8955);
or UO_1458 (O_1458,N_8661,N_9269);
or UO_1459 (O_1459,N_9024,N_9468);
and UO_1460 (O_1460,N_8168,N_8165);
or UO_1461 (O_1461,N_9730,N_9747);
and UO_1462 (O_1462,N_8377,N_8199);
and UO_1463 (O_1463,N_8085,N_9888);
xor UO_1464 (O_1464,N_8060,N_9129);
nor UO_1465 (O_1465,N_8186,N_9378);
nand UO_1466 (O_1466,N_8517,N_8047);
or UO_1467 (O_1467,N_9991,N_8469);
xnor UO_1468 (O_1468,N_9805,N_8667);
and UO_1469 (O_1469,N_9721,N_9815);
nand UO_1470 (O_1470,N_9475,N_9024);
or UO_1471 (O_1471,N_8822,N_9354);
nand UO_1472 (O_1472,N_9835,N_8515);
and UO_1473 (O_1473,N_8405,N_8318);
nor UO_1474 (O_1474,N_8026,N_8727);
or UO_1475 (O_1475,N_9678,N_9735);
or UO_1476 (O_1476,N_9381,N_9551);
and UO_1477 (O_1477,N_9659,N_8533);
nand UO_1478 (O_1478,N_8653,N_8376);
or UO_1479 (O_1479,N_9737,N_9987);
and UO_1480 (O_1480,N_8312,N_8701);
or UO_1481 (O_1481,N_9204,N_8703);
or UO_1482 (O_1482,N_8763,N_8355);
nor UO_1483 (O_1483,N_9422,N_8494);
nand UO_1484 (O_1484,N_8857,N_9147);
or UO_1485 (O_1485,N_8163,N_8761);
and UO_1486 (O_1486,N_9826,N_9893);
xnor UO_1487 (O_1487,N_9094,N_9071);
nor UO_1488 (O_1488,N_8380,N_9428);
nor UO_1489 (O_1489,N_8219,N_8270);
xor UO_1490 (O_1490,N_9527,N_9502);
nand UO_1491 (O_1491,N_9266,N_8918);
or UO_1492 (O_1492,N_9740,N_9737);
and UO_1493 (O_1493,N_9802,N_9093);
nor UO_1494 (O_1494,N_9711,N_8503);
nand UO_1495 (O_1495,N_9345,N_8419);
nand UO_1496 (O_1496,N_8195,N_9477);
nor UO_1497 (O_1497,N_8576,N_9471);
nor UO_1498 (O_1498,N_8248,N_9475);
nand UO_1499 (O_1499,N_8233,N_9573);
endmodule