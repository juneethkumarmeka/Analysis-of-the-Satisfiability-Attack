module basic_1500_15000_2000_60_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nor U0 (N_0,In_365,In_102);
xnor U1 (N_1,In_1468,In_1274);
or U2 (N_2,In_261,In_756);
or U3 (N_3,In_575,In_717);
xor U4 (N_4,In_672,In_948);
nor U5 (N_5,In_646,In_778);
nor U6 (N_6,In_1341,In_801);
or U7 (N_7,In_293,In_803);
xor U8 (N_8,In_1441,In_1267);
and U9 (N_9,In_306,In_14);
nor U10 (N_10,In_1297,In_219);
xor U11 (N_11,In_713,In_125);
xor U12 (N_12,In_602,In_1426);
and U13 (N_13,In_753,In_1);
xor U14 (N_14,In_1478,In_168);
nand U15 (N_15,In_60,In_483);
and U16 (N_16,In_586,In_104);
nand U17 (N_17,In_1256,In_820);
xnor U18 (N_18,In_360,In_204);
xor U19 (N_19,In_66,In_662);
nor U20 (N_20,In_1474,In_1170);
nor U21 (N_21,In_1043,In_487);
nand U22 (N_22,In_96,In_1449);
or U23 (N_23,In_550,In_1091);
xnor U24 (N_24,In_540,In_749);
or U25 (N_25,In_880,In_546);
and U26 (N_26,In_775,In_918);
nand U27 (N_27,In_0,In_827);
nand U28 (N_28,In_1015,In_526);
or U29 (N_29,In_908,In_997);
or U30 (N_30,In_859,In_659);
or U31 (N_31,In_989,In_9);
or U32 (N_32,In_971,In_1296);
nor U33 (N_33,In_448,In_1487);
nor U34 (N_34,In_75,In_1239);
xnor U35 (N_35,In_349,In_1044);
xor U36 (N_36,In_561,In_501);
nor U37 (N_37,In_435,In_1188);
or U38 (N_38,In_33,In_1032);
nor U39 (N_39,In_887,In_845);
nor U40 (N_40,In_1454,In_326);
xnor U41 (N_41,In_488,In_509);
and U42 (N_42,In_1158,In_32);
or U43 (N_43,In_673,In_267);
nor U44 (N_44,In_1068,In_245);
nor U45 (N_45,In_996,In_490);
or U46 (N_46,In_199,In_1038);
or U47 (N_47,In_1176,In_190);
nor U48 (N_48,In_1471,In_424);
xnor U49 (N_49,In_519,In_76);
xnor U50 (N_50,In_122,In_1412);
xnor U51 (N_51,In_22,In_171);
or U52 (N_52,In_841,In_1151);
or U53 (N_53,In_904,In_923);
and U54 (N_54,In_1258,In_825);
nand U55 (N_55,In_1271,In_158);
nor U56 (N_56,In_1185,In_534);
nor U57 (N_57,In_416,In_1499);
and U58 (N_58,In_977,In_998);
nand U59 (N_59,In_1241,In_543);
nand U60 (N_60,In_1086,In_1000);
xnor U61 (N_61,In_191,In_1458);
and U62 (N_62,In_731,In_1421);
nor U63 (N_63,In_1154,In_134);
nand U64 (N_64,In_1446,In_671);
xor U65 (N_65,In_352,In_1025);
xnor U66 (N_66,In_1228,In_1148);
nor U67 (N_67,In_276,In_517);
and U68 (N_68,In_186,In_185);
or U69 (N_69,In_447,In_231);
nand U70 (N_70,In_202,In_1214);
and U71 (N_71,In_955,In_625);
xnor U72 (N_72,In_115,In_356);
nand U73 (N_73,In_271,In_1269);
nand U74 (N_74,In_1378,In_761);
or U75 (N_75,In_425,In_1019);
or U76 (N_76,In_938,In_763);
nor U77 (N_77,In_111,In_421);
xnor U78 (N_78,In_1257,In_1098);
nand U79 (N_79,In_497,In_1428);
or U80 (N_80,In_1021,In_711);
nor U81 (N_81,In_117,In_1051);
xor U82 (N_82,In_994,In_402);
and U83 (N_83,In_610,In_751);
or U84 (N_84,In_1074,In_1444);
nand U85 (N_85,In_824,In_319);
and U86 (N_86,In_536,In_198);
xor U87 (N_87,In_605,In_1096);
nand U88 (N_88,In_640,In_1222);
or U89 (N_89,In_736,In_936);
and U90 (N_90,In_757,In_1358);
nor U91 (N_91,In_1295,In_817);
nor U92 (N_92,In_1122,In_462);
or U93 (N_93,In_655,In_1392);
and U94 (N_94,In_818,In_1160);
nand U95 (N_95,In_1276,In_995);
nor U96 (N_96,In_153,In_338);
xnor U97 (N_97,In_1009,In_1182);
and U98 (N_98,In_325,In_725);
nand U99 (N_99,In_544,In_706);
nand U100 (N_100,In_260,In_684);
or U101 (N_101,In_240,In_1340);
or U102 (N_102,In_792,In_24);
or U103 (N_103,In_1242,In_188);
xnor U104 (N_104,In_1356,In_1233);
nand U105 (N_105,In_742,In_892);
nor U106 (N_106,In_926,In_438);
and U107 (N_107,In_1061,In_676);
and U108 (N_108,In_558,In_595);
nor U109 (N_109,In_929,In_888);
nand U110 (N_110,In_906,In_836);
or U111 (N_111,In_1461,In_74);
nand U112 (N_112,In_1435,In_846);
nor U113 (N_113,In_1060,In_280);
and U114 (N_114,In_1005,In_133);
nand U115 (N_115,In_499,In_155);
or U116 (N_116,In_414,In_1328);
xnor U117 (N_117,In_300,In_291);
nand U118 (N_118,In_982,In_287);
nor U119 (N_119,In_807,In_463);
nor U120 (N_120,In_148,In_62);
nor U121 (N_121,In_745,In_1357);
or U122 (N_122,In_1490,In_848);
nand U123 (N_123,In_1157,In_468);
nand U124 (N_124,In_166,In_1101);
and U125 (N_125,In_677,In_537);
nand U126 (N_126,In_735,In_1393);
nor U127 (N_127,In_1293,In_1459);
nor U128 (N_128,In_697,In_522);
or U129 (N_129,In_406,In_1350);
and U130 (N_130,In_227,In_486);
xor U131 (N_131,In_1094,In_1429);
or U132 (N_132,In_780,In_964);
or U133 (N_133,In_1305,In_128);
or U134 (N_134,In_1013,In_195);
or U135 (N_135,In_738,In_1385);
xnor U136 (N_136,In_978,In_632);
nand U137 (N_137,In_683,In_8);
or U138 (N_138,In_312,In_376);
and U139 (N_139,In_1118,In_1354);
xor U140 (N_140,In_456,In_467);
xnor U141 (N_141,In_71,In_1466);
xnor U142 (N_142,In_296,In_1294);
nor U143 (N_143,In_216,In_135);
nor U144 (N_144,In_515,In_1221);
and U145 (N_145,In_867,In_965);
and U146 (N_146,In_787,In_1431);
or U147 (N_147,In_443,In_89);
or U148 (N_148,In_307,In_710);
nor U149 (N_149,In_579,In_1041);
nor U150 (N_150,In_180,In_855);
nor U151 (N_151,In_644,In_1273);
nor U152 (N_152,In_73,In_85);
nor U153 (N_153,In_510,In_1376);
and U154 (N_154,In_895,In_1367);
or U155 (N_155,In_1407,In_1310);
xor U156 (N_156,In_1093,In_112);
xnor U157 (N_157,In_136,In_350);
nand U158 (N_158,In_1187,In_1161);
nor U159 (N_159,In_728,In_65);
nor U160 (N_160,In_819,In_353);
nand U161 (N_161,In_1220,In_1488);
xor U162 (N_162,In_698,In_371);
nand U163 (N_163,In_653,In_516);
or U164 (N_164,In_1075,In_839);
and U165 (N_165,In_123,In_1402);
and U166 (N_166,In_35,In_194);
xor U167 (N_167,In_1083,In_680);
nand U168 (N_168,In_466,In_1362);
xor U169 (N_169,In_113,In_103);
and U170 (N_170,In_452,In_985);
nor U171 (N_171,In_1339,In_847);
nand U172 (N_172,In_1131,In_583);
nand U173 (N_173,In_740,In_1497);
or U174 (N_174,In_1252,In_1448);
xnor U175 (N_175,In_284,In_601);
nand U176 (N_176,In_1304,In_916);
xnor U177 (N_177,In_782,In_1189);
and U178 (N_178,In_802,In_1262);
and U179 (N_179,In_1453,In_1047);
xnor U180 (N_180,In_1349,In_54);
or U181 (N_181,In_562,In_1351);
nor U182 (N_182,In_105,In_866);
nand U183 (N_183,In_1120,In_1181);
or U184 (N_184,In_437,In_345);
nand U185 (N_185,In_1040,In_991);
xnor U186 (N_186,In_256,In_1134);
xor U187 (N_187,In_26,In_1240);
nand U188 (N_188,In_570,In_639);
and U189 (N_189,In_1218,In_962);
and U190 (N_190,In_243,In_531);
nand U191 (N_191,In_156,In_176);
and U192 (N_192,In_864,In_1482);
nor U193 (N_193,In_232,In_981);
nor U194 (N_194,In_367,In_1265);
xnor U195 (N_195,In_167,In_1494);
or U196 (N_196,In_603,In_715);
and U197 (N_197,In_477,In_741);
nand U198 (N_198,In_637,In_157);
and U199 (N_199,In_44,In_832);
or U200 (N_200,In_1192,In_934);
xor U201 (N_201,In_246,In_142);
xor U202 (N_202,In_795,In_804);
xnor U203 (N_203,In_1004,In_1145);
nand U204 (N_204,In_1206,In_210);
nand U205 (N_205,In_1484,In_82);
nand U206 (N_206,In_337,In_831);
nor U207 (N_207,In_1219,In_712);
xnor U208 (N_208,In_1470,In_1331);
xnor U209 (N_209,In_69,In_170);
nand U210 (N_210,In_828,In_652);
nor U211 (N_211,In_1066,In_752);
nand U212 (N_212,In_1398,In_449);
nand U213 (N_213,In_886,In_169);
or U214 (N_214,In_1423,In_1103);
nor U215 (N_215,In_1057,In_611);
and U216 (N_216,In_10,In_798);
nand U217 (N_217,In_389,In_29);
or U218 (N_218,In_301,In_410);
nor U219 (N_219,In_1390,In_619);
nand U220 (N_220,In_346,In_1442);
and U221 (N_221,In_907,In_242);
xnor U222 (N_222,In_399,In_254);
and U223 (N_223,In_21,In_333);
nand U224 (N_224,In_1493,In_1226);
or U225 (N_225,In_1389,In_784);
or U226 (N_226,In_173,In_891);
nand U227 (N_227,In_1266,In_1202);
xor U228 (N_228,In_568,In_302);
and U229 (N_229,In_485,In_1072);
and U230 (N_230,In_699,In_1410);
xnor U231 (N_231,In_623,In_1234);
nand U232 (N_232,In_496,In_1300);
nand U233 (N_233,In_1380,In_701);
nor U234 (N_234,In_723,In_77);
and U235 (N_235,In_951,In_705);
nand U236 (N_236,In_1236,In_1455);
nor U237 (N_237,In_1396,In_1095);
or U238 (N_238,In_110,In_282);
and U239 (N_239,In_471,In_53);
and U240 (N_240,In_1383,In_229);
and U241 (N_241,In_461,In_45);
nor U242 (N_242,In_631,In_61);
and U243 (N_243,In_1191,In_1472);
or U244 (N_244,In_734,In_643);
xnor U245 (N_245,In_1028,In_620);
nand U246 (N_246,In_1238,In_324);
or U247 (N_247,In_1143,In_283);
nor U248 (N_248,In_1321,In_944);
nor U249 (N_249,In_732,In_857);
nor U250 (N_250,N_103,In_249);
and U251 (N_251,In_1338,In_766);
nor U252 (N_252,N_210,In_132);
or U253 (N_253,In_1084,In_48);
or U254 (N_254,In_890,N_161);
xor U255 (N_255,In_590,In_1137);
or U256 (N_256,In_221,N_213);
nand U257 (N_257,N_187,In_392);
or U258 (N_258,In_812,In_862);
nor U259 (N_259,N_160,In_1116);
nor U260 (N_260,In_656,In_1058);
and U261 (N_261,N_104,N_232);
nor U262 (N_262,In_236,In_95);
nor U263 (N_263,In_1301,In_1159);
nand U264 (N_264,In_1400,In_174);
nor U265 (N_265,In_557,In_1204);
xor U266 (N_266,In_386,In_1011);
xnor U267 (N_267,N_229,N_102);
nor U268 (N_268,In_1250,In_149);
nor U269 (N_269,N_57,In_559);
and U270 (N_270,In_355,N_117);
or U271 (N_271,N_234,In_1078);
or U272 (N_272,N_167,In_1313);
or U273 (N_273,In_714,In_52);
and U274 (N_274,In_472,In_881);
nor U275 (N_275,In_1055,In_16);
xnor U276 (N_276,In_151,In_638);
and U277 (N_277,In_937,In_1409);
nand U278 (N_278,In_1169,In_469);
nor U279 (N_279,In_1209,N_189);
xnor U280 (N_280,N_84,In_813);
or U281 (N_281,In_618,N_176);
or U282 (N_282,In_913,N_190);
and U283 (N_283,In_838,In_413);
nor U284 (N_284,In_629,N_67);
or U285 (N_285,In_793,In_903);
nand U286 (N_286,In_492,In_373);
nor U287 (N_287,In_919,In_844);
or U288 (N_288,In_1018,In_459);
or U289 (N_289,N_123,In_422);
and U290 (N_290,In_315,In_730);
or U291 (N_291,In_806,In_834);
nor U292 (N_292,N_24,In_457);
xor U293 (N_293,In_564,In_313);
and U294 (N_294,In_107,In_237);
nor U295 (N_295,In_40,In_341);
or U296 (N_296,N_108,In_850);
xnor U297 (N_297,In_121,In_799);
xnor U298 (N_298,In_1016,In_1027);
nand U299 (N_299,In_874,In_1345);
or U300 (N_300,In_893,In_1439);
or U301 (N_301,In_476,In_815);
and U302 (N_302,In_87,In_984);
and U303 (N_303,N_72,In_896);
xor U304 (N_304,In_647,N_248);
nor U305 (N_305,In_184,In_733);
xor U306 (N_306,N_247,In_691);
and U307 (N_307,N_40,In_114);
xor U308 (N_308,In_130,In_1088);
and U309 (N_309,In_220,N_60);
and U310 (N_310,In_598,In_947);
nand U311 (N_311,N_159,In_1332);
nand U312 (N_312,In_327,N_86);
and U313 (N_313,In_1024,In_587);
and U314 (N_314,N_3,N_147);
nand U315 (N_315,In_608,In_56);
or U316 (N_316,N_240,N_95);
xnor U317 (N_317,In_1001,In_1397);
nand U318 (N_318,In_1081,In_750);
or U319 (N_319,In_1465,In_591);
xnor U320 (N_320,In_46,In_1405);
nor U321 (N_321,In_621,In_1141);
nand U322 (N_322,N_39,In_1142);
and U323 (N_323,In_1244,In_1417);
and U324 (N_324,N_99,In_606);
nor U325 (N_325,In_1387,In_525);
nand U326 (N_326,In_1285,In_484);
and U327 (N_327,In_574,In_1288);
nor U328 (N_328,In_318,N_74);
xor U329 (N_329,N_208,N_51);
or U330 (N_330,In_634,In_172);
xnor U331 (N_331,In_385,In_299);
xor U332 (N_332,In_1388,In_811);
nand U333 (N_333,In_147,In_1370);
nor U334 (N_334,N_46,In_573);
xor U335 (N_335,In_152,N_106);
xnor U336 (N_336,N_120,In_1291);
nand U337 (N_337,In_797,In_15);
or U338 (N_338,In_175,In_94);
or U339 (N_339,N_249,In_286);
xor U340 (N_340,N_219,In_718);
xnor U341 (N_341,In_1100,In_80);
nor U342 (N_342,In_661,In_900);
xor U343 (N_343,In_1379,In_1440);
xor U344 (N_344,In_1012,N_134);
and U345 (N_345,In_165,In_1309);
nor U346 (N_346,In_1199,N_90);
nor U347 (N_347,In_635,In_1007);
or U348 (N_348,N_56,In_1017);
nor U349 (N_349,In_1163,In_241);
xnor U350 (N_350,In_1064,In_569);
or U351 (N_351,N_12,N_127);
or U352 (N_352,In_1498,In_379);
or U353 (N_353,N_244,In_1030);
and U354 (N_354,In_571,In_143);
and U355 (N_355,In_1014,In_933);
and U356 (N_356,In_228,In_396);
nand U357 (N_357,N_76,In_342);
and U358 (N_358,N_54,In_1034);
and U359 (N_359,In_833,N_94);
or U360 (N_360,In_589,In_905);
and U361 (N_361,In_1133,N_170);
or U362 (N_362,N_9,N_111);
or U363 (N_363,N_88,In_1469);
or U364 (N_364,N_13,In_78);
and U365 (N_365,In_578,In_1196);
or U366 (N_366,In_1165,In_514);
and U367 (N_367,In_2,In_1418);
nor U368 (N_368,In_269,N_238);
and U369 (N_369,In_37,In_853);
nor U370 (N_370,In_952,In_975);
and U371 (N_371,In_511,In_1201);
xor U372 (N_372,In_144,In_303);
nand U373 (N_373,In_1261,N_156);
or U374 (N_374,In_791,In_1283);
xor U375 (N_375,In_1422,In_259);
or U376 (N_376,In_209,In_940);
and U377 (N_377,In_856,N_6);
xnor U378 (N_378,In_682,In_1205);
nand U379 (N_379,In_34,In_967);
or U380 (N_380,In_719,In_776);
and U381 (N_381,In_141,In_1114);
nand U382 (N_382,In_30,In_1436);
nand U383 (N_383,N_192,In_1255);
nand U384 (N_384,In_458,In_599);
or U385 (N_385,In_1290,In_1303);
and U386 (N_386,N_23,N_38);
or U387 (N_387,In_835,In_781);
and U388 (N_388,In_1085,In_860);
and U389 (N_389,In_320,In_547);
and U390 (N_390,In_902,N_124);
or U391 (N_391,In_138,In_555);
and U392 (N_392,N_169,N_145);
and U393 (N_393,N_175,In_116);
nand U394 (N_394,In_247,In_275);
and U395 (N_395,In_878,N_100);
nand U396 (N_396,In_108,In_678);
nor U397 (N_397,N_201,In_943);
and U398 (N_398,In_446,In_685);
and U399 (N_399,In_532,In_1366);
and U400 (N_400,In_1106,In_63);
or U401 (N_401,N_197,In_1144);
xnor U402 (N_402,In_1419,In_1113);
xnor U403 (N_403,In_145,In_378);
xor U404 (N_404,In_1208,In_362);
nand U405 (N_405,In_339,N_8);
xnor U406 (N_406,In_481,In_106);
xor U407 (N_407,In_401,In_411);
nand U408 (N_408,N_81,In_1438);
or U409 (N_409,N_158,N_27);
or U410 (N_410,In_794,In_179);
xor U411 (N_411,In_234,In_1045);
and U412 (N_412,In_716,In_1167);
or U413 (N_413,In_1171,In_1186);
or U414 (N_414,In_97,In_542);
and U415 (N_415,In_1275,In_358);
and U416 (N_416,In_1198,N_212);
xor U417 (N_417,N_153,In_201);
xor U418 (N_418,In_1399,In_1020);
nand U419 (N_419,In_1010,In_556);
and U420 (N_420,In_1391,N_30);
nand U421 (N_421,N_135,In_257);
and U422 (N_422,In_120,N_49);
and U423 (N_423,N_131,In_1053);
xor U424 (N_424,In_405,In_1483);
nor U425 (N_425,In_1077,In_1433);
or U426 (N_426,N_68,In_268);
nor U427 (N_427,In_36,N_214);
and U428 (N_428,In_1408,In_582);
or U429 (N_429,In_309,In_772);
and U430 (N_430,In_1427,In_505);
nand U431 (N_431,In_987,In_829);
xor U432 (N_432,In_205,N_75);
xor U433 (N_433,In_665,N_221);
and U434 (N_434,In_263,In_789);
or U435 (N_435,In_397,N_227);
xor U436 (N_436,In_1314,In_238);
and U437 (N_437,In_912,In_1336);
nor U438 (N_438,In_1126,In_876);
xor U439 (N_439,In_415,In_999);
and U440 (N_440,In_1462,N_196);
or U441 (N_441,In_533,In_1031);
nand U442 (N_442,N_186,In_921);
and U443 (N_443,In_504,N_15);
or U444 (N_444,In_1211,In_495);
nor U445 (N_445,N_47,In_861);
nor U446 (N_446,In_1212,In_1346);
nand U447 (N_447,In_1052,In_658);
nor U448 (N_448,N_91,In_764);
nand U449 (N_449,In_953,In_626);
nand U450 (N_450,In_1003,In_1215);
and U451 (N_451,In_946,In_1280);
and U452 (N_452,In_429,In_207);
and U453 (N_453,In_681,In_164);
xnor U454 (N_454,In_59,In_674);
and U455 (N_455,In_1002,In_910);
nor U456 (N_456,In_1386,In_1099);
or U457 (N_457,In_593,In_1177);
xnor U458 (N_458,N_33,In_90);
or U459 (N_459,N_178,In_651);
nand U460 (N_460,In_1235,In_774);
xor U461 (N_461,In_258,N_138);
nand U462 (N_462,In_351,In_576);
and U463 (N_463,In_885,In_394);
and U464 (N_464,In_884,In_1056);
nand U465 (N_465,In_1193,In_248);
or U466 (N_466,In_1225,In_99);
and U467 (N_467,In_251,N_226);
nor U468 (N_468,In_270,N_71);
or U469 (N_469,N_133,N_64);
and U470 (N_470,In_292,N_66);
nor U471 (N_471,In_1029,In_931);
nand U472 (N_472,N_115,In_1477);
nor U473 (N_473,In_1135,In_272);
nor U474 (N_474,In_354,In_57);
and U475 (N_475,In_1203,In_528);
xor U476 (N_476,N_207,In_225);
and U477 (N_477,In_668,In_870);
and U478 (N_478,In_18,N_151);
or U479 (N_479,In_928,In_1048);
nand U480 (N_480,In_79,In_1298);
and U481 (N_481,In_686,In_6);
or U482 (N_482,In_821,N_65);
nor U483 (N_483,In_1130,In_88);
nand U484 (N_484,N_10,In_849);
nor U485 (N_485,In_594,In_480);
nor U486 (N_486,In_539,In_398);
nand U487 (N_487,N_92,N_193);
nor U488 (N_488,In_1039,In_941);
nor U489 (N_489,In_1377,In_330);
nand U490 (N_490,In_428,N_183);
xor U491 (N_491,In_426,In_1050);
nor U492 (N_492,N_146,In_983);
or U493 (N_493,In_535,In_612);
nor U494 (N_494,N_137,In_19);
or U495 (N_495,N_7,In_67);
nor U496 (N_496,In_109,In_1432);
nand U497 (N_497,In_729,In_837);
and U498 (N_498,N_16,In_1138);
nand U499 (N_499,N_130,In_1481);
xor U500 (N_500,N_55,In_298);
nor U501 (N_501,In_968,N_465);
nand U502 (N_502,N_411,In_770);
or U503 (N_503,In_317,In_482);
and U504 (N_504,In_1026,In_150);
and U505 (N_505,In_596,In_92);
nor U506 (N_506,N_463,N_431);
xor U507 (N_507,In_622,N_163);
xor U508 (N_508,In_427,N_450);
xnor U509 (N_509,In_1425,N_185);
and U510 (N_510,N_417,In_633);
or U511 (N_511,In_181,N_181);
nor U512 (N_512,In_660,In_1125);
xor U513 (N_513,In_1452,N_306);
xor U514 (N_514,In_1069,In_25);
or U515 (N_515,N_314,In_1327);
xor U516 (N_516,N_492,N_370);
nand U517 (N_517,In_131,In_3);
and U518 (N_518,In_502,In_506);
nand U519 (N_519,In_359,N_343);
nand U520 (N_520,N_430,N_17);
xnor U521 (N_521,In_12,In_1174);
nand U522 (N_522,N_73,In_762);
or U523 (N_523,N_278,N_20);
nor U524 (N_524,In_988,In_830);
or U525 (N_525,N_225,N_474);
xor U526 (N_526,In_1485,In_1368);
nor U527 (N_527,In_1090,In_305);
and U528 (N_528,In_924,N_280);
xor U529 (N_529,N_195,N_171);
and U530 (N_530,In_1355,In_1284);
or U531 (N_531,In_852,N_270);
nand U532 (N_532,In_383,In_911);
or U533 (N_533,N_172,In_1263);
and U534 (N_534,N_263,N_89);
nor U535 (N_535,N_451,N_173);
nand U536 (N_536,In_1318,N_143);
nand U537 (N_537,N_174,In_613);
nand U538 (N_538,N_58,N_155);
xor U539 (N_539,In_974,N_310);
nand U540 (N_540,N_350,In_737);
xnor U541 (N_541,In_669,In_1360);
or U542 (N_542,N_0,N_144);
nor U543 (N_543,N_303,In_491);
or U544 (N_544,In_433,In_161);
xnor U545 (N_545,In_945,In_917);
nand U546 (N_546,In_577,In_1067);
xnor U547 (N_547,In_206,In_239);
and U548 (N_548,In_347,In_688);
nor U549 (N_549,In_391,N_479);
nand U550 (N_550,In_1123,In_1112);
xor U551 (N_551,In_1479,In_1375);
xor U552 (N_552,In_213,In_1374);
xor U553 (N_553,In_1382,In_786);
and U554 (N_554,In_439,N_45);
or U555 (N_555,In_523,In_43);
and U556 (N_556,In_790,In_1316);
nand U557 (N_557,In_1173,In_873);
nand U558 (N_558,In_879,In_768);
and U559 (N_559,In_530,N_475);
xnor U560 (N_560,In_1230,N_43);
or U561 (N_561,N_157,In_524);
xnor U562 (N_562,N_85,N_446);
nand U563 (N_563,N_152,N_347);
nor U564 (N_564,In_1080,In_1268);
nor U565 (N_565,In_580,N_11);
and U566 (N_566,N_481,In_1270);
nand U567 (N_567,N_467,In_666);
xor U568 (N_568,In_777,In_529);
or U569 (N_569,In_545,In_454);
or U570 (N_570,In_279,In_507);
or U571 (N_571,In_1243,In_636);
xnor U572 (N_572,N_373,In_17);
or U573 (N_573,In_494,In_1352);
xor U574 (N_574,In_217,In_865);
or U575 (N_575,N_35,In_1249);
and U576 (N_576,In_381,N_129);
or U577 (N_577,N_285,In_1348);
xor U578 (N_578,In_553,In_211);
or U579 (N_579,In_1333,In_1264);
xor U580 (N_580,In_973,In_563);
nand U581 (N_581,In_1248,In_1292);
nor U582 (N_582,N_447,In_192);
xnor U583 (N_583,In_869,N_426);
nand U584 (N_584,In_1254,In_473);
nor U585 (N_585,N_281,In_939);
and U586 (N_586,In_990,N_489);
xnor U587 (N_587,N_202,N_419);
and U588 (N_588,N_482,In_1330);
nor U589 (N_589,N_237,N_37);
nand U590 (N_590,In_343,In_722);
nor U591 (N_591,N_460,N_407);
nand U592 (N_592,In_538,In_645);
xor U593 (N_593,In_627,In_465);
xor U594 (N_594,N_259,In_597);
and U595 (N_595,In_868,In_445);
nand U596 (N_596,In_915,In_1115);
nor U597 (N_597,In_160,N_177);
nand U598 (N_598,N_220,N_387);
nor U599 (N_599,N_455,N_401);
xnor U600 (N_600,N_262,In_370);
xnor U601 (N_601,N_114,In_1092);
xor U602 (N_602,N_400,In_146);
or U603 (N_603,In_1184,In_255);
nor U604 (N_604,In_1152,N_142);
and U605 (N_605,In_475,In_288);
and U606 (N_606,N_434,In_289);
xnor U607 (N_607,In_1054,N_415);
and U608 (N_608,In_58,In_375);
and U609 (N_609,N_368,In_901);
nand U610 (N_610,In_440,N_253);
nand U611 (N_611,N_78,N_466);
xnor U612 (N_612,N_432,In_1178);
xnor U613 (N_613,N_141,In_233);
nand U614 (N_614,In_297,N_209);
nand U615 (N_615,In_177,In_5);
and U616 (N_616,N_199,N_485);
and U617 (N_617,In_1491,In_700);
or U618 (N_618,N_441,In_805);
nor U619 (N_619,In_1245,N_490);
xor U620 (N_620,N_437,In_387);
or U621 (N_621,In_1401,In_664);
or U622 (N_622,In_197,N_363);
xnor U623 (N_623,In_432,N_453);
nand U624 (N_624,N_325,In_969);
nand U625 (N_625,N_381,In_1087);
and U626 (N_626,In_1281,N_205);
and U627 (N_627,In_696,In_1227);
xor U628 (N_628,N_420,N_338);
nand U629 (N_629,N_28,N_473);
xnor U630 (N_630,N_452,In_70);
or U631 (N_631,In_1420,N_480);
or U632 (N_632,In_1162,N_397);
or U633 (N_633,In_28,In_521);
or U634 (N_634,N_298,N_274);
nand U635 (N_635,In_560,In_93);
or U636 (N_636,In_1287,In_163);
nand U637 (N_637,In_20,N_96);
or U638 (N_638,In_1247,N_255);
xor U639 (N_639,In_189,N_21);
xnor U640 (N_640,N_188,N_112);
nor U641 (N_641,In_614,In_453);
xor U642 (N_642,In_1463,In_1329);
or U643 (N_643,In_1149,N_366);
xor U644 (N_644,In_1299,In_64);
and U645 (N_645,In_384,N_1);
xor U646 (N_646,In_541,In_1172);
or U647 (N_647,N_69,In_823);
nand U648 (N_648,In_47,In_567);
or U649 (N_649,In_1246,In_409);
or U650 (N_650,In_518,In_1272);
xnor U651 (N_651,In_1415,In_551);
or U652 (N_652,N_440,N_311);
and U653 (N_653,In_1156,In_1073);
xor U654 (N_654,In_746,N_217);
nor U655 (N_655,In_1150,In_129);
and U656 (N_656,N_385,N_341);
xor U657 (N_657,In_720,In_760);
xnor U658 (N_658,In_1315,In_1207);
nand U659 (N_659,N_126,In_809);
nand U660 (N_660,In_970,In_281);
or U661 (N_661,In_1164,N_376);
or U662 (N_662,N_162,In_68);
and U663 (N_663,N_304,In_1046);
and U664 (N_664,In_212,N_486);
or U665 (N_665,In_657,N_287);
nor U666 (N_666,N_293,In_771);
and U667 (N_667,In_1217,N_326);
or U668 (N_668,In_316,N_353);
and U669 (N_669,N_251,In_1022);
xnor U670 (N_670,In_328,In_600);
xor U671 (N_671,In_294,In_956);
and U672 (N_672,In_581,N_369);
xor U673 (N_673,In_366,In_1059);
nor U674 (N_674,In_390,In_215);
or U675 (N_675,In_788,N_422);
nand U676 (N_676,In_565,N_318);
or U677 (N_677,N_433,N_200);
xnor U678 (N_678,N_125,N_301);
and U679 (N_679,In_278,N_395);
nand U680 (N_680,N_204,In_200);
nand U681 (N_681,N_61,In_882);
or U682 (N_682,N_121,In_464);
and U683 (N_683,N_53,N_360);
and U684 (N_684,In_140,In_773);
and U685 (N_685,In_1361,In_1146);
nor U686 (N_686,N_470,N_354);
xor U687 (N_687,N_436,In_1473);
or U688 (N_688,In_336,N_228);
xnor U689 (N_689,In_493,In_703);
xor U690 (N_690,In_223,In_1062);
and U691 (N_691,N_107,N_150);
nand U692 (N_692,In_500,In_1480);
xnor U693 (N_693,N_282,In_513);
nand U694 (N_694,N_498,In_549);
and U695 (N_695,N_297,N_269);
and U696 (N_696,In_1036,In_86);
nor U697 (N_697,In_512,N_462);
xnor U698 (N_698,In_400,N_59);
and U699 (N_699,N_423,In_162);
or U700 (N_700,In_690,In_455);
xor U701 (N_701,In_667,N_140);
nand U702 (N_702,N_488,In_214);
nor U703 (N_703,In_208,In_11);
or U704 (N_704,N_352,N_182);
nor U705 (N_705,In_408,In_1430);
xor U706 (N_706,In_1049,In_779);
nand U707 (N_707,In_1384,In_311);
xnor U708 (N_708,In_348,In_314);
or U709 (N_709,N_284,N_468);
or U710 (N_710,N_339,In_826);
and U711 (N_711,N_421,N_404);
and U712 (N_712,In_727,In_1307);
xor U713 (N_713,In_1129,N_50);
or U714 (N_714,In_266,In_1373);
nand U715 (N_715,In_1197,In_334);
xor U716 (N_716,In_81,N_403);
or U717 (N_717,In_1320,In_670);
nand U718 (N_718,N_427,N_317);
nand U719 (N_719,N_179,In_695);
xnor U720 (N_720,N_168,N_321);
and U721 (N_721,In_489,In_1065);
xor U722 (N_722,In_126,In_479);
xnor U723 (N_723,In_154,In_308);
and U724 (N_724,N_442,In_883);
or U725 (N_725,In_1364,In_1319);
and U726 (N_726,In_615,N_243);
xor U727 (N_727,N_384,In_654);
nand U728 (N_728,In_1132,In_986);
or U729 (N_729,In_407,N_216);
and U730 (N_730,In_1259,N_105);
nor U731 (N_731,In_274,In_863);
and U732 (N_732,In_843,In_755);
nand U733 (N_733,In_552,In_960);
or U734 (N_734,N_383,N_372);
nor U735 (N_735,In_1223,N_264);
nor U736 (N_736,In_1451,In_584);
xor U737 (N_737,In_1008,In_72);
and U738 (N_738,In_7,N_290);
nor U739 (N_739,N_180,In_585);
xnor U740 (N_740,N_409,In_1063);
and U741 (N_741,In_321,In_958);
nor U742 (N_742,In_675,In_335);
nor U743 (N_743,N_18,In_344);
nor U744 (N_744,N_355,In_470);
nor U745 (N_745,In_704,N_44);
and U746 (N_746,N_309,In_1347);
or U747 (N_747,N_241,In_816);
and U748 (N_748,N_279,N_359);
and U749 (N_749,N_258,N_41);
and U750 (N_750,In_1128,N_32);
nand U751 (N_751,N_300,N_110);
or U752 (N_752,In_1381,N_565);
xnor U753 (N_753,N_537,In_687);
xor U754 (N_754,N_697,N_495);
and U755 (N_755,In_759,N_266);
or U756 (N_756,N_624,In_357);
nor U757 (N_757,In_1033,N_654);
nand U758 (N_758,N_222,N_502);
xor U759 (N_759,In_1117,In_1070);
and U760 (N_760,In_708,In_1486);
nor U761 (N_761,N_231,In_412);
nand U762 (N_762,N_491,N_723);
nand U763 (N_763,N_681,In_420);
nand U764 (N_764,In_196,N_690);
xor U765 (N_765,In_898,N_398);
xor U766 (N_766,In_1102,In_119);
or U767 (N_767,N_554,N_223);
nor U768 (N_768,N_597,In_800);
xnor U769 (N_769,In_1403,N_203);
nand U770 (N_770,N_744,N_48);
and U771 (N_771,N_424,N_523);
xor U772 (N_772,N_276,N_261);
nor U773 (N_773,N_345,In_769);
and U774 (N_774,N_530,N_645);
xor U775 (N_775,N_655,In_957);
or U776 (N_776,N_493,N_598);
nand U777 (N_777,N_605,In_304);
or U778 (N_778,N_101,N_642);
xor U779 (N_779,N_603,In_972);
and U780 (N_780,N_459,N_418);
nor U781 (N_781,N_406,N_25);
and U782 (N_782,In_932,N_631);
xnor U783 (N_783,N_647,In_1079);
nor U784 (N_784,N_575,In_1119);
and U785 (N_785,N_2,N_508);
nor U786 (N_786,N_563,In_137);
xor U787 (N_787,In_42,In_13);
xnor U788 (N_788,N_472,In_1147);
nand U789 (N_789,In_607,N_630);
xor U790 (N_790,N_577,N_742);
or U791 (N_791,In_323,N_271);
xnor U792 (N_792,In_1168,In_765);
nand U793 (N_793,N_399,N_632);
xor U794 (N_794,In_1326,In_694);
and U795 (N_795,In_840,In_1324);
xor U796 (N_796,N_549,In_1213);
or U797 (N_797,In_922,In_592);
nor U798 (N_798,In_909,In_1289);
and U799 (N_799,In_1306,N_536);
nor U800 (N_800,In_39,In_980);
xor U801 (N_801,N_617,N_581);
and U802 (N_802,In_1179,N_334);
nor U803 (N_803,N_633,N_522);
and U804 (N_804,N_567,N_746);
nor U805 (N_805,In_624,N_307);
xnor U806 (N_806,N_476,N_734);
xor U807 (N_807,In_920,In_942);
and U808 (N_808,In_1359,N_611);
xnor U809 (N_809,N_22,N_573);
nor U810 (N_810,N_670,N_444);
or U811 (N_811,N_733,N_570);
or U812 (N_812,N_535,In_1424);
xnor U813 (N_813,In_527,N_149);
or U814 (N_814,N_583,N_532);
or U815 (N_815,N_717,N_588);
nand U816 (N_816,In_1342,In_285);
nor U817 (N_817,In_1111,N_740);
and U818 (N_818,N_402,N_337);
and U819 (N_819,N_728,In_329);
nand U820 (N_820,In_1121,In_1035);
nor U821 (N_821,N_607,N_692);
and U822 (N_822,In_949,N_273);
and U823 (N_823,N_629,In_1322);
or U824 (N_824,In_822,In_1136);
nand U825 (N_825,In_889,N_396);
nand U826 (N_826,In_743,In_395);
or U827 (N_827,N_672,N_405);
xnor U828 (N_828,N_571,N_561);
and U829 (N_829,In_1071,In_1175);
and U830 (N_830,In_100,In_1110);
nand U831 (N_831,In_1365,N_600);
nor U832 (N_832,In_851,In_182);
and U833 (N_833,N_709,N_574);
or U834 (N_834,In_1464,N_215);
nand U835 (N_835,N_564,N_729);
or U836 (N_836,In_91,In_340);
xnor U837 (N_837,N_568,N_429);
xor U838 (N_838,In_1194,N_79);
xnor U839 (N_839,N_164,In_709);
nor U840 (N_840,In_872,N_267);
or U841 (N_841,N_529,N_292);
xor U842 (N_842,In_23,In_663);
nand U843 (N_843,N_413,N_628);
or U844 (N_844,N_349,N_719);
xnor U845 (N_845,In_430,In_363);
xor U846 (N_846,In_1210,N_389);
and U847 (N_847,In_930,In_1437);
and U848 (N_848,N_516,N_665);
and U849 (N_849,In_739,In_290);
or U850 (N_850,N_722,N_721);
nor U851 (N_851,In_218,N_591);
or U852 (N_852,N_26,N_707);
nor U853 (N_853,N_394,N_428);
or U854 (N_854,In_642,N_477);
and U855 (N_855,N_745,In_899);
xor U856 (N_856,N_612,In_1183);
xor U857 (N_857,In_1253,N_622);
and U858 (N_858,In_858,In_1124);
nand U859 (N_859,N_286,N_636);
or U860 (N_860,N_289,N_252);
nor U861 (N_861,N_596,In_1406);
xnor U862 (N_862,In_554,N_712);
or U863 (N_863,In_1476,N_291);
and U864 (N_864,In_927,N_414);
and U865 (N_865,N_478,N_380);
and U866 (N_866,N_684,N_711);
and U867 (N_867,N_592,In_1445);
xor U868 (N_868,N_320,In_650);
xor U869 (N_869,N_461,N_517);
nor U870 (N_870,In_1371,In_796);
nand U871 (N_871,N_19,N_275);
or U872 (N_872,In_950,N_616);
xor U873 (N_873,In_1344,In_1302);
nor U874 (N_874,N_635,In_649);
xnor U875 (N_875,N_356,N_118);
and U876 (N_876,In_1139,N_327);
and U877 (N_877,N_332,N_294);
or U878 (N_878,N_312,N_699);
nand U879 (N_879,In_1190,N_313);
nor U880 (N_880,N_582,In_1434);
nand U881 (N_881,N_346,In_961);
xor U882 (N_882,In_1140,N_358);
nand U883 (N_883,In_810,N_98);
or U884 (N_884,In_877,N_627);
xor U885 (N_885,N_716,N_416);
nor U886 (N_886,N_547,N_504);
and U887 (N_887,N_374,N_747);
nand U888 (N_888,N_653,N_743);
xnor U889 (N_889,N_663,In_1395);
or U890 (N_890,N_718,N_708);
or U891 (N_891,N_685,N_83);
nor U892 (N_892,N_242,N_545);
and U893 (N_893,N_316,In_616);
and U894 (N_894,In_1335,N_578);
and U895 (N_895,In_1334,In_49);
nor U896 (N_896,N_551,In_101);
and U897 (N_897,N_542,In_630);
nand U898 (N_898,N_435,In_265);
xor U899 (N_899,N_524,N_675);
or U900 (N_900,N_621,In_1153);
and U901 (N_901,N_691,In_403);
xnor U902 (N_902,N_695,N_471);
nor U903 (N_903,N_661,In_628);
xor U904 (N_904,In_548,N_644);
xnor U905 (N_905,N_390,In_767);
xnor U906 (N_906,In_368,N_687);
and U907 (N_907,N_5,N_93);
nor U908 (N_908,In_264,N_594);
or U909 (N_909,N_272,N_483);
xor U910 (N_910,N_724,N_445);
nand U911 (N_911,N_335,N_500);
or U912 (N_912,In_1279,N_408);
xnor U913 (N_913,N_283,N_680);
xnor U914 (N_914,In_418,In_226);
or U915 (N_915,In_1456,N_494);
xnor U916 (N_916,N_748,In_31);
nand U917 (N_917,In_1492,In_914);
nor U918 (N_918,N_136,In_183);
nand U919 (N_919,N_501,In_1413);
and U920 (N_920,N_438,N_323);
nand U921 (N_921,In_442,N_132);
nand U922 (N_922,N_288,N_520);
nor U923 (N_923,In_871,N_727);
or U924 (N_924,In_1231,In_1286);
xnor U925 (N_925,N_375,N_348);
or U926 (N_926,N_589,N_693);
xnor U927 (N_927,N_87,In_382);
xnor U928 (N_928,N_557,N_638);
or U929 (N_929,N_513,In_954);
xor U930 (N_930,N_666,In_1042);
nor U931 (N_931,In_1277,In_1216);
nor U932 (N_932,In_277,N_4);
nor U933 (N_933,N_558,N_648);
xor U934 (N_934,In_372,N_656);
or U935 (N_935,In_959,In_252);
and U936 (N_936,N_556,N_572);
xor U937 (N_937,In_641,N_245);
nor U938 (N_938,N_365,N_510);
xor U939 (N_939,N_378,In_1312);
nor U940 (N_940,N_254,N_602);
nand U941 (N_941,N_609,N_730);
xor U942 (N_942,N_683,N_562);
xnor U943 (N_943,In_1353,N_623);
nor U944 (N_944,N_541,In_707);
nor U945 (N_945,In_1447,In_993);
and U946 (N_946,N_625,N_527);
and U947 (N_947,In_588,N_80);
and U948 (N_948,In_1323,N_299);
and U949 (N_949,N_14,N_660);
and U950 (N_950,N_82,N_555);
nand U951 (N_951,In_1363,N_379);
nor U952 (N_952,N_34,N_585);
and U953 (N_953,N_546,N_333);
and U954 (N_954,N_586,In_450);
and U955 (N_955,N_382,In_38);
or U956 (N_956,N_328,N_52);
nand U957 (N_957,N_507,N_550);
nor U958 (N_958,N_682,In_1311);
nand U959 (N_959,N_233,N_457);
xor U960 (N_960,In_178,In_159);
xor U961 (N_961,N_412,N_662);
nand U962 (N_962,N_698,N_340);
nor U963 (N_963,N_119,N_726);
nand U964 (N_964,In_250,In_193);
and U965 (N_965,In_322,In_4);
or U966 (N_966,In_431,N_651);
nor U967 (N_967,In_566,N_62);
and U968 (N_968,In_702,N_512);
or U969 (N_969,N_579,N_511);
or U970 (N_970,In_222,In_253);
nand U971 (N_971,In_1104,N_449);
nor U972 (N_972,In_648,N_330);
and U973 (N_973,In_503,N_701);
nor U974 (N_974,In_84,In_1076);
nand U975 (N_975,In_854,N_235);
or U976 (N_976,In_224,N_109);
nor U977 (N_977,N_531,In_1037);
or U978 (N_978,N_230,In_1443);
nor U979 (N_979,In_273,In_604);
xor U980 (N_980,In_1414,In_976);
xor U981 (N_981,N_464,N_643);
nand U982 (N_982,N_533,N_626);
xnor U983 (N_983,In_1180,In_1107);
or U984 (N_984,N_580,N_166);
nor U985 (N_985,N_618,In_295);
and U986 (N_986,N_236,N_319);
or U987 (N_987,In_724,N_599);
xnor U988 (N_988,In_692,In_27);
and U989 (N_989,N_668,In_754);
xnor U990 (N_990,In_1394,In_1372);
and U991 (N_991,N_497,N_148);
and U992 (N_992,N_329,N_539);
nand U993 (N_993,N_637,In_434);
or U994 (N_994,N_639,In_1343);
nand U995 (N_995,In_203,N_528);
or U996 (N_996,In_417,N_518);
nand U997 (N_997,In_331,In_139);
xor U998 (N_998,N_391,In_244);
nor U999 (N_999,N_165,In_1489);
nand U1000 (N_1000,N_544,N_469);
nor U1001 (N_1001,N_975,N_154);
or U1002 (N_1002,N_905,N_357);
or U1003 (N_1003,In_572,N_895);
or U1004 (N_1004,In_992,N_849);
or U1005 (N_1005,N_590,N_634);
and U1006 (N_1006,N_935,N_559);
nand U1007 (N_1007,N_509,N_976);
and U1008 (N_1008,N_206,N_649);
xor U1009 (N_1009,N_678,N_751);
nor U1010 (N_1010,N_641,N_833);
or U1011 (N_1011,N_425,N_946);
and U1012 (N_1012,In_1237,N_981);
nand U1013 (N_1013,N_198,In_478);
nand U1014 (N_1014,N_970,N_783);
or U1015 (N_1015,In_508,N_871);
and U1016 (N_1016,In_310,N_732);
and U1017 (N_1017,N_851,N_484);
and U1018 (N_1018,N_939,N_63);
xnor U1019 (N_1019,In_1278,N_42);
xnor U1020 (N_1020,In_127,N_818);
or U1021 (N_1021,N_36,N_812);
and U1022 (N_1022,N_773,N_386);
xnor U1023 (N_1023,N_657,N_29);
nand U1024 (N_1024,N_947,N_963);
xnor U1025 (N_1025,In_230,In_98);
and U1026 (N_1026,N_926,N_911);
or U1027 (N_1027,In_498,N_113);
xnor U1028 (N_1028,N_752,N_828);
nor U1029 (N_1029,N_615,N_587);
and U1030 (N_1030,N_704,N_936);
nand U1031 (N_1031,N_614,N_854);
xor U1032 (N_1032,N_919,N_538);
nor U1033 (N_1033,N_897,In_842);
nor U1034 (N_1034,In_1260,N_785);
nand U1035 (N_1035,N_367,In_332);
xor U1036 (N_1036,N_246,N_861);
or U1037 (N_1037,N_769,N_943);
or U1038 (N_1038,N_852,In_1006);
xnor U1039 (N_1039,N_706,N_601);
and U1040 (N_1040,N_806,N_922);
and U1041 (N_1041,N_902,In_451);
xor U1042 (N_1042,N_184,N_765);
nand U1043 (N_1043,N_505,N_908);
or U1044 (N_1044,In_361,N_696);
and U1045 (N_1045,N_874,N_817);
nor U1046 (N_1046,N_351,In_744);
nand U1047 (N_1047,N_990,N_856);
and U1048 (N_1048,N_810,N_31);
and U1049 (N_1049,N_454,N_841);
and U1050 (N_1050,In_814,N_713);
xor U1051 (N_1051,In_388,N_980);
and U1052 (N_1052,N_993,N_791);
and U1053 (N_1053,In_1450,N_260);
xor U1054 (N_1054,N_888,N_868);
nor U1055 (N_1055,N_771,N_77);
xnor U1056 (N_1056,N_967,N_604);
or U1057 (N_1057,In_444,N_362);
nor U1058 (N_1058,N_987,N_296);
xor U1059 (N_1059,In_1224,N_881);
or U1060 (N_1060,In_1317,N_929);
nor U1061 (N_1061,N_945,In_808);
nand U1062 (N_1062,N_829,N_764);
or U1063 (N_1063,N_839,N_850);
xnor U1064 (N_1064,N_128,N_974);
xnor U1065 (N_1065,N_676,N_277);
xnor U1066 (N_1066,In_51,N_97);
nor U1067 (N_1067,N_918,N_754);
and U1068 (N_1068,N_239,N_688);
nor U1069 (N_1069,N_741,N_997);
or U1070 (N_1070,In_1404,N_731);
xnor U1071 (N_1071,In_894,N_801);
xnor U1072 (N_1072,N_766,N_928);
and U1073 (N_1073,N_342,N_965);
xnor U1074 (N_1074,N_650,In_364);
and U1075 (N_1075,N_224,N_789);
nor U1076 (N_1076,N_816,N_857);
or U1077 (N_1077,In_124,N_308);
or U1078 (N_1078,N_912,N_797);
xor U1079 (N_1079,N_755,N_659);
nor U1080 (N_1080,In_726,N_904);
nor U1081 (N_1081,N_879,N_843);
nand U1082 (N_1082,N_664,N_799);
and U1083 (N_1083,N_959,N_956);
or U1084 (N_1084,N_576,N_827);
and U1085 (N_1085,N_925,N_860);
nand U1086 (N_1086,N_896,In_966);
nand U1087 (N_1087,In_1166,N_914);
or U1088 (N_1088,N_844,N_950);
nor U1089 (N_1089,N_923,N_821);
xor U1090 (N_1090,In_369,N_620);
xnor U1091 (N_1091,In_1232,N_772);
nor U1092 (N_1092,N_410,N_377);
nand U1093 (N_1093,In_748,N_986);
xnor U1094 (N_1094,N_322,N_813);
xnor U1095 (N_1095,N_364,N_870);
nand U1096 (N_1096,N_762,N_738);
and U1097 (N_1097,N_606,In_1200);
or U1098 (N_1098,In_83,In_963);
or U1099 (N_1099,N_953,N_758);
or U1100 (N_1100,N_873,N_983);
or U1101 (N_1101,N_800,N_777);
xor U1102 (N_1102,In_118,N_503);
nor U1103 (N_1103,N_703,In_1416);
xor U1104 (N_1104,N_526,N_855);
nand U1105 (N_1105,N_331,N_811);
nor U1106 (N_1106,N_915,N_646);
xnor U1107 (N_1107,N_753,N_802);
or U1108 (N_1108,N_776,In_1089);
or U1109 (N_1109,N_265,N_969);
or U1110 (N_1110,N_891,N_566);
and U1111 (N_1111,N_548,N_191);
nor U1112 (N_1112,In_374,N_679);
or U1113 (N_1113,N_866,In_1251);
nand U1114 (N_1114,In_897,N_819);
xnor U1115 (N_1115,N_894,N_836);
nor U1116 (N_1116,In_423,N_991);
nand U1117 (N_1117,N_885,In_1467);
nor U1118 (N_1118,In_1282,In_1229);
or U1119 (N_1119,N_814,N_996);
xnor U1120 (N_1120,In_1023,N_864);
or U1121 (N_1121,In_758,N_877);
nand U1122 (N_1122,N_948,N_790);
nor U1123 (N_1123,In_783,N_705);
nand U1124 (N_1124,N_979,N_940);
nand U1125 (N_1125,N_780,N_552);
nand U1126 (N_1126,N_985,N_784);
nor U1127 (N_1127,N_998,N_736);
nor U1128 (N_1128,In_50,In_979);
xnor U1129 (N_1129,N_957,N_977);
or U1130 (N_1130,N_834,N_853);
or U1131 (N_1131,In_41,N_781);
and U1132 (N_1132,N_70,In_609);
nand U1133 (N_1133,N_796,N_982);
and U1134 (N_1134,N_971,N_737);
nand U1135 (N_1135,N_906,N_194);
nand U1136 (N_1136,N_815,N_702);
nor U1137 (N_1137,N_250,N_933);
and U1138 (N_1138,N_921,N_984);
nor U1139 (N_1139,N_506,N_989);
nand U1140 (N_1140,N_305,N_139);
xor U1141 (N_1141,N_824,N_934);
or U1142 (N_1142,N_898,N_955);
and U1143 (N_1143,N_610,N_994);
and U1144 (N_1144,In_679,N_710);
or U1145 (N_1145,N_838,N_122);
or U1146 (N_1146,In_235,N_809);
nand U1147 (N_1147,N_768,N_295);
nor U1148 (N_1148,N_907,In_419);
nand U1149 (N_1149,In_520,N_962);
or U1150 (N_1150,N_960,N_593);
nor U1151 (N_1151,N_689,N_525);
xnor U1152 (N_1152,N_931,N_954);
and U1153 (N_1153,In_1155,In_187);
nor U1154 (N_1154,N_514,N_978);
or U1155 (N_1155,N_792,N_835);
xnor U1156 (N_1156,N_880,N_913);
xor U1157 (N_1157,N_826,N_336);
and U1158 (N_1158,N_820,N_951);
nor U1159 (N_1159,N_900,N_927);
and U1160 (N_1160,N_519,N_756);
or U1161 (N_1161,In_1325,In_441);
and U1162 (N_1162,N_787,In_474);
nor U1163 (N_1163,N_878,N_218);
nand U1164 (N_1164,N_456,N_393);
xor U1165 (N_1165,N_640,N_392);
and U1166 (N_1166,N_916,N_673);
nand U1167 (N_1167,N_257,N_757);
xnor U1168 (N_1168,N_760,N_608);
nand U1169 (N_1169,N_788,N_886);
xor U1170 (N_1170,In_55,N_268);
or U1171 (N_1171,In_380,N_863);
nor U1172 (N_1172,N_859,N_862);
or U1173 (N_1173,N_830,N_941);
or U1174 (N_1174,N_763,N_669);
nand U1175 (N_1175,In_377,N_823);
nor U1176 (N_1176,N_804,N_899);
nand U1177 (N_1177,N_770,N_793);
or U1178 (N_1178,N_942,In_617);
nand U1179 (N_1179,N_371,In_689);
nor U1180 (N_1180,N_761,In_1337);
xor U1181 (N_1181,In_1460,N_840);
xnor U1182 (N_1182,N_890,In_721);
or U1183 (N_1183,N_917,N_778);
and U1184 (N_1184,N_924,N_324);
xnor U1185 (N_1185,In_785,N_938);
nand U1186 (N_1186,N_903,N_920);
or U1187 (N_1187,N_694,N_499);
xnor U1188 (N_1188,N_443,N_973);
nor U1189 (N_1189,N_759,N_652);
or U1190 (N_1190,N_116,N_782);
xnor U1191 (N_1191,In_1195,N_775);
nor U1192 (N_1192,N_677,N_803);
xor U1193 (N_1193,N_725,N_798);
nor U1194 (N_1194,N_540,In_875);
or U1195 (N_1195,In_393,N_786);
xor U1196 (N_1196,In_935,N_584);
nor U1197 (N_1197,N_992,N_858);
nor U1198 (N_1198,In_1457,N_560);
xor U1199 (N_1199,N_845,N_961);
nor U1200 (N_1200,In_925,In_1105);
nor U1201 (N_1201,N_750,In_747);
xor U1202 (N_1202,N_865,N_361);
nand U1203 (N_1203,N_807,N_883);
or U1204 (N_1204,In_1082,N_876);
and U1205 (N_1205,N_930,N_869);
nor U1206 (N_1206,In_460,N_831);
or U1207 (N_1207,N_521,N_968);
or U1208 (N_1208,N_884,In_1097);
nand U1209 (N_1209,N_779,In_262);
nand U1210 (N_1210,N_739,N_972);
nor U1211 (N_1211,In_1127,N_872);
nand U1212 (N_1212,In_1369,In_1475);
or U1213 (N_1213,N_749,N_910);
and U1214 (N_1214,N_837,N_256);
nand U1215 (N_1215,N_999,N_553);
nor U1216 (N_1216,N_882,N_932);
nor U1217 (N_1217,N_686,N_715);
nand U1218 (N_1218,N_613,N_487);
nor U1219 (N_1219,N_619,N_892);
nand U1220 (N_1220,N_595,N_767);
nor U1221 (N_1221,N_889,In_404);
or U1222 (N_1222,N_808,In_1411);
xnor U1223 (N_1223,N_995,N_958);
and U1224 (N_1224,N_966,N_515);
and U1225 (N_1225,In_1308,N_720);
and U1226 (N_1226,N_774,N_822);
xnor U1227 (N_1227,N_944,N_667);
nand U1228 (N_1228,N_543,N_658);
and U1229 (N_1229,N_671,N_847);
and U1230 (N_1230,N_909,N_846);
and U1231 (N_1231,N_458,N_388);
nand U1232 (N_1232,N_496,N_937);
nand U1233 (N_1233,In_1496,N_805);
nor U1234 (N_1234,N_848,N_211);
xor U1235 (N_1235,N_735,In_1495);
xnor U1236 (N_1236,In_1108,N_344);
and U1237 (N_1237,N_794,In_693);
or U1238 (N_1238,N_893,N_949);
nor U1239 (N_1239,N_825,N_964);
and U1240 (N_1240,N_534,N_795);
nor U1241 (N_1241,N_988,N_867);
or U1242 (N_1242,N_315,N_302);
or U1243 (N_1243,N_842,N_714);
nor U1244 (N_1244,N_875,N_439);
or U1245 (N_1245,N_901,N_569);
nor U1246 (N_1246,N_887,In_436);
nand U1247 (N_1247,N_674,N_952);
nand U1248 (N_1248,N_832,In_1109);
and U1249 (N_1249,N_448,N_700);
nor U1250 (N_1250,N_1063,N_1231);
nand U1251 (N_1251,N_1094,N_1237);
nor U1252 (N_1252,N_1124,N_1229);
and U1253 (N_1253,N_1088,N_1238);
nand U1254 (N_1254,N_1188,N_1008);
nand U1255 (N_1255,N_1058,N_1097);
or U1256 (N_1256,N_1148,N_1033);
or U1257 (N_1257,N_1143,N_1043);
nand U1258 (N_1258,N_1120,N_1089);
or U1259 (N_1259,N_1056,N_1163);
and U1260 (N_1260,N_1187,N_1005);
or U1261 (N_1261,N_1227,N_1152);
nor U1262 (N_1262,N_1192,N_1181);
nand U1263 (N_1263,N_1007,N_1159);
or U1264 (N_1264,N_1109,N_1233);
and U1265 (N_1265,N_1145,N_1015);
nor U1266 (N_1266,N_1217,N_1203);
xor U1267 (N_1267,N_1074,N_1240);
nor U1268 (N_1268,N_1023,N_1161);
and U1269 (N_1269,N_1000,N_1084);
and U1270 (N_1270,N_1006,N_1234);
nand U1271 (N_1271,N_1073,N_1025);
and U1272 (N_1272,N_1051,N_1222);
nand U1273 (N_1273,N_1052,N_1134);
nand U1274 (N_1274,N_1127,N_1042);
nor U1275 (N_1275,N_1218,N_1106);
or U1276 (N_1276,N_1072,N_1001);
nand U1277 (N_1277,N_1016,N_1102);
xnor U1278 (N_1278,N_1012,N_1021);
and U1279 (N_1279,N_1093,N_1128);
nor U1280 (N_1280,N_1223,N_1244);
and U1281 (N_1281,N_1071,N_1209);
nand U1282 (N_1282,N_1154,N_1009);
and U1283 (N_1283,N_1100,N_1091);
and U1284 (N_1284,N_1156,N_1049);
nor U1285 (N_1285,N_1060,N_1064);
and U1286 (N_1286,N_1096,N_1018);
nand U1287 (N_1287,N_1135,N_1151);
xnor U1288 (N_1288,N_1214,N_1020);
xnor U1289 (N_1289,N_1057,N_1220);
nor U1290 (N_1290,N_1228,N_1131);
nand U1291 (N_1291,N_1062,N_1150);
xnor U1292 (N_1292,N_1067,N_1139);
xor U1293 (N_1293,N_1078,N_1160);
or U1294 (N_1294,N_1115,N_1235);
nand U1295 (N_1295,N_1004,N_1123);
nand U1296 (N_1296,N_1061,N_1153);
xnor U1297 (N_1297,N_1162,N_1213);
xor U1298 (N_1298,N_1095,N_1101);
nor U1299 (N_1299,N_1149,N_1204);
and U1300 (N_1300,N_1076,N_1069);
xor U1301 (N_1301,N_1122,N_1036);
and U1302 (N_1302,N_1142,N_1247);
nor U1303 (N_1303,N_1175,N_1011);
xnor U1304 (N_1304,N_1208,N_1199);
nand U1305 (N_1305,N_1184,N_1226);
nand U1306 (N_1306,N_1243,N_1099);
nor U1307 (N_1307,N_1138,N_1136);
or U1308 (N_1308,N_1083,N_1144);
nor U1309 (N_1309,N_1080,N_1191);
or U1310 (N_1310,N_1180,N_1044);
or U1311 (N_1311,N_1040,N_1190);
or U1312 (N_1312,N_1249,N_1157);
or U1313 (N_1313,N_1114,N_1194);
or U1314 (N_1314,N_1225,N_1130);
or U1315 (N_1315,N_1118,N_1119);
nand U1316 (N_1316,N_1116,N_1206);
and U1317 (N_1317,N_1068,N_1079);
nand U1318 (N_1318,N_1167,N_1183);
or U1319 (N_1319,N_1082,N_1010);
nor U1320 (N_1320,N_1087,N_1186);
nand U1321 (N_1321,N_1105,N_1028);
nand U1322 (N_1322,N_1041,N_1179);
or U1323 (N_1323,N_1147,N_1117);
nor U1324 (N_1324,N_1155,N_1216);
and U1325 (N_1325,N_1129,N_1248);
nand U1326 (N_1326,N_1221,N_1030);
and U1327 (N_1327,N_1031,N_1230);
nand U1328 (N_1328,N_1113,N_1107);
and U1329 (N_1329,N_1165,N_1133);
or U1330 (N_1330,N_1164,N_1121);
xnor U1331 (N_1331,N_1171,N_1224);
xnor U1332 (N_1332,N_1108,N_1207);
and U1333 (N_1333,N_1137,N_1195);
xor U1334 (N_1334,N_1053,N_1200);
or U1335 (N_1335,N_1189,N_1193);
nand U1336 (N_1336,N_1059,N_1172);
or U1337 (N_1337,N_1054,N_1174);
nand U1338 (N_1338,N_1092,N_1066);
xor U1339 (N_1339,N_1019,N_1046);
nand U1340 (N_1340,N_1081,N_1048);
or U1341 (N_1341,N_1196,N_1166);
xor U1342 (N_1342,N_1236,N_1038);
or U1343 (N_1343,N_1034,N_1246);
nand U1344 (N_1344,N_1176,N_1065);
or U1345 (N_1345,N_1178,N_1245);
xnor U1346 (N_1346,N_1242,N_1141);
xnor U1347 (N_1347,N_1098,N_1132);
xor U1348 (N_1348,N_1212,N_1050);
and U1349 (N_1349,N_1182,N_1070);
and U1350 (N_1350,N_1197,N_1103);
or U1351 (N_1351,N_1013,N_1185);
nand U1352 (N_1352,N_1241,N_1027);
xor U1353 (N_1353,N_1075,N_1039);
xnor U1354 (N_1354,N_1173,N_1239);
or U1355 (N_1355,N_1022,N_1125);
or U1356 (N_1356,N_1002,N_1205);
nor U1357 (N_1357,N_1110,N_1085);
or U1358 (N_1358,N_1170,N_1090);
nor U1359 (N_1359,N_1024,N_1045);
nor U1360 (N_1360,N_1232,N_1037);
or U1361 (N_1361,N_1032,N_1219);
or U1362 (N_1362,N_1126,N_1112);
nand U1363 (N_1363,N_1169,N_1146);
and U1364 (N_1364,N_1003,N_1198);
nor U1365 (N_1365,N_1026,N_1168);
nand U1366 (N_1366,N_1077,N_1014);
and U1367 (N_1367,N_1140,N_1211);
and U1368 (N_1368,N_1104,N_1210);
nand U1369 (N_1369,N_1035,N_1086);
or U1370 (N_1370,N_1017,N_1158);
nand U1371 (N_1371,N_1202,N_1201);
or U1372 (N_1372,N_1029,N_1111);
nor U1373 (N_1373,N_1215,N_1047);
nor U1374 (N_1374,N_1177,N_1055);
and U1375 (N_1375,N_1225,N_1010);
or U1376 (N_1376,N_1197,N_1117);
xor U1377 (N_1377,N_1242,N_1024);
nor U1378 (N_1378,N_1101,N_1075);
xor U1379 (N_1379,N_1161,N_1050);
nor U1380 (N_1380,N_1172,N_1198);
nand U1381 (N_1381,N_1022,N_1240);
nor U1382 (N_1382,N_1065,N_1164);
nand U1383 (N_1383,N_1142,N_1168);
nor U1384 (N_1384,N_1157,N_1145);
or U1385 (N_1385,N_1065,N_1017);
and U1386 (N_1386,N_1053,N_1172);
nand U1387 (N_1387,N_1093,N_1039);
or U1388 (N_1388,N_1208,N_1206);
or U1389 (N_1389,N_1248,N_1083);
and U1390 (N_1390,N_1135,N_1011);
nand U1391 (N_1391,N_1190,N_1149);
and U1392 (N_1392,N_1229,N_1100);
or U1393 (N_1393,N_1190,N_1095);
nor U1394 (N_1394,N_1036,N_1229);
or U1395 (N_1395,N_1091,N_1185);
nor U1396 (N_1396,N_1114,N_1035);
nand U1397 (N_1397,N_1163,N_1192);
and U1398 (N_1398,N_1071,N_1216);
nor U1399 (N_1399,N_1035,N_1196);
nand U1400 (N_1400,N_1162,N_1225);
and U1401 (N_1401,N_1025,N_1213);
xnor U1402 (N_1402,N_1179,N_1135);
nand U1403 (N_1403,N_1153,N_1103);
nor U1404 (N_1404,N_1024,N_1176);
nand U1405 (N_1405,N_1178,N_1099);
or U1406 (N_1406,N_1098,N_1033);
or U1407 (N_1407,N_1046,N_1009);
or U1408 (N_1408,N_1206,N_1218);
nor U1409 (N_1409,N_1074,N_1021);
xnor U1410 (N_1410,N_1142,N_1054);
or U1411 (N_1411,N_1197,N_1045);
and U1412 (N_1412,N_1153,N_1191);
nand U1413 (N_1413,N_1114,N_1019);
xor U1414 (N_1414,N_1073,N_1229);
or U1415 (N_1415,N_1089,N_1075);
nor U1416 (N_1416,N_1050,N_1058);
nand U1417 (N_1417,N_1061,N_1149);
xnor U1418 (N_1418,N_1135,N_1063);
nor U1419 (N_1419,N_1098,N_1035);
or U1420 (N_1420,N_1004,N_1005);
xnor U1421 (N_1421,N_1028,N_1231);
xor U1422 (N_1422,N_1110,N_1080);
xor U1423 (N_1423,N_1078,N_1164);
nand U1424 (N_1424,N_1118,N_1135);
and U1425 (N_1425,N_1243,N_1183);
nand U1426 (N_1426,N_1106,N_1203);
nand U1427 (N_1427,N_1195,N_1077);
and U1428 (N_1428,N_1087,N_1148);
nand U1429 (N_1429,N_1170,N_1197);
nand U1430 (N_1430,N_1163,N_1147);
or U1431 (N_1431,N_1126,N_1105);
and U1432 (N_1432,N_1247,N_1185);
or U1433 (N_1433,N_1002,N_1192);
and U1434 (N_1434,N_1068,N_1075);
nand U1435 (N_1435,N_1152,N_1161);
or U1436 (N_1436,N_1028,N_1034);
and U1437 (N_1437,N_1026,N_1217);
xnor U1438 (N_1438,N_1042,N_1148);
nor U1439 (N_1439,N_1101,N_1165);
xor U1440 (N_1440,N_1237,N_1027);
nor U1441 (N_1441,N_1217,N_1072);
or U1442 (N_1442,N_1207,N_1161);
nor U1443 (N_1443,N_1009,N_1130);
or U1444 (N_1444,N_1008,N_1237);
or U1445 (N_1445,N_1180,N_1155);
nand U1446 (N_1446,N_1083,N_1244);
and U1447 (N_1447,N_1143,N_1049);
and U1448 (N_1448,N_1012,N_1115);
and U1449 (N_1449,N_1083,N_1077);
nand U1450 (N_1450,N_1031,N_1142);
nand U1451 (N_1451,N_1055,N_1114);
nand U1452 (N_1452,N_1084,N_1143);
nand U1453 (N_1453,N_1064,N_1209);
or U1454 (N_1454,N_1017,N_1068);
xor U1455 (N_1455,N_1152,N_1102);
xnor U1456 (N_1456,N_1038,N_1210);
nor U1457 (N_1457,N_1054,N_1238);
or U1458 (N_1458,N_1171,N_1117);
nor U1459 (N_1459,N_1196,N_1150);
or U1460 (N_1460,N_1218,N_1023);
or U1461 (N_1461,N_1208,N_1033);
nand U1462 (N_1462,N_1228,N_1121);
xnor U1463 (N_1463,N_1023,N_1242);
nand U1464 (N_1464,N_1174,N_1048);
nor U1465 (N_1465,N_1100,N_1026);
and U1466 (N_1466,N_1071,N_1156);
nand U1467 (N_1467,N_1031,N_1005);
nand U1468 (N_1468,N_1247,N_1019);
nand U1469 (N_1469,N_1082,N_1230);
or U1470 (N_1470,N_1146,N_1189);
xor U1471 (N_1471,N_1095,N_1116);
nor U1472 (N_1472,N_1123,N_1119);
and U1473 (N_1473,N_1243,N_1125);
nand U1474 (N_1474,N_1102,N_1077);
or U1475 (N_1475,N_1110,N_1238);
or U1476 (N_1476,N_1135,N_1188);
nand U1477 (N_1477,N_1083,N_1223);
or U1478 (N_1478,N_1106,N_1023);
nand U1479 (N_1479,N_1208,N_1212);
xnor U1480 (N_1480,N_1157,N_1072);
nor U1481 (N_1481,N_1247,N_1178);
nand U1482 (N_1482,N_1228,N_1100);
xnor U1483 (N_1483,N_1098,N_1151);
and U1484 (N_1484,N_1146,N_1043);
or U1485 (N_1485,N_1062,N_1098);
xor U1486 (N_1486,N_1214,N_1057);
nand U1487 (N_1487,N_1025,N_1212);
and U1488 (N_1488,N_1090,N_1144);
nor U1489 (N_1489,N_1208,N_1247);
nand U1490 (N_1490,N_1100,N_1174);
or U1491 (N_1491,N_1066,N_1125);
and U1492 (N_1492,N_1087,N_1191);
nand U1493 (N_1493,N_1051,N_1057);
and U1494 (N_1494,N_1067,N_1025);
nor U1495 (N_1495,N_1199,N_1016);
xnor U1496 (N_1496,N_1069,N_1124);
or U1497 (N_1497,N_1117,N_1227);
nor U1498 (N_1498,N_1152,N_1222);
and U1499 (N_1499,N_1090,N_1165);
nand U1500 (N_1500,N_1258,N_1453);
nor U1501 (N_1501,N_1434,N_1382);
nand U1502 (N_1502,N_1479,N_1406);
nor U1503 (N_1503,N_1441,N_1271);
nor U1504 (N_1504,N_1426,N_1357);
nor U1505 (N_1505,N_1279,N_1308);
and U1506 (N_1506,N_1262,N_1338);
nor U1507 (N_1507,N_1335,N_1344);
and U1508 (N_1508,N_1389,N_1469);
nor U1509 (N_1509,N_1294,N_1260);
nor U1510 (N_1510,N_1359,N_1325);
xnor U1511 (N_1511,N_1440,N_1489);
xor U1512 (N_1512,N_1435,N_1473);
or U1513 (N_1513,N_1345,N_1298);
xnor U1514 (N_1514,N_1418,N_1485);
and U1515 (N_1515,N_1276,N_1466);
or U1516 (N_1516,N_1456,N_1307);
and U1517 (N_1517,N_1468,N_1402);
xnor U1518 (N_1518,N_1495,N_1322);
or U1519 (N_1519,N_1302,N_1459);
nand U1520 (N_1520,N_1331,N_1347);
or U1521 (N_1521,N_1269,N_1285);
nor U1522 (N_1522,N_1481,N_1482);
nor U1523 (N_1523,N_1278,N_1341);
or U1524 (N_1524,N_1484,N_1442);
or U1525 (N_1525,N_1405,N_1305);
nand U1526 (N_1526,N_1490,N_1355);
nor U1527 (N_1527,N_1300,N_1493);
or U1528 (N_1528,N_1461,N_1398);
nor U1529 (N_1529,N_1358,N_1403);
xnor U1530 (N_1530,N_1264,N_1324);
nor U1531 (N_1531,N_1304,N_1366);
nand U1532 (N_1532,N_1370,N_1392);
or U1533 (N_1533,N_1457,N_1272);
and U1534 (N_1534,N_1429,N_1374);
or U1535 (N_1535,N_1477,N_1250);
xor U1536 (N_1536,N_1399,N_1404);
or U1537 (N_1537,N_1474,N_1417);
or U1538 (N_1538,N_1336,N_1386);
or U1539 (N_1539,N_1314,N_1467);
nor U1540 (N_1540,N_1444,N_1446);
and U1541 (N_1541,N_1257,N_1369);
or U1542 (N_1542,N_1259,N_1261);
nand U1543 (N_1543,N_1497,N_1330);
nand U1544 (N_1544,N_1373,N_1313);
xnor U1545 (N_1545,N_1408,N_1372);
or U1546 (N_1546,N_1309,N_1475);
or U1547 (N_1547,N_1430,N_1470);
xor U1548 (N_1548,N_1351,N_1471);
xnor U1549 (N_1549,N_1480,N_1385);
or U1550 (N_1550,N_1329,N_1353);
or U1551 (N_1551,N_1312,N_1360);
nand U1552 (N_1552,N_1340,N_1422);
nand U1553 (N_1553,N_1281,N_1303);
and U1554 (N_1554,N_1296,N_1295);
nand U1555 (N_1555,N_1381,N_1445);
and U1556 (N_1556,N_1299,N_1428);
xor U1557 (N_1557,N_1443,N_1253);
xor U1558 (N_1558,N_1297,N_1301);
nor U1559 (N_1559,N_1454,N_1394);
or U1560 (N_1560,N_1488,N_1432);
and U1561 (N_1561,N_1458,N_1275);
nor U1562 (N_1562,N_1496,N_1363);
xor U1563 (N_1563,N_1286,N_1375);
nor U1564 (N_1564,N_1319,N_1327);
or U1565 (N_1565,N_1362,N_1255);
nand U1566 (N_1566,N_1395,N_1317);
or U1567 (N_1567,N_1437,N_1499);
nand U1568 (N_1568,N_1332,N_1265);
and U1569 (N_1569,N_1311,N_1333);
nand U1570 (N_1570,N_1256,N_1465);
and U1571 (N_1571,N_1483,N_1449);
or U1572 (N_1572,N_1321,N_1411);
nand U1573 (N_1573,N_1414,N_1326);
nand U1574 (N_1574,N_1270,N_1419);
or U1575 (N_1575,N_1284,N_1424);
or U1576 (N_1576,N_1288,N_1439);
or U1577 (N_1577,N_1415,N_1455);
or U1578 (N_1578,N_1486,N_1320);
xnor U1579 (N_1579,N_1447,N_1282);
nand U1580 (N_1580,N_1409,N_1384);
xor U1581 (N_1581,N_1252,N_1268);
nand U1582 (N_1582,N_1462,N_1316);
or U1583 (N_1583,N_1431,N_1400);
and U1584 (N_1584,N_1361,N_1349);
and U1585 (N_1585,N_1451,N_1263);
or U1586 (N_1586,N_1342,N_1254);
and U1587 (N_1587,N_1354,N_1396);
or U1588 (N_1588,N_1464,N_1387);
and U1589 (N_1589,N_1380,N_1390);
nand U1590 (N_1590,N_1352,N_1339);
or U1591 (N_1591,N_1377,N_1448);
and U1592 (N_1592,N_1425,N_1472);
xor U1593 (N_1593,N_1476,N_1371);
nand U1594 (N_1594,N_1498,N_1343);
or U1595 (N_1595,N_1350,N_1287);
nor U1596 (N_1596,N_1289,N_1266);
or U1597 (N_1597,N_1436,N_1397);
or U1598 (N_1598,N_1376,N_1412);
or U1599 (N_1599,N_1334,N_1492);
xnor U1600 (N_1600,N_1267,N_1423);
and U1601 (N_1601,N_1478,N_1416);
xnor U1602 (N_1602,N_1348,N_1291);
nor U1603 (N_1603,N_1420,N_1421);
and U1604 (N_1604,N_1251,N_1337);
nor U1605 (N_1605,N_1410,N_1310);
xnor U1606 (N_1606,N_1401,N_1407);
xor U1607 (N_1607,N_1323,N_1346);
nand U1608 (N_1608,N_1438,N_1487);
and U1609 (N_1609,N_1315,N_1463);
or U1610 (N_1610,N_1433,N_1283);
nand U1611 (N_1611,N_1367,N_1452);
or U1612 (N_1612,N_1318,N_1388);
nand U1613 (N_1613,N_1274,N_1450);
or U1614 (N_1614,N_1273,N_1306);
or U1615 (N_1615,N_1328,N_1292);
nor U1616 (N_1616,N_1460,N_1378);
nor U1617 (N_1617,N_1494,N_1491);
xor U1618 (N_1618,N_1280,N_1393);
xnor U1619 (N_1619,N_1290,N_1365);
and U1620 (N_1620,N_1293,N_1391);
and U1621 (N_1621,N_1356,N_1364);
nor U1622 (N_1622,N_1379,N_1427);
or U1623 (N_1623,N_1277,N_1413);
and U1624 (N_1624,N_1368,N_1383);
nand U1625 (N_1625,N_1258,N_1403);
and U1626 (N_1626,N_1321,N_1387);
xor U1627 (N_1627,N_1394,N_1483);
and U1628 (N_1628,N_1302,N_1404);
nand U1629 (N_1629,N_1329,N_1449);
xnor U1630 (N_1630,N_1313,N_1333);
xor U1631 (N_1631,N_1297,N_1381);
nor U1632 (N_1632,N_1321,N_1384);
and U1633 (N_1633,N_1252,N_1491);
nor U1634 (N_1634,N_1419,N_1338);
nand U1635 (N_1635,N_1279,N_1415);
or U1636 (N_1636,N_1254,N_1279);
nand U1637 (N_1637,N_1299,N_1467);
nand U1638 (N_1638,N_1474,N_1351);
nor U1639 (N_1639,N_1281,N_1256);
nor U1640 (N_1640,N_1432,N_1359);
or U1641 (N_1641,N_1349,N_1325);
or U1642 (N_1642,N_1271,N_1367);
and U1643 (N_1643,N_1306,N_1439);
nand U1644 (N_1644,N_1321,N_1296);
nand U1645 (N_1645,N_1488,N_1407);
xnor U1646 (N_1646,N_1348,N_1487);
nand U1647 (N_1647,N_1286,N_1449);
nand U1648 (N_1648,N_1458,N_1392);
xor U1649 (N_1649,N_1276,N_1421);
xnor U1650 (N_1650,N_1403,N_1332);
or U1651 (N_1651,N_1304,N_1484);
nand U1652 (N_1652,N_1457,N_1437);
nor U1653 (N_1653,N_1310,N_1265);
or U1654 (N_1654,N_1278,N_1340);
nand U1655 (N_1655,N_1303,N_1360);
or U1656 (N_1656,N_1422,N_1342);
or U1657 (N_1657,N_1250,N_1292);
nand U1658 (N_1658,N_1397,N_1475);
nor U1659 (N_1659,N_1452,N_1336);
xnor U1660 (N_1660,N_1436,N_1359);
and U1661 (N_1661,N_1343,N_1385);
and U1662 (N_1662,N_1373,N_1455);
or U1663 (N_1663,N_1352,N_1357);
xnor U1664 (N_1664,N_1309,N_1448);
nor U1665 (N_1665,N_1429,N_1306);
xnor U1666 (N_1666,N_1311,N_1451);
nand U1667 (N_1667,N_1250,N_1367);
nand U1668 (N_1668,N_1397,N_1371);
or U1669 (N_1669,N_1338,N_1325);
or U1670 (N_1670,N_1496,N_1464);
and U1671 (N_1671,N_1496,N_1259);
and U1672 (N_1672,N_1367,N_1279);
nand U1673 (N_1673,N_1483,N_1406);
nand U1674 (N_1674,N_1448,N_1404);
nor U1675 (N_1675,N_1256,N_1287);
nor U1676 (N_1676,N_1369,N_1382);
nor U1677 (N_1677,N_1496,N_1492);
nand U1678 (N_1678,N_1270,N_1303);
nor U1679 (N_1679,N_1330,N_1325);
nand U1680 (N_1680,N_1380,N_1271);
nand U1681 (N_1681,N_1495,N_1288);
or U1682 (N_1682,N_1379,N_1393);
and U1683 (N_1683,N_1259,N_1443);
and U1684 (N_1684,N_1445,N_1376);
nor U1685 (N_1685,N_1357,N_1348);
xor U1686 (N_1686,N_1392,N_1386);
nand U1687 (N_1687,N_1299,N_1400);
nand U1688 (N_1688,N_1294,N_1495);
nor U1689 (N_1689,N_1431,N_1368);
and U1690 (N_1690,N_1303,N_1462);
or U1691 (N_1691,N_1495,N_1463);
or U1692 (N_1692,N_1491,N_1400);
or U1693 (N_1693,N_1490,N_1385);
or U1694 (N_1694,N_1351,N_1316);
nor U1695 (N_1695,N_1272,N_1296);
and U1696 (N_1696,N_1394,N_1411);
xnor U1697 (N_1697,N_1376,N_1341);
nand U1698 (N_1698,N_1437,N_1468);
and U1699 (N_1699,N_1316,N_1420);
xor U1700 (N_1700,N_1371,N_1387);
or U1701 (N_1701,N_1468,N_1317);
nand U1702 (N_1702,N_1286,N_1281);
nand U1703 (N_1703,N_1311,N_1385);
nand U1704 (N_1704,N_1349,N_1271);
or U1705 (N_1705,N_1375,N_1305);
nor U1706 (N_1706,N_1266,N_1421);
or U1707 (N_1707,N_1354,N_1494);
nor U1708 (N_1708,N_1392,N_1423);
or U1709 (N_1709,N_1442,N_1318);
nor U1710 (N_1710,N_1258,N_1288);
or U1711 (N_1711,N_1267,N_1379);
xnor U1712 (N_1712,N_1469,N_1387);
xor U1713 (N_1713,N_1292,N_1374);
xor U1714 (N_1714,N_1364,N_1346);
and U1715 (N_1715,N_1380,N_1440);
nand U1716 (N_1716,N_1321,N_1252);
and U1717 (N_1717,N_1345,N_1432);
nor U1718 (N_1718,N_1289,N_1307);
nor U1719 (N_1719,N_1489,N_1465);
xor U1720 (N_1720,N_1459,N_1425);
or U1721 (N_1721,N_1498,N_1415);
and U1722 (N_1722,N_1372,N_1303);
and U1723 (N_1723,N_1484,N_1319);
or U1724 (N_1724,N_1270,N_1499);
nand U1725 (N_1725,N_1422,N_1486);
and U1726 (N_1726,N_1253,N_1400);
and U1727 (N_1727,N_1367,N_1381);
or U1728 (N_1728,N_1455,N_1436);
or U1729 (N_1729,N_1265,N_1489);
or U1730 (N_1730,N_1439,N_1265);
nand U1731 (N_1731,N_1469,N_1485);
or U1732 (N_1732,N_1436,N_1403);
or U1733 (N_1733,N_1458,N_1370);
xnor U1734 (N_1734,N_1452,N_1371);
and U1735 (N_1735,N_1361,N_1442);
xor U1736 (N_1736,N_1321,N_1351);
nor U1737 (N_1737,N_1253,N_1380);
nor U1738 (N_1738,N_1295,N_1491);
nor U1739 (N_1739,N_1301,N_1265);
or U1740 (N_1740,N_1293,N_1468);
or U1741 (N_1741,N_1370,N_1343);
and U1742 (N_1742,N_1435,N_1267);
and U1743 (N_1743,N_1277,N_1454);
xnor U1744 (N_1744,N_1260,N_1308);
nand U1745 (N_1745,N_1390,N_1394);
xor U1746 (N_1746,N_1357,N_1345);
nand U1747 (N_1747,N_1299,N_1436);
xor U1748 (N_1748,N_1405,N_1359);
and U1749 (N_1749,N_1285,N_1340);
nor U1750 (N_1750,N_1675,N_1524);
and U1751 (N_1751,N_1585,N_1501);
nor U1752 (N_1752,N_1632,N_1694);
nand U1753 (N_1753,N_1627,N_1701);
nand U1754 (N_1754,N_1713,N_1527);
nor U1755 (N_1755,N_1715,N_1615);
and U1756 (N_1756,N_1595,N_1546);
or U1757 (N_1757,N_1616,N_1558);
or U1758 (N_1758,N_1673,N_1730);
xnor U1759 (N_1759,N_1676,N_1657);
or U1760 (N_1760,N_1606,N_1552);
or U1761 (N_1761,N_1709,N_1555);
nand U1762 (N_1762,N_1681,N_1742);
xor U1763 (N_1763,N_1559,N_1581);
or U1764 (N_1764,N_1579,N_1703);
nand U1765 (N_1765,N_1593,N_1688);
nor U1766 (N_1766,N_1622,N_1652);
nor U1767 (N_1767,N_1729,N_1698);
and U1768 (N_1768,N_1537,N_1726);
nand U1769 (N_1769,N_1695,N_1665);
or U1770 (N_1770,N_1594,N_1566);
xor U1771 (N_1771,N_1692,N_1656);
and U1772 (N_1772,N_1533,N_1690);
nor U1773 (N_1773,N_1516,N_1658);
and U1774 (N_1774,N_1597,N_1560);
nand U1775 (N_1775,N_1663,N_1738);
and U1776 (N_1776,N_1633,N_1635);
xnor U1777 (N_1777,N_1746,N_1519);
or U1778 (N_1778,N_1741,N_1564);
and U1779 (N_1779,N_1568,N_1655);
or U1780 (N_1780,N_1509,N_1605);
or U1781 (N_1781,N_1708,N_1562);
nor U1782 (N_1782,N_1611,N_1721);
or U1783 (N_1783,N_1569,N_1660);
nand U1784 (N_1784,N_1506,N_1630);
nor U1785 (N_1785,N_1667,N_1666);
nand U1786 (N_1786,N_1526,N_1674);
xnor U1787 (N_1787,N_1700,N_1522);
nor U1788 (N_1788,N_1542,N_1580);
nand U1789 (N_1789,N_1511,N_1531);
and U1790 (N_1790,N_1724,N_1710);
nand U1791 (N_1791,N_1685,N_1554);
and U1792 (N_1792,N_1601,N_1696);
or U1793 (N_1793,N_1647,N_1587);
xnor U1794 (N_1794,N_1716,N_1736);
nand U1795 (N_1795,N_1661,N_1548);
nand U1796 (N_1796,N_1590,N_1505);
and U1797 (N_1797,N_1515,N_1586);
nor U1798 (N_1798,N_1639,N_1550);
xnor U1799 (N_1799,N_1651,N_1598);
or U1800 (N_1800,N_1603,N_1504);
xor U1801 (N_1801,N_1722,N_1677);
or U1802 (N_1802,N_1507,N_1572);
and U1803 (N_1803,N_1679,N_1536);
nand U1804 (N_1804,N_1547,N_1529);
xnor U1805 (N_1805,N_1743,N_1592);
nor U1806 (N_1806,N_1517,N_1664);
or U1807 (N_1807,N_1570,N_1620);
nor U1808 (N_1808,N_1723,N_1596);
and U1809 (N_1809,N_1749,N_1699);
xnor U1810 (N_1810,N_1577,N_1539);
or U1811 (N_1811,N_1640,N_1512);
xnor U1812 (N_1812,N_1538,N_1565);
nor U1813 (N_1813,N_1563,N_1528);
or U1814 (N_1814,N_1520,N_1574);
and U1815 (N_1815,N_1613,N_1745);
nand U1816 (N_1816,N_1602,N_1544);
and U1817 (N_1817,N_1588,N_1582);
nor U1818 (N_1818,N_1553,N_1631);
xnor U1819 (N_1819,N_1567,N_1600);
or U1820 (N_1820,N_1648,N_1521);
and U1821 (N_1821,N_1735,N_1610);
or U1822 (N_1822,N_1625,N_1671);
nor U1823 (N_1823,N_1619,N_1670);
xor U1824 (N_1824,N_1662,N_1518);
or U1825 (N_1825,N_1530,N_1689);
xnor U1826 (N_1826,N_1669,N_1556);
xnor U1827 (N_1827,N_1653,N_1624);
nor U1828 (N_1828,N_1514,N_1734);
or U1829 (N_1829,N_1604,N_1683);
nor U1830 (N_1830,N_1628,N_1584);
and U1831 (N_1831,N_1644,N_1634);
nor U1832 (N_1832,N_1659,N_1702);
and U1833 (N_1833,N_1682,N_1589);
and U1834 (N_1834,N_1740,N_1561);
and U1835 (N_1835,N_1733,N_1711);
and U1836 (N_1836,N_1502,N_1575);
nand U1837 (N_1837,N_1571,N_1618);
and U1838 (N_1838,N_1557,N_1599);
and U1839 (N_1839,N_1612,N_1614);
and U1840 (N_1840,N_1646,N_1532);
or U1841 (N_1841,N_1525,N_1649);
nor U1842 (N_1842,N_1500,N_1642);
nor U1843 (N_1843,N_1744,N_1576);
xnor U1844 (N_1844,N_1704,N_1629);
xor U1845 (N_1845,N_1551,N_1684);
or U1846 (N_1846,N_1678,N_1541);
or U1847 (N_1847,N_1617,N_1672);
or U1848 (N_1848,N_1623,N_1712);
nand U1849 (N_1849,N_1641,N_1643);
nand U1850 (N_1850,N_1707,N_1697);
and U1851 (N_1851,N_1705,N_1645);
nor U1852 (N_1852,N_1719,N_1739);
nand U1853 (N_1853,N_1510,N_1732);
or U1854 (N_1854,N_1731,N_1609);
xnor U1855 (N_1855,N_1728,N_1540);
nand U1856 (N_1856,N_1687,N_1654);
nor U1857 (N_1857,N_1714,N_1718);
nor U1858 (N_1858,N_1650,N_1573);
or U1859 (N_1859,N_1534,N_1513);
nor U1860 (N_1860,N_1578,N_1747);
or U1861 (N_1861,N_1638,N_1636);
xor U1862 (N_1862,N_1748,N_1717);
nor U1863 (N_1863,N_1680,N_1686);
nand U1864 (N_1864,N_1545,N_1591);
or U1865 (N_1865,N_1583,N_1737);
or U1866 (N_1866,N_1727,N_1508);
and U1867 (N_1867,N_1549,N_1668);
nor U1868 (N_1868,N_1535,N_1720);
nand U1869 (N_1869,N_1608,N_1691);
nand U1870 (N_1870,N_1706,N_1607);
or U1871 (N_1871,N_1725,N_1503);
xor U1872 (N_1872,N_1626,N_1621);
nor U1873 (N_1873,N_1693,N_1637);
xnor U1874 (N_1874,N_1523,N_1543);
nand U1875 (N_1875,N_1703,N_1586);
and U1876 (N_1876,N_1745,N_1674);
xor U1877 (N_1877,N_1608,N_1702);
xor U1878 (N_1878,N_1607,N_1709);
or U1879 (N_1879,N_1632,N_1512);
and U1880 (N_1880,N_1604,N_1503);
and U1881 (N_1881,N_1506,N_1558);
or U1882 (N_1882,N_1548,N_1646);
nor U1883 (N_1883,N_1506,N_1697);
nand U1884 (N_1884,N_1504,N_1661);
or U1885 (N_1885,N_1500,N_1532);
or U1886 (N_1886,N_1708,N_1726);
xor U1887 (N_1887,N_1732,N_1672);
xor U1888 (N_1888,N_1589,N_1725);
nor U1889 (N_1889,N_1614,N_1693);
or U1890 (N_1890,N_1703,N_1523);
and U1891 (N_1891,N_1588,N_1722);
and U1892 (N_1892,N_1661,N_1512);
or U1893 (N_1893,N_1601,N_1654);
xor U1894 (N_1894,N_1649,N_1504);
nor U1895 (N_1895,N_1657,N_1542);
or U1896 (N_1896,N_1732,N_1500);
nand U1897 (N_1897,N_1666,N_1712);
and U1898 (N_1898,N_1735,N_1646);
or U1899 (N_1899,N_1563,N_1660);
and U1900 (N_1900,N_1630,N_1667);
nor U1901 (N_1901,N_1545,N_1568);
xor U1902 (N_1902,N_1603,N_1676);
and U1903 (N_1903,N_1710,N_1536);
nor U1904 (N_1904,N_1733,N_1742);
nor U1905 (N_1905,N_1571,N_1739);
nand U1906 (N_1906,N_1501,N_1644);
and U1907 (N_1907,N_1628,N_1509);
nor U1908 (N_1908,N_1547,N_1749);
nor U1909 (N_1909,N_1724,N_1545);
xnor U1910 (N_1910,N_1659,N_1559);
xor U1911 (N_1911,N_1695,N_1529);
nand U1912 (N_1912,N_1513,N_1665);
nor U1913 (N_1913,N_1682,N_1618);
xnor U1914 (N_1914,N_1670,N_1623);
or U1915 (N_1915,N_1714,N_1570);
xnor U1916 (N_1916,N_1631,N_1516);
nand U1917 (N_1917,N_1747,N_1719);
or U1918 (N_1918,N_1584,N_1581);
and U1919 (N_1919,N_1576,N_1746);
nand U1920 (N_1920,N_1618,N_1653);
nor U1921 (N_1921,N_1744,N_1537);
and U1922 (N_1922,N_1500,N_1573);
or U1923 (N_1923,N_1669,N_1628);
and U1924 (N_1924,N_1671,N_1602);
and U1925 (N_1925,N_1626,N_1530);
xnor U1926 (N_1926,N_1663,N_1591);
nand U1927 (N_1927,N_1642,N_1530);
and U1928 (N_1928,N_1549,N_1584);
nor U1929 (N_1929,N_1622,N_1694);
or U1930 (N_1930,N_1677,N_1608);
and U1931 (N_1931,N_1746,N_1653);
xor U1932 (N_1932,N_1701,N_1706);
nor U1933 (N_1933,N_1711,N_1652);
xnor U1934 (N_1934,N_1603,N_1746);
or U1935 (N_1935,N_1744,N_1669);
nand U1936 (N_1936,N_1530,N_1578);
nor U1937 (N_1937,N_1638,N_1513);
nor U1938 (N_1938,N_1505,N_1642);
nand U1939 (N_1939,N_1547,N_1510);
nand U1940 (N_1940,N_1636,N_1669);
xor U1941 (N_1941,N_1583,N_1649);
nor U1942 (N_1942,N_1511,N_1674);
nand U1943 (N_1943,N_1504,N_1552);
nand U1944 (N_1944,N_1699,N_1589);
nor U1945 (N_1945,N_1569,N_1525);
nand U1946 (N_1946,N_1690,N_1542);
nand U1947 (N_1947,N_1684,N_1742);
or U1948 (N_1948,N_1615,N_1633);
or U1949 (N_1949,N_1635,N_1544);
or U1950 (N_1950,N_1668,N_1652);
and U1951 (N_1951,N_1522,N_1650);
nor U1952 (N_1952,N_1697,N_1621);
xnor U1953 (N_1953,N_1563,N_1531);
nand U1954 (N_1954,N_1618,N_1737);
nor U1955 (N_1955,N_1661,N_1547);
or U1956 (N_1956,N_1743,N_1633);
nor U1957 (N_1957,N_1620,N_1679);
nor U1958 (N_1958,N_1539,N_1519);
nand U1959 (N_1959,N_1673,N_1728);
and U1960 (N_1960,N_1619,N_1667);
or U1961 (N_1961,N_1617,N_1599);
nor U1962 (N_1962,N_1698,N_1681);
xor U1963 (N_1963,N_1513,N_1714);
nand U1964 (N_1964,N_1693,N_1570);
nand U1965 (N_1965,N_1730,N_1522);
xnor U1966 (N_1966,N_1631,N_1704);
and U1967 (N_1967,N_1520,N_1666);
and U1968 (N_1968,N_1729,N_1689);
or U1969 (N_1969,N_1708,N_1727);
nor U1970 (N_1970,N_1608,N_1693);
xor U1971 (N_1971,N_1741,N_1610);
and U1972 (N_1972,N_1717,N_1702);
or U1973 (N_1973,N_1704,N_1650);
or U1974 (N_1974,N_1548,N_1522);
and U1975 (N_1975,N_1557,N_1646);
xnor U1976 (N_1976,N_1553,N_1534);
nand U1977 (N_1977,N_1504,N_1503);
nor U1978 (N_1978,N_1670,N_1569);
or U1979 (N_1979,N_1626,N_1680);
nor U1980 (N_1980,N_1633,N_1737);
xnor U1981 (N_1981,N_1640,N_1502);
xnor U1982 (N_1982,N_1678,N_1591);
or U1983 (N_1983,N_1501,N_1615);
nand U1984 (N_1984,N_1733,N_1503);
nor U1985 (N_1985,N_1518,N_1575);
and U1986 (N_1986,N_1518,N_1550);
or U1987 (N_1987,N_1601,N_1569);
or U1988 (N_1988,N_1638,N_1640);
or U1989 (N_1989,N_1692,N_1740);
or U1990 (N_1990,N_1724,N_1675);
nand U1991 (N_1991,N_1589,N_1646);
nor U1992 (N_1992,N_1577,N_1529);
nand U1993 (N_1993,N_1628,N_1524);
nand U1994 (N_1994,N_1662,N_1591);
nand U1995 (N_1995,N_1598,N_1589);
and U1996 (N_1996,N_1640,N_1716);
nand U1997 (N_1997,N_1513,N_1724);
and U1998 (N_1998,N_1542,N_1724);
nand U1999 (N_1999,N_1657,N_1643);
nor U2000 (N_2000,N_1999,N_1804);
and U2001 (N_2001,N_1900,N_1887);
nand U2002 (N_2002,N_1920,N_1873);
xor U2003 (N_2003,N_1846,N_1946);
xnor U2004 (N_2004,N_1784,N_1943);
nand U2005 (N_2005,N_1826,N_1782);
nor U2006 (N_2006,N_1908,N_1811);
or U2007 (N_2007,N_1903,N_1750);
xnor U2008 (N_2008,N_1914,N_1842);
xnor U2009 (N_2009,N_1978,N_1785);
xor U2010 (N_2010,N_1951,N_1921);
nor U2011 (N_2011,N_1995,N_1828);
xor U2012 (N_2012,N_1917,N_1923);
nor U2013 (N_2013,N_1896,N_1849);
and U2014 (N_2014,N_1988,N_1947);
and U2015 (N_2015,N_1948,N_1837);
or U2016 (N_2016,N_1961,N_1981);
xnor U2017 (N_2017,N_1845,N_1895);
nand U2018 (N_2018,N_1971,N_1833);
xnor U2019 (N_2019,N_1765,N_1994);
nand U2020 (N_2020,N_1788,N_1777);
nor U2021 (N_2021,N_1773,N_1862);
xor U2022 (N_2022,N_1958,N_1997);
nor U2023 (N_2023,N_1753,N_1752);
nand U2024 (N_2024,N_1930,N_1793);
or U2025 (N_2025,N_1822,N_1913);
or U2026 (N_2026,N_1912,N_1816);
and U2027 (N_2027,N_1883,N_1976);
nor U2028 (N_2028,N_1910,N_1904);
nor U2029 (N_2029,N_1852,N_1808);
or U2030 (N_2030,N_1843,N_1969);
nor U2031 (N_2031,N_1933,N_1834);
xor U2032 (N_2032,N_1878,N_1998);
or U2033 (N_2033,N_1757,N_1957);
or U2034 (N_2034,N_1906,N_1877);
nor U2035 (N_2035,N_1956,N_1886);
and U2036 (N_2036,N_1876,N_1861);
and U2037 (N_2037,N_1963,N_1893);
and U2038 (N_2038,N_1848,N_1991);
or U2039 (N_2039,N_1954,N_1823);
and U2040 (N_2040,N_1813,N_1966);
xnor U2041 (N_2041,N_1818,N_1984);
or U2042 (N_2042,N_1800,N_1891);
nand U2043 (N_2043,N_1875,N_1760);
nand U2044 (N_2044,N_1856,N_1769);
or U2045 (N_2045,N_1858,N_1841);
and U2046 (N_2046,N_1840,N_1980);
or U2047 (N_2047,N_1795,N_1829);
nand U2048 (N_2048,N_1927,N_1867);
nor U2049 (N_2049,N_1938,N_1815);
nand U2050 (N_2050,N_1871,N_1766);
and U2051 (N_2051,N_1780,N_1960);
nor U2052 (N_2052,N_1870,N_1844);
xnor U2053 (N_2053,N_1874,N_1770);
or U2054 (N_2054,N_1803,N_1909);
and U2055 (N_2055,N_1790,N_1810);
nor U2056 (N_2056,N_1789,N_1787);
nand U2057 (N_2057,N_1799,N_1935);
nor U2058 (N_2058,N_1907,N_1776);
nand U2059 (N_2059,N_1827,N_1945);
xor U2060 (N_2060,N_1940,N_1755);
or U2061 (N_2061,N_1854,N_1899);
nor U2062 (N_2062,N_1764,N_1898);
xnor U2063 (N_2063,N_1949,N_1855);
nor U2064 (N_2064,N_1791,N_1825);
or U2065 (N_2065,N_1996,N_1866);
nor U2066 (N_2066,N_1953,N_1754);
and U2067 (N_2067,N_1925,N_1761);
nor U2068 (N_2068,N_1993,N_1889);
and U2069 (N_2069,N_1865,N_1763);
nor U2070 (N_2070,N_1794,N_1892);
xor U2071 (N_2071,N_1885,N_1836);
nand U2072 (N_2072,N_1894,N_1902);
or U2073 (N_2073,N_1942,N_1879);
nand U2074 (N_2074,N_1857,N_1934);
nand U2075 (N_2075,N_1916,N_1937);
nand U2076 (N_2076,N_1897,N_1905);
xnor U2077 (N_2077,N_1987,N_1758);
xor U2078 (N_2078,N_1944,N_1767);
xnor U2079 (N_2079,N_1792,N_1964);
or U2080 (N_2080,N_1973,N_1809);
nand U2081 (N_2081,N_1779,N_1989);
or U2082 (N_2082,N_1839,N_1796);
xnor U2083 (N_2083,N_1983,N_1962);
xor U2084 (N_2084,N_1884,N_1819);
nand U2085 (N_2085,N_1932,N_1778);
xnor U2086 (N_2086,N_1814,N_1798);
nand U2087 (N_2087,N_1880,N_1941);
nor U2088 (N_2088,N_1919,N_1952);
nor U2089 (N_2089,N_1824,N_1847);
nand U2090 (N_2090,N_1982,N_1979);
or U2091 (N_2091,N_1859,N_1901);
nand U2092 (N_2092,N_1939,N_1911);
nor U2093 (N_2093,N_1805,N_1801);
xor U2094 (N_2094,N_1924,N_1967);
nand U2095 (N_2095,N_1812,N_1781);
and U2096 (N_2096,N_1955,N_1950);
and U2097 (N_2097,N_1817,N_1918);
nand U2098 (N_2098,N_1835,N_1868);
nand U2099 (N_2099,N_1970,N_1882);
and U2100 (N_2100,N_1931,N_1863);
xnor U2101 (N_2101,N_1965,N_1771);
nor U2102 (N_2102,N_1797,N_1890);
nor U2103 (N_2103,N_1775,N_1972);
xor U2104 (N_2104,N_1802,N_1977);
and U2105 (N_2105,N_1990,N_1928);
xor U2106 (N_2106,N_1915,N_1831);
or U2107 (N_2107,N_1986,N_1807);
xor U2108 (N_2108,N_1783,N_1772);
xnor U2109 (N_2109,N_1968,N_1830);
nand U2110 (N_2110,N_1926,N_1992);
xnor U2111 (N_2111,N_1936,N_1860);
xnor U2112 (N_2112,N_1864,N_1806);
and U2113 (N_2113,N_1959,N_1768);
or U2114 (N_2114,N_1985,N_1869);
and U2115 (N_2115,N_1888,N_1759);
xnor U2116 (N_2116,N_1821,N_1872);
xor U2117 (N_2117,N_1832,N_1929);
xor U2118 (N_2118,N_1851,N_1881);
nand U2119 (N_2119,N_1756,N_1922);
nor U2120 (N_2120,N_1838,N_1975);
nand U2121 (N_2121,N_1762,N_1774);
or U2122 (N_2122,N_1974,N_1853);
or U2123 (N_2123,N_1786,N_1850);
nor U2124 (N_2124,N_1820,N_1751);
nor U2125 (N_2125,N_1932,N_1798);
nand U2126 (N_2126,N_1922,N_1961);
xor U2127 (N_2127,N_1848,N_1795);
and U2128 (N_2128,N_1977,N_1891);
xnor U2129 (N_2129,N_1903,N_1822);
nor U2130 (N_2130,N_1925,N_1764);
xnor U2131 (N_2131,N_1964,N_1829);
and U2132 (N_2132,N_1917,N_1857);
nand U2133 (N_2133,N_1822,N_1809);
nor U2134 (N_2134,N_1915,N_1842);
or U2135 (N_2135,N_1771,N_1765);
and U2136 (N_2136,N_1785,N_1933);
nor U2137 (N_2137,N_1899,N_1809);
or U2138 (N_2138,N_1867,N_1928);
or U2139 (N_2139,N_1809,N_1984);
and U2140 (N_2140,N_1776,N_1796);
nor U2141 (N_2141,N_1841,N_1856);
or U2142 (N_2142,N_1852,N_1999);
nor U2143 (N_2143,N_1879,N_1888);
nand U2144 (N_2144,N_1940,N_1793);
nor U2145 (N_2145,N_1994,N_1774);
nand U2146 (N_2146,N_1998,N_1874);
or U2147 (N_2147,N_1850,N_1900);
or U2148 (N_2148,N_1804,N_1850);
and U2149 (N_2149,N_1968,N_1831);
xor U2150 (N_2150,N_1916,N_1817);
nand U2151 (N_2151,N_1853,N_1885);
nor U2152 (N_2152,N_1799,N_1758);
or U2153 (N_2153,N_1844,N_1951);
nor U2154 (N_2154,N_1957,N_1804);
or U2155 (N_2155,N_1941,N_1836);
nor U2156 (N_2156,N_1783,N_1889);
nand U2157 (N_2157,N_1878,N_1983);
or U2158 (N_2158,N_1857,N_1778);
xnor U2159 (N_2159,N_1824,N_1821);
nand U2160 (N_2160,N_1890,N_1880);
nand U2161 (N_2161,N_1901,N_1868);
nor U2162 (N_2162,N_1858,N_1994);
xnor U2163 (N_2163,N_1844,N_1949);
and U2164 (N_2164,N_1761,N_1880);
nand U2165 (N_2165,N_1842,N_1840);
xor U2166 (N_2166,N_1971,N_1938);
or U2167 (N_2167,N_1823,N_1898);
and U2168 (N_2168,N_1928,N_1994);
or U2169 (N_2169,N_1905,N_1855);
or U2170 (N_2170,N_1846,N_1795);
nor U2171 (N_2171,N_1869,N_1759);
or U2172 (N_2172,N_1828,N_1933);
nand U2173 (N_2173,N_1875,N_1904);
xnor U2174 (N_2174,N_1845,N_1833);
nor U2175 (N_2175,N_1913,N_1904);
xnor U2176 (N_2176,N_1854,N_1792);
xor U2177 (N_2177,N_1764,N_1909);
xnor U2178 (N_2178,N_1897,N_1777);
xor U2179 (N_2179,N_1952,N_1899);
and U2180 (N_2180,N_1952,N_1867);
or U2181 (N_2181,N_1796,N_1909);
or U2182 (N_2182,N_1817,N_1771);
nor U2183 (N_2183,N_1824,N_1826);
nor U2184 (N_2184,N_1825,N_1997);
or U2185 (N_2185,N_1769,N_1854);
xor U2186 (N_2186,N_1823,N_1811);
and U2187 (N_2187,N_1998,N_1976);
xnor U2188 (N_2188,N_1937,N_1925);
or U2189 (N_2189,N_1905,N_1951);
xnor U2190 (N_2190,N_1896,N_1899);
xnor U2191 (N_2191,N_1835,N_1946);
nand U2192 (N_2192,N_1940,N_1988);
nand U2193 (N_2193,N_1771,N_1883);
and U2194 (N_2194,N_1841,N_1862);
nor U2195 (N_2195,N_1784,N_1967);
xor U2196 (N_2196,N_1784,N_1762);
nand U2197 (N_2197,N_1978,N_1923);
nand U2198 (N_2198,N_1987,N_1996);
or U2199 (N_2199,N_1759,N_1798);
and U2200 (N_2200,N_1999,N_1966);
or U2201 (N_2201,N_1946,N_1776);
nor U2202 (N_2202,N_1754,N_1752);
and U2203 (N_2203,N_1970,N_1760);
nor U2204 (N_2204,N_1856,N_1793);
nor U2205 (N_2205,N_1787,N_1954);
xnor U2206 (N_2206,N_1980,N_1954);
and U2207 (N_2207,N_1869,N_1979);
and U2208 (N_2208,N_1966,N_1894);
and U2209 (N_2209,N_1972,N_1760);
nand U2210 (N_2210,N_1996,N_1925);
nor U2211 (N_2211,N_1868,N_1780);
xnor U2212 (N_2212,N_1847,N_1999);
nor U2213 (N_2213,N_1955,N_1990);
xnor U2214 (N_2214,N_1987,N_1787);
nand U2215 (N_2215,N_1786,N_1834);
or U2216 (N_2216,N_1890,N_1838);
or U2217 (N_2217,N_1955,N_1803);
and U2218 (N_2218,N_1929,N_1988);
and U2219 (N_2219,N_1923,N_1803);
nand U2220 (N_2220,N_1808,N_1833);
xor U2221 (N_2221,N_1833,N_1967);
and U2222 (N_2222,N_1842,N_1841);
xor U2223 (N_2223,N_1751,N_1844);
xnor U2224 (N_2224,N_1966,N_1914);
or U2225 (N_2225,N_1927,N_1760);
or U2226 (N_2226,N_1990,N_1849);
or U2227 (N_2227,N_1879,N_1775);
nand U2228 (N_2228,N_1962,N_1836);
nand U2229 (N_2229,N_1910,N_1765);
or U2230 (N_2230,N_1830,N_1864);
and U2231 (N_2231,N_1824,N_1778);
xnor U2232 (N_2232,N_1809,N_1943);
nor U2233 (N_2233,N_1847,N_1806);
or U2234 (N_2234,N_1928,N_1815);
and U2235 (N_2235,N_1854,N_1816);
and U2236 (N_2236,N_1822,N_1828);
and U2237 (N_2237,N_1776,N_1982);
nand U2238 (N_2238,N_1826,N_1752);
nor U2239 (N_2239,N_1935,N_1994);
nor U2240 (N_2240,N_1843,N_1858);
and U2241 (N_2241,N_1912,N_1795);
nand U2242 (N_2242,N_1905,N_1879);
or U2243 (N_2243,N_1781,N_1910);
and U2244 (N_2244,N_1803,N_1833);
or U2245 (N_2245,N_1861,N_1862);
nand U2246 (N_2246,N_1955,N_1769);
and U2247 (N_2247,N_1763,N_1762);
nand U2248 (N_2248,N_1973,N_1986);
xnor U2249 (N_2249,N_1791,N_1844);
or U2250 (N_2250,N_2210,N_2051);
nor U2251 (N_2251,N_2037,N_2108);
and U2252 (N_2252,N_2234,N_2199);
nor U2253 (N_2253,N_2084,N_2160);
or U2254 (N_2254,N_2066,N_2131);
or U2255 (N_2255,N_2033,N_2224);
or U2256 (N_2256,N_2101,N_2045);
xor U2257 (N_2257,N_2161,N_2061);
and U2258 (N_2258,N_2163,N_2046);
xor U2259 (N_2259,N_2026,N_2188);
nor U2260 (N_2260,N_2135,N_2152);
and U2261 (N_2261,N_2057,N_2203);
nand U2262 (N_2262,N_2170,N_2103);
nor U2263 (N_2263,N_2179,N_2047);
nand U2264 (N_2264,N_2154,N_2235);
xor U2265 (N_2265,N_2071,N_2102);
nor U2266 (N_2266,N_2001,N_2124);
nand U2267 (N_2267,N_2090,N_2095);
xnor U2268 (N_2268,N_2132,N_2014);
or U2269 (N_2269,N_2139,N_2231);
xor U2270 (N_2270,N_2200,N_2127);
nor U2271 (N_2271,N_2216,N_2169);
nor U2272 (N_2272,N_2162,N_2120);
nor U2273 (N_2273,N_2064,N_2155);
xnor U2274 (N_2274,N_2085,N_2016);
or U2275 (N_2275,N_2219,N_2242);
nand U2276 (N_2276,N_2146,N_2073);
nor U2277 (N_2277,N_2144,N_2067);
nand U2278 (N_2278,N_2094,N_2214);
nor U2279 (N_2279,N_2236,N_2070);
nand U2280 (N_2280,N_2043,N_2012);
xnor U2281 (N_2281,N_2056,N_2195);
nor U2282 (N_2282,N_2083,N_2055);
and U2283 (N_2283,N_2075,N_2029);
and U2284 (N_2284,N_2137,N_2237);
xor U2285 (N_2285,N_2206,N_2157);
nor U2286 (N_2286,N_2228,N_2192);
nand U2287 (N_2287,N_2211,N_2181);
nor U2288 (N_2288,N_2226,N_2099);
xnor U2289 (N_2289,N_2038,N_2238);
and U2290 (N_2290,N_2180,N_2118);
xor U2291 (N_2291,N_2027,N_2150);
nor U2292 (N_2292,N_2246,N_2105);
or U2293 (N_2293,N_2044,N_2185);
and U2294 (N_2294,N_2054,N_2194);
and U2295 (N_2295,N_2184,N_2215);
and U2296 (N_2296,N_2092,N_2187);
and U2297 (N_2297,N_2111,N_2114);
nand U2298 (N_2298,N_2119,N_2109);
nand U2299 (N_2299,N_2138,N_2060);
and U2300 (N_2300,N_2177,N_2230);
or U2301 (N_2301,N_2244,N_2098);
or U2302 (N_2302,N_2130,N_2148);
and U2303 (N_2303,N_2158,N_2010);
nand U2304 (N_2304,N_2086,N_2225);
xor U2305 (N_2305,N_2196,N_2023);
or U2306 (N_2306,N_2233,N_2053);
xor U2307 (N_2307,N_2036,N_2243);
nand U2308 (N_2308,N_2201,N_2112);
or U2309 (N_2309,N_2204,N_2167);
nand U2310 (N_2310,N_2025,N_2168);
or U2311 (N_2311,N_2142,N_2147);
xor U2312 (N_2312,N_2091,N_2072);
nor U2313 (N_2313,N_2006,N_2207);
xor U2314 (N_2314,N_2197,N_2013);
nor U2315 (N_2315,N_2082,N_2175);
and U2316 (N_2316,N_2133,N_2129);
or U2317 (N_2317,N_2136,N_2209);
xor U2318 (N_2318,N_2165,N_2050);
nand U2319 (N_2319,N_2134,N_2208);
nand U2320 (N_2320,N_2110,N_2052);
and U2321 (N_2321,N_2116,N_2007);
nor U2322 (N_2322,N_2240,N_2032);
and U2323 (N_2323,N_2106,N_2193);
xnor U2324 (N_2324,N_2232,N_2122);
or U2325 (N_2325,N_2079,N_2113);
or U2326 (N_2326,N_2004,N_2097);
xor U2327 (N_2327,N_2081,N_2182);
xnor U2328 (N_2328,N_2034,N_2140);
xnor U2329 (N_2329,N_2176,N_2218);
and U2330 (N_2330,N_2076,N_2009);
nand U2331 (N_2331,N_2121,N_2049);
nor U2332 (N_2332,N_2178,N_2171);
and U2333 (N_2333,N_2048,N_2190);
and U2334 (N_2334,N_2117,N_2145);
and U2335 (N_2335,N_2149,N_2183);
nand U2336 (N_2336,N_2123,N_2000);
nor U2337 (N_2337,N_2035,N_2041);
nor U2338 (N_2338,N_2151,N_2068);
nor U2339 (N_2339,N_2141,N_2078);
and U2340 (N_2340,N_2126,N_2104);
nor U2341 (N_2341,N_2017,N_2005);
xor U2342 (N_2342,N_2011,N_2040);
or U2343 (N_2343,N_2059,N_2028);
or U2344 (N_2344,N_2241,N_2003);
and U2345 (N_2345,N_2173,N_2143);
or U2346 (N_2346,N_2227,N_2096);
nor U2347 (N_2347,N_2249,N_2223);
or U2348 (N_2348,N_2074,N_2062);
and U2349 (N_2349,N_2202,N_2008);
nor U2350 (N_2350,N_2015,N_2089);
nor U2351 (N_2351,N_2125,N_2205);
nor U2352 (N_2352,N_2217,N_2248);
xnor U2353 (N_2353,N_2022,N_2020);
xnor U2354 (N_2354,N_2063,N_2247);
nand U2355 (N_2355,N_2164,N_2002);
nand U2356 (N_2356,N_2128,N_2031);
and U2357 (N_2357,N_2222,N_2030);
nor U2358 (N_2358,N_2087,N_2174);
nand U2359 (N_2359,N_2100,N_2019);
nand U2360 (N_2360,N_2159,N_2080);
and U2361 (N_2361,N_2115,N_2239);
and U2362 (N_2362,N_2021,N_2213);
and U2363 (N_2363,N_2156,N_2191);
nor U2364 (N_2364,N_2189,N_2088);
xnor U2365 (N_2365,N_2065,N_2069);
xor U2366 (N_2366,N_2198,N_2212);
nor U2367 (N_2367,N_2042,N_2172);
nand U2368 (N_2368,N_2039,N_2186);
nor U2369 (N_2369,N_2245,N_2018);
nand U2370 (N_2370,N_2093,N_2058);
nor U2371 (N_2371,N_2220,N_2024);
nand U2372 (N_2372,N_2077,N_2166);
nand U2373 (N_2373,N_2153,N_2107);
and U2374 (N_2374,N_2221,N_2229);
nand U2375 (N_2375,N_2046,N_2224);
nor U2376 (N_2376,N_2058,N_2218);
nand U2377 (N_2377,N_2194,N_2080);
or U2378 (N_2378,N_2175,N_2193);
nand U2379 (N_2379,N_2230,N_2009);
or U2380 (N_2380,N_2229,N_2213);
or U2381 (N_2381,N_2085,N_2044);
nor U2382 (N_2382,N_2236,N_2079);
nor U2383 (N_2383,N_2013,N_2189);
nor U2384 (N_2384,N_2117,N_2096);
xor U2385 (N_2385,N_2120,N_2113);
and U2386 (N_2386,N_2160,N_2153);
and U2387 (N_2387,N_2083,N_2110);
or U2388 (N_2388,N_2138,N_2177);
and U2389 (N_2389,N_2055,N_2149);
or U2390 (N_2390,N_2004,N_2134);
nor U2391 (N_2391,N_2095,N_2185);
or U2392 (N_2392,N_2144,N_2065);
xor U2393 (N_2393,N_2069,N_2249);
and U2394 (N_2394,N_2135,N_2118);
nor U2395 (N_2395,N_2232,N_2115);
or U2396 (N_2396,N_2167,N_2129);
nor U2397 (N_2397,N_2189,N_2195);
nand U2398 (N_2398,N_2248,N_2235);
or U2399 (N_2399,N_2017,N_2201);
xor U2400 (N_2400,N_2077,N_2198);
nand U2401 (N_2401,N_2144,N_2049);
or U2402 (N_2402,N_2115,N_2005);
xor U2403 (N_2403,N_2108,N_2024);
or U2404 (N_2404,N_2237,N_2244);
or U2405 (N_2405,N_2168,N_2230);
xor U2406 (N_2406,N_2027,N_2026);
or U2407 (N_2407,N_2103,N_2019);
xor U2408 (N_2408,N_2110,N_2193);
nor U2409 (N_2409,N_2152,N_2064);
or U2410 (N_2410,N_2049,N_2076);
or U2411 (N_2411,N_2102,N_2021);
nor U2412 (N_2412,N_2172,N_2219);
nand U2413 (N_2413,N_2033,N_2092);
nand U2414 (N_2414,N_2230,N_2103);
nand U2415 (N_2415,N_2130,N_2020);
or U2416 (N_2416,N_2066,N_2175);
xor U2417 (N_2417,N_2209,N_2239);
nor U2418 (N_2418,N_2133,N_2176);
and U2419 (N_2419,N_2235,N_2160);
or U2420 (N_2420,N_2227,N_2234);
nor U2421 (N_2421,N_2226,N_2027);
nand U2422 (N_2422,N_2017,N_2062);
xnor U2423 (N_2423,N_2248,N_2156);
xor U2424 (N_2424,N_2217,N_2246);
and U2425 (N_2425,N_2227,N_2239);
or U2426 (N_2426,N_2025,N_2013);
and U2427 (N_2427,N_2037,N_2110);
or U2428 (N_2428,N_2011,N_2051);
nand U2429 (N_2429,N_2157,N_2247);
nor U2430 (N_2430,N_2012,N_2069);
xnor U2431 (N_2431,N_2171,N_2092);
xnor U2432 (N_2432,N_2105,N_2181);
nor U2433 (N_2433,N_2247,N_2242);
and U2434 (N_2434,N_2170,N_2094);
nand U2435 (N_2435,N_2228,N_2062);
or U2436 (N_2436,N_2115,N_2144);
nand U2437 (N_2437,N_2157,N_2080);
or U2438 (N_2438,N_2012,N_2034);
nor U2439 (N_2439,N_2079,N_2227);
and U2440 (N_2440,N_2184,N_2070);
nor U2441 (N_2441,N_2241,N_2236);
xor U2442 (N_2442,N_2114,N_2011);
nor U2443 (N_2443,N_2119,N_2194);
or U2444 (N_2444,N_2073,N_2052);
and U2445 (N_2445,N_2128,N_2127);
xor U2446 (N_2446,N_2060,N_2041);
or U2447 (N_2447,N_2065,N_2129);
and U2448 (N_2448,N_2000,N_2067);
and U2449 (N_2449,N_2083,N_2024);
nand U2450 (N_2450,N_2189,N_2012);
and U2451 (N_2451,N_2098,N_2073);
or U2452 (N_2452,N_2203,N_2129);
or U2453 (N_2453,N_2066,N_2112);
nor U2454 (N_2454,N_2192,N_2016);
and U2455 (N_2455,N_2042,N_2085);
and U2456 (N_2456,N_2146,N_2231);
nand U2457 (N_2457,N_2162,N_2174);
and U2458 (N_2458,N_2249,N_2045);
xor U2459 (N_2459,N_2001,N_2074);
and U2460 (N_2460,N_2172,N_2030);
xor U2461 (N_2461,N_2133,N_2222);
xnor U2462 (N_2462,N_2148,N_2021);
nand U2463 (N_2463,N_2198,N_2169);
and U2464 (N_2464,N_2055,N_2075);
xnor U2465 (N_2465,N_2152,N_2115);
and U2466 (N_2466,N_2052,N_2120);
nor U2467 (N_2467,N_2218,N_2106);
and U2468 (N_2468,N_2118,N_2083);
or U2469 (N_2469,N_2173,N_2185);
nor U2470 (N_2470,N_2207,N_2030);
nand U2471 (N_2471,N_2056,N_2128);
and U2472 (N_2472,N_2021,N_2052);
nor U2473 (N_2473,N_2154,N_2018);
nand U2474 (N_2474,N_2114,N_2080);
nor U2475 (N_2475,N_2059,N_2044);
nor U2476 (N_2476,N_2199,N_2024);
nand U2477 (N_2477,N_2101,N_2088);
and U2478 (N_2478,N_2139,N_2163);
nand U2479 (N_2479,N_2092,N_2190);
xnor U2480 (N_2480,N_2035,N_2173);
and U2481 (N_2481,N_2016,N_2149);
nor U2482 (N_2482,N_2214,N_2033);
nor U2483 (N_2483,N_2123,N_2087);
nand U2484 (N_2484,N_2174,N_2204);
nand U2485 (N_2485,N_2035,N_2121);
nand U2486 (N_2486,N_2015,N_2133);
and U2487 (N_2487,N_2182,N_2207);
nor U2488 (N_2488,N_2160,N_2180);
nor U2489 (N_2489,N_2176,N_2141);
nand U2490 (N_2490,N_2012,N_2066);
nand U2491 (N_2491,N_2209,N_2131);
and U2492 (N_2492,N_2074,N_2005);
nand U2493 (N_2493,N_2229,N_2171);
and U2494 (N_2494,N_2135,N_2050);
nand U2495 (N_2495,N_2224,N_2167);
xnor U2496 (N_2496,N_2227,N_2229);
nor U2497 (N_2497,N_2231,N_2172);
nand U2498 (N_2498,N_2029,N_2117);
nand U2499 (N_2499,N_2219,N_2218);
and U2500 (N_2500,N_2461,N_2492);
nand U2501 (N_2501,N_2337,N_2280);
and U2502 (N_2502,N_2316,N_2325);
nor U2503 (N_2503,N_2304,N_2297);
nand U2504 (N_2504,N_2386,N_2342);
xor U2505 (N_2505,N_2318,N_2407);
or U2506 (N_2506,N_2430,N_2414);
xor U2507 (N_2507,N_2479,N_2260);
xnor U2508 (N_2508,N_2463,N_2438);
nor U2509 (N_2509,N_2499,N_2268);
nor U2510 (N_2510,N_2370,N_2271);
xnor U2511 (N_2511,N_2364,N_2340);
and U2512 (N_2512,N_2313,N_2419);
or U2513 (N_2513,N_2397,N_2354);
xnor U2514 (N_2514,N_2376,N_2345);
xor U2515 (N_2515,N_2487,N_2338);
nor U2516 (N_2516,N_2323,N_2331);
nand U2517 (N_2517,N_2418,N_2333);
xor U2518 (N_2518,N_2305,N_2366);
nand U2519 (N_2519,N_2347,N_2399);
and U2520 (N_2520,N_2413,N_2393);
xor U2521 (N_2521,N_2263,N_2484);
or U2522 (N_2522,N_2285,N_2434);
xnor U2523 (N_2523,N_2468,N_2350);
xor U2524 (N_2524,N_2450,N_2277);
and U2525 (N_2525,N_2358,N_2469);
nor U2526 (N_2526,N_2289,N_2330);
or U2527 (N_2527,N_2357,N_2429);
nand U2528 (N_2528,N_2381,N_2483);
nand U2529 (N_2529,N_2497,N_2290);
xor U2530 (N_2530,N_2395,N_2267);
or U2531 (N_2531,N_2281,N_2328);
nand U2532 (N_2532,N_2329,N_2459);
nor U2533 (N_2533,N_2384,N_2346);
or U2534 (N_2534,N_2390,N_2261);
xor U2535 (N_2535,N_2435,N_2476);
or U2536 (N_2536,N_2437,N_2380);
or U2537 (N_2537,N_2389,N_2482);
and U2538 (N_2538,N_2415,N_2465);
nand U2539 (N_2539,N_2258,N_2440);
nor U2540 (N_2540,N_2439,N_2427);
nand U2541 (N_2541,N_2335,N_2428);
nor U2542 (N_2542,N_2455,N_2474);
or U2543 (N_2543,N_2443,N_2262);
or U2544 (N_2544,N_2276,N_2495);
xor U2545 (N_2545,N_2284,N_2489);
nand U2546 (N_2546,N_2367,N_2272);
or U2547 (N_2547,N_2256,N_2308);
xor U2548 (N_2548,N_2259,N_2255);
or U2549 (N_2549,N_2472,N_2447);
or U2550 (N_2550,N_2486,N_2360);
nor U2551 (N_2551,N_2475,N_2425);
nor U2552 (N_2552,N_2394,N_2311);
xnor U2553 (N_2553,N_2396,N_2303);
or U2554 (N_2554,N_2266,N_2403);
and U2555 (N_2555,N_2462,N_2453);
xor U2556 (N_2556,N_2250,N_2336);
or U2557 (N_2557,N_2377,N_2426);
nor U2558 (N_2558,N_2400,N_2321);
or U2559 (N_2559,N_2375,N_2398);
and U2560 (N_2560,N_2464,N_2362);
nand U2561 (N_2561,N_2471,N_2294);
nand U2562 (N_2562,N_2436,N_2298);
and U2563 (N_2563,N_2454,N_2320);
xnor U2564 (N_2564,N_2349,N_2273);
and U2565 (N_2565,N_2301,N_2287);
or U2566 (N_2566,N_2456,N_2490);
nand U2567 (N_2567,N_2296,N_2442);
or U2568 (N_2568,N_2401,N_2293);
and U2569 (N_2569,N_2352,N_2310);
or U2570 (N_2570,N_2449,N_2339);
xor U2571 (N_2571,N_2411,N_2373);
nand U2572 (N_2572,N_2312,N_2275);
nor U2573 (N_2573,N_2417,N_2319);
nand U2574 (N_2574,N_2446,N_2416);
nand U2575 (N_2575,N_2433,N_2452);
xnor U2576 (N_2576,N_2405,N_2374);
xor U2577 (N_2577,N_2404,N_2420);
xnor U2578 (N_2578,N_2302,N_2361);
nand U2579 (N_2579,N_2291,N_2444);
or U2580 (N_2580,N_2286,N_2431);
and U2581 (N_2581,N_2481,N_2314);
nor U2582 (N_2582,N_2441,N_2423);
and U2583 (N_2583,N_2251,N_2382);
nor U2584 (N_2584,N_2283,N_2480);
xnor U2585 (N_2585,N_2460,N_2363);
or U2586 (N_2586,N_2478,N_2493);
or U2587 (N_2587,N_2424,N_2343);
nor U2588 (N_2588,N_2445,N_2356);
or U2589 (N_2589,N_2332,N_2409);
and U2590 (N_2590,N_2326,N_2494);
nand U2591 (N_2591,N_2451,N_2369);
xnor U2592 (N_2592,N_2278,N_2353);
nand U2593 (N_2593,N_2300,N_2288);
nor U2594 (N_2594,N_2448,N_2269);
and U2595 (N_2595,N_2412,N_2334);
xor U2596 (N_2596,N_2477,N_2327);
nor U2597 (N_2597,N_2351,N_2292);
nor U2598 (N_2598,N_2299,N_2378);
nand U2599 (N_2599,N_2348,N_2470);
and U2600 (N_2600,N_2406,N_2315);
or U2601 (N_2601,N_2322,N_2392);
and U2602 (N_2602,N_2391,N_2496);
nor U2603 (N_2603,N_2421,N_2307);
and U2604 (N_2604,N_2274,N_2402);
xnor U2605 (N_2605,N_2295,N_2408);
and U2606 (N_2606,N_2355,N_2368);
nand U2607 (N_2607,N_2254,N_2488);
or U2608 (N_2608,N_2279,N_2270);
nor U2609 (N_2609,N_2252,N_2344);
or U2610 (N_2610,N_2458,N_2264);
and U2611 (N_2611,N_2467,N_2422);
and U2612 (N_2612,N_2317,N_2341);
and U2613 (N_2613,N_2485,N_2387);
nor U2614 (N_2614,N_2371,N_2498);
nor U2615 (N_2615,N_2306,N_2253);
xnor U2616 (N_2616,N_2379,N_2257);
or U2617 (N_2617,N_2410,N_2473);
xnor U2618 (N_2618,N_2383,N_2359);
or U2619 (N_2619,N_2372,N_2265);
and U2620 (N_2620,N_2385,N_2365);
or U2621 (N_2621,N_2324,N_2309);
nand U2622 (N_2622,N_2388,N_2466);
nand U2623 (N_2623,N_2491,N_2457);
and U2624 (N_2624,N_2282,N_2432);
nor U2625 (N_2625,N_2414,N_2345);
xnor U2626 (N_2626,N_2366,N_2431);
or U2627 (N_2627,N_2403,N_2413);
xor U2628 (N_2628,N_2457,N_2424);
or U2629 (N_2629,N_2295,N_2453);
nor U2630 (N_2630,N_2448,N_2439);
and U2631 (N_2631,N_2381,N_2336);
or U2632 (N_2632,N_2341,N_2461);
xnor U2633 (N_2633,N_2469,N_2277);
or U2634 (N_2634,N_2296,N_2330);
nand U2635 (N_2635,N_2449,N_2350);
and U2636 (N_2636,N_2400,N_2367);
and U2637 (N_2637,N_2384,N_2413);
xor U2638 (N_2638,N_2396,N_2314);
xnor U2639 (N_2639,N_2456,N_2432);
nor U2640 (N_2640,N_2489,N_2482);
nor U2641 (N_2641,N_2472,N_2250);
nor U2642 (N_2642,N_2259,N_2334);
or U2643 (N_2643,N_2335,N_2346);
or U2644 (N_2644,N_2338,N_2309);
nor U2645 (N_2645,N_2433,N_2412);
xnor U2646 (N_2646,N_2495,N_2280);
nand U2647 (N_2647,N_2374,N_2274);
nand U2648 (N_2648,N_2478,N_2442);
and U2649 (N_2649,N_2274,N_2293);
or U2650 (N_2650,N_2296,N_2481);
nor U2651 (N_2651,N_2485,N_2322);
nand U2652 (N_2652,N_2455,N_2497);
xnor U2653 (N_2653,N_2498,N_2478);
or U2654 (N_2654,N_2371,N_2334);
xor U2655 (N_2655,N_2294,N_2410);
xor U2656 (N_2656,N_2283,N_2394);
nand U2657 (N_2657,N_2325,N_2296);
xnor U2658 (N_2658,N_2263,N_2476);
or U2659 (N_2659,N_2413,N_2498);
or U2660 (N_2660,N_2417,N_2290);
xnor U2661 (N_2661,N_2475,N_2490);
xnor U2662 (N_2662,N_2387,N_2444);
or U2663 (N_2663,N_2390,N_2334);
or U2664 (N_2664,N_2401,N_2265);
xnor U2665 (N_2665,N_2443,N_2307);
or U2666 (N_2666,N_2491,N_2349);
and U2667 (N_2667,N_2267,N_2251);
or U2668 (N_2668,N_2395,N_2285);
or U2669 (N_2669,N_2369,N_2359);
nand U2670 (N_2670,N_2309,N_2473);
or U2671 (N_2671,N_2479,N_2452);
xnor U2672 (N_2672,N_2440,N_2393);
and U2673 (N_2673,N_2297,N_2429);
nor U2674 (N_2674,N_2261,N_2329);
nor U2675 (N_2675,N_2431,N_2415);
or U2676 (N_2676,N_2429,N_2471);
or U2677 (N_2677,N_2400,N_2498);
nor U2678 (N_2678,N_2343,N_2456);
nor U2679 (N_2679,N_2385,N_2495);
xor U2680 (N_2680,N_2277,N_2302);
nor U2681 (N_2681,N_2396,N_2452);
and U2682 (N_2682,N_2493,N_2336);
and U2683 (N_2683,N_2496,N_2354);
or U2684 (N_2684,N_2387,N_2406);
or U2685 (N_2685,N_2377,N_2423);
nand U2686 (N_2686,N_2325,N_2343);
or U2687 (N_2687,N_2381,N_2375);
nand U2688 (N_2688,N_2473,N_2374);
or U2689 (N_2689,N_2293,N_2406);
and U2690 (N_2690,N_2380,N_2263);
and U2691 (N_2691,N_2316,N_2332);
xor U2692 (N_2692,N_2484,N_2482);
nor U2693 (N_2693,N_2296,N_2444);
or U2694 (N_2694,N_2497,N_2382);
nand U2695 (N_2695,N_2307,N_2260);
and U2696 (N_2696,N_2417,N_2351);
and U2697 (N_2697,N_2485,N_2486);
or U2698 (N_2698,N_2262,N_2380);
or U2699 (N_2699,N_2337,N_2372);
xor U2700 (N_2700,N_2451,N_2353);
xnor U2701 (N_2701,N_2482,N_2289);
or U2702 (N_2702,N_2448,N_2340);
or U2703 (N_2703,N_2277,N_2299);
nand U2704 (N_2704,N_2300,N_2409);
and U2705 (N_2705,N_2480,N_2353);
xor U2706 (N_2706,N_2373,N_2394);
xor U2707 (N_2707,N_2491,N_2264);
and U2708 (N_2708,N_2426,N_2466);
xnor U2709 (N_2709,N_2373,N_2495);
nand U2710 (N_2710,N_2323,N_2282);
nand U2711 (N_2711,N_2471,N_2308);
xnor U2712 (N_2712,N_2361,N_2480);
and U2713 (N_2713,N_2322,N_2453);
nand U2714 (N_2714,N_2265,N_2479);
and U2715 (N_2715,N_2313,N_2468);
nor U2716 (N_2716,N_2425,N_2494);
and U2717 (N_2717,N_2348,N_2341);
and U2718 (N_2718,N_2254,N_2454);
nand U2719 (N_2719,N_2350,N_2464);
or U2720 (N_2720,N_2451,N_2467);
xor U2721 (N_2721,N_2290,N_2419);
or U2722 (N_2722,N_2407,N_2468);
and U2723 (N_2723,N_2419,N_2434);
and U2724 (N_2724,N_2288,N_2340);
or U2725 (N_2725,N_2412,N_2406);
or U2726 (N_2726,N_2486,N_2299);
and U2727 (N_2727,N_2333,N_2354);
nor U2728 (N_2728,N_2304,N_2411);
xor U2729 (N_2729,N_2430,N_2464);
nor U2730 (N_2730,N_2361,N_2307);
nand U2731 (N_2731,N_2496,N_2278);
and U2732 (N_2732,N_2317,N_2303);
nor U2733 (N_2733,N_2374,N_2399);
nand U2734 (N_2734,N_2426,N_2385);
or U2735 (N_2735,N_2284,N_2288);
or U2736 (N_2736,N_2393,N_2448);
xnor U2737 (N_2737,N_2367,N_2297);
nor U2738 (N_2738,N_2496,N_2285);
and U2739 (N_2739,N_2437,N_2300);
xnor U2740 (N_2740,N_2316,N_2295);
or U2741 (N_2741,N_2387,N_2329);
and U2742 (N_2742,N_2397,N_2468);
nor U2743 (N_2743,N_2425,N_2451);
nor U2744 (N_2744,N_2387,N_2466);
or U2745 (N_2745,N_2283,N_2426);
xor U2746 (N_2746,N_2344,N_2337);
nor U2747 (N_2747,N_2464,N_2361);
nand U2748 (N_2748,N_2377,N_2321);
nand U2749 (N_2749,N_2346,N_2487);
or U2750 (N_2750,N_2725,N_2737);
nor U2751 (N_2751,N_2646,N_2558);
and U2752 (N_2752,N_2667,N_2680);
or U2753 (N_2753,N_2615,N_2693);
or U2754 (N_2754,N_2559,N_2566);
and U2755 (N_2755,N_2735,N_2729);
or U2756 (N_2756,N_2565,N_2658);
nor U2757 (N_2757,N_2652,N_2673);
or U2758 (N_2758,N_2719,N_2604);
nor U2759 (N_2759,N_2746,N_2718);
nor U2760 (N_2760,N_2589,N_2659);
nand U2761 (N_2761,N_2630,N_2510);
or U2762 (N_2762,N_2650,N_2583);
xor U2763 (N_2763,N_2522,N_2526);
nand U2764 (N_2764,N_2597,N_2561);
nor U2765 (N_2765,N_2520,N_2633);
and U2766 (N_2766,N_2519,N_2517);
or U2767 (N_2767,N_2696,N_2608);
xor U2768 (N_2768,N_2654,N_2628);
xnor U2769 (N_2769,N_2582,N_2535);
or U2770 (N_2770,N_2656,N_2541);
nand U2771 (N_2771,N_2500,N_2647);
xor U2772 (N_2772,N_2699,N_2689);
and U2773 (N_2773,N_2660,N_2592);
and U2774 (N_2774,N_2664,N_2730);
nand U2775 (N_2775,N_2570,N_2532);
nand U2776 (N_2776,N_2666,N_2528);
nand U2777 (N_2777,N_2578,N_2703);
or U2778 (N_2778,N_2545,N_2739);
nand U2779 (N_2779,N_2555,N_2643);
and U2780 (N_2780,N_2724,N_2749);
and U2781 (N_2781,N_2648,N_2713);
xor U2782 (N_2782,N_2537,N_2672);
nor U2783 (N_2783,N_2540,N_2538);
xnor U2784 (N_2784,N_2549,N_2586);
nor U2785 (N_2785,N_2716,N_2641);
and U2786 (N_2786,N_2695,N_2547);
nand U2787 (N_2787,N_2553,N_2694);
or U2788 (N_2788,N_2710,N_2601);
xor U2789 (N_2789,N_2571,N_2590);
nand U2790 (N_2790,N_2536,N_2705);
or U2791 (N_2791,N_2539,N_2620);
xor U2792 (N_2792,N_2594,N_2697);
or U2793 (N_2793,N_2550,N_2613);
or U2794 (N_2794,N_2564,N_2611);
nand U2795 (N_2795,N_2744,N_2501);
nand U2796 (N_2796,N_2677,N_2584);
and U2797 (N_2797,N_2707,N_2577);
or U2798 (N_2798,N_2605,N_2568);
and U2799 (N_2799,N_2627,N_2513);
xor U2800 (N_2800,N_2554,N_2657);
xor U2801 (N_2801,N_2642,N_2665);
nand U2802 (N_2802,N_2684,N_2567);
or U2803 (N_2803,N_2552,N_2534);
xor U2804 (N_2804,N_2669,N_2575);
or U2805 (N_2805,N_2653,N_2511);
and U2806 (N_2806,N_2527,N_2557);
nor U2807 (N_2807,N_2624,N_2506);
or U2808 (N_2808,N_2728,N_2626);
xor U2809 (N_2809,N_2533,N_2629);
nor U2810 (N_2810,N_2574,N_2742);
xor U2811 (N_2811,N_2674,N_2682);
nand U2812 (N_2812,N_2748,N_2731);
or U2813 (N_2813,N_2637,N_2610);
and U2814 (N_2814,N_2727,N_2720);
or U2815 (N_2815,N_2717,N_2544);
and U2816 (N_2816,N_2618,N_2638);
or U2817 (N_2817,N_2560,N_2607);
or U2818 (N_2818,N_2521,N_2688);
and U2819 (N_2819,N_2747,N_2603);
and U2820 (N_2820,N_2745,N_2702);
or U2821 (N_2821,N_2606,N_2736);
and U2822 (N_2822,N_2675,N_2640);
nand U2823 (N_2823,N_2609,N_2681);
xor U2824 (N_2824,N_2639,N_2644);
nor U2825 (N_2825,N_2556,N_2580);
nand U2826 (N_2826,N_2595,N_2734);
nand U2827 (N_2827,N_2531,N_2635);
nor U2828 (N_2828,N_2581,N_2712);
or U2829 (N_2829,N_2631,N_2542);
or U2830 (N_2830,N_2701,N_2546);
or U2831 (N_2831,N_2598,N_2525);
nor U2832 (N_2832,N_2503,N_2562);
nand U2833 (N_2833,N_2543,N_2508);
nor U2834 (N_2834,N_2679,N_2661);
or U2835 (N_2835,N_2516,N_2706);
and U2836 (N_2836,N_2723,N_2588);
nor U2837 (N_2837,N_2708,N_2502);
xnor U2838 (N_2838,N_2504,N_2722);
nand U2839 (N_2839,N_2569,N_2683);
nand U2840 (N_2840,N_2671,N_2600);
xnor U2841 (N_2841,N_2616,N_2632);
or U2842 (N_2842,N_2548,N_2617);
xnor U2843 (N_2843,N_2602,N_2507);
nor U2844 (N_2844,N_2738,N_2523);
xnor U2845 (N_2845,N_2515,N_2663);
and U2846 (N_2846,N_2576,N_2691);
xnor U2847 (N_2847,N_2714,N_2668);
and U2848 (N_2848,N_2692,N_2678);
xnor U2849 (N_2849,N_2625,N_2614);
nand U2850 (N_2850,N_2529,N_2709);
and U2851 (N_2851,N_2741,N_2686);
nand U2852 (N_2852,N_2573,N_2670);
xnor U2853 (N_2853,N_2698,N_2524);
nor U2854 (N_2854,N_2645,N_2662);
and U2855 (N_2855,N_2530,N_2587);
xor U2856 (N_2856,N_2711,N_2721);
nand U2857 (N_2857,N_2551,N_2649);
and U2858 (N_2858,N_2505,N_2512);
xnor U2859 (N_2859,N_2740,N_2518);
and U2860 (N_2860,N_2599,N_2655);
nor U2861 (N_2861,N_2676,N_2572);
or U2862 (N_2862,N_2619,N_2636);
nor U2863 (N_2863,N_2596,N_2715);
or U2864 (N_2864,N_2726,N_2563);
nor U2865 (N_2865,N_2687,N_2579);
xnor U2866 (N_2866,N_2634,N_2612);
and U2867 (N_2867,N_2743,N_2622);
nor U2868 (N_2868,N_2509,N_2651);
or U2869 (N_2869,N_2732,N_2585);
nand U2870 (N_2870,N_2685,N_2733);
or U2871 (N_2871,N_2593,N_2621);
and U2872 (N_2872,N_2704,N_2514);
nor U2873 (N_2873,N_2690,N_2700);
xnor U2874 (N_2874,N_2591,N_2623);
nor U2875 (N_2875,N_2671,N_2720);
nor U2876 (N_2876,N_2546,N_2698);
xor U2877 (N_2877,N_2610,N_2535);
nor U2878 (N_2878,N_2690,N_2667);
or U2879 (N_2879,N_2706,N_2564);
and U2880 (N_2880,N_2689,N_2561);
xor U2881 (N_2881,N_2747,N_2598);
nand U2882 (N_2882,N_2688,N_2646);
xnor U2883 (N_2883,N_2603,N_2507);
nor U2884 (N_2884,N_2657,N_2603);
nand U2885 (N_2885,N_2600,N_2617);
and U2886 (N_2886,N_2679,N_2630);
nand U2887 (N_2887,N_2508,N_2717);
or U2888 (N_2888,N_2654,N_2524);
and U2889 (N_2889,N_2657,N_2615);
nor U2890 (N_2890,N_2573,N_2593);
nand U2891 (N_2891,N_2607,N_2549);
and U2892 (N_2892,N_2571,N_2561);
nand U2893 (N_2893,N_2690,N_2675);
and U2894 (N_2894,N_2679,N_2722);
or U2895 (N_2895,N_2625,N_2518);
xnor U2896 (N_2896,N_2621,N_2651);
nand U2897 (N_2897,N_2719,N_2525);
or U2898 (N_2898,N_2630,N_2597);
nor U2899 (N_2899,N_2528,N_2698);
xor U2900 (N_2900,N_2670,N_2649);
xnor U2901 (N_2901,N_2708,N_2734);
nand U2902 (N_2902,N_2728,N_2647);
nand U2903 (N_2903,N_2688,N_2725);
and U2904 (N_2904,N_2646,N_2674);
nand U2905 (N_2905,N_2719,N_2648);
xnor U2906 (N_2906,N_2677,N_2542);
xnor U2907 (N_2907,N_2723,N_2710);
nor U2908 (N_2908,N_2512,N_2664);
or U2909 (N_2909,N_2552,N_2617);
xor U2910 (N_2910,N_2506,N_2628);
xnor U2911 (N_2911,N_2681,N_2674);
or U2912 (N_2912,N_2564,N_2738);
or U2913 (N_2913,N_2640,N_2631);
nor U2914 (N_2914,N_2670,N_2507);
nor U2915 (N_2915,N_2559,N_2672);
nor U2916 (N_2916,N_2500,N_2639);
or U2917 (N_2917,N_2669,N_2626);
xor U2918 (N_2918,N_2671,N_2645);
nor U2919 (N_2919,N_2700,N_2745);
or U2920 (N_2920,N_2674,N_2624);
and U2921 (N_2921,N_2676,N_2721);
and U2922 (N_2922,N_2630,N_2544);
nor U2923 (N_2923,N_2533,N_2692);
nor U2924 (N_2924,N_2545,N_2649);
xnor U2925 (N_2925,N_2610,N_2620);
or U2926 (N_2926,N_2709,N_2639);
nor U2927 (N_2927,N_2554,N_2655);
and U2928 (N_2928,N_2673,N_2747);
nor U2929 (N_2929,N_2598,N_2696);
nand U2930 (N_2930,N_2724,N_2685);
or U2931 (N_2931,N_2641,N_2690);
nand U2932 (N_2932,N_2669,N_2625);
and U2933 (N_2933,N_2735,N_2669);
xor U2934 (N_2934,N_2646,N_2719);
and U2935 (N_2935,N_2539,N_2704);
nand U2936 (N_2936,N_2517,N_2595);
and U2937 (N_2937,N_2663,N_2574);
nor U2938 (N_2938,N_2633,N_2559);
or U2939 (N_2939,N_2602,N_2749);
and U2940 (N_2940,N_2502,N_2682);
and U2941 (N_2941,N_2581,N_2666);
or U2942 (N_2942,N_2665,N_2520);
nor U2943 (N_2943,N_2570,N_2510);
nor U2944 (N_2944,N_2624,N_2501);
and U2945 (N_2945,N_2652,N_2711);
nand U2946 (N_2946,N_2723,N_2546);
nor U2947 (N_2947,N_2706,N_2674);
and U2948 (N_2948,N_2636,N_2736);
and U2949 (N_2949,N_2628,N_2732);
nor U2950 (N_2950,N_2598,N_2679);
or U2951 (N_2951,N_2748,N_2596);
nand U2952 (N_2952,N_2570,N_2723);
or U2953 (N_2953,N_2688,N_2644);
nor U2954 (N_2954,N_2516,N_2530);
or U2955 (N_2955,N_2646,N_2607);
or U2956 (N_2956,N_2590,N_2632);
nor U2957 (N_2957,N_2742,N_2730);
xnor U2958 (N_2958,N_2579,N_2635);
nand U2959 (N_2959,N_2501,N_2530);
and U2960 (N_2960,N_2531,N_2693);
xnor U2961 (N_2961,N_2553,N_2558);
nor U2962 (N_2962,N_2686,N_2625);
nand U2963 (N_2963,N_2643,N_2743);
and U2964 (N_2964,N_2558,N_2541);
xnor U2965 (N_2965,N_2690,N_2591);
nor U2966 (N_2966,N_2504,N_2634);
and U2967 (N_2967,N_2560,N_2684);
or U2968 (N_2968,N_2578,N_2716);
or U2969 (N_2969,N_2690,N_2523);
nor U2970 (N_2970,N_2535,N_2596);
nand U2971 (N_2971,N_2749,N_2673);
and U2972 (N_2972,N_2516,N_2695);
or U2973 (N_2973,N_2681,N_2749);
xnor U2974 (N_2974,N_2516,N_2548);
xnor U2975 (N_2975,N_2535,N_2747);
nor U2976 (N_2976,N_2625,N_2667);
nand U2977 (N_2977,N_2635,N_2570);
nand U2978 (N_2978,N_2592,N_2707);
or U2979 (N_2979,N_2526,N_2747);
and U2980 (N_2980,N_2713,N_2613);
nor U2981 (N_2981,N_2578,N_2609);
or U2982 (N_2982,N_2538,N_2524);
nand U2983 (N_2983,N_2695,N_2624);
and U2984 (N_2984,N_2661,N_2502);
or U2985 (N_2985,N_2635,N_2518);
and U2986 (N_2986,N_2680,N_2560);
nor U2987 (N_2987,N_2561,N_2542);
or U2988 (N_2988,N_2549,N_2712);
nor U2989 (N_2989,N_2739,N_2504);
nor U2990 (N_2990,N_2700,N_2554);
nor U2991 (N_2991,N_2705,N_2563);
or U2992 (N_2992,N_2527,N_2506);
nor U2993 (N_2993,N_2721,N_2658);
or U2994 (N_2994,N_2536,N_2558);
nand U2995 (N_2995,N_2566,N_2663);
nor U2996 (N_2996,N_2600,N_2638);
nand U2997 (N_2997,N_2748,N_2572);
or U2998 (N_2998,N_2622,N_2502);
or U2999 (N_2999,N_2660,N_2504);
or U3000 (N_3000,N_2864,N_2952);
or U3001 (N_3001,N_2910,N_2931);
xnor U3002 (N_3002,N_2989,N_2858);
and U3003 (N_3003,N_2774,N_2871);
nand U3004 (N_3004,N_2885,N_2894);
nor U3005 (N_3005,N_2821,N_2769);
nand U3006 (N_3006,N_2817,N_2980);
or U3007 (N_3007,N_2761,N_2920);
nor U3008 (N_3008,N_2843,N_2969);
nor U3009 (N_3009,N_2831,N_2791);
and U3010 (N_3010,N_2878,N_2919);
or U3011 (N_3011,N_2766,N_2890);
nor U3012 (N_3012,N_2900,N_2868);
or U3013 (N_3013,N_2923,N_2767);
and U3014 (N_3014,N_2782,N_2916);
nor U3015 (N_3015,N_2880,N_2865);
or U3016 (N_3016,N_2903,N_2771);
xnor U3017 (N_3017,N_2962,N_2902);
nand U3018 (N_3018,N_2828,N_2854);
xor U3019 (N_3019,N_2979,N_2976);
xor U3020 (N_3020,N_2847,N_2863);
nor U3021 (N_3021,N_2837,N_2841);
or U3022 (N_3022,N_2888,N_2783);
or U3023 (N_3023,N_2895,N_2812);
nand U3024 (N_3024,N_2948,N_2951);
or U3025 (N_3025,N_2772,N_2794);
and U3026 (N_3026,N_2852,N_2891);
and U3027 (N_3027,N_2950,N_2877);
nand U3028 (N_3028,N_2855,N_2915);
or U3029 (N_3029,N_2781,N_2998);
nand U3030 (N_3030,N_2760,N_2874);
nand U3031 (N_3031,N_2779,N_2941);
nor U3032 (N_3032,N_2896,N_2913);
or U3033 (N_3033,N_2964,N_2882);
nor U3034 (N_3034,N_2924,N_2929);
xnor U3035 (N_3035,N_2972,N_2912);
xnor U3036 (N_3036,N_2974,N_2961);
xnor U3037 (N_3037,N_2869,N_2893);
and U3038 (N_3038,N_2884,N_2826);
or U3039 (N_3039,N_2862,N_2849);
or U3040 (N_3040,N_2856,N_2938);
nand U3041 (N_3041,N_2802,N_2773);
and U3042 (N_3042,N_2955,N_2925);
or U3043 (N_3043,N_2993,N_2755);
or U3044 (N_3044,N_2759,N_2887);
nor U3045 (N_3045,N_2906,N_2753);
nand U3046 (N_3046,N_2844,N_2751);
nand U3047 (N_3047,N_2807,N_2795);
and U3048 (N_3048,N_2822,N_2968);
or U3049 (N_3049,N_2987,N_2805);
xor U3050 (N_3050,N_2940,N_2965);
nor U3051 (N_3051,N_2909,N_2872);
and U3052 (N_3052,N_2978,N_2997);
and U3053 (N_3053,N_2918,N_2780);
and U3054 (N_3054,N_2975,N_2823);
or U3055 (N_3055,N_2834,N_2765);
xnor U3056 (N_3056,N_2889,N_2928);
nor U3057 (N_3057,N_2934,N_2776);
xnor U3058 (N_3058,N_2775,N_2992);
or U3059 (N_3059,N_2984,N_2908);
or U3060 (N_3060,N_2901,N_2846);
nand U3061 (N_3061,N_2991,N_2827);
nor U3062 (N_3062,N_2792,N_2947);
nand U3063 (N_3063,N_2957,N_2801);
and U3064 (N_3064,N_2944,N_2754);
nand U3065 (N_3065,N_2879,N_2939);
nand U3066 (N_3066,N_2845,N_2914);
or U3067 (N_3067,N_2756,N_2803);
xor U3068 (N_3068,N_2777,N_2936);
or U3069 (N_3069,N_2994,N_2830);
or U3070 (N_3070,N_2922,N_2850);
or U3071 (N_3071,N_2857,N_2829);
xnor U3072 (N_3072,N_2866,N_2860);
xor U3073 (N_3073,N_2876,N_2945);
and U3074 (N_3074,N_2764,N_2935);
nand U3075 (N_3075,N_2977,N_2832);
nor U3076 (N_3076,N_2995,N_2971);
or U3077 (N_3077,N_2806,N_2959);
nand U3078 (N_3078,N_2785,N_2799);
xor U3079 (N_3079,N_2768,N_2953);
nor U3080 (N_3080,N_2946,N_2958);
xor U3081 (N_3081,N_2808,N_2796);
nor U3082 (N_3082,N_2937,N_2790);
or U3083 (N_3083,N_2851,N_2824);
nor U3084 (N_3084,N_2983,N_2836);
xnor U3085 (N_3085,N_2839,N_2750);
or U3086 (N_3086,N_2942,N_2907);
and U3087 (N_3087,N_2981,N_2752);
and U3088 (N_3088,N_2949,N_2873);
xnor U3089 (N_3089,N_2954,N_2818);
nor U3090 (N_3090,N_2786,N_2911);
or U3091 (N_3091,N_2933,N_2897);
nand U3092 (N_3092,N_2886,N_2820);
nor U3093 (N_3093,N_2905,N_2838);
or U3094 (N_3094,N_2809,N_2917);
and U3095 (N_3095,N_2784,N_2793);
and U3096 (N_3096,N_2788,N_2800);
or U3097 (N_3097,N_2932,N_2787);
nand U3098 (N_3098,N_2970,N_2899);
or U3099 (N_3099,N_2757,N_2892);
xnor U3100 (N_3100,N_2921,N_2778);
xor U3101 (N_3101,N_2999,N_2835);
nor U3102 (N_3102,N_2943,N_2811);
xor U3103 (N_3103,N_2813,N_2797);
nand U3104 (N_3104,N_2758,N_2926);
nand U3105 (N_3105,N_2762,N_2842);
and U3106 (N_3106,N_2982,N_2815);
nor U3107 (N_3107,N_2985,N_2804);
or U3108 (N_3108,N_2881,N_2853);
nor U3109 (N_3109,N_2898,N_2840);
nor U3110 (N_3110,N_2927,N_2904);
xor U3111 (N_3111,N_2996,N_2798);
and U3112 (N_3112,N_2967,N_2960);
nand U3113 (N_3113,N_2966,N_2986);
nand U3114 (N_3114,N_2867,N_2833);
nand U3115 (N_3115,N_2810,N_2848);
nor U3116 (N_3116,N_2816,N_2990);
or U3117 (N_3117,N_2988,N_2861);
or U3118 (N_3118,N_2789,N_2770);
xor U3119 (N_3119,N_2870,N_2956);
and U3120 (N_3120,N_2973,N_2814);
nor U3121 (N_3121,N_2763,N_2963);
xor U3122 (N_3122,N_2875,N_2825);
xnor U3123 (N_3123,N_2883,N_2930);
or U3124 (N_3124,N_2859,N_2819);
xor U3125 (N_3125,N_2827,N_2882);
and U3126 (N_3126,N_2909,N_2838);
nand U3127 (N_3127,N_2852,N_2986);
and U3128 (N_3128,N_2946,N_2938);
nor U3129 (N_3129,N_2898,N_2886);
nor U3130 (N_3130,N_2787,N_2865);
nand U3131 (N_3131,N_2951,N_2845);
or U3132 (N_3132,N_2802,N_2975);
nor U3133 (N_3133,N_2837,N_2844);
or U3134 (N_3134,N_2898,N_2954);
or U3135 (N_3135,N_2979,N_2773);
nor U3136 (N_3136,N_2876,N_2821);
and U3137 (N_3137,N_2938,N_2806);
or U3138 (N_3138,N_2903,N_2884);
and U3139 (N_3139,N_2800,N_2907);
nand U3140 (N_3140,N_2956,N_2811);
xnor U3141 (N_3141,N_2887,N_2753);
nand U3142 (N_3142,N_2967,N_2892);
nand U3143 (N_3143,N_2975,N_2767);
nand U3144 (N_3144,N_2767,N_2795);
nand U3145 (N_3145,N_2907,N_2999);
nor U3146 (N_3146,N_2770,N_2818);
and U3147 (N_3147,N_2883,N_2802);
or U3148 (N_3148,N_2924,N_2753);
or U3149 (N_3149,N_2895,N_2921);
or U3150 (N_3150,N_2952,N_2849);
or U3151 (N_3151,N_2837,N_2981);
and U3152 (N_3152,N_2901,N_2800);
and U3153 (N_3153,N_2972,N_2889);
and U3154 (N_3154,N_2953,N_2990);
or U3155 (N_3155,N_2784,N_2755);
xnor U3156 (N_3156,N_2975,N_2769);
xnor U3157 (N_3157,N_2800,N_2751);
or U3158 (N_3158,N_2939,N_2752);
and U3159 (N_3159,N_2865,N_2899);
or U3160 (N_3160,N_2799,N_2806);
nor U3161 (N_3161,N_2835,N_2898);
xor U3162 (N_3162,N_2923,N_2761);
nand U3163 (N_3163,N_2858,N_2999);
or U3164 (N_3164,N_2840,N_2892);
or U3165 (N_3165,N_2870,N_2940);
nand U3166 (N_3166,N_2830,N_2821);
or U3167 (N_3167,N_2810,N_2816);
or U3168 (N_3168,N_2778,N_2822);
xor U3169 (N_3169,N_2957,N_2910);
nand U3170 (N_3170,N_2974,N_2907);
and U3171 (N_3171,N_2903,N_2956);
xnor U3172 (N_3172,N_2837,N_2927);
nor U3173 (N_3173,N_2899,N_2806);
or U3174 (N_3174,N_2907,N_2875);
or U3175 (N_3175,N_2888,N_2794);
and U3176 (N_3176,N_2787,N_2937);
xor U3177 (N_3177,N_2820,N_2866);
or U3178 (N_3178,N_2946,N_2869);
nand U3179 (N_3179,N_2971,N_2951);
nor U3180 (N_3180,N_2939,N_2819);
nor U3181 (N_3181,N_2824,N_2959);
xor U3182 (N_3182,N_2902,N_2869);
nand U3183 (N_3183,N_2865,N_2759);
nor U3184 (N_3184,N_2930,N_2858);
nor U3185 (N_3185,N_2833,N_2751);
xor U3186 (N_3186,N_2867,N_2804);
xor U3187 (N_3187,N_2929,N_2766);
nor U3188 (N_3188,N_2764,N_2769);
xor U3189 (N_3189,N_2912,N_2751);
or U3190 (N_3190,N_2979,N_2993);
nor U3191 (N_3191,N_2941,N_2963);
nand U3192 (N_3192,N_2804,N_2752);
and U3193 (N_3193,N_2862,N_2987);
and U3194 (N_3194,N_2917,N_2838);
nor U3195 (N_3195,N_2876,N_2844);
nand U3196 (N_3196,N_2825,N_2908);
and U3197 (N_3197,N_2944,N_2780);
xor U3198 (N_3198,N_2869,N_2774);
nand U3199 (N_3199,N_2768,N_2862);
nand U3200 (N_3200,N_2761,N_2839);
nand U3201 (N_3201,N_2784,N_2781);
nand U3202 (N_3202,N_2896,N_2758);
nand U3203 (N_3203,N_2909,N_2820);
xnor U3204 (N_3204,N_2905,N_2785);
nand U3205 (N_3205,N_2888,N_2927);
or U3206 (N_3206,N_2916,N_2877);
nand U3207 (N_3207,N_2900,N_2796);
xnor U3208 (N_3208,N_2975,N_2954);
nor U3209 (N_3209,N_2958,N_2954);
and U3210 (N_3210,N_2957,N_2917);
or U3211 (N_3211,N_2750,N_2930);
and U3212 (N_3212,N_2996,N_2938);
or U3213 (N_3213,N_2908,N_2928);
nand U3214 (N_3214,N_2842,N_2787);
xnor U3215 (N_3215,N_2950,N_2890);
or U3216 (N_3216,N_2780,N_2940);
nor U3217 (N_3217,N_2900,N_2947);
or U3218 (N_3218,N_2768,N_2811);
or U3219 (N_3219,N_2776,N_2769);
nor U3220 (N_3220,N_2810,N_2808);
or U3221 (N_3221,N_2894,N_2996);
and U3222 (N_3222,N_2895,N_2759);
xor U3223 (N_3223,N_2752,N_2763);
nor U3224 (N_3224,N_2963,N_2962);
and U3225 (N_3225,N_2757,N_2785);
nor U3226 (N_3226,N_2940,N_2803);
nor U3227 (N_3227,N_2785,N_2831);
nor U3228 (N_3228,N_2781,N_2803);
nand U3229 (N_3229,N_2889,N_2943);
xor U3230 (N_3230,N_2962,N_2978);
nor U3231 (N_3231,N_2829,N_2782);
or U3232 (N_3232,N_2907,N_2983);
or U3233 (N_3233,N_2864,N_2765);
or U3234 (N_3234,N_2893,N_2954);
and U3235 (N_3235,N_2963,N_2764);
and U3236 (N_3236,N_2971,N_2984);
nand U3237 (N_3237,N_2873,N_2921);
nor U3238 (N_3238,N_2799,N_2844);
nand U3239 (N_3239,N_2968,N_2871);
nor U3240 (N_3240,N_2892,N_2924);
xnor U3241 (N_3241,N_2847,N_2853);
or U3242 (N_3242,N_2896,N_2807);
and U3243 (N_3243,N_2806,N_2997);
xnor U3244 (N_3244,N_2786,N_2887);
xnor U3245 (N_3245,N_2835,N_2983);
xor U3246 (N_3246,N_2862,N_2878);
and U3247 (N_3247,N_2941,N_2899);
or U3248 (N_3248,N_2891,N_2887);
nand U3249 (N_3249,N_2785,N_2847);
nor U3250 (N_3250,N_3188,N_3233);
and U3251 (N_3251,N_3198,N_3076);
or U3252 (N_3252,N_3115,N_3124);
or U3253 (N_3253,N_3005,N_3003);
nand U3254 (N_3254,N_3236,N_3037);
and U3255 (N_3255,N_3052,N_3117);
nand U3256 (N_3256,N_3237,N_3174);
nor U3257 (N_3257,N_3066,N_3130);
nand U3258 (N_3258,N_3069,N_3009);
or U3259 (N_3259,N_3216,N_3012);
and U3260 (N_3260,N_3050,N_3245);
and U3261 (N_3261,N_3224,N_3008);
nor U3262 (N_3262,N_3205,N_3067);
xnor U3263 (N_3263,N_3144,N_3157);
nand U3264 (N_3264,N_3092,N_3112);
and U3265 (N_3265,N_3156,N_3019);
xor U3266 (N_3266,N_3183,N_3129);
and U3267 (N_3267,N_3047,N_3091);
or U3268 (N_3268,N_3154,N_3201);
nand U3269 (N_3269,N_3170,N_3192);
nor U3270 (N_3270,N_3095,N_3122);
xnor U3271 (N_3271,N_3014,N_3049);
nand U3272 (N_3272,N_3246,N_3006);
nand U3273 (N_3273,N_3149,N_3186);
and U3274 (N_3274,N_3102,N_3202);
nor U3275 (N_3275,N_3025,N_3203);
nor U3276 (N_3276,N_3045,N_3204);
nand U3277 (N_3277,N_3165,N_3247);
xnor U3278 (N_3278,N_3036,N_3041);
nand U3279 (N_3279,N_3029,N_3075);
xor U3280 (N_3280,N_3150,N_3086);
nand U3281 (N_3281,N_3125,N_3176);
or U3282 (N_3282,N_3042,N_3128);
nor U3283 (N_3283,N_3032,N_3051);
and U3284 (N_3284,N_3013,N_3134);
or U3285 (N_3285,N_3072,N_3127);
nor U3286 (N_3286,N_3242,N_3104);
and U3287 (N_3287,N_3038,N_3173);
nor U3288 (N_3288,N_3081,N_3161);
nand U3289 (N_3289,N_3147,N_3004);
or U3290 (N_3290,N_3145,N_3109);
nand U3291 (N_3291,N_3024,N_3087);
nand U3292 (N_3292,N_3189,N_3158);
nand U3293 (N_3293,N_3044,N_3133);
nor U3294 (N_3294,N_3151,N_3214);
nand U3295 (N_3295,N_3120,N_3230);
and U3296 (N_3296,N_3055,N_3022);
or U3297 (N_3297,N_3135,N_3167);
and U3298 (N_3298,N_3184,N_3221);
and U3299 (N_3299,N_3121,N_3043);
xnor U3300 (N_3300,N_3153,N_3116);
xor U3301 (N_3301,N_3046,N_3181);
nand U3302 (N_3302,N_3064,N_3061);
nand U3303 (N_3303,N_3199,N_3108);
or U3304 (N_3304,N_3168,N_3232);
xnor U3305 (N_3305,N_3023,N_3059);
or U3306 (N_3306,N_3088,N_3131);
nand U3307 (N_3307,N_3197,N_3175);
nor U3308 (N_3308,N_3090,N_3239);
or U3309 (N_3309,N_3039,N_3063);
nor U3310 (N_3310,N_3096,N_3136);
or U3311 (N_3311,N_3169,N_3082);
nor U3312 (N_3312,N_3099,N_3140);
or U3313 (N_3313,N_3021,N_3123);
and U3314 (N_3314,N_3240,N_3195);
nand U3315 (N_3315,N_3103,N_3077);
nor U3316 (N_3316,N_3097,N_3200);
xnor U3317 (N_3317,N_3190,N_3011);
xor U3318 (N_3318,N_3163,N_3015);
nand U3319 (N_3319,N_3060,N_3068);
xnor U3320 (N_3320,N_3000,N_3223);
and U3321 (N_3321,N_3016,N_3118);
and U3322 (N_3322,N_3146,N_3179);
and U3323 (N_3323,N_3018,N_3126);
nand U3324 (N_3324,N_3027,N_3178);
nor U3325 (N_3325,N_3152,N_3110);
and U3326 (N_3326,N_3079,N_3002);
xnor U3327 (N_3327,N_3074,N_3148);
nor U3328 (N_3328,N_3028,N_3248);
and U3329 (N_3329,N_3159,N_3107);
xnor U3330 (N_3330,N_3111,N_3155);
nor U3331 (N_3331,N_3139,N_3225);
xnor U3332 (N_3332,N_3211,N_3244);
or U3333 (N_3333,N_3114,N_3053);
xor U3334 (N_3334,N_3085,N_3058);
and U3335 (N_3335,N_3222,N_3007);
and U3336 (N_3336,N_3171,N_3185);
nand U3337 (N_3337,N_3071,N_3084);
xnor U3338 (N_3338,N_3057,N_3056);
nor U3339 (N_3339,N_3243,N_3017);
xnor U3340 (N_3340,N_3106,N_3166);
nand U3341 (N_3341,N_3217,N_3241);
xor U3342 (N_3342,N_3101,N_3209);
nor U3343 (N_3343,N_3048,N_3132);
and U3344 (N_3344,N_3080,N_3020);
nor U3345 (N_3345,N_3113,N_3034);
or U3346 (N_3346,N_3215,N_3070);
or U3347 (N_3347,N_3162,N_3073);
or U3348 (N_3348,N_3227,N_3083);
nor U3349 (N_3349,N_3119,N_3035);
xor U3350 (N_3350,N_3105,N_3226);
nand U3351 (N_3351,N_3031,N_3194);
or U3352 (N_3352,N_3098,N_3141);
xnor U3353 (N_3353,N_3177,N_3010);
xor U3354 (N_3354,N_3208,N_3182);
nor U3355 (N_3355,N_3193,N_3054);
and U3356 (N_3356,N_3218,N_3030);
xnor U3357 (N_3357,N_3219,N_3229);
and U3358 (N_3358,N_3228,N_3160);
nor U3359 (N_3359,N_3033,N_3094);
nor U3360 (N_3360,N_3206,N_3210);
nand U3361 (N_3361,N_3220,N_3093);
or U3362 (N_3362,N_3191,N_3164);
nor U3363 (N_3363,N_3065,N_3231);
nor U3364 (N_3364,N_3143,N_3040);
or U3365 (N_3365,N_3213,N_3172);
and U3366 (N_3366,N_3249,N_3187);
and U3367 (N_3367,N_3212,N_3196);
xnor U3368 (N_3368,N_3001,N_3089);
xor U3369 (N_3369,N_3137,N_3234);
xnor U3370 (N_3370,N_3180,N_3138);
nor U3371 (N_3371,N_3100,N_3142);
nor U3372 (N_3372,N_3026,N_3207);
nand U3373 (N_3373,N_3078,N_3238);
and U3374 (N_3374,N_3062,N_3235);
nand U3375 (N_3375,N_3025,N_3003);
nand U3376 (N_3376,N_3129,N_3072);
nand U3377 (N_3377,N_3232,N_3002);
xor U3378 (N_3378,N_3224,N_3217);
nand U3379 (N_3379,N_3058,N_3144);
nor U3380 (N_3380,N_3226,N_3191);
nor U3381 (N_3381,N_3161,N_3119);
nor U3382 (N_3382,N_3182,N_3159);
xor U3383 (N_3383,N_3192,N_3123);
nand U3384 (N_3384,N_3043,N_3042);
nand U3385 (N_3385,N_3153,N_3210);
xor U3386 (N_3386,N_3153,N_3183);
or U3387 (N_3387,N_3050,N_3004);
and U3388 (N_3388,N_3192,N_3186);
nand U3389 (N_3389,N_3225,N_3223);
or U3390 (N_3390,N_3029,N_3177);
nand U3391 (N_3391,N_3137,N_3249);
xnor U3392 (N_3392,N_3105,N_3215);
xnor U3393 (N_3393,N_3249,N_3100);
nand U3394 (N_3394,N_3220,N_3154);
xor U3395 (N_3395,N_3094,N_3066);
nand U3396 (N_3396,N_3066,N_3078);
nor U3397 (N_3397,N_3146,N_3024);
nor U3398 (N_3398,N_3154,N_3212);
nor U3399 (N_3399,N_3143,N_3190);
or U3400 (N_3400,N_3129,N_3101);
and U3401 (N_3401,N_3223,N_3058);
or U3402 (N_3402,N_3107,N_3100);
nand U3403 (N_3403,N_3015,N_3179);
xnor U3404 (N_3404,N_3201,N_3033);
nand U3405 (N_3405,N_3193,N_3021);
xnor U3406 (N_3406,N_3025,N_3218);
or U3407 (N_3407,N_3105,N_3197);
and U3408 (N_3408,N_3225,N_3076);
xor U3409 (N_3409,N_3241,N_3144);
xnor U3410 (N_3410,N_3178,N_3164);
or U3411 (N_3411,N_3142,N_3234);
nor U3412 (N_3412,N_3154,N_3012);
nor U3413 (N_3413,N_3150,N_3145);
xnor U3414 (N_3414,N_3204,N_3210);
nor U3415 (N_3415,N_3011,N_3128);
xnor U3416 (N_3416,N_3077,N_3045);
and U3417 (N_3417,N_3073,N_3044);
and U3418 (N_3418,N_3240,N_3001);
nor U3419 (N_3419,N_3100,N_3027);
nand U3420 (N_3420,N_3127,N_3168);
and U3421 (N_3421,N_3012,N_3099);
nor U3422 (N_3422,N_3028,N_3060);
nand U3423 (N_3423,N_3202,N_3002);
xnor U3424 (N_3424,N_3165,N_3220);
xnor U3425 (N_3425,N_3221,N_3063);
xor U3426 (N_3426,N_3243,N_3095);
or U3427 (N_3427,N_3019,N_3239);
xor U3428 (N_3428,N_3005,N_3007);
nor U3429 (N_3429,N_3023,N_3107);
or U3430 (N_3430,N_3228,N_3060);
nor U3431 (N_3431,N_3071,N_3125);
nor U3432 (N_3432,N_3012,N_3091);
xor U3433 (N_3433,N_3019,N_3035);
or U3434 (N_3434,N_3050,N_3088);
or U3435 (N_3435,N_3119,N_3078);
or U3436 (N_3436,N_3202,N_3103);
nor U3437 (N_3437,N_3046,N_3142);
xor U3438 (N_3438,N_3076,N_3183);
nand U3439 (N_3439,N_3116,N_3205);
xor U3440 (N_3440,N_3227,N_3058);
or U3441 (N_3441,N_3075,N_3091);
xnor U3442 (N_3442,N_3155,N_3006);
xnor U3443 (N_3443,N_3143,N_3012);
nand U3444 (N_3444,N_3216,N_3169);
nor U3445 (N_3445,N_3209,N_3231);
or U3446 (N_3446,N_3118,N_3060);
xor U3447 (N_3447,N_3174,N_3172);
and U3448 (N_3448,N_3175,N_3159);
nor U3449 (N_3449,N_3173,N_3166);
or U3450 (N_3450,N_3053,N_3234);
nand U3451 (N_3451,N_3108,N_3219);
or U3452 (N_3452,N_3145,N_3094);
or U3453 (N_3453,N_3042,N_3017);
xor U3454 (N_3454,N_3001,N_3138);
and U3455 (N_3455,N_3214,N_3226);
xor U3456 (N_3456,N_3223,N_3014);
nand U3457 (N_3457,N_3169,N_3119);
and U3458 (N_3458,N_3136,N_3083);
nand U3459 (N_3459,N_3145,N_3002);
and U3460 (N_3460,N_3083,N_3128);
nand U3461 (N_3461,N_3075,N_3198);
and U3462 (N_3462,N_3114,N_3183);
xor U3463 (N_3463,N_3128,N_3166);
or U3464 (N_3464,N_3207,N_3017);
xnor U3465 (N_3465,N_3175,N_3036);
nor U3466 (N_3466,N_3022,N_3094);
and U3467 (N_3467,N_3041,N_3203);
or U3468 (N_3468,N_3208,N_3144);
nor U3469 (N_3469,N_3110,N_3022);
nand U3470 (N_3470,N_3028,N_3023);
xor U3471 (N_3471,N_3170,N_3070);
or U3472 (N_3472,N_3083,N_3066);
or U3473 (N_3473,N_3107,N_3240);
xnor U3474 (N_3474,N_3034,N_3103);
or U3475 (N_3475,N_3030,N_3177);
xnor U3476 (N_3476,N_3218,N_3094);
or U3477 (N_3477,N_3023,N_3140);
xnor U3478 (N_3478,N_3149,N_3242);
xnor U3479 (N_3479,N_3029,N_3160);
and U3480 (N_3480,N_3029,N_3125);
xor U3481 (N_3481,N_3217,N_3165);
xnor U3482 (N_3482,N_3044,N_3147);
xor U3483 (N_3483,N_3185,N_3168);
or U3484 (N_3484,N_3215,N_3038);
nand U3485 (N_3485,N_3074,N_3032);
and U3486 (N_3486,N_3047,N_3192);
xor U3487 (N_3487,N_3209,N_3243);
nor U3488 (N_3488,N_3163,N_3239);
or U3489 (N_3489,N_3236,N_3206);
xor U3490 (N_3490,N_3194,N_3207);
and U3491 (N_3491,N_3164,N_3151);
and U3492 (N_3492,N_3130,N_3068);
or U3493 (N_3493,N_3067,N_3021);
nand U3494 (N_3494,N_3169,N_3019);
nor U3495 (N_3495,N_3130,N_3231);
or U3496 (N_3496,N_3027,N_3126);
or U3497 (N_3497,N_3143,N_3031);
or U3498 (N_3498,N_3238,N_3113);
or U3499 (N_3499,N_3119,N_3249);
xor U3500 (N_3500,N_3397,N_3408);
and U3501 (N_3501,N_3368,N_3470);
nor U3502 (N_3502,N_3262,N_3399);
xnor U3503 (N_3503,N_3425,N_3442);
nor U3504 (N_3504,N_3317,N_3440);
nor U3505 (N_3505,N_3272,N_3328);
and U3506 (N_3506,N_3324,N_3452);
and U3507 (N_3507,N_3251,N_3486);
xnor U3508 (N_3508,N_3257,N_3363);
nand U3509 (N_3509,N_3323,N_3358);
nor U3510 (N_3510,N_3403,N_3285);
nand U3511 (N_3511,N_3493,N_3499);
nor U3512 (N_3512,N_3299,N_3335);
or U3513 (N_3513,N_3436,N_3427);
xnor U3514 (N_3514,N_3406,N_3396);
and U3515 (N_3515,N_3401,N_3482);
xor U3516 (N_3516,N_3333,N_3441);
nor U3517 (N_3517,N_3289,N_3264);
or U3518 (N_3518,N_3355,N_3402);
or U3519 (N_3519,N_3428,N_3437);
xor U3520 (N_3520,N_3426,N_3495);
xor U3521 (N_3521,N_3250,N_3263);
or U3522 (N_3522,N_3458,N_3271);
xnor U3523 (N_3523,N_3438,N_3258);
nor U3524 (N_3524,N_3477,N_3287);
and U3525 (N_3525,N_3460,N_3383);
and U3526 (N_3526,N_3261,N_3356);
nor U3527 (N_3527,N_3412,N_3365);
or U3528 (N_3528,N_3471,N_3390);
xor U3529 (N_3529,N_3337,N_3453);
nor U3530 (N_3530,N_3419,N_3349);
nor U3531 (N_3531,N_3488,N_3445);
or U3532 (N_3532,N_3252,N_3463);
or U3533 (N_3533,N_3306,N_3353);
nor U3534 (N_3534,N_3344,N_3431);
nand U3535 (N_3535,N_3290,N_3494);
xor U3536 (N_3536,N_3283,N_3320);
and U3537 (N_3537,N_3280,N_3256);
or U3538 (N_3538,N_3322,N_3313);
and U3539 (N_3539,N_3366,N_3465);
nand U3540 (N_3540,N_3370,N_3449);
nand U3541 (N_3541,N_3475,N_3298);
nand U3542 (N_3542,N_3443,N_3255);
nor U3543 (N_3543,N_3297,N_3336);
and U3544 (N_3544,N_3469,N_3325);
xnor U3545 (N_3545,N_3367,N_3480);
xnor U3546 (N_3546,N_3373,N_3372);
and U3547 (N_3547,N_3421,N_3351);
nand U3548 (N_3548,N_3318,N_3360);
nand U3549 (N_3549,N_3339,N_3434);
or U3550 (N_3550,N_3269,N_3378);
nor U3551 (N_3551,N_3316,N_3352);
nor U3552 (N_3552,N_3418,N_3489);
nor U3553 (N_3553,N_3393,N_3468);
xnor U3554 (N_3554,N_3310,N_3295);
or U3555 (N_3555,N_3332,N_3304);
and U3556 (N_3556,N_3301,N_3330);
nand U3557 (N_3557,N_3415,N_3305);
or U3558 (N_3558,N_3476,N_3432);
nor U3559 (N_3559,N_3260,N_3292);
nand U3560 (N_3560,N_3398,N_3446);
nor U3561 (N_3561,N_3341,N_3478);
xor U3562 (N_3562,N_3448,N_3424);
xor U3563 (N_3563,N_3490,N_3496);
and U3564 (N_3564,N_3491,N_3409);
and U3565 (N_3565,N_3479,N_3314);
and U3566 (N_3566,N_3410,N_3347);
and U3567 (N_3567,N_3277,N_3362);
or U3568 (N_3568,N_3411,N_3492);
or U3569 (N_3569,N_3481,N_3273);
and U3570 (N_3570,N_3414,N_3451);
and U3571 (N_3571,N_3423,N_3276);
xnor U3572 (N_3572,N_3361,N_3384);
nor U3573 (N_3573,N_3498,N_3312);
xor U3574 (N_3574,N_3359,N_3319);
nor U3575 (N_3575,N_3422,N_3435);
or U3576 (N_3576,N_3382,N_3266);
nand U3577 (N_3577,N_3392,N_3288);
xnor U3578 (N_3578,N_3400,N_3279);
xor U3579 (N_3579,N_3385,N_3278);
and U3580 (N_3580,N_3429,N_3308);
nor U3581 (N_3581,N_3459,N_3375);
xnor U3582 (N_3582,N_3315,N_3270);
xor U3583 (N_3583,N_3387,N_3329);
or U3584 (N_3584,N_3473,N_3291);
or U3585 (N_3585,N_3267,N_3294);
nand U3586 (N_3586,N_3274,N_3405);
and U3587 (N_3587,N_3379,N_3430);
nand U3588 (N_3588,N_3487,N_3450);
xnor U3589 (N_3589,N_3377,N_3388);
xnor U3590 (N_3590,N_3455,N_3342);
nand U3591 (N_3591,N_3462,N_3281);
nand U3592 (N_3592,N_3282,N_3474);
nand U3593 (N_3593,N_3369,N_3254);
and U3594 (N_3594,N_3300,N_3311);
nand U3595 (N_3595,N_3253,N_3374);
and U3596 (N_3596,N_3334,N_3338);
nor U3597 (N_3597,N_3293,N_3381);
nor U3598 (N_3598,N_3497,N_3484);
nand U3599 (N_3599,N_3302,N_3457);
xor U3600 (N_3600,N_3268,N_3454);
nor U3601 (N_3601,N_3346,N_3485);
or U3602 (N_3602,N_3466,N_3307);
nand U3603 (N_3603,N_3364,N_3340);
or U3604 (N_3604,N_3354,N_3321);
or U3605 (N_3605,N_3357,N_3309);
nand U3606 (N_3606,N_3326,N_3447);
or U3607 (N_3607,N_3343,N_3284);
or U3608 (N_3608,N_3286,N_3404);
xor U3609 (N_3609,N_3296,N_3371);
and U3610 (N_3610,N_3395,N_3259);
xor U3611 (N_3611,N_3407,N_3391);
nand U3612 (N_3612,N_3413,N_3439);
nand U3613 (N_3613,N_3464,N_3265);
xnor U3614 (N_3614,N_3433,N_3376);
and U3615 (N_3615,N_3444,N_3380);
xnor U3616 (N_3616,N_3416,N_3394);
xnor U3617 (N_3617,N_3472,N_3461);
nand U3618 (N_3618,N_3350,N_3483);
or U3619 (N_3619,N_3345,N_3331);
and U3620 (N_3620,N_3456,N_3386);
nor U3621 (N_3621,N_3417,N_3327);
xnor U3622 (N_3622,N_3467,N_3275);
nor U3623 (N_3623,N_3420,N_3303);
and U3624 (N_3624,N_3348,N_3389);
xor U3625 (N_3625,N_3300,N_3401);
nand U3626 (N_3626,N_3288,N_3475);
nor U3627 (N_3627,N_3298,N_3275);
nand U3628 (N_3628,N_3448,N_3376);
nor U3629 (N_3629,N_3414,N_3286);
nand U3630 (N_3630,N_3490,N_3449);
or U3631 (N_3631,N_3250,N_3408);
nand U3632 (N_3632,N_3293,N_3403);
xor U3633 (N_3633,N_3373,N_3290);
xnor U3634 (N_3634,N_3367,N_3453);
nor U3635 (N_3635,N_3385,N_3368);
nand U3636 (N_3636,N_3302,N_3465);
and U3637 (N_3637,N_3385,N_3440);
nand U3638 (N_3638,N_3414,N_3357);
xor U3639 (N_3639,N_3327,N_3477);
and U3640 (N_3640,N_3459,N_3452);
and U3641 (N_3641,N_3411,N_3398);
and U3642 (N_3642,N_3414,N_3346);
and U3643 (N_3643,N_3292,N_3325);
nand U3644 (N_3644,N_3448,N_3282);
xnor U3645 (N_3645,N_3474,N_3255);
xnor U3646 (N_3646,N_3297,N_3493);
nand U3647 (N_3647,N_3390,N_3278);
or U3648 (N_3648,N_3401,N_3396);
and U3649 (N_3649,N_3266,N_3297);
nand U3650 (N_3650,N_3467,N_3379);
xor U3651 (N_3651,N_3315,N_3453);
nor U3652 (N_3652,N_3392,N_3265);
nor U3653 (N_3653,N_3407,N_3323);
nand U3654 (N_3654,N_3376,N_3425);
nor U3655 (N_3655,N_3406,N_3262);
nor U3656 (N_3656,N_3461,N_3251);
nor U3657 (N_3657,N_3373,N_3475);
nand U3658 (N_3658,N_3293,N_3256);
nor U3659 (N_3659,N_3357,N_3298);
or U3660 (N_3660,N_3383,N_3255);
and U3661 (N_3661,N_3383,N_3430);
or U3662 (N_3662,N_3371,N_3291);
and U3663 (N_3663,N_3281,N_3383);
nand U3664 (N_3664,N_3292,N_3357);
or U3665 (N_3665,N_3477,N_3275);
nor U3666 (N_3666,N_3282,N_3280);
and U3667 (N_3667,N_3294,N_3355);
nor U3668 (N_3668,N_3365,N_3369);
xor U3669 (N_3669,N_3471,N_3288);
nor U3670 (N_3670,N_3472,N_3325);
nor U3671 (N_3671,N_3460,N_3421);
nor U3672 (N_3672,N_3261,N_3355);
or U3673 (N_3673,N_3383,N_3442);
and U3674 (N_3674,N_3257,N_3306);
or U3675 (N_3675,N_3486,N_3288);
nor U3676 (N_3676,N_3400,N_3458);
nor U3677 (N_3677,N_3442,N_3307);
nor U3678 (N_3678,N_3443,N_3317);
nor U3679 (N_3679,N_3281,N_3455);
nor U3680 (N_3680,N_3251,N_3469);
and U3681 (N_3681,N_3495,N_3470);
xnor U3682 (N_3682,N_3344,N_3490);
nand U3683 (N_3683,N_3491,N_3306);
or U3684 (N_3684,N_3401,N_3385);
and U3685 (N_3685,N_3356,N_3426);
xnor U3686 (N_3686,N_3271,N_3330);
nand U3687 (N_3687,N_3287,N_3360);
nand U3688 (N_3688,N_3263,N_3494);
and U3689 (N_3689,N_3407,N_3359);
xnor U3690 (N_3690,N_3382,N_3355);
or U3691 (N_3691,N_3334,N_3454);
or U3692 (N_3692,N_3365,N_3385);
nand U3693 (N_3693,N_3488,N_3290);
xnor U3694 (N_3694,N_3374,N_3271);
xor U3695 (N_3695,N_3267,N_3462);
nor U3696 (N_3696,N_3328,N_3271);
nor U3697 (N_3697,N_3415,N_3324);
nor U3698 (N_3698,N_3339,N_3403);
and U3699 (N_3699,N_3483,N_3428);
nor U3700 (N_3700,N_3416,N_3328);
and U3701 (N_3701,N_3402,N_3460);
xor U3702 (N_3702,N_3253,N_3311);
xnor U3703 (N_3703,N_3414,N_3252);
or U3704 (N_3704,N_3462,N_3365);
nor U3705 (N_3705,N_3416,N_3432);
nand U3706 (N_3706,N_3314,N_3342);
or U3707 (N_3707,N_3323,N_3313);
or U3708 (N_3708,N_3339,N_3313);
or U3709 (N_3709,N_3412,N_3396);
xor U3710 (N_3710,N_3477,N_3467);
xor U3711 (N_3711,N_3258,N_3338);
nand U3712 (N_3712,N_3332,N_3301);
nand U3713 (N_3713,N_3398,N_3272);
nor U3714 (N_3714,N_3379,N_3342);
or U3715 (N_3715,N_3387,N_3440);
nand U3716 (N_3716,N_3281,N_3356);
or U3717 (N_3717,N_3459,N_3282);
xor U3718 (N_3718,N_3418,N_3389);
xor U3719 (N_3719,N_3267,N_3346);
nand U3720 (N_3720,N_3288,N_3476);
nor U3721 (N_3721,N_3376,N_3288);
and U3722 (N_3722,N_3289,N_3460);
or U3723 (N_3723,N_3355,N_3299);
and U3724 (N_3724,N_3260,N_3323);
nand U3725 (N_3725,N_3374,N_3285);
or U3726 (N_3726,N_3300,N_3383);
xnor U3727 (N_3727,N_3354,N_3462);
or U3728 (N_3728,N_3475,N_3387);
nand U3729 (N_3729,N_3361,N_3391);
xor U3730 (N_3730,N_3343,N_3312);
or U3731 (N_3731,N_3318,N_3390);
and U3732 (N_3732,N_3482,N_3278);
nor U3733 (N_3733,N_3416,N_3454);
and U3734 (N_3734,N_3352,N_3427);
or U3735 (N_3735,N_3404,N_3317);
or U3736 (N_3736,N_3309,N_3356);
and U3737 (N_3737,N_3300,N_3270);
or U3738 (N_3738,N_3262,N_3424);
nand U3739 (N_3739,N_3493,N_3341);
nor U3740 (N_3740,N_3404,N_3365);
or U3741 (N_3741,N_3484,N_3436);
and U3742 (N_3742,N_3430,N_3488);
or U3743 (N_3743,N_3338,N_3438);
nor U3744 (N_3744,N_3302,N_3393);
and U3745 (N_3745,N_3462,N_3490);
nor U3746 (N_3746,N_3475,N_3394);
nor U3747 (N_3747,N_3392,N_3376);
nand U3748 (N_3748,N_3444,N_3276);
and U3749 (N_3749,N_3480,N_3407);
nor U3750 (N_3750,N_3724,N_3519);
or U3751 (N_3751,N_3664,N_3518);
or U3752 (N_3752,N_3731,N_3744);
xnor U3753 (N_3753,N_3659,N_3588);
xnor U3754 (N_3754,N_3748,N_3740);
nand U3755 (N_3755,N_3680,N_3749);
nand U3756 (N_3756,N_3662,N_3728);
xnor U3757 (N_3757,N_3642,N_3734);
nand U3758 (N_3758,N_3556,N_3729);
and U3759 (N_3759,N_3550,N_3658);
or U3760 (N_3760,N_3527,N_3632);
and U3761 (N_3761,N_3657,N_3617);
nand U3762 (N_3762,N_3538,N_3641);
and U3763 (N_3763,N_3597,N_3705);
and U3764 (N_3764,N_3548,N_3513);
nand U3765 (N_3765,N_3634,N_3512);
nor U3766 (N_3766,N_3741,N_3521);
xor U3767 (N_3767,N_3569,N_3541);
xor U3768 (N_3768,N_3733,N_3544);
nand U3769 (N_3769,N_3668,N_3665);
xor U3770 (N_3770,N_3502,N_3675);
nand U3771 (N_3771,N_3537,N_3577);
nand U3772 (N_3772,N_3511,N_3661);
nand U3773 (N_3773,N_3655,N_3506);
nand U3774 (N_3774,N_3633,N_3670);
and U3775 (N_3775,N_3643,N_3745);
or U3776 (N_3776,N_3702,N_3660);
and U3777 (N_3777,N_3639,N_3534);
nor U3778 (N_3778,N_3644,N_3703);
nand U3779 (N_3779,N_3601,N_3524);
nand U3780 (N_3780,N_3585,N_3715);
and U3781 (N_3781,N_3546,N_3504);
nor U3782 (N_3782,N_3674,N_3507);
xor U3783 (N_3783,N_3543,N_3536);
nand U3784 (N_3784,N_3640,N_3626);
and U3785 (N_3785,N_3718,N_3528);
nor U3786 (N_3786,N_3720,N_3688);
and U3787 (N_3787,N_3686,N_3631);
and U3788 (N_3788,N_3553,N_3586);
nor U3789 (N_3789,N_3532,N_3619);
nand U3790 (N_3790,N_3738,N_3737);
nor U3791 (N_3791,N_3709,N_3630);
nand U3792 (N_3792,N_3520,N_3576);
xnor U3793 (N_3793,N_3522,N_3501);
xor U3794 (N_3794,N_3691,N_3531);
or U3795 (N_3795,N_3627,N_3578);
and U3796 (N_3796,N_3628,N_3525);
xor U3797 (N_3797,N_3547,N_3612);
xor U3798 (N_3798,N_3725,N_3567);
or U3799 (N_3799,N_3559,N_3594);
nand U3800 (N_3800,N_3574,N_3719);
xnor U3801 (N_3801,N_3678,N_3713);
xor U3802 (N_3802,N_3676,N_3746);
nor U3803 (N_3803,N_3714,N_3510);
or U3804 (N_3804,N_3539,N_3614);
and U3805 (N_3805,N_3560,N_3618);
xnor U3806 (N_3806,N_3636,N_3726);
and U3807 (N_3807,N_3505,N_3599);
and U3808 (N_3808,N_3698,N_3598);
or U3809 (N_3809,N_3591,N_3727);
and U3810 (N_3810,N_3516,N_3723);
or U3811 (N_3811,N_3517,N_3575);
nand U3812 (N_3812,N_3610,N_3721);
and U3813 (N_3813,N_3666,N_3672);
nor U3814 (N_3814,N_3566,N_3654);
nor U3815 (N_3815,N_3635,N_3595);
or U3816 (N_3816,N_3535,N_3604);
and U3817 (N_3817,N_3708,N_3616);
nand U3818 (N_3818,N_3648,N_3558);
nor U3819 (N_3819,N_3608,N_3609);
nor U3820 (N_3820,N_3707,N_3573);
and U3821 (N_3821,N_3596,N_3580);
xor U3822 (N_3822,N_3551,N_3603);
nand U3823 (N_3823,N_3572,N_3582);
xnor U3824 (N_3824,N_3717,N_3514);
and U3825 (N_3825,N_3523,N_3689);
xor U3826 (N_3826,N_3637,N_3568);
nand U3827 (N_3827,N_3682,N_3646);
and U3828 (N_3828,N_3623,N_3581);
nor U3829 (N_3829,N_3704,N_3681);
or U3830 (N_3830,N_3711,N_3621);
nand U3831 (N_3831,N_3656,N_3557);
xnor U3832 (N_3832,N_3542,N_3555);
nand U3833 (N_3833,N_3685,N_3700);
nand U3834 (N_3834,N_3692,N_3673);
nor U3835 (N_3835,N_3699,N_3683);
or U3836 (N_3836,N_3706,N_3624);
xor U3837 (N_3837,N_3684,N_3565);
nor U3838 (N_3838,N_3671,N_3590);
xnor U3839 (N_3839,N_3554,N_3645);
or U3840 (N_3840,N_3564,N_3722);
or U3841 (N_3841,N_3561,N_3697);
and U3842 (N_3842,N_3625,N_3562);
nor U3843 (N_3843,N_3508,N_3730);
xor U3844 (N_3844,N_3552,N_3739);
or U3845 (N_3845,N_3651,N_3742);
nand U3846 (N_3846,N_3736,N_3606);
xnor U3847 (N_3847,N_3607,N_3587);
and U3848 (N_3848,N_3638,N_3710);
nand U3849 (N_3849,N_3735,N_3500);
xor U3850 (N_3850,N_3600,N_3592);
nand U3851 (N_3851,N_3743,N_3677);
or U3852 (N_3852,N_3694,N_3696);
or U3853 (N_3853,N_3732,N_3622);
or U3854 (N_3854,N_3545,N_3563);
nor U3855 (N_3855,N_3652,N_3602);
or U3856 (N_3856,N_3613,N_3571);
or U3857 (N_3857,N_3515,N_3526);
xnor U3858 (N_3858,N_3570,N_3663);
and U3859 (N_3859,N_3647,N_3649);
nand U3860 (N_3860,N_3605,N_3687);
nor U3861 (N_3861,N_3579,N_3669);
and U3862 (N_3862,N_3667,N_3540);
xnor U3863 (N_3863,N_3693,N_3533);
xnor U3864 (N_3864,N_3629,N_3716);
or U3865 (N_3865,N_3615,N_3589);
or U3866 (N_3866,N_3701,N_3690);
xor U3867 (N_3867,N_3650,N_3530);
or U3868 (N_3868,N_3679,N_3549);
nand U3869 (N_3869,N_3503,N_3695);
nand U3870 (N_3870,N_3620,N_3584);
nand U3871 (N_3871,N_3593,N_3611);
nand U3872 (N_3872,N_3747,N_3509);
nand U3873 (N_3873,N_3529,N_3583);
nand U3874 (N_3874,N_3653,N_3712);
and U3875 (N_3875,N_3537,N_3665);
or U3876 (N_3876,N_3701,N_3625);
or U3877 (N_3877,N_3638,N_3728);
nand U3878 (N_3878,N_3691,N_3547);
or U3879 (N_3879,N_3718,N_3624);
xnor U3880 (N_3880,N_3736,N_3538);
and U3881 (N_3881,N_3712,N_3636);
and U3882 (N_3882,N_3520,N_3723);
or U3883 (N_3883,N_3714,N_3657);
nand U3884 (N_3884,N_3636,N_3717);
xor U3885 (N_3885,N_3727,N_3662);
xnor U3886 (N_3886,N_3504,N_3501);
xor U3887 (N_3887,N_3619,N_3544);
xnor U3888 (N_3888,N_3564,N_3529);
and U3889 (N_3889,N_3684,N_3524);
xor U3890 (N_3890,N_3525,N_3606);
or U3891 (N_3891,N_3560,N_3519);
or U3892 (N_3892,N_3743,N_3689);
nand U3893 (N_3893,N_3592,N_3528);
nand U3894 (N_3894,N_3603,N_3660);
nand U3895 (N_3895,N_3629,N_3538);
and U3896 (N_3896,N_3667,N_3725);
nor U3897 (N_3897,N_3610,N_3639);
nand U3898 (N_3898,N_3664,N_3643);
nand U3899 (N_3899,N_3668,N_3634);
nor U3900 (N_3900,N_3527,N_3728);
nor U3901 (N_3901,N_3746,N_3686);
nor U3902 (N_3902,N_3555,N_3503);
or U3903 (N_3903,N_3522,N_3520);
and U3904 (N_3904,N_3531,N_3551);
nand U3905 (N_3905,N_3631,N_3620);
nand U3906 (N_3906,N_3700,N_3741);
nor U3907 (N_3907,N_3551,N_3729);
xor U3908 (N_3908,N_3514,N_3553);
xor U3909 (N_3909,N_3500,N_3515);
or U3910 (N_3910,N_3585,N_3695);
xor U3911 (N_3911,N_3596,N_3682);
nor U3912 (N_3912,N_3576,N_3551);
and U3913 (N_3913,N_3549,N_3574);
or U3914 (N_3914,N_3570,N_3743);
or U3915 (N_3915,N_3542,N_3509);
xnor U3916 (N_3916,N_3632,N_3639);
nand U3917 (N_3917,N_3558,N_3566);
xor U3918 (N_3918,N_3570,N_3615);
or U3919 (N_3919,N_3584,N_3678);
nand U3920 (N_3920,N_3707,N_3562);
xnor U3921 (N_3921,N_3691,N_3533);
nor U3922 (N_3922,N_3705,N_3716);
xor U3923 (N_3923,N_3635,N_3535);
nor U3924 (N_3924,N_3568,N_3679);
nand U3925 (N_3925,N_3521,N_3608);
xnor U3926 (N_3926,N_3578,N_3620);
xnor U3927 (N_3927,N_3737,N_3715);
nor U3928 (N_3928,N_3725,N_3620);
nor U3929 (N_3929,N_3507,N_3579);
xnor U3930 (N_3930,N_3516,N_3520);
nor U3931 (N_3931,N_3501,N_3634);
or U3932 (N_3932,N_3621,N_3598);
or U3933 (N_3933,N_3734,N_3605);
nor U3934 (N_3934,N_3580,N_3599);
or U3935 (N_3935,N_3616,N_3683);
xnor U3936 (N_3936,N_3511,N_3538);
nor U3937 (N_3937,N_3632,N_3572);
nor U3938 (N_3938,N_3656,N_3548);
or U3939 (N_3939,N_3566,N_3530);
nand U3940 (N_3940,N_3627,N_3629);
or U3941 (N_3941,N_3713,N_3643);
and U3942 (N_3942,N_3722,N_3535);
or U3943 (N_3943,N_3513,N_3523);
nor U3944 (N_3944,N_3541,N_3553);
nor U3945 (N_3945,N_3546,N_3621);
nand U3946 (N_3946,N_3509,N_3684);
xnor U3947 (N_3947,N_3629,N_3534);
nand U3948 (N_3948,N_3518,N_3717);
nand U3949 (N_3949,N_3654,N_3641);
or U3950 (N_3950,N_3748,N_3545);
or U3951 (N_3951,N_3713,N_3542);
nand U3952 (N_3952,N_3562,N_3744);
nand U3953 (N_3953,N_3539,N_3660);
nand U3954 (N_3954,N_3501,N_3631);
nor U3955 (N_3955,N_3663,N_3742);
nand U3956 (N_3956,N_3551,N_3644);
nor U3957 (N_3957,N_3547,N_3645);
nand U3958 (N_3958,N_3616,N_3719);
or U3959 (N_3959,N_3512,N_3581);
nor U3960 (N_3960,N_3571,N_3668);
nand U3961 (N_3961,N_3744,N_3662);
or U3962 (N_3962,N_3616,N_3699);
and U3963 (N_3963,N_3613,N_3584);
nand U3964 (N_3964,N_3575,N_3620);
and U3965 (N_3965,N_3573,N_3675);
nand U3966 (N_3966,N_3673,N_3586);
or U3967 (N_3967,N_3538,N_3661);
nor U3968 (N_3968,N_3647,N_3730);
xor U3969 (N_3969,N_3648,N_3708);
nand U3970 (N_3970,N_3572,N_3681);
or U3971 (N_3971,N_3687,N_3512);
nand U3972 (N_3972,N_3634,N_3656);
or U3973 (N_3973,N_3692,N_3509);
nor U3974 (N_3974,N_3712,N_3713);
xnor U3975 (N_3975,N_3641,N_3514);
nor U3976 (N_3976,N_3730,N_3646);
nor U3977 (N_3977,N_3718,N_3546);
xnor U3978 (N_3978,N_3648,N_3582);
nor U3979 (N_3979,N_3565,N_3525);
nand U3980 (N_3980,N_3646,N_3684);
xor U3981 (N_3981,N_3502,N_3580);
nor U3982 (N_3982,N_3689,N_3727);
nor U3983 (N_3983,N_3674,N_3648);
and U3984 (N_3984,N_3567,N_3502);
and U3985 (N_3985,N_3653,N_3607);
xor U3986 (N_3986,N_3611,N_3646);
nand U3987 (N_3987,N_3633,N_3658);
or U3988 (N_3988,N_3690,N_3653);
xnor U3989 (N_3989,N_3547,N_3550);
and U3990 (N_3990,N_3674,N_3562);
or U3991 (N_3991,N_3654,N_3680);
xnor U3992 (N_3992,N_3623,N_3542);
and U3993 (N_3993,N_3675,N_3552);
and U3994 (N_3994,N_3522,N_3574);
or U3995 (N_3995,N_3572,N_3540);
or U3996 (N_3996,N_3617,N_3565);
or U3997 (N_3997,N_3515,N_3720);
or U3998 (N_3998,N_3515,N_3646);
nor U3999 (N_3999,N_3742,N_3563);
nand U4000 (N_4000,N_3803,N_3753);
nor U4001 (N_4001,N_3926,N_3777);
and U4002 (N_4002,N_3922,N_3770);
and U4003 (N_4003,N_3795,N_3906);
and U4004 (N_4004,N_3780,N_3824);
xor U4005 (N_4005,N_3932,N_3915);
nor U4006 (N_4006,N_3917,N_3785);
or U4007 (N_4007,N_3907,N_3869);
nand U4008 (N_4008,N_3769,N_3884);
and U4009 (N_4009,N_3923,N_3788);
or U4010 (N_4010,N_3796,N_3874);
nand U4011 (N_4011,N_3924,N_3763);
xnor U4012 (N_4012,N_3976,N_3837);
nor U4013 (N_4013,N_3895,N_3980);
or U4014 (N_4014,N_3776,N_3904);
or U4015 (N_4015,N_3896,N_3850);
xnor U4016 (N_4016,N_3921,N_3849);
or U4017 (N_4017,N_3998,N_3820);
xor U4018 (N_4018,N_3938,N_3978);
and U4019 (N_4019,N_3944,N_3897);
xnor U4020 (N_4020,N_3844,N_3819);
nor U4021 (N_4021,N_3965,N_3758);
and U4022 (N_4022,N_3905,N_3971);
or U4023 (N_4023,N_3989,N_3766);
and U4024 (N_4024,N_3969,N_3784);
nand U4025 (N_4025,N_3892,N_3867);
nor U4026 (N_4026,N_3960,N_3790);
nor U4027 (N_4027,N_3822,N_3750);
xnor U4028 (N_4028,N_3848,N_3950);
xnor U4029 (N_4029,N_3979,N_3830);
and U4030 (N_4030,N_3833,N_3885);
nor U4031 (N_4031,N_3811,N_3786);
xnor U4032 (N_4032,N_3875,N_3845);
and U4033 (N_4033,N_3759,N_3829);
nor U4034 (N_4034,N_3988,N_3768);
or U4035 (N_4035,N_3911,N_3963);
nor U4036 (N_4036,N_3870,N_3956);
xnor U4037 (N_4037,N_3983,N_3909);
and U4038 (N_4038,N_3787,N_3982);
nor U4039 (N_4039,N_3972,N_3990);
or U4040 (N_4040,N_3992,N_3903);
nor U4041 (N_4041,N_3826,N_3958);
nor U4042 (N_4042,N_3832,N_3880);
nor U4043 (N_4043,N_3818,N_3898);
and U4044 (N_4044,N_3856,N_3968);
and U4045 (N_4045,N_3952,N_3970);
or U4046 (N_4046,N_3984,N_3839);
or U4047 (N_4047,N_3751,N_3894);
and U4048 (N_4048,N_3806,N_3815);
nor U4049 (N_4049,N_3914,N_3858);
and U4050 (N_4050,N_3857,N_3912);
nor U4051 (N_4051,N_3812,N_3995);
nand U4052 (N_4052,N_3893,N_3999);
nand U4053 (N_4053,N_3836,N_3821);
nor U4054 (N_4054,N_3834,N_3800);
nand U4055 (N_4055,N_3953,N_3878);
or U4056 (N_4056,N_3919,N_3946);
nand U4057 (N_4057,N_3752,N_3765);
or U4058 (N_4058,N_3910,N_3762);
xor U4059 (N_4059,N_3756,N_3781);
nor U4060 (N_4060,N_3957,N_3817);
nand U4061 (N_4061,N_3846,N_3805);
nand U4062 (N_4062,N_3838,N_3901);
nand U4063 (N_4063,N_3929,N_3835);
xnor U4064 (N_4064,N_3890,N_3961);
nand U4065 (N_4065,N_3987,N_3948);
and U4066 (N_4066,N_3888,N_3927);
and U4067 (N_4067,N_3964,N_3852);
or U4068 (N_4068,N_3967,N_3810);
nand U4069 (N_4069,N_3775,N_3862);
nor U4070 (N_4070,N_3802,N_3936);
and U4071 (N_4071,N_3986,N_3974);
or U4072 (N_4072,N_3789,N_3814);
nand U4073 (N_4073,N_3851,N_3761);
and U4074 (N_4074,N_3935,N_3886);
and U4075 (N_4075,N_3954,N_3985);
nor U4076 (N_4076,N_3942,N_3782);
nor U4077 (N_4077,N_3792,N_3997);
nand U4078 (N_4078,N_3843,N_3823);
nand U4079 (N_4079,N_3783,N_3865);
xnor U4080 (N_4080,N_3757,N_3793);
and U4081 (N_4081,N_3841,N_3925);
or U4082 (N_4082,N_3881,N_3854);
nand U4083 (N_4083,N_3920,N_3827);
nor U4084 (N_4084,N_3930,N_3807);
or U4085 (N_4085,N_3861,N_3918);
nor U4086 (N_4086,N_3916,N_3873);
nand U4087 (N_4087,N_3872,N_3991);
nand U4088 (N_4088,N_3816,N_3764);
nand U4089 (N_4089,N_3864,N_3799);
nor U4090 (N_4090,N_3966,N_3772);
xor U4091 (N_4091,N_3859,N_3778);
and U4092 (N_4092,N_3801,N_3868);
xnor U4093 (N_4093,N_3931,N_3913);
and U4094 (N_4094,N_3853,N_3809);
and U4095 (N_4095,N_3900,N_3831);
nor U4096 (N_4096,N_3755,N_3804);
nand U4097 (N_4097,N_3949,N_3860);
and U4098 (N_4098,N_3975,N_3808);
nor U4099 (N_4099,N_3981,N_3933);
or U4100 (N_4100,N_3791,N_3876);
and U4101 (N_4101,N_3959,N_3899);
and U4102 (N_4102,N_3994,N_3891);
and U4103 (N_4103,N_3879,N_3940);
or U4104 (N_4104,N_3798,N_3908);
xnor U4105 (N_4105,N_3855,N_3828);
or U4106 (N_4106,N_3840,N_3794);
nor U4107 (N_4107,N_3902,N_3847);
and U4108 (N_4108,N_3797,N_3996);
and U4109 (N_4109,N_3973,N_3882);
nand U4110 (N_4110,N_3813,N_3887);
nor U4111 (N_4111,N_3866,N_3773);
or U4112 (N_4112,N_3928,N_3825);
nor U4113 (N_4113,N_3760,N_3754);
or U4114 (N_4114,N_3945,N_3962);
xor U4115 (N_4115,N_3955,N_3871);
nand U4116 (N_4116,N_3842,N_3771);
or U4117 (N_4117,N_3977,N_3947);
xor U4118 (N_4118,N_3934,N_3774);
nor U4119 (N_4119,N_3943,N_3883);
or U4120 (N_4120,N_3863,N_3937);
nor U4121 (N_4121,N_3993,N_3767);
xor U4122 (N_4122,N_3941,N_3889);
and U4123 (N_4123,N_3951,N_3779);
xnor U4124 (N_4124,N_3877,N_3939);
nand U4125 (N_4125,N_3922,N_3889);
xnor U4126 (N_4126,N_3965,N_3925);
and U4127 (N_4127,N_3850,N_3777);
nand U4128 (N_4128,N_3797,N_3803);
or U4129 (N_4129,N_3894,N_3856);
xnor U4130 (N_4130,N_3850,N_3763);
xor U4131 (N_4131,N_3962,N_3787);
xnor U4132 (N_4132,N_3777,N_3880);
nand U4133 (N_4133,N_3865,N_3790);
nor U4134 (N_4134,N_3910,N_3828);
nor U4135 (N_4135,N_3764,N_3939);
nand U4136 (N_4136,N_3972,N_3891);
or U4137 (N_4137,N_3760,N_3932);
nand U4138 (N_4138,N_3780,N_3808);
nand U4139 (N_4139,N_3897,N_3988);
and U4140 (N_4140,N_3891,N_3776);
or U4141 (N_4141,N_3974,N_3834);
or U4142 (N_4142,N_3846,N_3971);
and U4143 (N_4143,N_3931,N_3927);
or U4144 (N_4144,N_3901,N_3947);
nor U4145 (N_4145,N_3808,N_3902);
and U4146 (N_4146,N_3889,N_3912);
nor U4147 (N_4147,N_3801,N_3927);
nor U4148 (N_4148,N_3939,N_3927);
or U4149 (N_4149,N_3798,N_3863);
nor U4150 (N_4150,N_3862,N_3848);
nand U4151 (N_4151,N_3901,N_3762);
nor U4152 (N_4152,N_3753,N_3995);
and U4153 (N_4153,N_3835,N_3897);
and U4154 (N_4154,N_3758,N_3942);
or U4155 (N_4155,N_3922,N_3921);
or U4156 (N_4156,N_3761,N_3854);
nor U4157 (N_4157,N_3795,N_3944);
xor U4158 (N_4158,N_3924,N_3750);
nor U4159 (N_4159,N_3933,N_3954);
nand U4160 (N_4160,N_3754,N_3772);
xor U4161 (N_4161,N_3860,N_3841);
nor U4162 (N_4162,N_3808,N_3870);
nand U4163 (N_4163,N_3852,N_3814);
nor U4164 (N_4164,N_3985,N_3865);
or U4165 (N_4165,N_3837,N_3886);
nand U4166 (N_4166,N_3785,N_3912);
nand U4167 (N_4167,N_3822,N_3930);
or U4168 (N_4168,N_3996,N_3756);
or U4169 (N_4169,N_3849,N_3913);
nand U4170 (N_4170,N_3984,N_3791);
or U4171 (N_4171,N_3799,N_3833);
xor U4172 (N_4172,N_3909,N_3966);
and U4173 (N_4173,N_3887,N_3928);
nand U4174 (N_4174,N_3819,N_3890);
or U4175 (N_4175,N_3843,N_3947);
and U4176 (N_4176,N_3977,N_3915);
and U4177 (N_4177,N_3865,N_3769);
nor U4178 (N_4178,N_3848,N_3767);
or U4179 (N_4179,N_3875,N_3847);
nand U4180 (N_4180,N_3799,N_3922);
xor U4181 (N_4181,N_3797,N_3852);
nand U4182 (N_4182,N_3968,N_3877);
xnor U4183 (N_4183,N_3848,N_3986);
nand U4184 (N_4184,N_3919,N_3893);
xnor U4185 (N_4185,N_3938,N_3799);
or U4186 (N_4186,N_3878,N_3879);
and U4187 (N_4187,N_3984,N_3983);
and U4188 (N_4188,N_3886,N_3802);
nor U4189 (N_4189,N_3968,N_3997);
and U4190 (N_4190,N_3824,N_3802);
xor U4191 (N_4191,N_3784,N_3974);
and U4192 (N_4192,N_3893,N_3924);
xnor U4193 (N_4193,N_3773,N_3777);
xnor U4194 (N_4194,N_3952,N_3763);
nand U4195 (N_4195,N_3768,N_3949);
nand U4196 (N_4196,N_3768,N_3806);
nand U4197 (N_4197,N_3939,N_3780);
or U4198 (N_4198,N_3837,N_3991);
nor U4199 (N_4199,N_3918,N_3929);
nand U4200 (N_4200,N_3796,N_3821);
nand U4201 (N_4201,N_3847,N_3873);
or U4202 (N_4202,N_3873,N_3988);
and U4203 (N_4203,N_3769,N_3764);
nor U4204 (N_4204,N_3837,N_3863);
nor U4205 (N_4205,N_3922,N_3805);
or U4206 (N_4206,N_3763,N_3843);
nand U4207 (N_4207,N_3972,N_3957);
or U4208 (N_4208,N_3986,N_3909);
nor U4209 (N_4209,N_3767,N_3904);
or U4210 (N_4210,N_3995,N_3867);
nor U4211 (N_4211,N_3808,N_3772);
and U4212 (N_4212,N_3932,N_3862);
xor U4213 (N_4213,N_3758,N_3825);
nor U4214 (N_4214,N_3813,N_3904);
nor U4215 (N_4215,N_3955,N_3944);
or U4216 (N_4216,N_3810,N_3751);
or U4217 (N_4217,N_3938,N_3939);
nand U4218 (N_4218,N_3822,N_3862);
nand U4219 (N_4219,N_3844,N_3823);
nor U4220 (N_4220,N_3804,N_3995);
nor U4221 (N_4221,N_3906,N_3902);
xnor U4222 (N_4222,N_3891,N_3934);
nor U4223 (N_4223,N_3838,N_3916);
or U4224 (N_4224,N_3751,N_3762);
xnor U4225 (N_4225,N_3902,N_3838);
nor U4226 (N_4226,N_3994,N_3786);
and U4227 (N_4227,N_3752,N_3851);
or U4228 (N_4228,N_3842,N_3825);
and U4229 (N_4229,N_3880,N_3811);
nor U4230 (N_4230,N_3829,N_3873);
xnor U4231 (N_4231,N_3905,N_3763);
xor U4232 (N_4232,N_3934,N_3903);
nand U4233 (N_4233,N_3775,N_3932);
and U4234 (N_4234,N_3978,N_3804);
or U4235 (N_4235,N_3909,N_3836);
nor U4236 (N_4236,N_3877,N_3936);
nor U4237 (N_4237,N_3872,N_3804);
nand U4238 (N_4238,N_3807,N_3972);
and U4239 (N_4239,N_3964,N_3832);
nor U4240 (N_4240,N_3843,N_3876);
xnor U4241 (N_4241,N_3766,N_3851);
or U4242 (N_4242,N_3779,N_3766);
xor U4243 (N_4243,N_3865,N_3931);
nand U4244 (N_4244,N_3894,N_3780);
or U4245 (N_4245,N_3773,N_3781);
xnor U4246 (N_4246,N_3985,N_3908);
xor U4247 (N_4247,N_3832,N_3888);
or U4248 (N_4248,N_3888,N_3942);
nand U4249 (N_4249,N_3767,N_3837);
xnor U4250 (N_4250,N_4154,N_4235);
or U4251 (N_4251,N_4170,N_4055);
xnor U4252 (N_4252,N_4041,N_4056);
nor U4253 (N_4253,N_4140,N_4087);
and U4254 (N_4254,N_4149,N_4122);
or U4255 (N_4255,N_4010,N_4133);
nor U4256 (N_4256,N_4228,N_4023);
xnor U4257 (N_4257,N_4031,N_4136);
nand U4258 (N_4258,N_4244,N_4129);
and U4259 (N_4259,N_4179,N_4134);
or U4260 (N_4260,N_4232,N_4245);
and U4261 (N_4261,N_4003,N_4025);
nand U4262 (N_4262,N_4126,N_4046);
or U4263 (N_4263,N_4247,N_4182);
or U4264 (N_4264,N_4231,N_4117);
nor U4265 (N_4265,N_4180,N_4081);
and U4266 (N_4266,N_4050,N_4106);
nand U4267 (N_4267,N_4135,N_4205);
nor U4268 (N_4268,N_4236,N_4116);
xor U4269 (N_4269,N_4045,N_4004);
nor U4270 (N_4270,N_4162,N_4193);
nand U4271 (N_4271,N_4167,N_4014);
and U4272 (N_4272,N_4013,N_4137);
nand U4273 (N_4273,N_4121,N_4070);
xnor U4274 (N_4274,N_4184,N_4053);
nand U4275 (N_4275,N_4217,N_4212);
nor U4276 (N_4276,N_4157,N_4216);
nand U4277 (N_4277,N_4049,N_4108);
nor U4278 (N_4278,N_4089,N_4197);
xor U4279 (N_4279,N_4145,N_4096);
and U4280 (N_4280,N_4099,N_4102);
and U4281 (N_4281,N_4153,N_4227);
xor U4282 (N_4282,N_4033,N_4036);
nand U4283 (N_4283,N_4171,N_4202);
and U4284 (N_4284,N_4026,N_4011);
and U4285 (N_4285,N_4063,N_4047);
or U4286 (N_4286,N_4000,N_4176);
and U4287 (N_4287,N_4206,N_4187);
and U4288 (N_4288,N_4175,N_4163);
nand U4289 (N_4289,N_4118,N_4028);
or U4290 (N_4290,N_4119,N_4148);
nand U4291 (N_4291,N_4172,N_4141);
or U4292 (N_4292,N_4181,N_4060);
nor U4293 (N_4293,N_4094,N_4083);
or U4294 (N_4294,N_4128,N_4072);
xor U4295 (N_4295,N_4224,N_4146);
nor U4296 (N_4296,N_4085,N_4188);
nor U4297 (N_4297,N_4071,N_4018);
xor U4298 (N_4298,N_4221,N_4169);
xor U4299 (N_4299,N_4009,N_4067);
and U4300 (N_4300,N_4032,N_4204);
and U4301 (N_4301,N_4142,N_4074);
nand U4302 (N_4302,N_4120,N_4064);
xnor U4303 (N_4303,N_4103,N_4022);
or U4304 (N_4304,N_4203,N_4002);
nand U4305 (N_4305,N_4138,N_4243);
xor U4306 (N_4306,N_4210,N_4185);
nor U4307 (N_4307,N_4090,N_4048);
nand U4308 (N_4308,N_4143,N_4226);
or U4309 (N_4309,N_4068,N_4110);
xnor U4310 (N_4310,N_4211,N_4069);
xnor U4311 (N_4311,N_4194,N_4017);
and U4312 (N_4312,N_4218,N_4214);
or U4313 (N_4313,N_4127,N_4076);
nand U4314 (N_4314,N_4015,N_4132);
xnor U4315 (N_4315,N_4125,N_4209);
or U4316 (N_4316,N_4101,N_4020);
nand U4317 (N_4317,N_4091,N_4215);
and U4318 (N_4318,N_4173,N_4238);
and U4319 (N_4319,N_4156,N_4027);
nor U4320 (N_4320,N_4054,N_4016);
and U4321 (N_4321,N_4177,N_4174);
nand U4322 (N_4322,N_4240,N_4124);
or U4323 (N_4323,N_4104,N_4159);
nand U4324 (N_4324,N_4233,N_4196);
nor U4325 (N_4325,N_4065,N_4021);
and U4326 (N_4326,N_4160,N_4201);
xor U4327 (N_4327,N_4168,N_4225);
and U4328 (N_4328,N_4086,N_4029);
xor U4329 (N_4329,N_4079,N_4165);
or U4330 (N_4330,N_4005,N_4001);
nor U4331 (N_4331,N_4114,N_4057);
or U4332 (N_4332,N_4088,N_4246);
and U4333 (N_4333,N_4111,N_4190);
xnor U4334 (N_4334,N_4062,N_4147);
xor U4335 (N_4335,N_4078,N_4199);
or U4336 (N_4336,N_4059,N_4130);
nand U4337 (N_4337,N_4248,N_4024);
and U4338 (N_4338,N_4234,N_4042);
nand U4339 (N_4339,N_4229,N_4075);
nand U4340 (N_4340,N_4151,N_4166);
nand U4341 (N_4341,N_4223,N_4100);
or U4342 (N_4342,N_4112,N_4038);
nor U4343 (N_4343,N_4139,N_4061);
and U4344 (N_4344,N_4150,N_4186);
nand U4345 (N_4345,N_4035,N_4249);
and U4346 (N_4346,N_4030,N_4113);
nor U4347 (N_4347,N_4008,N_4207);
or U4348 (N_4348,N_4123,N_4158);
or U4349 (N_4349,N_4222,N_4080);
nor U4350 (N_4350,N_4107,N_4084);
xor U4351 (N_4351,N_4052,N_4043);
and U4352 (N_4352,N_4237,N_4098);
nor U4353 (N_4353,N_4093,N_4208);
nand U4354 (N_4354,N_4155,N_4044);
nor U4355 (N_4355,N_4242,N_4007);
xor U4356 (N_4356,N_4039,N_4239);
nor U4357 (N_4357,N_4241,N_4037);
and U4358 (N_4358,N_4066,N_4012);
or U4359 (N_4359,N_4095,N_4097);
and U4360 (N_4360,N_4115,N_4152);
xor U4361 (N_4361,N_4073,N_4161);
nand U4362 (N_4362,N_4191,N_4105);
or U4363 (N_4363,N_4198,N_4131);
or U4364 (N_4364,N_4183,N_4219);
nand U4365 (N_4365,N_4164,N_4178);
nand U4366 (N_4366,N_4058,N_4077);
and U4367 (N_4367,N_4034,N_4230);
and U4368 (N_4368,N_4051,N_4040);
nor U4369 (N_4369,N_4082,N_4144);
or U4370 (N_4370,N_4220,N_4006);
or U4371 (N_4371,N_4192,N_4195);
nor U4372 (N_4372,N_4092,N_4200);
xor U4373 (N_4373,N_4213,N_4189);
nand U4374 (N_4374,N_4109,N_4019);
nand U4375 (N_4375,N_4021,N_4177);
nand U4376 (N_4376,N_4030,N_4012);
and U4377 (N_4377,N_4110,N_4092);
or U4378 (N_4378,N_4197,N_4153);
or U4379 (N_4379,N_4072,N_4249);
xor U4380 (N_4380,N_4050,N_4113);
xnor U4381 (N_4381,N_4006,N_4120);
or U4382 (N_4382,N_4193,N_4054);
nor U4383 (N_4383,N_4184,N_4234);
or U4384 (N_4384,N_4146,N_4093);
xor U4385 (N_4385,N_4129,N_4064);
xnor U4386 (N_4386,N_4197,N_4208);
xnor U4387 (N_4387,N_4224,N_4227);
or U4388 (N_4388,N_4076,N_4114);
and U4389 (N_4389,N_4116,N_4168);
or U4390 (N_4390,N_4009,N_4228);
nand U4391 (N_4391,N_4202,N_4016);
and U4392 (N_4392,N_4083,N_4169);
or U4393 (N_4393,N_4235,N_4017);
and U4394 (N_4394,N_4048,N_4040);
xnor U4395 (N_4395,N_4131,N_4105);
or U4396 (N_4396,N_4122,N_4040);
xor U4397 (N_4397,N_4194,N_4248);
or U4398 (N_4398,N_4145,N_4161);
nand U4399 (N_4399,N_4182,N_4020);
nand U4400 (N_4400,N_4008,N_4173);
and U4401 (N_4401,N_4227,N_4209);
or U4402 (N_4402,N_4018,N_4202);
nor U4403 (N_4403,N_4088,N_4221);
or U4404 (N_4404,N_4040,N_4191);
and U4405 (N_4405,N_4098,N_4093);
and U4406 (N_4406,N_4152,N_4008);
xor U4407 (N_4407,N_4007,N_4146);
or U4408 (N_4408,N_4001,N_4015);
nor U4409 (N_4409,N_4088,N_4117);
or U4410 (N_4410,N_4140,N_4040);
xnor U4411 (N_4411,N_4003,N_4204);
and U4412 (N_4412,N_4139,N_4052);
and U4413 (N_4413,N_4035,N_4203);
and U4414 (N_4414,N_4113,N_4159);
or U4415 (N_4415,N_4173,N_4201);
xnor U4416 (N_4416,N_4116,N_4079);
nor U4417 (N_4417,N_4064,N_4160);
and U4418 (N_4418,N_4034,N_4141);
xnor U4419 (N_4419,N_4161,N_4166);
nand U4420 (N_4420,N_4054,N_4164);
or U4421 (N_4421,N_4005,N_4162);
and U4422 (N_4422,N_4239,N_4181);
nor U4423 (N_4423,N_4105,N_4189);
nor U4424 (N_4424,N_4235,N_4099);
and U4425 (N_4425,N_4191,N_4161);
nand U4426 (N_4426,N_4165,N_4166);
or U4427 (N_4427,N_4110,N_4186);
or U4428 (N_4428,N_4164,N_4225);
or U4429 (N_4429,N_4133,N_4190);
or U4430 (N_4430,N_4245,N_4021);
and U4431 (N_4431,N_4202,N_4088);
nor U4432 (N_4432,N_4057,N_4081);
xnor U4433 (N_4433,N_4078,N_4054);
and U4434 (N_4434,N_4152,N_4229);
or U4435 (N_4435,N_4201,N_4197);
or U4436 (N_4436,N_4150,N_4026);
nand U4437 (N_4437,N_4018,N_4168);
nand U4438 (N_4438,N_4115,N_4093);
xor U4439 (N_4439,N_4216,N_4224);
xor U4440 (N_4440,N_4241,N_4176);
and U4441 (N_4441,N_4020,N_4183);
xor U4442 (N_4442,N_4237,N_4162);
xor U4443 (N_4443,N_4107,N_4141);
or U4444 (N_4444,N_4071,N_4069);
or U4445 (N_4445,N_4207,N_4209);
nand U4446 (N_4446,N_4175,N_4184);
nor U4447 (N_4447,N_4247,N_4125);
and U4448 (N_4448,N_4019,N_4164);
nor U4449 (N_4449,N_4100,N_4180);
nor U4450 (N_4450,N_4176,N_4069);
and U4451 (N_4451,N_4020,N_4238);
nor U4452 (N_4452,N_4197,N_4085);
and U4453 (N_4453,N_4170,N_4116);
nand U4454 (N_4454,N_4153,N_4008);
and U4455 (N_4455,N_4242,N_4194);
and U4456 (N_4456,N_4210,N_4234);
xnor U4457 (N_4457,N_4193,N_4036);
nor U4458 (N_4458,N_4138,N_4054);
xnor U4459 (N_4459,N_4088,N_4190);
nor U4460 (N_4460,N_4122,N_4073);
and U4461 (N_4461,N_4203,N_4094);
nand U4462 (N_4462,N_4042,N_4075);
nor U4463 (N_4463,N_4007,N_4038);
nor U4464 (N_4464,N_4203,N_4162);
xor U4465 (N_4465,N_4190,N_4028);
xnor U4466 (N_4466,N_4025,N_4036);
nand U4467 (N_4467,N_4012,N_4028);
nand U4468 (N_4468,N_4090,N_4124);
nor U4469 (N_4469,N_4138,N_4115);
xor U4470 (N_4470,N_4093,N_4210);
and U4471 (N_4471,N_4132,N_4106);
and U4472 (N_4472,N_4054,N_4022);
nor U4473 (N_4473,N_4053,N_4162);
nor U4474 (N_4474,N_4078,N_4060);
or U4475 (N_4475,N_4038,N_4034);
nor U4476 (N_4476,N_4121,N_4194);
xor U4477 (N_4477,N_4055,N_4076);
xnor U4478 (N_4478,N_4222,N_4238);
nor U4479 (N_4479,N_4154,N_4125);
xnor U4480 (N_4480,N_4053,N_4231);
or U4481 (N_4481,N_4013,N_4123);
or U4482 (N_4482,N_4171,N_4096);
nand U4483 (N_4483,N_4191,N_4073);
nand U4484 (N_4484,N_4139,N_4124);
and U4485 (N_4485,N_4159,N_4093);
and U4486 (N_4486,N_4075,N_4048);
xnor U4487 (N_4487,N_4065,N_4004);
nand U4488 (N_4488,N_4061,N_4195);
and U4489 (N_4489,N_4038,N_4105);
xor U4490 (N_4490,N_4245,N_4045);
or U4491 (N_4491,N_4138,N_4045);
nor U4492 (N_4492,N_4227,N_4066);
nand U4493 (N_4493,N_4180,N_4201);
nor U4494 (N_4494,N_4012,N_4074);
nor U4495 (N_4495,N_4013,N_4191);
or U4496 (N_4496,N_4008,N_4076);
xnor U4497 (N_4497,N_4030,N_4045);
nand U4498 (N_4498,N_4032,N_4097);
nor U4499 (N_4499,N_4004,N_4019);
nor U4500 (N_4500,N_4494,N_4330);
xor U4501 (N_4501,N_4322,N_4477);
and U4502 (N_4502,N_4482,N_4470);
or U4503 (N_4503,N_4343,N_4369);
xnor U4504 (N_4504,N_4462,N_4487);
or U4505 (N_4505,N_4284,N_4434);
and U4506 (N_4506,N_4303,N_4358);
nor U4507 (N_4507,N_4262,N_4307);
xor U4508 (N_4508,N_4421,N_4376);
nand U4509 (N_4509,N_4313,N_4292);
or U4510 (N_4510,N_4269,N_4472);
and U4511 (N_4511,N_4306,N_4280);
and U4512 (N_4512,N_4281,N_4252);
nand U4513 (N_4513,N_4475,N_4411);
xor U4514 (N_4514,N_4394,N_4282);
nor U4515 (N_4515,N_4366,N_4398);
nor U4516 (N_4516,N_4317,N_4427);
nand U4517 (N_4517,N_4342,N_4350);
and U4518 (N_4518,N_4412,N_4444);
nor U4519 (N_4519,N_4495,N_4327);
and U4520 (N_4520,N_4288,N_4498);
xnor U4521 (N_4521,N_4432,N_4254);
xnor U4522 (N_4522,N_4344,N_4459);
nor U4523 (N_4523,N_4298,N_4290);
xnor U4524 (N_4524,N_4296,N_4471);
and U4525 (N_4525,N_4304,N_4357);
nand U4526 (N_4526,N_4389,N_4493);
xor U4527 (N_4527,N_4251,N_4364);
nand U4528 (N_4528,N_4271,N_4361);
or U4529 (N_4529,N_4287,N_4491);
and U4530 (N_4530,N_4426,N_4429);
xor U4531 (N_4531,N_4450,N_4309);
and U4532 (N_4532,N_4333,N_4469);
xnor U4533 (N_4533,N_4323,N_4331);
or U4534 (N_4534,N_4305,N_4410);
nor U4535 (N_4535,N_4338,N_4279);
nor U4536 (N_4536,N_4413,N_4285);
nand U4537 (N_4537,N_4250,N_4291);
nand U4538 (N_4538,N_4463,N_4419);
xnor U4539 (N_4539,N_4461,N_4267);
and U4540 (N_4540,N_4355,N_4422);
or U4541 (N_4541,N_4383,N_4439);
or U4542 (N_4542,N_4467,N_4380);
nor U4543 (N_4543,N_4485,N_4457);
nor U4544 (N_4544,N_4446,N_4480);
and U4545 (N_4545,N_4395,N_4295);
and U4546 (N_4546,N_4321,N_4385);
and U4547 (N_4547,N_4418,N_4393);
nand U4548 (N_4548,N_4356,N_4397);
or U4549 (N_4549,N_4415,N_4403);
or U4550 (N_4550,N_4399,N_4449);
nor U4551 (N_4551,N_4367,N_4371);
nand U4552 (N_4552,N_4276,N_4324);
and U4553 (N_4553,N_4318,N_4340);
xnor U4554 (N_4554,N_4489,N_4261);
nor U4555 (N_4555,N_4263,N_4320);
xnor U4556 (N_4556,N_4428,N_4479);
nor U4557 (N_4557,N_4414,N_4440);
nor U4558 (N_4558,N_4417,N_4329);
nand U4559 (N_4559,N_4497,N_4359);
and U4560 (N_4560,N_4386,N_4454);
and U4561 (N_4561,N_4264,N_4272);
nor U4562 (N_4562,N_4265,N_4373);
and U4563 (N_4563,N_4390,N_4260);
nor U4564 (N_4564,N_4308,N_4448);
nand U4565 (N_4565,N_4468,N_4409);
and U4566 (N_4566,N_4488,N_4314);
nand U4567 (N_4567,N_4381,N_4336);
nor U4568 (N_4568,N_4348,N_4388);
or U4569 (N_4569,N_4337,N_4431);
nor U4570 (N_4570,N_4266,N_4425);
nor U4571 (N_4571,N_4352,N_4456);
or U4572 (N_4572,N_4382,N_4401);
nand U4573 (N_4573,N_4496,N_4453);
nor U4574 (N_4574,N_4378,N_4402);
nand U4575 (N_4575,N_4436,N_4297);
nand U4576 (N_4576,N_4465,N_4377);
nand U4577 (N_4577,N_4408,N_4257);
nor U4578 (N_4578,N_4258,N_4283);
nor U4579 (N_4579,N_4384,N_4458);
xor U4580 (N_4580,N_4300,N_4286);
xor U4581 (N_4581,N_4325,N_4312);
or U4582 (N_4582,N_4478,N_4407);
or U4583 (N_4583,N_4430,N_4315);
or U4584 (N_4584,N_4374,N_4341);
and U4585 (N_4585,N_4435,N_4363);
nand U4586 (N_4586,N_4391,N_4351);
nor U4587 (N_4587,N_4289,N_4476);
nand U4588 (N_4588,N_4445,N_4362);
nor U4589 (N_4589,N_4474,N_4452);
and U4590 (N_4590,N_4311,N_4437);
or U4591 (N_4591,N_4372,N_4392);
or U4592 (N_4592,N_4259,N_4473);
nor U4593 (N_4593,N_4294,N_4379);
xor U4594 (N_4594,N_4438,N_4274);
nor U4595 (N_4595,N_4416,N_4433);
and U4596 (N_4596,N_4484,N_4332);
or U4597 (N_4597,N_4370,N_4443);
nand U4598 (N_4598,N_4277,N_4256);
nor U4599 (N_4599,N_4339,N_4483);
and U4600 (N_4600,N_4375,N_4404);
xnor U4601 (N_4601,N_4368,N_4451);
xnor U4602 (N_4602,N_4481,N_4420);
xnor U4603 (N_4603,N_4268,N_4400);
and U4604 (N_4604,N_4466,N_4405);
nor U4605 (N_4605,N_4492,N_4486);
xnor U4606 (N_4606,N_4302,N_4293);
or U4607 (N_4607,N_4353,N_4354);
nor U4608 (N_4608,N_4346,N_4441);
nand U4609 (N_4609,N_4406,N_4328);
nand U4610 (N_4610,N_4360,N_4334);
or U4611 (N_4611,N_4278,N_4255);
nand U4612 (N_4612,N_4316,N_4464);
nor U4613 (N_4613,N_4270,N_4455);
nor U4614 (N_4614,N_4447,N_4273);
and U4615 (N_4615,N_4345,N_4424);
or U4616 (N_4616,N_4460,N_4387);
or U4617 (N_4617,N_4253,N_4442);
nor U4618 (N_4618,N_4396,N_4310);
nor U4619 (N_4619,N_4326,N_4349);
nor U4620 (N_4620,N_4299,N_4275);
nand U4621 (N_4621,N_4347,N_4365);
xnor U4622 (N_4622,N_4499,N_4335);
and U4623 (N_4623,N_4319,N_4490);
and U4624 (N_4624,N_4423,N_4301);
or U4625 (N_4625,N_4357,N_4312);
or U4626 (N_4626,N_4497,N_4403);
xor U4627 (N_4627,N_4432,N_4357);
nor U4628 (N_4628,N_4273,N_4394);
nand U4629 (N_4629,N_4334,N_4374);
nor U4630 (N_4630,N_4483,N_4395);
xnor U4631 (N_4631,N_4440,N_4404);
or U4632 (N_4632,N_4406,N_4367);
and U4633 (N_4633,N_4458,N_4405);
and U4634 (N_4634,N_4448,N_4262);
nor U4635 (N_4635,N_4438,N_4320);
nor U4636 (N_4636,N_4422,N_4282);
and U4637 (N_4637,N_4456,N_4419);
nand U4638 (N_4638,N_4263,N_4276);
or U4639 (N_4639,N_4400,N_4445);
or U4640 (N_4640,N_4426,N_4255);
nand U4641 (N_4641,N_4483,N_4340);
and U4642 (N_4642,N_4337,N_4439);
nor U4643 (N_4643,N_4360,N_4353);
nor U4644 (N_4644,N_4334,N_4366);
xnor U4645 (N_4645,N_4467,N_4343);
or U4646 (N_4646,N_4264,N_4490);
xnor U4647 (N_4647,N_4288,N_4381);
xnor U4648 (N_4648,N_4356,N_4323);
nor U4649 (N_4649,N_4460,N_4266);
or U4650 (N_4650,N_4341,N_4464);
nor U4651 (N_4651,N_4388,N_4281);
and U4652 (N_4652,N_4438,N_4491);
nand U4653 (N_4653,N_4481,N_4456);
xnor U4654 (N_4654,N_4274,N_4383);
nand U4655 (N_4655,N_4392,N_4278);
and U4656 (N_4656,N_4306,N_4367);
nand U4657 (N_4657,N_4309,N_4381);
nand U4658 (N_4658,N_4258,N_4422);
or U4659 (N_4659,N_4410,N_4253);
xnor U4660 (N_4660,N_4412,N_4339);
or U4661 (N_4661,N_4398,N_4365);
and U4662 (N_4662,N_4325,N_4418);
nand U4663 (N_4663,N_4355,N_4414);
and U4664 (N_4664,N_4485,N_4260);
xor U4665 (N_4665,N_4394,N_4429);
and U4666 (N_4666,N_4492,N_4398);
or U4667 (N_4667,N_4332,N_4302);
nor U4668 (N_4668,N_4496,N_4385);
xnor U4669 (N_4669,N_4329,N_4355);
xnor U4670 (N_4670,N_4270,N_4360);
or U4671 (N_4671,N_4440,N_4441);
or U4672 (N_4672,N_4425,N_4418);
or U4673 (N_4673,N_4379,N_4409);
nand U4674 (N_4674,N_4481,N_4295);
nor U4675 (N_4675,N_4410,N_4283);
nor U4676 (N_4676,N_4491,N_4294);
nand U4677 (N_4677,N_4444,N_4331);
and U4678 (N_4678,N_4432,N_4343);
nor U4679 (N_4679,N_4447,N_4351);
or U4680 (N_4680,N_4464,N_4313);
xor U4681 (N_4681,N_4466,N_4397);
xor U4682 (N_4682,N_4255,N_4350);
xnor U4683 (N_4683,N_4323,N_4395);
nand U4684 (N_4684,N_4251,N_4270);
nand U4685 (N_4685,N_4461,N_4306);
xnor U4686 (N_4686,N_4363,N_4250);
nor U4687 (N_4687,N_4264,N_4346);
nand U4688 (N_4688,N_4373,N_4372);
xnor U4689 (N_4689,N_4361,N_4324);
and U4690 (N_4690,N_4411,N_4363);
or U4691 (N_4691,N_4270,N_4408);
nand U4692 (N_4692,N_4328,N_4277);
or U4693 (N_4693,N_4410,N_4465);
nor U4694 (N_4694,N_4254,N_4461);
and U4695 (N_4695,N_4305,N_4466);
xor U4696 (N_4696,N_4252,N_4337);
or U4697 (N_4697,N_4488,N_4382);
xor U4698 (N_4698,N_4365,N_4340);
xnor U4699 (N_4699,N_4482,N_4403);
and U4700 (N_4700,N_4384,N_4282);
xor U4701 (N_4701,N_4369,N_4494);
nor U4702 (N_4702,N_4262,N_4326);
nor U4703 (N_4703,N_4458,N_4481);
or U4704 (N_4704,N_4267,N_4302);
nand U4705 (N_4705,N_4362,N_4275);
or U4706 (N_4706,N_4393,N_4421);
nand U4707 (N_4707,N_4483,N_4325);
xor U4708 (N_4708,N_4342,N_4382);
nand U4709 (N_4709,N_4344,N_4418);
nand U4710 (N_4710,N_4325,N_4397);
or U4711 (N_4711,N_4490,N_4303);
nor U4712 (N_4712,N_4360,N_4454);
xor U4713 (N_4713,N_4256,N_4386);
or U4714 (N_4714,N_4400,N_4494);
or U4715 (N_4715,N_4460,N_4319);
or U4716 (N_4716,N_4430,N_4420);
and U4717 (N_4717,N_4307,N_4298);
and U4718 (N_4718,N_4424,N_4480);
nand U4719 (N_4719,N_4489,N_4288);
or U4720 (N_4720,N_4367,N_4352);
xor U4721 (N_4721,N_4383,N_4422);
nor U4722 (N_4722,N_4373,N_4381);
or U4723 (N_4723,N_4330,N_4437);
nor U4724 (N_4724,N_4260,N_4357);
nor U4725 (N_4725,N_4447,N_4300);
or U4726 (N_4726,N_4487,N_4370);
or U4727 (N_4727,N_4493,N_4268);
nor U4728 (N_4728,N_4332,N_4395);
xnor U4729 (N_4729,N_4368,N_4349);
nand U4730 (N_4730,N_4295,N_4463);
xnor U4731 (N_4731,N_4434,N_4382);
and U4732 (N_4732,N_4488,N_4446);
and U4733 (N_4733,N_4277,N_4331);
or U4734 (N_4734,N_4475,N_4466);
or U4735 (N_4735,N_4478,N_4356);
and U4736 (N_4736,N_4267,N_4293);
or U4737 (N_4737,N_4349,N_4313);
nor U4738 (N_4738,N_4479,N_4319);
xor U4739 (N_4739,N_4337,N_4497);
nor U4740 (N_4740,N_4325,N_4407);
nand U4741 (N_4741,N_4306,N_4499);
xnor U4742 (N_4742,N_4392,N_4477);
or U4743 (N_4743,N_4490,N_4431);
nand U4744 (N_4744,N_4473,N_4274);
xnor U4745 (N_4745,N_4261,N_4492);
nand U4746 (N_4746,N_4256,N_4475);
and U4747 (N_4747,N_4396,N_4252);
and U4748 (N_4748,N_4458,N_4273);
or U4749 (N_4749,N_4486,N_4461);
or U4750 (N_4750,N_4567,N_4712);
or U4751 (N_4751,N_4585,N_4557);
nor U4752 (N_4752,N_4556,N_4688);
and U4753 (N_4753,N_4690,N_4631);
nand U4754 (N_4754,N_4629,N_4543);
or U4755 (N_4755,N_4608,N_4583);
and U4756 (N_4756,N_4637,N_4587);
nand U4757 (N_4757,N_4730,N_4715);
or U4758 (N_4758,N_4737,N_4569);
or U4759 (N_4759,N_4521,N_4524);
or U4760 (N_4760,N_4577,N_4705);
xor U4761 (N_4761,N_4596,N_4736);
nand U4762 (N_4762,N_4536,N_4500);
xnor U4763 (N_4763,N_4575,N_4564);
and U4764 (N_4764,N_4535,N_4719);
xnor U4765 (N_4765,N_4619,N_4503);
xor U4766 (N_4766,N_4698,N_4630);
nand U4767 (N_4767,N_4611,N_4668);
nand U4768 (N_4768,N_4566,N_4646);
xor U4769 (N_4769,N_4592,N_4553);
or U4770 (N_4770,N_4538,N_4679);
and U4771 (N_4771,N_4732,N_4729);
xor U4772 (N_4772,N_4655,N_4509);
nand U4773 (N_4773,N_4501,N_4584);
xor U4774 (N_4774,N_4708,N_4692);
and U4775 (N_4775,N_4635,N_4512);
or U4776 (N_4776,N_4643,N_4505);
or U4777 (N_4777,N_4517,N_4714);
or U4778 (N_4778,N_4740,N_4595);
and U4779 (N_4779,N_4588,N_4523);
nand U4780 (N_4780,N_4573,N_4527);
xor U4781 (N_4781,N_4609,N_4651);
xor U4782 (N_4782,N_4615,N_4665);
or U4783 (N_4783,N_4604,N_4599);
nand U4784 (N_4784,N_4676,N_4534);
nand U4785 (N_4785,N_4576,N_4638);
nand U4786 (N_4786,N_4547,N_4673);
nor U4787 (N_4787,N_4516,N_4513);
nor U4788 (N_4788,N_4677,N_4626);
or U4789 (N_4789,N_4636,N_4649);
xor U4790 (N_4790,N_4525,N_4682);
and U4791 (N_4791,N_4519,N_4544);
or U4792 (N_4792,N_4614,N_4693);
or U4793 (N_4793,N_4537,N_4597);
xnor U4794 (N_4794,N_4617,N_4645);
nand U4795 (N_4795,N_4545,N_4733);
and U4796 (N_4796,N_4713,N_4704);
nand U4797 (N_4797,N_4650,N_4506);
and U4798 (N_4798,N_4647,N_4669);
xor U4799 (N_4799,N_4749,N_4558);
nor U4800 (N_4800,N_4685,N_4671);
nor U4801 (N_4801,N_4747,N_4510);
nand U4802 (N_4802,N_4548,N_4724);
and U4803 (N_4803,N_4530,N_4504);
xnor U4804 (N_4804,N_4582,N_4574);
and U4805 (N_4805,N_4533,N_4554);
nor U4806 (N_4806,N_4551,N_4623);
xor U4807 (N_4807,N_4628,N_4743);
or U4808 (N_4808,N_4586,N_4672);
or U4809 (N_4809,N_4684,N_4641);
and U4810 (N_4810,N_4546,N_4696);
xnor U4811 (N_4811,N_4687,N_4571);
and U4812 (N_4812,N_4560,N_4662);
or U4813 (N_4813,N_4702,N_4642);
or U4814 (N_4814,N_4520,N_4699);
nand U4815 (N_4815,N_4598,N_4689);
xnor U4816 (N_4816,N_4658,N_4652);
nand U4817 (N_4817,N_4578,N_4620);
nand U4818 (N_4818,N_4691,N_4694);
nor U4819 (N_4819,N_4541,N_4745);
and U4820 (N_4820,N_4563,N_4528);
and U4821 (N_4821,N_4559,N_4707);
xor U4822 (N_4822,N_4591,N_4674);
xnor U4823 (N_4823,N_4718,N_4744);
nor U4824 (N_4824,N_4640,N_4581);
xor U4825 (N_4825,N_4602,N_4670);
nand U4826 (N_4826,N_4697,N_4663);
nor U4827 (N_4827,N_4657,N_4700);
and U4828 (N_4828,N_4656,N_4717);
and U4829 (N_4829,N_4644,N_4526);
xor U4830 (N_4830,N_4661,N_4667);
xor U4831 (N_4831,N_4728,N_4675);
nor U4832 (N_4832,N_4603,N_4709);
and U4833 (N_4833,N_4622,N_4726);
or U4834 (N_4834,N_4561,N_4746);
nand U4835 (N_4835,N_4735,N_4706);
or U4836 (N_4836,N_4522,N_4727);
and U4837 (N_4837,N_4701,N_4664);
and U4838 (N_4838,N_4725,N_4508);
nand U4839 (N_4839,N_4552,N_4711);
and U4840 (N_4840,N_4632,N_4565);
nand U4841 (N_4841,N_4739,N_4678);
nor U4842 (N_4842,N_4593,N_4748);
or U4843 (N_4843,N_4531,N_4594);
nor U4844 (N_4844,N_4600,N_4666);
or U4845 (N_4845,N_4627,N_4514);
nor U4846 (N_4846,N_4741,N_4654);
or U4847 (N_4847,N_4634,N_4731);
and U4848 (N_4848,N_4695,N_4710);
nor U4849 (N_4849,N_4579,N_4555);
nand U4850 (N_4850,N_4625,N_4605);
and U4851 (N_4851,N_4721,N_4539);
nor U4852 (N_4852,N_4529,N_4502);
or U4853 (N_4853,N_4621,N_4624);
or U4854 (N_4854,N_4686,N_4590);
nand U4855 (N_4855,N_4703,N_4518);
nand U4856 (N_4856,N_4610,N_4738);
and U4857 (N_4857,N_4606,N_4681);
nor U4858 (N_4858,N_4580,N_4542);
xnor U4859 (N_4859,N_4601,N_4734);
xnor U4860 (N_4860,N_4723,N_4659);
xnor U4861 (N_4861,N_4633,N_4653);
nor U4862 (N_4862,N_4680,N_4618);
nor U4863 (N_4863,N_4683,N_4515);
nand U4864 (N_4864,N_4613,N_4607);
nor U4865 (N_4865,N_4722,N_4570);
nor U4866 (N_4866,N_4532,N_4568);
and U4867 (N_4867,N_4562,N_4549);
xor U4868 (N_4868,N_4720,N_4616);
nor U4869 (N_4869,N_4511,N_4540);
nor U4870 (N_4870,N_4660,N_4612);
xor U4871 (N_4871,N_4648,N_4716);
nor U4872 (N_4872,N_4742,N_4589);
nand U4873 (N_4873,N_4550,N_4572);
xor U4874 (N_4874,N_4507,N_4639);
xor U4875 (N_4875,N_4572,N_4694);
nor U4876 (N_4876,N_4621,N_4665);
or U4877 (N_4877,N_4724,N_4744);
nand U4878 (N_4878,N_4599,N_4520);
nand U4879 (N_4879,N_4636,N_4618);
and U4880 (N_4880,N_4519,N_4507);
xnor U4881 (N_4881,N_4640,N_4503);
nor U4882 (N_4882,N_4502,N_4743);
or U4883 (N_4883,N_4600,N_4735);
nand U4884 (N_4884,N_4522,N_4569);
nand U4885 (N_4885,N_4593,N_4555);
xor U4886 (N_4886,N_4677,N_4697);
and U4887 (N_4887,N_4674,N_4556);
nor U4888 (N_4888,N_4641,N_4661);
or U4889 (N_4889,N_4505,N_4728);
or U4890 (N_4890,N_4578,N_4676);
and U4891 (N_4891,N_4737,N_4655);
nor U4892 (N_4892,N_4649,N_4618);
nor U4893 (N_4893,N_4614,N_4507);
or U4894 (N_4894,N_4623,N_4648);
nor U4895 (N_4895,N_4600,N_4650);
nand U4896 (N_4896,N_4704,N_4722);
and U4897 (N_4897,N_4518,N_4563);
xnor U4898 (N_4898,N_4519,N_4590);
nand U4899 (N_4899,N_4689,N_4621);
or U4900 (N_4900,N_4634,N_4708);
xnor U4901 (N_4901,N_4704,N_4573);
nor U4902 (N_4902,N_4569,N_4666);
xnor U4903 (N_4903,N_4741,N_4674);
nand U4904 (N_4904,N_4549,N_4708);
or U4905 (N_4905,N_4577,N_4668);
nand U4906 (N_4906,N_4674,N_4748);
nand U4907 (N_4907,N_4747,N_4544);
nor U4908 (N_4908,N_4608,N_4743);
xnor U4909 (N_4909,N_4649,N_4537);
nand U4910 (N_4910,N_4558,N_4739);
and U4911 (N_4911,N_4547,N_4524);
nand U4912 (N_4912,N_4518,N_4599);
nand U4913 (N_4913,N_4629,N_4647);
or U4914 (N_4914,N_4665,N_4631);
or U4915 (N_4915,N_4522,N_4517);
or U4916 (N_4916,N_4707,N_4736);
and U4917 (N_4917,N_4626,N_4584);
nand U4918 (N_4918,N_4621,N_4625);
nor U4919 (N_4919,N_4509,N_4732);
and U4920 (N_4920,N_4697,N_4664);
or U4921 (N_4921,N_4743,N_4567);
nor U4922 (N_4922,N_4568,N_4577);
xnor U4923 (N_4923,N_4721,N_4660);
nor U4924 (N_4924,N_4664,N_4555);
or U4925 (N_4925,N_4571,N_4679);
xnor U4926 (N_4926,N_4720,N_4623);
or U4927 (N_4927,N_4707,N_4731);
nand U4928 (N_4928,N_4696,N_4712);
nand U4929 (N_4929,N_4573,N_4548);
or U4930 (N_4930,N_4681,N_4686);
nor U4931 (N_4931,N_4634,N_4584);
xnor U4932 (N_4932,N_4722,N_4628);
or U4933 (N_4933,N_4580,N_4738);
xor U4934 (N_4934,N_4587,N_4721);
nor U4935 (N_4935,N_4583,N_4691);
xnor U4936 (N_4936,N_4607,N_4503);
or U4937 (N_4937,N_4525,N_4610);
nor U4938 (N_4938,N_4698,N_4689);
xor U4939 (N_4939,N_4643,N_4539);
xnor U4940 (N_4940,N_4672,N_4532);
xor U4941 (N_4941,N_4605,N_4697);
or U4942 (N_4942,N_4725,N_4685);
or U4943 (N_4943,N_4702,N_4609);
or U4944 (N_4944,N_4501,N_4680);
and U4945 (N_4945,N_4642,N_4667);
and U4946 (N_4946,N_4653,N_4730);
or U4947 (N_4947,N_4639,N_4571);
xnor U4948 (N_4948,N_4525,N_4706);
or U4949 (N_4949,N_4632,N_4543);
nor U4950 (N_4950,N_4563,N_4708);
or U4951 (N_4951,N_4516,N_4540);
or U4952 (N_4952,N_4661,N_4558);
nand U4953 (N_4953,N_4519,N_4648);
and U4954 (N_4954,N_4594,N_4532);
nor U4955 (N_4955,N_4607,N_4501);
nand U4956 (N_4956,N_4590,N_4622);
nor U4957 (N_4957,N_4556,N_4516);
or U4958 (N_4958,N_4511,N_4711);
or U4959 (N_4959,N_4582,N_4549);
nor U4960 (N_4960,N_4549,N_4534);
nand U4961 (N_4961,N_4591,N_4640);
xnor U4962 (N_4962,N_4667,N_4626);
xor U4963 (N_4963,N_4529,N_4503);
or U4964 (N_4964,N_4603,N_4570);
or U4965 (N_4965,N_4584,N_4514);
xnor U4966 (N_4966,N_4540,N_4682);
nand U4967 (N_4967,N_4668,N_4736);
nand U4968 (N_4968,N_4511,N_4746);
or U4969 (N_4969,N_4619,N_4540);
and U4970 (N_4970,N_4554,N_4640);
nand U4971 (N_4971,N_4567,N_4605);
or U4972 (N_4972,N_4633,N_4739);
and U4973 (N_4973,N_4652,N_4700);
or U4974 (N_4974,N_4723,N_4748);
nand U4975 (N_4975,N_4645,N_4548);
nand U4976 (N_4976,N_4571,N_4699);
nand U4977 (N_4977,N_4712,N_4589);
nand U4978 (N_4978,N_4724,N_4523);
xor U4979 (N_4979,N_4626,N_4601);
xnor U4980 (N_4980,N_4672,N_4623);
nand U4981 (N_4981,N_4689,N_4601);
and U4982 (N_4982,N_4644,N_4586);
xor U4983 (N_4983,N_4569,N_4640);
xor U4984 (N_4984,N_4524,N_4541);
nand U4985 (N_4985,N_4508,N_4653);
or U4986 (N_4986,N_4514,N_4617);
nand U4987 (N_4987,N_4728,N_4560);
nand U4988 (N_4988,N_4730,N_4705);
and U4989 (N_4989,N_4630,N_4530);
nor U4990 (N_4990,N_4726,N_4576);
xnor U4991 (N_4991,N_4617,N_4505);
xnor U4992 (N_4992,N_4546,N_4716);
xor U4993 (N_4993,N_4726,N_4647);
or U4994 (N_4994,N_4538,N_4646);
nor U4995 (N_4995,N_4573,N_4639);
nor U4996 (N_4996,N_4622,N_4730);
and U4997 (N_4997,N_4577,N_4537);
nand U4998 (N_4998,N_4594,N_4502);
or U4999 (N_4999,N_4560,N_4683);
or U5000 (N_5000,N_4758,N_4930);
or U5001 (N_5001,N_4885,N_4760);
nor U5002 (N_5002,N_4899,N_4856);
nor U5003 (N_5003,N_4996,N_4862);
and U5004 (N_5004,N_4986,N_4750);
nand U5005 (N_5005,N_4827,N_4910);
xnor U5006 (N_5006,N_4824,N_4890);
xor U5007 (N_5007,N_4975,N_4840);
nand U5008 (N_5008,N_4917,N_4880);
nand U5009 (N_5009,N_4847,N_4763);
xnor U5010 (N_5010,N_4764,N_4867);
nand U5011 (N_5011,N_4762,N_4883);
xnor U5012 (N_5012,N_4989,N_4962);
or U5013 (N_5013,N_4804,N_4871);
nand U5014 (N_5014,N_4904,N_4822);
and U5015 (N_5015,N_4948,N_4855);
or U5016 (N_5016,N_4797,N_4935);
or U5017 (N_5017,N_4898,N_4915);
or U5018 (N_5018,N_4753,N_4994);
or U5019 (N_5019,N_4921,N_4909);
nand U5020 (N_5020,N_4928,N_4842);
and U5021 (N_5021,N_4980,N_4990);
or U5022 (N_5022,N_4852,N_4756);
or U5023 (N_5023,N_4821,N_4775);
xnor U5024 (N_5024,N_4950,N_4783);
nor U5025 (N_5025,N_4985,N_4901);
nand U5026 (N_5026,N_4944,N_4997);
or U5027 (N_5027,N_4964,N_4794);
nand U5028 (N_5028,N_4957,N_4864);
and U5029 (N_5029,N_4843,N_4854);
and U5030 (N_5030,N_4916,N_4933);
nor U5031 (N_5031,N_4981,N_4960);
and U5032 (N_5032,N_4979,N_4970);
xor U5033 (N_5033,N_4926,N_4788);
or U5034 (N_5034,N_4776,N_4959);
or U5035 (N_5035,N_4778,N_4799);
or U5036 (N_5036,N_4971,N_4768);
and U5037 (N_5037,N_4813,N_4936);
xnor U5038 (N_5038,N_4808,N_4995);
nand U5039 (N_5039,N_4943,N_4984);
xor U5040 (N_5040,N_4832,N_4913);
and U5041 (N_5041,N_4912,N_4868);
nor U5042 (N_5042,N_4789,N_4850);
and U5043 (N_5043,N_4825,N_4836);
and U5044 (N_5044,N_4860,N_4818);
and U5045 (N_5045,N_4781,N_4774);
nand U5046 (N_5046,N_4873,N_4896);
and U5047 (N_5047,N_4817,N_4988);
nand U5048 (N_5048,N_4844,N_4866);
or U5049 (N_5049,N_4881,N_4830);
and U5050 (N_5050,N_4805,N_4958);
nor U5051 (N_5051,N_4816,N_4888);
nand U5052 (N_5052,N_4780,N_4978);
nor U5053 (N_5053,N_4894,N_4861);
xnor U5054 (N_5054,N_4998,N_4754);
xor U5055 (N_5055,N_4870,N_4823);
nand U5056 (N_5056,N_4863,N_4982);
nand U5057 (N_5057,N_4927,N_4974);
nand U5058 (N_5058,N_4886,N_4908);
xnor U5059 (N_5059,N_4968,N_4769);
xnor U5060 (N_5060,N_4869,N_4900);
or U5061 (N_5061,N_4973,N_4963);
nor U5062 (N_5062,N_4892,N_4798);
nor U5063 (N_5063,N_4807,N_4949);
nor U5064 (N_5064,N_4846,N_4952);
nor U5065 (N_5065,N_4801,N_4879);
and U5066 (N_5066,N_4977,N_4993);
xor U5067 (N_5067,N_4777,N_4940);
and U5068 (N_5068,N_4865,N_4939);
nor U5069 (N_5069,N_4831,N_4945);
nand U5070 (N_5070,N_4877,N_4857);
xor U5071 (N_5071,N_4853,N_4884);
xor U5072 (N_5072,N_4755,N_4765);
nor U5073 (N_5073,N_4837,N_4903);
xnor U5074 (N_5074,N_4876,N_4923);
or U5075 (N_5075,N_4809,N_4951);
and U5076 (N_5076,N_4812,N_4925);
or U5077 (N_5077,N_4875,N_4829);
and U5078 (N_5078,N_4773,N_4838);
xor U5079 (N_5079,N_4793,N_4800);
nand U5080 (N_5080,N_4779,N_4999);
and U5081 (N_5081,N_4914,N_4972);
nand U5082 (N_5082,N_4924,N_4932);
or U5083 (N_5083,N_4992,N_4803);
nand U5084 (N_5084,N_4782,N_4893);
xor U5085 (N_5085,N_4983,N_4770);
and U5086 (N_5086,N_4859,N_4802);
and U5087 (N_5087,N_4839,N_4761);
xnor U5088 (N_5088,N_4759,N_4820);
nor U5089 (N_5089,N_4787,N_4810);
nor U5090 (N_5090,N_4791,N_4965);
or U5091 (N_5091,N_4766,N_4967);
or U5092 (N_5092,N_4889,N_4815);
nor U5093 (N_5093,N_4934,N_4772);
and U5094 (N_5094,N_4833,N_4796);
xnor U5095 (N_5095,N_4858,N_4942);
or U5096 (N_5096,N_4784,N_4874);
xor U5097 (N_5097,N_4969,N_4941);
and U5098 (N_5098,N_4991,N_4849);
or U5099 (N_5099,N_4786,N_4966);
and U5100 (N_5100,N_4757,N_4811);
or U5101 (N_5101,N_4938,N_4878);
nor U5102 (N_5102,N_4911,N_4851);
nand U5103 (N_5103,N_4918,N_4895);
nand U5104 (N_5104,N_4826,N_4835);
or U5105 (N_5105,N_4931,N_4887);
and U5106 (N_5106,N_4953,N_4905);
xnor U5107 (N_5107,N_4976,N_4897);
nor U5108 (N_5108,N_4767,N_4828);
xnor U5109 (N_5109,N_4961,N_4841);
xnor U5110 (N_5110,N_4906,N_4954);
nand U5111 (N_5111,N_4956,N_4790);
and U5112 (N_5112,N_4834,N_4920);
and U5113 (N_5113,N_4785,N_4882);
xor U5114 (N_5114,N_4922,N_4771);
or U5115 (N_5115,N_4891,N_4872);
and U5116 (N_5116,N_4929,N_4902);
nand U5117 (N_5117,N_4919,N_4955);
nand U5118 (N_5118,N_4845,N_4806);
xor U5119 (N_5119,N_4819,N_4848);
nand U5120 (N_5120,N_4792,N_4987);
or U5121 (N_5121,N_4946,N_4752);
nor U5122 (N_5122,N_4814,N_4947);
or U5123 (N_5123,N_4907,N_4937);
or U5124 (N_5124,N_4795,N_4751);
and U5125 (N_5125,N_4761,N_4949);
and U5126 (N_5126,N_4907,N_4757);
or U5127 (N_5127,N_4937,N_4974);
or U5128 (N_5128,N_4879,N_4883);
xnor U5129 (N_5129,N_4970,N_4791);
and U5130 (N_5130,N_4842,N_4853);
nor U5131 (N_5131,N_4862,N_4758);
xor U5132 (N_5132,N_4794,N_4847);
nand U5133 (N_5133,N_4923,N_4830);
xnor U5134 (N_5134,N_4864,N_4892);
nor U5135 (N_5135,N_4775,N_4913);
nand U5136 (N_5136,N_4808,N_4960);
xor U5137 (N_5137,N_4972,N_4970);
nand U5138 (N_5138,N_4799,N_4763);
and U5139 (N_5139,N_4753,N_4936);
xnor U5140 (N_5140,N_4906,N_4811);
nor U5141 (N_5141,N_4956,N_4847);
or U5142 (N_5142,N_4909,N_4858);
or U5143 (N_5143,N_4846,N_4894);
xor U5144 (N_5144,N_4987,N_4875);
nand U5145 (N_5145,N_4883,N_4761);
nor U5146 (N_5146,N_4879,N_4825);
and U5147 (N_5147,N_4781,N_4910);
xor U5148 (N_5148,N_4882,N_4915);
xnor U5149 (N_5149,N_4832,N_4940);
nand U5150 (N_5150,N_4851,N_4896);
xor U5151 (N_5151,N_4753,N_4832);
and U5152 (N_5152,N_4943,N_4989);
nor U5153 (N_5153,N_4805,N_4867);
and U5154 (N_5154,N_4897,N_4802);
nor U5155 (N_5155,N_4872,N_4835);
or U5156 (N_5156,N_4820,N_4914);
nand U5157 (N_5157,N_4964,N_4774);
nor U5158 (N_5158,N_4945,N_4916);
nor U5159 (N_5159,N_4884,N_4848);
xnor U5160 (N_5160,N_4885,N_4838);
nand U5161 (N_5161,N_4996,N_4999);
or U5162 (N_5162,N_4768,N_4983);
nor U5163 (N_5163,N_4883,N_4804);
nor U5164 (N_5164,N_4890,N_4915);
or U5165 (N_5165,N_4771,N_4797);
or U5166 (N_5166,N_4908,N_4888);
nor U5167 (N_5167,N_4894,N_4797);
nand U5168 (N_5168,N_4828,N_4927);
and U5169 (N_5169,N_4780,N_4775);
xor U5170 (N_5170,N_4955,N_4982);
nand U5171 (N_5171,N_4864,N_4803);
nand U5172 (N_5172,N_4845,N_4989);
and U5173 (N_5173,N_4940,N_4838);
and U5174 (N_5174,N_4958,N_4891);
nor U5175 (N_5175,N_4758,N_4871);
or U5176 (N_5176,N_4983,N_4930);
nand U5177 (N_5177,N_4970,N_4805);
nand U5178 (N_5178,N_4921,N_4764);
xnor U5179 (N_5179,N_4929,N_4759);
nand U5180 (N_5180,N_4928,N_4835);
and U5181 (N_5181,N_4801,N_4867);
and U5182 (N_5182,N_4845,N_4778);
nor U5183 (N_5183,N_4842,N_4891);
nor U5184 (N_5184,N_4794,N_4854);
xor U5185 (N_5185,N_4985,N_4832);
nand U5186 (N_5186,N_4929,N_4775);
and U5187 (N_5187,N_4769,N_4942);
nand U5188 (N_5188,N_4983,N_4912);
nor U5189 (N_5189,N_4968,N_4998);
xor U5190 (N_5190,N_4959,N_4894);
xnor U5191 (N_5191,N_4834,N_4977);
and U5192 (N_5192,N_4782,N_4960);
nand U5193 (N_5193,N_4917,N_4953);
and U5194 (N_5194,N_4922,N_4795);
and U5195 (N_5195,N_4758,N_4887);
nand U5196 (N_5196,N_4998,N_4927);
xor U5197 (N_5197,N_4792,N_4906);
or U5198 (N_5198,N_4998,N_4828);
nor U5199 (N_5199,N_4884,N_4891);
nand U5200 (N_5200,N_4881,N_4841);
and U5201 (N_5201,N_4864,N_4819);
nor U5202 (N_5202,N_4992,N_4936);
xnor U5203 (N_5203,N_4851,N_4752);
nand U5204 (N_5204,N_4923,N_4823);
xor U5205 (N_5205,N_4937,N_4829);
and U5206 (N_5206,N_4818,N_4890);
and U5207 (N_5207,N_4972,N_4792);
nand U5208 (N_5208,N_4988,N_4822);
nor U5209 (N_5209,N_4851,N_4964);
nor U5210 (N_5210,N_4793,N_4920);
xor U5211 (N_5211,N_4769,N_4912);
xor U5212 (N_5212,N_4820,N_4844);
nor U5213 (N_5213,N_4822,N_4986);
nor U5214 (N_5214,N_4923,N_4814);
and U5215 (N_5215,N_4837,N_4808);
nor U5216 (N_5216,N_4768,N_4905);
nand U5217 (N_5217,N_4825,N_4754);
and U5218 (N_5218,N_4780,N_4893);
nand U5219 (N_5219,N_4766,N_4781);
and U5220 (N_5220,N_4805,N_4952);
and U5221 (N_5221,N_4991,N_4915);
xor U5222 (N_5222,N_4795,N_4798);
nor U5223 (N_5223,N_4805,N_4964);
nand U5224 (N_5224,N_4973,N_4872);
xnor U5225 (N_5225,N_4891,N_4919);
and U5226 (N_5226,N_4926,N_4915);
nand U5227 (N_5227,N_4970,N_4775);
nand U5228 (N_5228,N_4855,N_4922);
nand U5229 (N_5229,N_4841,N_4957);
nor U5230 (N_5230,N_4950,N_4895);
nand U5231 (N_5231,N_4760,N_4889);
nand U5232 (N_5232,N_4842,N_4954);
nor U5233 (N_5233,N_4850,N_4906);
xor U5234 (N_5234,N_4981,N_4916);
xnor U5235 (N_5235,N_4894,N_4926);
nor U5236 (N_5236,N_4986,N_4782);
xor U5237 (N_5237,N_4961,N_4826);
nor U5238 (N_5238,N_4796,N_4765);
or U5239 (N_5239,N_4844,N_4767);
xor U5240 (N_5240,N_4957,N_4842);
and U5241 (N_5241,N_4860,N_4975);
nand U5242 (N_5242,N_4772,N_4840);
and U5243 (N_5243,N_4907,N_4941);
or U5244 (N_5244,N_4829,N_4838);
nand U5245 (N_5245,N_4794,N_4753);
or U5246 (N_5246,N_4927,N_4997);
or U5247 (N_5247,N_4837,N_4751);
or U5248 (N_5248,N_4788,N_4929);
xor U5249 (N_5249,N_4912,N_4956);
nor U5250 (N_5250,N_5111,N_5040);
and U5251 (N_5251,N_5159,N_5233);
and U5252 (N_5252,N_5082,N_5246);
nand U5253 (N_5253,N_5003,N_5012);
xnor U5254 (N_5254,N_5002,N_5187);
or U5255 (N_5255,N_5054,N_5090);
xor U5256 (N_5256,N_5170,N_5141);
xor U5257 (N_5257,N_5195,N_5125);
nand U5258 (N_5258,N_5210,N_5249);
and U5259 (N_5259,N_5147,N_5184);
or U5260 (N_5260,N_5023,N_5154);
or U5261 (N_5261,N_5069,N_5005);
and U5262 (N_5262,N_5174,N_5096);
or U5263 (N_5263,N_5139,N_5214);
nor U5264 (N_5264,N_5104,N_5133);
nand U5265 (N_5265,N_5025,N_5213);
and U5266 (N_5266,N_5020,N_5227);
xor U5267 (N_5267,N_5240,N_5135);
nand U5268 (N_5268,N_5228,N_5206);
nor U5269 (N_5269,N_5085,N_5065);
or U5270 (N_5270,N_5120,N_5110);
xor U5271 (N_5271,N_5118,N_5115);
and U5272 (N_5272,N_5089,N_5225);
xnor U5273 (N_5273,N_5245,N_5045);
nor U5274 (N_5274,N_5145,N_5030);
or U5275 (N_5275,N_5243,N_5209);
or U5276 (N_5276,N_5211,N_5168);
or U5277 (N_5277,N_5155,N_5208);
or U5278 (N_5278,N_5226,N_5117);
or U5279 (N_5279,N_5193,N_5015);
nor U5280 (N_5280,N_5018,N_5083);
nor U5281 (N_5281,N_5244,N_5132);
and U5282 (N_5282,N_5248,N_5217);
and U5283 (N_5283,N_5212,N_5163);
or U5284 (N_5284,N_5029,N_5199);
nor U5285 (N_5285,N_5241,N_5197);
or U5286 (N_5286,N_5027,N_5239);
or U5287 (N_5287,N_5032,N_5144);
xor U5288 (N_5288,N_5162,N_5181);
or U5289 (N_5289,N_5156,N_5143);
and U5290 (N_5290,N_5000,N_5234);
or U5291 (N_5291,N_5222,N_5112);
and U5292 (N_5292,N_5161,N_5024);
xor U5293 (N_5293,N_5176,N_5060);
nor U5294 (N_5294,N_5216,N_5014);
and U5295 (N_5295,N_5007,N_5198);
and U5296 (N_5296,N_5042,N_5073);
nand U5297 (N_5297,N_5140,N_5077);
or U5298 (N_5298,N_5131,N_5055);
xor U5299 (N_5299,N_5093,N_5021);
nor U5300 (N_5300,N_5220,N_5178);
nand U5301 (N_5301,N_5050,N_5201);
or U5302 (N_5302,N_5041,N_5231);
and U5303 (N_5303,N_5072,N_5011);
nand U5304 (N_5304,N_5238,N_5019);
nor U5305 (N_5305,N_5043,N_5204);
and U5306 (N_5306,N_5128,N_5049);
nand U5307 (N_5307,N_5129,N_5136);
and U5308 (N_5308,N_5190,N_5114);
nand U5309 (N_5309,N_5086,N_5183);
or U5310 (N_5310,N_5189,N_5048);
or U5311 (N_5311,N_5173,N_5009);
or U5312 (N_5312,N_5242,N_5106);
and U5313 (N_5313,N_5097,N_5013);
and U5314 (N_5314,N_5033,N_5078);
nor U5315 (N_5315,N_5022,N_5094);
and U5316 (N_5316,N_5108,N_5175);
or U5317 (N_5317,N_5230,N_5116);
and U5318 (N_5318,N_5063,N_5235);
and U5319 (N_5319,N_5105,N_5061);
nand U5320 (N_5320,N_5223,N_5130);
or U5321 (N_5321,N_5122,N_5107);
and U5322 (N_5322,N_5150,N_5177);
nand U5323 (N_5323,N_5124,N_5121);
xor U5324 (N_5324,N_5091,N_5188);
xor U5325 (N_5325,N_5057,N_5229);
or U5326 (N_5326,N_5098,N_5001);
nor U5327 (N_5327,N_5016,N_5102);
xor U5328 (N_5328,N_5010,N_5053);
and U5329 (N_5329,N_5247,N_5034);
nand U5330 (N_5330,N_5221,N_5182);
nor U5331 (N_5331,N_5171,N_5205);
nand U5332 (N_5332,N_5075,N_5166);
and U5333 (N_5333,N_5236,N_5200);
and U5334 (N_5334,N_5160,N_5026);
xnor U5335 (N_5335,N_5099,N_5064);
and U5336 (N_5336,N_5215,N_5056);
nand U5337 (N_5337,N_5169,N_5037);
or U5338 (N_5338,N_5146,N_5058);
xnor U5339 (N_5339,N_5047,N_5180);
xor U5340 (N_5340,N_5172,N_5237);
nand U5341 (N_5341,N_5192,N_5088);
nand U5342 (N_5342,N_5006,N_5028);
nor U5343 (N_5343,N_5036,N_5167);
or U5344 (N_5344,N_5157,N_5087);
xor U5345 (N_5345,N_5202,N_5185);
xnor U5346 (N_5346,N_5071,N_5126);
nand U5347 (N_5347,N_5046,N_5207);
nand U5348 (N_5348,N_5070,N_5044);
nor U5349 (N_5349,N_5059,N_5052);
nor U5350 (N_5350,N_5232,N_5138);
nand U5351 (N_5351,N_5031,N_5113);
nand U5352 (N_5352,N_5038,N_5151);
and U5353 (N_5353,N_5074,N_5039);
xnor U5354 (N_5354,N_5084,N_5165);
or U5355 (N_5355,N_5092,N_5080);
nand U5356 (N_5356,N_5123,N_5142);
xor U5357 (N_5357,N_5158,N_5008);
nor U5358 (N_5358,N_5004,N_5062);
or U5359 (N_5359,N_5219,N_5079);
or U5360 (N_5360,N_5153,N_5100);
xor U5361 (N_5361,N_5164,N_5218);
and U5362 (N_5362,N_5017,N_5196);
and U5363 (N_5363,N_5186,N_5149);
nand U5364 (N_5364,N_5127,N_5076);
and U5365 (N_5365,N_5148,N_5134);
nor U5366 (N_5366,N_5191,N_5119);
nor U5367 (N_5367,N_5152,N_5103);
xnor U5368 (N_5368,N_5203,N_5067);
xor U5369 (N_5369,N_5137,N_5101);
nand U5370 (N_5370,N_5095,N_5194);
nand U5371 (N_5371,N_5081,N_5179);
nor U5372 (N_5372,N_5035,N_5051);
or U5373 (N_5373,N_5068,N_5224);
xnor U5374 (N_5374,N_5109,N_5066);
nand U5375 (N_5375,N_5143,N_5162);
or U5376 (N_5376,N_5120,N_5149);
and U5377 (N_5377,N_5155,N_5224);
and U5378 (N_5378,N_5108,N_5133);
nand U5379 (N_5379,N_5166,N_5069);
nand U5380 (N_5380,N_5141,N_5126);
nand U5381 (N_5381,N_5193,N_5013);
or U5382 (N_5382,N_5228,N_5045);
nand U5383 (N_5383,N_5245,N_5226);
nor U5384 (N_5384,N_5224,N_5150);
xnor U5385 (N_5385,N_5049,N_5183);
or U5386 (N_5386,N_5027,N_5142);
and U5387 (N_5387,N_5172,N_5090);
and U5388 (N_5388,N_5079,N_5100);
xor U5389 (N_5389,N_5073,N_5086);
xor U5390 (N_5390,N_5224,N_5035);
xor U5391 (N_5391,N_5055,N_5051);
xnor U5392 (N_5392,N_5089,N_5109);
and U5393 (N_5393,N_5143,N_5075);
nor U5394 (N_5394,N_5088,N_5184);
nor U5395 (N_5395,N_5098,N_5141);
or U5396 (N_5396,N_5074,N_5246);
or U5397 (N_5397,N_5226,N_5081);
and U5398 (N_5398,N_5003,N_5217);
xnor U5399 (N_5399,N_5121,N_5042);
xnor U5400 (N_5400,N_5144,N_5228);
nand U5401 (N_5401,N_5029,N_5027);
or U5402 (N_5402,N_5204,N_5078);
nor U5403 (N_5403,N_5096,N_5145);
nor U5404 (N_5404,N_5185,N_5003);
or U5405 (N_5405,N_5088,N_5183);
and U5406 (N_5406,N_5237,N_5055);
nand U5407 (N_5407,N_5242,N_5176);
or U5408 (N_5408,N_5035,N_5210);
or U5409 (N_5409,N_5015,N_5070);
nor U5410 (N_5410,N_5084,N_5233);
xor U5411 (N_5411,N_5168,N_5130);
nand U5412 (N_5412,N_5174,N_5133);
or U5413 (N_5413,N_5134,N_5140);
or U5414 (N_5414,N_5094,N_5226);
or U5415 (N_5415,N_5013,N_5195);
or U5416 (N_5416,N_5163,N_5226);
or U5417 (N_5417,N_5137,N_5157);
xnor U5418 (N_5418,N_5157,N_5213);
xor U5419 (N_5419,N_5240,N_5136);
and U5420 (N_5420,N_5157,N_5210);
xor U5421 (N_5421,N_5180,N_5225);
or U5422 (N_5422,N_5007,N_5052);
or U5423 (N_5423,N_5238,N_5049);
or U5424 (N_5424,N_5211,N_5196);
or U5425 (N_5425,N_5131,N_5080);
nand U5426 (N_5426,N_5144,N_5148);
and U5427 (N_5427,N_5158,N_5014);
xor U5428 (N_5428,N_5075,N_5196);
nand U5429 (N_5429,N_5047,N_5087);
or U5430 (N_5430,N_5206,N_5019);
nor U5431 (N_5431,N_5139,N_5042);
nand U5432 (N_5432,N_5015,N_5146);
nor U5433 (N_5433,N_5173,N_5001);
and U5434 (N_5434,N_5070,N_5047);
nand U5435 (N_5435,N_5054,N_5240);
or U5436 (N_5436,N_5097,N_5049);
nor U5437 (N_5437,N_5147,N_5139);
or U5438 (N_5438,N_5157,N_5083);
or U5439 (N_5439,N_5061,N_5239);
or U5440 (N_5440,N_5156,N_5083);
or U5441 (N_5441,N_5124,N_5029);
or U5442 (N_5442,N_5147,N_5030);
xor U5443 (N_5443,N_5212,N_5174);
nor U5444 (N_5444,N_5074,N_5015);
or U5445 (N_5445,N_5054,N_5091);
nand U5446 (N_5446,N_5100,N_5166);
or U5447 (N_5447,N_5161,N_5158);
nor U5448 (N_5448,N_5239,N_5127);
nor U5449 (N_5449,N_5195,N_5050);
and U5450 (N_5450,N_5103,N_5109);
xor U5451 (N_5451,N_5191,N_5207);
xor U5452 (N_5452,N_5066,N_5222);
nor U5453 (N_5453,N_5233,N_5239);
nand U5454 (N_5454,N_5237,N_5247);
and U5455 (N_5455,N_5244,N_5228);
or U5456 (N_5456,N_5005,N_5105);
nand U5457 (N_5457,N_5033,N_5208);
xnor U5458 (N_5458,N_5203,N_5232);
and U5459 (N_5459,N_5004,N_5240);
and U5460 (N_5460,N_5208,N_5066);
or U5461 (N_5461,N_5161,N_5169);
or U5462 (N_5462,N_5003,N_5191);
xnor U5463 (N_5463,N_5017,N_5135);
nor U5464 (N_5464,N_5200,N_5179);
and U5465 (N_5465,N_5004,N_5108);
or U5466 (N_5466,N_5198,N_5095);
and U5467 (N_5467,N_5240,N_5043);
or U5468 (N_5468,N_5018,N_5148);
or U5469 (N_5469,N_5113,N_5207);
nor U5470 (N_5470,N_5074,N_5038);
xnor U5471 (N_5471,N_5131,N_5208);
or U5472 (N_5472,N_5226,N_5058);
nand U5473 (N_5473,N_5108,N_5186);
nand U5474 (N_5474,N_5172,N_5044);
nor U5475 (N_5475,N_5049,N_5161);
nor U5476 (N_5476,N_5075,N_5047);
or U5477 (N_5477,N_5237,N_5204);
or U5478 (N_5478,N_5119,N_5052);
nor U5479 (N_5479,N_5009,N_5147);
nand U5480 (N_5480,N_5208,N_5085);
xnor U5481 (N_5481,N_5202,N_5239);
xor U5482 (N_5482,N_5056,N_5203);
and U5483 (N_5483,N_5222,N_5180);
nand U5484 (N_5484,N_5173,N_5021);
or U5485 (N_5485,N_5215,N_5196);
nand U5486 (N_5486,N_5087,N_5046);
or U5487 (N_5487,N_5204,N_5123);
and U5488 (N_5488,N_5173,N_5108);
nor U5489 (N_5489,N_5092,N_5106);
nor U5490 (N_5490,N_5088,N_5042);
nand U5491 (N_5491,N_5219,N_5247);
or U5492 (N_5492,N_5215,N_5158);
xnor U5493 (N_5493,N_5197,N_5037);
and U5494 (N_5494,N_5170,N_5209);
xor U5495 (N_5495,N_5106,N_5043);
and U5496 (N_5496,N_5172,N_5098);
or U5497 (N_5497,N_5072,N_5026);
nor U5498 (N_5498,N_5011,N_5120);
xnor U5499 (N_5499,N_5127,N_5175);
or U5500 (N_5500,N_5261,N_5291);
xor U5501 (N_5501,N_5479,N_5497);
xor U5502 (N_5502,N_5401,N_5483);
xor U5503 (N_5503,N_5388,N_5443);
nor U5504 (N_5504,N_5438,N_5287);
and U5505 (N_5505,N_5278,N_5263);
and U5506 (N_5506,N_5283,N_5412);
nor U5507 (N_5507,N_5459,N_5432);
and U5508 (N_5508,N_5361,N_5471);
or U5509 (N_5509,N_5267,N_5450);
or U5510 (N_5510,N_5262,N_5408);
nand U5511 (N_5511,N_5323,N_5341);
or U5512 (N_5512,N_5436,N_5256);
or U5513 (N_5513,N_5268,N_5328);
xor U5514 (N_5514,N_5442,N_5290);
xor U5515 (N_5515,N_5304,N_5319);
xnor U5516 (N_5516,N_5332,N_5269);
nor U5517 (N_5517,N_5253,N_5416);
nor U5518 (N_5518,N_5277,N_5313);
xor U5519 (N_5519,N_5371,N_5308);
nor U5520 (N_5520,N_5469,N_5409);
nand U5521 (N_5521,N_5484,N_5357);
nand U5522 (N_5522,N_5329,N_5317);
and U5523 (N_5523,N_5399,N_5318);
nand U5524 (N_5524,N_5407,N_5423);
nand U5525 (N_5525,N_5372,N_5411);
xor U5526 (N_5526,N_5305,N_5280);
nand U5527 (N_5527,N_5316,N_5440);
xnor U5528 (N_5528,N_5380,N_5467);
nand U5529 (N_5529,N_5455,N_5474);
nand U5530 (N_5530,N_5499,N_5491);
nor U5531 (N_5531,N_5468,N_5314);
nor U5532 (N_5532,N_5342,N_5299);
xor U5533 (N_5533,N_5362,N_5393);
or U5534 (N_5534,N_5274,N_5335);
xor U5535 (N_5535,N_5338,N_5377);
nor U5536 (N_5536,N_5462,N_5494);
nand U5537 (N_5537,N_5309,N_5289);
nand U5538 (N_5538,N_5322,N_5394);
nor U5539 (N_5539,N_5281,N_5385);
and U5540 (N_5540,N_5360,N_5356);
or U5541 (N_5541,N_5434,N_5303);
or U5542 (N_5542,N_5458,N_5464);
nand U5543 (N_5543,N_5485,N_5252);
or U5544 (N_5544,N_5369,N_5365);
nand U5545 (N_5545,N_5441,N_5325);
nand U5546 (N_5546,N_5301,N_5446);
xor U5547 (N_5547,N_5279,N_5398);
or U5548 (N_5548,N_5306,N_5286);
nor U5549 (N_5549,N_5255,N_5363);
nor U5550 (N_5550,N_5354,N_5482);
nand U5551 (N_5551,N_5296,N_5430);
or U5552 (N_5552,N_5327,N_5344);
xor U5553 (N_5553,N_5271,N_5449);
nor U5554 (N_5554,N_5375,N_5498);
nor U5555 (N_5555,N_5366,N_5417);
or U5556 (N_5556,N_5295,N_5444);
and U5557 (N_5557,N_5374,N_5376);
xnor U5558 (N_5558,N_5367,N_5257);
nand U5559 (N_5559,N_5359,N_5390);
nand U5560 (N_5560,N_5452,N_5425);
or U5561 (N_5561,N_5473,N_5282);
and U5562 (N_5562,N_5272,N_5378);
nor U5563 (N_5563,N_5454,N_5493);
nand U5564 (N_5564,N_5403,N_5413);
or U5565 (N_5565,N_5463,N_5400);
nor U5566 (N_5566,N_5405,N_5324);
nand U5567 (N_5567,N_5448,N_5364);
nand U5568 (N_5568,N_5288,N_5495);
nor U5569 (N_5569,N_5435,N_5381);
or U5570 (N_5570,N_5476,N_5294);
nand U5571 (N_5571,N_5265,N_5461);
or U5572 (N_5572,N_5402,N_5336);
or U5573 (N_5573,N_5460,N_5453);
and U5574 (N_5574,N_5389,N_5297);
nand U5575 (N_5575,N_5259,N_5472);
and U5576 (N_5576,N_5445,N_5486);
nand U5577 (N_5577,N_5351,N_5475);
nor U5578 (N_5578,N_5273,N_5421);
and U5579 (N_5579,N_5391,N_5307);
and U5580 (N_5580,N_5312,N_5428);
xor U5581 (N_5581,N_5457,N_5422);
or U5582 (N_5582,N_5420,N_5370);
or U5583 (N_5583,N_5478,N_5410);
nand U5584 (N_5584,N_5333,N_5345);
nand U5585 (N_5585,N_5311,N_5386);
xnor U5586 (N_5586,N_5373,N_5431);
xnor U5587 (N_5587,N_5433,N_5418);
nand U5588 (N_5588,N_5326,N_5415);
xor U5589 (N_5589,N_5480,N_5260);
nor U5590 (N_5590,N_5368,N_5350);
or U5591 (N_5591,N_5488,N_5395);
or U5592 (N_5592,N_5315,N_5406);
or U5593 (N_5593,N_5258,N_5481);
nor U5594 (N_5594,N_5387,N_5320);
xor U5595 (N_5595,N_5451,N_5470);
xor U5596 (N_5596,N_5447,N_5264);
xnor U5597 (N_5597,N_5437,N_5339);
xor U5598 (N_5598,N_5419,N_5337);
nor U5599 (N_5599,N_5477,N_5250);
nand U5600 (N_5600,N_5358,N_5384);
nor U5601 (N_5601,N_5466,N_5404);
nor U5602 (N_5602,N_5284,N_5347);
nor U5603 (N_5603,N_5427,N_5348);
or U5604 (N_5604,N_5254,N_5275);
nand U5605 (N_5605,N_5396,N_5355);
nand U5606 (N_5606,N_5302,N_5382);
and U5607 (N_5607,N_5496,N_5349);
nand U5608 (N_5608,N_5353,N_5383);
or U5609 (N_5609,N_5492,N_5379);
nand U5610 (N_5610,N_5334,N_5340);
and U5611 (N_5611,N_5414,N_5392);
xor U5612 (N_5612,N_5270,N_5292);
or U5613 (N_5613,N_5352,N_5439);
and U5614 (N_5614,N_5266,N_5465);
nand U5615 (N_5615,N_5429,N_5487);
nand U5616 (N_5616,N_5298,N_5346);
or U5617 (N_5617,N_5343,N_5489);
xor U5618 (N_5618,N_5251,N_5397);
nor U5619 (N_5619,N_5456,N_5321);
nand U5620 (N_5620,N_5300,N_5490);
and U5621 (N_5621,N_5331,N_5293);
nor U5622 (N_5622,N_5426,N_5276);
nor U5623 (N_5623,N_5330,N_5285);
or U5624 (N_5624,N_5310,N_5424);
xnor U5625 (N_5625,N_5457,N_5414);
xnor U5626 (N_5626,N_5464,N_5296);
nand U5627 (N_5627,N_5348,N_5263);
nor U5628 (N_5628,N_5430,N_5363);
or U5629 (N_5629,N_5425,N_5318);
nand U5630 (N_5630,N_5425,N_5471);
xnor U5631 (N_5631,N_5304,N_5445);
or U5632 (N_5632,N_5451,N_5302);
nor U5633 (N_5633,N_5495,N_5289);
xor U5634 (N_5634,N_5464,N_5403);
and U5635 (N_5635,N_5289,N_5464);
nor U5636 (N_5636,N_5251,N_5279);
nor U5637 (N_5637,N_5439,N_5367);
or U5638 (N_5638,N_5311,N_5432);
or U5639 (N_5639,N_5452,N_5437);
xor U5640 (N_5640,N_5471,N_5426);
xnor U5641 (N_5641,N_5282,N_5272);
xor U5642 (N_5642,N_5415,N_5315);
nor U5643 (N_5643,N_5412,N_5288);
or U5644 (N_5644,N_5349,N_5294);
or U5645 (N_5645,N_5374,N_5488);
nand U5646 (N_5646,N_5484,N_5386);
xnor U5647 (N_5647,N_5460,N_5294);
and U5648 (N_5648,N_5350,N_5396);
and U5649 (N_5649,N_5427,N_5379);
and U5650 (N_5650,N_5380,N_5311);
nor U5651 (N_5651,N_5408,N_5281);
nor U5652 (N_5652,N_5396,N_5314);
xor U5653 (N_5653,N_5400,N_5446);
or U5654 (N_5654,N_5426,N_5457);
xnor U5655 (N_5655,N_5489,N_5367);
nor U5656 (N_5656,N_5425,N_5330);
nor U5657 (N_5657,N_5487,N_5355);
and U5658 (N_5658,N_5480,N_5368);
nor U5659 (N_5659,N_5312,N_5395);
and U5660 (N_5660,N_5262,N_5293);
nand U5661 (N_5661,N_5299,N_5325);
and U5662 (N_5662,N_5325,N_5300);
nor U5663 (N_5663,N_5432,N_5357);
nor U5664 (N_5664,N_5390,N_5377);
xnor U5665 (N_5665,N_5430,N_5288);
nor U5666 (N_5666,N_5472,N_5456);
and U5667 (N_5667,N_5447,N_5260);
or U5668 (N_5668,N_5394,N_5386);
nand U5669 (N_5669,N_5329,N_5255);
xor U5670 (N_5670,N_5317,N_5320);
xor U5671 (N_5671,N_5321,N_5490);
and U5672 (N_5672,N_5446,N_5324);
nand U5673 (N_5673,N_5338,N_5372);
nor U5674 (N_5674,N_5451,N_5358);
nor U5675 (N_5675,N_5360,N_5326);
and U5676 (N_5676,N_5429,N_5377);
nor U5677 (N_5677,N_5264,N_5381);
or U5678 (N_5678,N_5465,N_5337);
nand U5679 (N_5679,N_5305,N_5343);
nor U5680 (N_5680,N_5271,N_5496);
nor U5681 (N_5681,N_5418,N_5323);
or U5682 (N_5682,N_5458,N_5495);
nand U5683 (N_5683,N_5341,N_5335);
and U5684 (N_5684,N_5250,N_5342);
nor U5685 (N_5685,N_5397,N_5254);
and U5686 (N_5686,N_5473,N_5439);
or U5687 (N_5687,N_5309,N_5339);
xor U5688 (N_5688,N_5473,N_5336);
xor U5689 (N_5689,N_5358,N_5429);
xnor U5690 (N_5690,N_5440,N_5300);
and U5691 (N_5691,N_5378,N_5355);
or U5692 (N_5692,N_5393,N_5419);
and U5693 (N_5693,N_5276,N_5416);
xnor U5694 (N_5694,N_5466,N_5426);
nor U5695 (N_5695,N_5334,N_5288);
xor U5696 (N_5696,N_5309,N_5376);
or U5697 (N_5697,N_5472,N_5355);
nor U5698 (N_5698,N_5251,N_5398);
xor U5699 (N_5699,N_5339,N_5399);
nor U5700 (N_5700,N_5300,N_5452);
nand U5701 (N_5701,N_5348,N_5284);
xor U5702 (N_5702,N_5342,N_5270);
nand U5703 (N_5703,N_5469,N_5252);
xor U5704 (N_5704,N_5395,N_5435);
xor U5705 (N_5705,N_5398,N_5397);
xnor U5706 (N_5706,N_5281,N_5318);
xor U5707 (N_5707,N_5358,N_5269);
xor U5708 (N_5708,N_5362,N_5301);
xnor U5709 (N_5709,N_5351,N_5358);
and U5710 (N_5710,N_5296,N_5329);
and U5711 (N_5711,N_5263,N_5496);
and U5712 (N_5712,N_5486,N_5404);
nand U5713 (N_5713,N_5428,N_5305);
and U5714 (N_5714,N_5294,N_5497);
or U5715 (N_5715,N_5429,N_5431);
nor U5716 (N_5716,N_5321,N_5375);
xnor U5717 (N_5717,N_5314,N_5485);
nor U5718 (N_5718,N_5365,N_5371);
xnor U5719 (N_5719,N_5278,N_5266);
nor U5720 (N_5720,N_5430,N_5303);
and U5721 (N_5721,N_5336,N_5463);
xor U5722 (N_5722,N_5472,N_5345);
and U5723 (N_5723,N_5345,N_5349);
xnor U5724 (N_5724,N_5420,N_5462);
nor U5725 (N_5725,N_5330,N_5347);
xnor U5726 (N_5726,N_5474,N_5263);
nand U5727 (N_5727,N_5399,N_5451);
xnor U5728 (N_5728,N_5310,N_5290);
or U5729 (N_5729,N_5374,N_5493);
nor U5730 (N_5730,N_5282,N_5333);
and U5731 (N_5731,N_5270,N_5269);
nand U5732 (N_5732,N_5466,N_5398);
nor U5733 (N_5733,N_5369,N_5330);
and U5734 (N_5734,N_5482,N_5466);
or U5735 (N_5735,N_5469,N_5256);
nand U5736 (N_5736,N_5408,N_5295);
and U5737 (N_5737,N_5305,N_5273);
or U5738 (N_5738,N_5386,N_5422);
or U5739 (N_5739,N_5437,N_5350);
xor U5740 (N_5740,N_5461,N_5470);
nand U5741 (N_5741,N_5414,N_5399);
xnor U5742 (N_5742,N_5301,N_5478);
nor U5743 (N_5743,N_5488,N_5490);
nand U5744 (N_5744,N_5301,N_5273);
nand U5745 (N_5745,N_5346,N_5285);
nand U5746 (N_5746,N_5341,N_5356);
nor U5747 (N_5747,N_5473,N_5497);
nand U5748 (N_5748,N_5473,N_5338);
nand U5749 (N_5749,N_5259,N_5291);
and U5750 (N_5750,N_5618,N_5616);
xor U5751 (N_5751,N_5647,N_5668);
xor U5752 (N_5752,N_5586,N_5690);
nand U5753 (N_5753,N_5638,N_5521);
or U5754 (N_5754,N_5503,N_5508);
nor U5755 (N_5755,N_5667,N_5517);
or U5756 (N_5756,N_5661,N_5673);
nand U5757 (N_5757,N_5505,N_5604);
nand U5758 (N_5758,N_5737,N_5624);
xnor U5759 (N_5759,N_5590,N_5547);
or U5760 (N_5760,N_5636,N_5655);
xor U5761 (N_5761,N_5523,N_5736);
or U5762 (N_5762,N_5528,N_5657);
nand U5763 (N_5763,N_5536,N_5634);
or U5764 (N_5764,N_5645,N_5642);
nor U5765 (N_5765,N_5703,N_5600);
xnor U5766 (N_5766,N_5659,N_5622);
and U5767 (N_5767,N_5555,N_5591);
nor U5768 (N_5768,N_5646,N_5694);
xnor U5769 (N_5769,N_5734,N_5733);
and U5770 (N_5770,N_5565,N_5578);
or U5771 (N_5771,N_5558,N_5545);
and U5772 (N_5772,N_5715,N_5643);
nand U5773 (N_5773,N_5700,N_5705);
nand U5774 (N_5774,N_5524,N_5671);
nand U5775 (N_5775,N_5585,N_5619);
or U5776 (N_5776,N_5711,N_5731);
and U5777 (N_5777,N_5710,N_5539);
or U5778 (N_5778,N_5511,N_5682);
nor U5779 (N_5779,N_5632,N_5507);
nor U5780 (N_5780,N_5628,N_5670);
xnor U5781 (N_5781,N_5567,N_5575);
nand U5782 (N_5782,N_5743,N_5637);
nand U5783 (N_5783,N_5741,N_5656);
nor U5784 (N_5784,N_5553,N_5510);
nand U5785 (N_5785,N_5516,N_5685);
nand U5786 (N_5786,N_5641,N_5602);
or U5787 (N_5787,N_5698,N_5650);
xnor U5788 (N_5788,N_5720,N_5589);
nand U5789 (N_5789,N_5654,N_5688);
nand U5790 (N_5790,N_5631,N_5687);
or U5791 (N_5791,N_5635,N_5504);
nor U5792 (N_5792,N_5538,N_5730);
xor U5793 (N_5793,N_5615,N_5727);
xnor U5794 (N_5794,N_5546,N_5570);
nor U5795 (N_5795,N_5625,N_5584);
or U5796 (N_5796,N_5620,N_5571);
nand U5797 (N_5797,N_5531,N_5745);
xnor U5798 (N_5798,N_5725,N_5587);
nor U5799 (N_5799,N_5612,N_5593);
nor U5800 (N_5800,N_5562,N_5506);
nand U5801 (N_5801,N_5696,N_5701);
and U5802 (N_5802,N_5684,N_5629);
or U5803 (N_5803,N_5551,N_5563);
and U5804 (N_5804,N_5686,N_5706);
and U5805 (N_5805,N_5614,N_5648);
nor U5806 (N_5806,N_5713,N_5522);
nand U5807 (N_5807,N_5588,N_5738);
nor U5808 (N_5808,N_5535,N_5714);
and U5809 (N_5809,N_5679,N_5518);
xnor U5810 (N_5810,N_5735,N_5746);
nor U5811 (N_5811,N_5728,N_5542);
nor U5812 (N_5812,N_5739,N_5662);
nor U5813 (N_5813,N_5640,N_5515);
nand U5814 (N_5814,N_5644,N_5651);
xnor U5815 (N_5815,N_5717,N_5674);
nand U5816 (N_5816,N_5525,N_5649);
nor U5817 (N_5817,N_5676,N_5580);
or U5818 (N_5818,N_5729,N_5500);
and U5819 (N_5819,N_5557,N_5537);
nor U5820 (N_5820,N_5660,N_5617);
or U5821 (N_5821,N_5594,N_5527);
and U5822 (N_5822,N_5724,N_5675);
xor U5823 (N_5823,N_5598,N_5663);
nor U5824 (N_5824,N_5716,N_5672);
nor U5825 (N_5825,N_5561,N_5599);
xor U5826 (N_5826,N_5695,N_5573);
xor U5827 (N_5827,N_5549,N_5718);
or U5828 (N_5828,N_5689,N_5574);
xor U5829 (N_5829,N_5610,N_5582);
and U5830 (N_5830,N_5606,N_5566);
xnor U5831 (N_5831,N_5702,N_5568);
xnor U5832 (N_5832,N_5732,N_5658);
or U5833 (N_5833,N_5621,N_5595);
and U5834 (N_5834,N_5678,N_5577);
and U5835 (N_5835,N_5608,N_5550);
or U5836 (N_5836,N_5512,N_5699);
and U5837 (N_5837,N_5552,N_5559);
xnor U5838 (N_5838,N_5526,N_5747);
xor U5839 (N_5839,N_5540,N_5697);
nor U5840 (N_5840,N_5704,N_5677);
or U5841 (N_5841,N_5607,N_5601);
or U5842 (N_5842,N_5633,N_5722);
and U5843 (N_5843,N_5605,N_5592);
nor U5844 (N_5844,N_5639,N_5630);
nand U5845 (N_5845,N_5652,N_5581);
nand U5846 (N_5846,N_5572,N_5603);
and U5847 (N_5847,N_5556,N_5532);
nand U5848 (N_5848,N_5749,N_5583);
xnor U5849 (N_5849,N_5692,N_5613);
nor U5850 (N_5850,N_5740,N_5554);
or U5851 (N_5851,N_5627,N_5665);
nor U5852 (N_5852,N_5530,N_5712);
or U5853 (N_5853,N_5691,N_5534);
nor U5854 (N_5854,N_5707,N_5681);
nand U5855 (N_5855,N_5744,N_5723);
xnor U5856 (N_5856,N_5509,N_5569);
and U5857 (N_5857,N_5666,N_5560);
and U5858 (N_5858,N_5693,N_5683);
xor U5859 (N_5859,N_5721,N_5564);
and U5860 (N_5860,N_5519,N_5579);
xor U5861 (N_5861,N_5544,N_5596);
nand U5862 (N_5862,N_5576,N_5726);
nor U5863 (N_5863,N_5529,N_5541);
and U5864 (N_5864,N_5719,N_5520);
or U5865 (N_5865,N_5502,N_5623);
or U5866 (N_5866,N_5680,N_5611);
xor U5867 (N_5867,N_5742,N_5501);
nand U5868 (N_5868,N_5533,N_5653);
or U5869 (N_5869,N_5708,N_5664);
nand U5870 (N_5870,N_5669,N_5548);
nor U5871 (N_5871,N_5626,N_5597);
xor U5872 (N_5872,N_5514,N_5748);
and U5873 (N_5873,N_5543,N_5609);
nor U5874 (N_5874,N_5709,N_5513);
or U5875 (N_5875,N_5721,N_5728);
or U5876 (N_5876,N_5548,N_5510);
nand U5877 (N_5877,N_5688,N_5678);
nor U5878 (N_5878,N_5581,N_5692);
or U5879 (N_5879,N_5743,N_5725);
or U5880 (N_5880,N_5610,N_5638);
or U5881 (N_5881,N_5531,N_5722);
and U5882 (N_5882,N_5541,N_5548);
nor U5883 (N_5883,N_5527,N_5679);
nor U5884 (N_5884,N_5534,N_5546);
nand U5885 (N_5885,N_5740,N_5715);
xnor U5886 (N_5886,N_5697,N_5514);
xor U5887 (N_5887,N_5645,N_5550);
xnor U5888 (N_5888,N_5697,N_5691);
or U5889 (N_5889,N_5590,N_5533);
nand U5890 (N_5890,N_5723,N_5697);
and U5891 (N_5891,N_5675,N_5586);
nor U5892 (N_5892,N_5521,N_5660);
nand U5893 (N_5893,N_5732,N_5606);
xnor U5894 (N_5894,N_5611,N_5647);
and U5895 (N_5895,N_5631,N_5633);
and U5896 (N_5896,N_5619,N_5518);
nor U5897 (N_5897,N_5671,N_5537);
nor U5898 (N_5898,N_5681,N_5691);
nand U5899 (N_5899,N_5508,N_5674);
or U5900 (N_5900,N_5583,N_5745);
nand U5901 (N_5901,N_5729,N_5670);
and U5902 (N_5902,N_5513,N_5663);
and U5903 (N_5903,N_5524,N_5554);
and U5904 (N_5904,N_5713,N_5637);
nand U5905 (N_5905,N_5515,N_5596);
and U5906 (N_5906,N_5638,N_5702);
nor U5907 (N_5907,N_5556,N_5521);
and U5908 (N_5908,N_5635,N_5587);
nand U5909 (N_5909,N_5596,N_5608);
or U5910 (N_5910,N_5559,N_5694);
nand U5911 (N_5911,N_5616,N_5529);
nand U5912 (N_5912,N_5680,N_5523);
nor U5913 (N_5913,N_5653,N_5598);
xor U5914 (N_5914,N_5730,N_5548);
or U5915 (N_5915,N_5733,N_5710);
nand U5916 (N_5916,N_5696,N_5618);
xnor U5917 (N_5917,N_5635,N_5562);
xnor U5918 (N_5918,N_5503,N_5597);
and U5919 (N_5919,N_5509,N_5695);
or U5920 (N_5920,N_5584,N_5667);
xor U5921 (N_5921,N_5531,N_5717);
nand U5922 (N_5922,N_5704,N_5676);
nor U5923 (N_5923,N_5705,N_5659);
or U5924 (N_5924,N_5517,N_5706);
and U5925 (N_5925,N_5546,N_5619);
nand U5926 (N_5926,N_5612,N_5536);
nor U5927 (N_5927,N_5736,N_5532);
xnor U5928 (N_5928,N_5609,N_5584);
nor U5929 (N_5929,N_5697,N_5714);
and U5930 (N_5930,N_5713,N_5656);
nor U5931 (N_5931,N_5587,N_5650);
nor U5932 (N_5932,N_5688,N_5740);
nand U5933 (N_5933,N_5506,N_5567);
and U5934 (N_5934,N_5567,N_5570);
nand U5935 (N_5935,N_5539,N_5555);
nor U5936 (N_5936,N_5671,N_5644);
nand U5937 (N_5937,N_5524,N_5737);
and U5938 (N_5938,N_5609,N_5512);
or U5939 (N_5939,N_5676,N_5579);
nor U5940 (N_5940,N_5639,N_5562);
xnor U5941 (N_5941,N_5645,N_5655);
xnor U5942 (N_5942,N_5635,N_5577);
nor U5943 (N_5943,N_5580,N_5504);
nand U5944 (N_5944,N_5535,N_5591);
and U5945 (N_5945,N_5738,N_5506);
and U5946 (N_5946,N_5546,N_5605);
and U5947 (N_5947,N_5629,N_5590);
xor U5948 (N_5948,N_5538,N_5633);
nor U5949 (N_5949,N_5731,N_5633);
and U5950 (N_5950,N_5560,N_5502);
xnor U5951 (N_5951,N_5705,N_5729);
nand U5952 (N_5952,N_5628,N_5570);
xor U5953 (N_5953,N_5722,N_5661);
nor U5954 (N_5954,N_5554,N_5648);
or U5955 (N_5955,N_5618,N_5579);
and U5956 (N_5956,N_5654,N_5516);
nor U5957 (N_5957,N_5535,N_5583);
and U5958 (N_5958,N_5553,N_5722);
xnor U5959 (N_5959,N_5668,N_5625);
nor U5960 (N_5960,N_5611,N_5746);
and U5961 (N_5961,N_5654,N_5655);
nor U5962 (N_5962,N_5604,N_5652);
or U5963 (N_5963,N_5606,N_5730);
or U5964 (N_5964,N_5628,N_5505);
and U5965 (N_5965,N_5712,N_5721);
or U5966 (N_5966,N_5545,N_5717);
or U5967 (N_5967,N_5621,N_5725);
or U5968 (N_5968,N_5534,N_5662);
and U5969 (N_5969,N_5689,N_5675);
nand U5970 (N_5970,N_5675,N_5696);
or U5971 (N_5971,N_5669,N_5719);
nor U5972 (N_5972,N_5738,N_5746);
nand U5973 (N_5973,N_5747,N_5623);
nor U5974 (N_5974,N_5622,N_5575);
or U5975 (N_5975,N_5637,N_5664);
xor U5976 (N_5976,N_5623,N_5694);
xnor U5977 (N_5977,N_5557,N_5525);
xnor U5978 (N_5978,N_5506,N_5746);
xnor U5979 (N_5979,N_5628,N_5736);
nand U5980 (N_5980,N_5641,N_5617);
xor U5981 (N_5981,N_5682,N_5652);
xnor U5982 (N_5982,N_5627,N_5683);
or U5983 (N_5983,N_5561,N_5725);
xnor U5984 (N_5984,N_5525,N_5679);
xor U5985 (N_5985,N_5597,N_5669);
nor U5986 (N_5986,N_5549,N_5664);
or U5987 (N_5987,N_5740,N_5590);
nor U5988 (N_5988,N_5627,N_5522);
nor U5989 (N_5989,N_5724,N_5596);
and U5990 (N_5990,N_5679,N_5575);
nor U5991 (N_5991,N_5676,N_5571);
nor U5992 (N_5992,N_5593,N_5607);
nand U5993 (N_5993,N_5749,N_5676);
and U5994 (N_5994,N_5694,N_5569);
nor U5995 (N_5995,N_5625,N_5678);
and U5996 (N_5996,N_5721,N_5664);
nor U5997 (N_5997,N_5715,N_5648);
nand U5998 (N_5998,N_5736,N_5667);
xor U5999 (N_5999,N_5678,N_5557);
or U6000 (N_6000,N_5977,N_5963);
and U6001 (N_6001,N_5823,N_5979);
or U6002 (N_6002,N_5813,N_5885);
nand U6003 (N_6003,N_5850,N_5815);
nand U6004 (N_6004,N_5757,N_5770);
nor U6005 (N_6005,N_5990,N_5951);
nor U6006 (N_6006,N_5777,N_5988);
nor U6007 (N_6007,N_5836,N_5771);
and U6008 (N_6008,N_5843,N_5928);
xnor U6009 (N_6009,N_5837,N_5825);
nor U6010 (N_6010,N_5874,N_5911);
nand U6011 (N_6011,N_5931,N_5962);
nor U6012 (N_6012,N_5958,N_5844);
nand U6013 (N_6013,N_5792,N_5884);
and U6014 (N_6014,N_5966,N_5896);
or U6015 (N_6015,N_5876,N_5855);
and U6016 (N_6016,N_5760,N_5942);
nand U6017 (N_6017,N_5886,N_5801);
xnor U6018 (N_6018,N_5926,N_5915);
nand U6019 (N_6019,N_5961,N_5812);
nor U6020 (N_6020,N_5806,N_5793);
nand U6021 (N_6021,N_5953,N_5831);
and U6022 (N_6022,N_5819,N_5780);
and U6023 (N_6023,N_5754,N_5758);
and U6024 (N_6024,N_5827,N_5893);
nor U6025 (N_6025,N_5950,N_5860);
xnor U6026 (N_6026,N_5820,N_5755);
nand U6027 (N_6027,N_5762,N_5955);
or U6028 (N_6028,N_5790,N_5952);
or U6029 (N_6029,N_5861,N_5798);
or U6030 (N_6030,N_5808,N_5883);
nand U6031 (N_6031,N_5982,N_5769);
or U6032 (N_6032,N_5872,N_5787);
and U6033 (N_6033,N_5995,N_5975);
or U6034 (N_6034,N_5985,N_5869);
or U6035 (N_6035,N_5940,N_5935);
and U6036 (N_6036,N_5853,N_5878);
xnor U6037 (N_6037,N_5981,N_5903);
xor U6038 (N_6038,N_5774,N_5829);
nor U6039 (N_6039,N_5840,N_5773);
nand U6040 (N_6040,N_5752,N_5765);
nor U6041 (N_6041,N_5897,N_5838);
nand U6042 (N_6042,N_5857,N_5980);
xor U6043 (N_6043,N_5764,N_5870);
xnor U6044 (N_6044,N_5851,N_5889);
or U6045 (N_6045,N_5919,N_5892);
nand U6046 (N_6046,N_5946,N_5904);
nand U6047 (N_6047,N_5994,N_5880);
and U6048 (N_6048,N_5841,N_5927);
xnor U6049 (N_6049,N_5863,N_5772);
nand U6050 (N_6050,N_5879,N_5932);
or U6051 (N_6051,N_5828,N_5906);
or U6052 (N_6052,N_5751,N_5921);
nand U6053 (N_6053,N_5888,N_5865);
nor U6054 (N_6054,N_5845,N_5891);
nor U6055 (N_6055,N_5895,N_5766);
or U6056 (N_6056,N_5759,N_5991);
or U6057 (N_6057,N_5875,N_5978);
and U6058 (N_6058,N_5778,N_5954);
nor U6059 (N_6059,N_5924,N_5968);
nand U6060 (N_6060,N_5803,N_5934);
xor U6061 (N_6061,N_5923,N_5856);
nand U6062 (N_6062,N_5913,N_5937);
xnor U6063 (N_6063,N_5941,N_5871);
and U6064 (N_6064,N_5842,N_5796);
and U6065 (N_6065,N_5816,N_5784);
and U6066 (N_6066,N_5900,N_5914);
nand U6067 (N_6067,N_5992,N_5908);
nand U6068 (N_6068,N_5918,N_5789);
or U6069 (N_6069,N_5750,N_5993);
xor U6070 (N_6070,N_5902,N_5998);
nor U6071 (N_6071,N_5916,N_5894);
or U6072 (N_6072,N_5810,N_5852);
nand U6073 (N_6073,N_5881,N_5887);
or U6074 (N_6074,N_5948,N_5939);
xor U6075 (N_6075,N_5868,N_5910);
and U6076 (N_6076,N_5821,N_5965);
nor U6077 (N_6077,N_5767,N_5756);
xor U6078 (N_6078,N_5971,N_5936);
nand U6079 (N_6079,N_5802,N_5818);
nand U6080 (N_6080,N_5804,N_5817);
nor U6081 (N_6081,N_5768,N_5967);
xnor U6082 (N_6082,N_5794,N_5786);
and U6083 (N_6083,N_5989,N_5890);
nand U6084 (N_6084,N_5848,N_5944);
and U6085 (N_6085,N_5996,N_5933);
and U6086 (N_6086,N_5969,N_5938);
or U6087 (N_6087,N_5866,N_5877);
and U6088 (N_6088,N_5912,N_5864);
xnor U6089 (N_6089,N_5970,N_5800);
and U6090 (N_6090,N_5846,N_5832);
nor U6091 (N_6091,N_5809,N_5972);
or U6092 (N_6092,N_5779,N_5959);
xnor U6093 (N_6093,N_5834,N_5943);
nand U6094 (N_6094,N_5826,N_5882);
xor U6095 (N_6095,N_5781,N_5901);
xor U6096 (N_6096,N_5805,N_5899);
and U6097 (N_6097,N_5945,N_5814);
nand U6098 (N_6098,N_5983,N_5999);
nand U6099 (N_6099,N_5775,N_5947);
xor U6100 (N_6100,N_5930,N_5822);
nor U6101 (N_6101,N_5763,N_5839);
and U6102 (N_6102,N_5974,N_5791);
xnor U6103 (N_6103,N_5835,N_5811);
nor U6104 (N_6104,N_5905,N_5795);
xor U6105 (N_6105,N_5753,N_5956);
xor U6106 (N_6106,N_5907,N_5922);
or U6107 (N_6107,N_5929,N_5783);
xor U6108 (N_6108,N_5964,N_5854);
and U6109 (N_6109,N_5973,N_5785);
or U6110 (N_6110,N_5830,N_5782);
or U6111 (N_6111,N_5984,N_5824);
xor U6112 (N_6112,N_5960,N_5976);
xor U6113 (N_6113,N_5920,N_5862);
nand U6114 (N_6114,N_5761,N_5858);
nor U6115 (N_6115,N_5917,N_5957);
nand U6116 (N_6116,N_5833,N_5873);
and U6117 (N_6117,N_5847,N_5925);
nand U6118 (N_6118,N_5807,N_5849);
nor U6119 (N_6119,N_5986,N_5949);
and U6120 (N_6120,N_5776,N_5797);
nor U6121 (N_6121,N_5788,N_5909);
nand U6122 (N_6122,N_5859,N_5997);
and U6123 (N_6123,N_5867,N_5987);
or U6124 (N_6124,N_5799,N_5898);
or U6125 (N_6125,N_5774,N_5892);
or U6126 (N_6126,N_5881,N_5989);
xor U6127 (N_6127,N_5914,N_5898);
xor U6128 (N_6128,N_5761,N_5885);
nand U6129 (N_6129,N_5965,N_5931);
or U6130 (N_6130,N_5750,N_5904);
and U6131 (N_6131,N_5760,N_5754);
or U6132 (N_6132,N_5990,N_5817);
or U6133 (N_6133,N_5903,N_5805);
nor U6134 (N_6134,N_5776,N_5813);
and U6135 (N_6135,N_5794,N_5791);
nand U6136 (N_6136,N_5755,N_5860);
or U6137 (N_6137,N_5910,N_5802);
nor U6138 (N_6138,N_5924,N_5953);
and U6139 (N_6139,N_5885,N_5942);
xor U6140 (N_6140,N_5800,N_5804);
nand U6141 (N_6141,N_5806,N_5828);
nand U6142 (N_6142,N_5766,N_5893);
xor U6143 (N_6143,N_5779,N_5851);
xnor U6144 (N_6144,N_5888,N_5866);
nand U6145 (N_6145,N_5977,N_5878);
or U6146 (N_6146,N_5860,N_5764);
or U6147 (N_6147,N_5810,N_5995);
and U6148 (N_6148,N_5856,N_5823);
nand U6149 (N_6149,N_5761,N_5897);
nor U6150 (N_6150,N_5783,N_5840);
or U6151 (N_6151,N_5818,N_5855);
nand U6152 (N_6152,N_5988,N_5818);
nand U6153 (N_6153,N_5783,N_5996);
or U6154 (N_6154,N_5758,N_5808);
and U6155 (N_6155,N_5757,N_5999);
xor U6156 (N_6156,N_5792,N_5812);
xnor U6157 (N_6157,N_5973,N_5859);
nand U6158 (N_6158,N_5788,N_5805);
nor U6159 (N_6159,N_5936,N_5856);
nand U6160 (N_6160,N_5933,N_5764);
nand U6161 (N_6161,N_5782,N_5828);
nand U6162 (N_6162,N_5931,N_5752);
nor U6163 (N_6163,N_5871,N_5775);
nor U6164 (N_6164,N_5849,N_5806);
and U6165 (N_6165,N_5776,N_5854);
xnor U6166 (N_6166,N_5992,N_5993);
and U6167 (N_6167,N_5843,N_5923);
and U6168 (N_6168,N_5947,N_5776);
xnor U6169 (N_6169,N_5786,N_5918);
or U6170 (N_6170,N_5840,N_5907);
or U6171 (N_6171,N_5868,N_5805);
and U6172 (N_6172,N_5817,N_5848);
xor U6173 (N_6173,N_5951,N_5804);
and U6174 (N_6174,N_5934,N_5921);
or U6175 (N_6175,N_5853,N_5938);
nand U6176 (N_6176,N_5797,N_5936);
and U6177 (N_6177,N_5909,N_5997);
nand U6178 (N_6178,N_5989,N_5770);
xnor U6179 (N_6179,N_5916,N_5951);
nand U6180 (N_6180,N_5836,N_5982);
nor U6181 (N_6181,N_5904,N_5781);
or U6182 (N_6182,N_5847,N_5903);
or U6183 (N_6183,N_5811,N_5934);
nand U6184 (N_6184,N_5919,N_5917);
or U6185 (N_6185,N_5913,N_5798);
and U6186 (N_6186,N_5890,N_5759);
nand U6187 (N_6187,N_5929,N_5847);
nand U6188 (N_6188,N_5801,N_5990);
and U6189 (N_6189,N_5898,N_5920);
nor U6190 (N_6190,N_5813,N_5893);
nand U6191 (N_6191,N_5865,N_5872);
and U6192 (N_6192,N_5920,N_5844);
nand U6193 (N_6193,N_5927,N_5838);
nand U6194 (N_6194,N_5759,N_5840);
nor U6195 (N_6195,N_5897,N_5755);
or U6196 (N_6196,N_5910,N_5906);
xnor U6197 (N_6197,N_5960,N_5910);
or U6198 (N_6198,N_5786,N_5905);
xnor U6199 (N_6199,N_5999,N_5893);
xnor U6200 (N_6200,N_5826,N_5920);
and U6201 (N_6201,N_5779,N_5952);
nor U6202 (N_6202,N_5953,N_5751);
nor U6203 (N_6203,N_5819,N_5856);
and U6204 (N_6204,N_5955,N_5791);
nor U6205 (N_6205,N_5860,N_5822);
or U6206 (N_6206,N_5997,N_5949);
nor U6207 (N_6207,N_5856,N_5913);
xnor U6208 (N_6208,N_5782,N_5951);
nand U6209 (N_6209,N_5823,N_5957);
nor U6210 (N_6210,N_5808,N_5958);
and U6211 (N_6211,N_5782,N_5950);
nor U6212 (N_6212,N_5909,N_5999);
and U6213 (N_6213,N_5955,N_5895);
or U6214 (N_6214,N_5949,N_5775);
nor U6215 (N_6215,N_5954,N_5878);
xor U6216 (N_6216,N_5862,N_5797);
xor U6217 (N_6217,N_5998,N_5794);
or U6218 (N_6218,N_5855,N_5785);
nand U6219 (N_6219,N_5832,N_5963);
nor U6220 (N_6220,N_5804,N_5947);
nand U6221 (N_6221,N_5786,N_5882);
or U6222 (N_6222,N_5915,N_5752);
nand U6223 (N_6223,N_5995,N_5920);
or U6224 (N_6224,N_5939,N_5884);
xnor U6225 (N_6225,N_5902,N_5912);
nand U6226 (N_6226,N_5947,N_5982);
or U6227 (N_6227,N_5887,N_5815);
or U6228 (N_6228,N_5892,N_5794);
xnor U6229 (N_6229,N_5956,N_5770);
nor U6230 (N_6230,N_5846,N_5823);
nand U6231 (N_6231,N_5881,N_5921);
nand U6232 (N_6232,N_5849,N_5949);
xnor U6233 (N_6233,N_5818,N_5809);
nand U6234 (N_6234,N_5915,N_5978);
xnor U6235 (N_6235,N_5959,N_5795);
or U6236 (N_6236,N_5921,N_5913);
nand U6237 (N_6237,N_5857,N_5939);
nand U6238 (N_6238,N_5768,N_5865);
xnor U6239 (N_6239,N_5774,N_5950);
or U6240 (N_6240,N_5903,N_5961);
nor U6241 (N_6241,N_5885,N_5811);
and U6242 (N_6242,N_5785,N_5762);
nand U6243 (N_6243,N_5781,N_5835);
nand U6244 (N_6244,N_5822,N_5790);
nand U6245 (N_6245,N_5775,N_5785);
nor U6246 (N_6246,N_5894,N_5856);
or U6247 (N_6247,N_5973,N_5783);
nor U6248 (N_6248,N_5966,N_5785);
or U6249 (N_6249,N_5762,N_5807);
nand U6250 (N_6250,N_6033,N_6143);
nand U6251 (N_6251,N_6059,N_6189);
nand U6252 (N_6252,N_6003,N_6045);
and U6253 (N_6253,N_6244,N_6175);
xnor U6254 (N_6254,N_6069,N_6150);
and U6255 (N_6255,N_6158,N_6099);
nor U6256 (N_6256,N_6162,N_6134);
xnor U6257 (N_6257,N_6040,N_6064);
xor U6258 (N_6258,N_6186,N_6226);
and U6259 (N_6259,N_6246,N_6047);
nand U6260 (N_6260,N_6085,N_6007);
and U6261 (N_6261,N_6093,N_6027);
nand U6262 (N_6262,N_6185,N_6001);
or U6263 (N_6263,N_6243,N_6133);
nor U6264 (N_6264,N_6196,N_6234);
or U6265 (N_6265,N_6044,N_6124);
or U6266 (N_6266,N_6160,N_6097);
or U6267 (N_6267,N_6023,N_6213);
nand U6268 (N_6268,N_6232,N_6063);
nand U6269 (N_6269,N_6238,N_6089);
and U6270 (N_6270,N_6177,N_6173);
nor U6271 (N_6271,N_6168,N_6169);
or U6272 (N_6272,N_6154,N_6030);
or U6273 (N_6273,N_6037,N_6049);
or U6274 (N_6274,N_6181,N_6114);
nand U6275 (N_6275,N_6212,N_6237);
or U6276 (N_6276,N_6245,N_6071);
or U6277 (N_6277,N_6151,N_6068);
nor U6278 (N_6278,N_6078,N_6241);
xnor U6279 (N_6279,N_6225,N_6176);
and U6280 (N_6280,N_6190,N_6054);
nand U6281 (N_6281,N_6077,N_6102);
or U6282 (N_6282,N_6180,N_6012);
xor U6283 (N_6283,N_6005,N_6022);
nor U6284 (N_6284,N_6126,N_6062);
nor U6285 (N_6285,N_6018,N_6248);
nor U6286 (N_6286,N_6163,N_6046);
and U6287 (N_6287,N_6067,N_6026);
or U6288 (N_6288,N_6110,N_6210);
or U6289 (N_6289,N_6036,N_6032);
xnor U6290 (N_6290,N_6011,N_6056);
xnor U6291 (N_6291,N_6184,N_6136);
xor U6292 (N_6292,N_6187,N_6205);
xor U6293 (N_6293,N_6122,N_6132);
xnor U6294 (N_6294,N_6195,N_6209);
or U6295 (N_6295,N_6082,N_6129);
nor U6296 (N_6296,N_6020,N_6161);
nor U6297 (N_6297,N_6025,N_6084);
nor U6298 (N_6298,N_6021,N_6038);
xor U6299 (N_6299,N_6066,N_6247);
and U6300 (N_6300,N_6029,N_6142);
nor U6301 (N_6301,N_6157,N_6172);
and U6302 (N_6302,N_6174,N_6211);
nand U6303 (N_6303,N_6206,N_6095);
nor U6304 (N_6304,N_6140,N_6204);
xor U6305 (N_6305,N_6115,N_6164);
and U6306 (N_6306,N_6149,N_6106);
and U6307 (N_6307,N_6188,N_6017);
nand U6308 (N_6308,N_6070,N_6087);
nand U6309 (N_6309,N_6167,N_6192);
and U6310 (N_6310,N_6166,N_6178);
or U6311 (N_6311,N_6222,N_6135);
nand U6312 (N_6312,N_6165,N_6112);
xnor U6313 (N_6313,N_6083,N_6145);
or U6314 (N_6314,N_6052,N_6117);
xnor U6315 (N_6315,N_6235,N_6239);
nand U6316 (N_6316,N_6220,N_6240);
nor U6317 (N_6317,N_6197,N_6128);
and U6318 (N_6318,N_6050,N_6219);
nand U6319 (N_6319,N_6016,N_6086);
and U6320 (N_6320,N_6091,N_6061);
or U6321 (N_6321,N_6221,N_6171);
or U6322 (N_6322,N_6002,N_6101);
nand U6323 (N_6323,N_6155,N_6242);
nand U6324 (N_6324,N_6073,N_6138);
and U6325 (N_6325,N_6193,N_6121);
or U6326 (N_6326,N_6113,N_6207);
and U6327 (N_6327,N_6053,N_6229);
and U6328 (N_6328,N_6183,N_6152);
nor U6329 (N_6329,N_6014,N_6105);
nor U6330 (N_6330,N_6060,N_6081);
and U6331 (N_6331,N_6182,N_6057);
nand U6332 (N_6332,N_6228,N_6043);
nor U6333 (N_6333,N_6146,N_6088);
nand U6334 (N_6334,N_6058,N_6216);
xnor U6335 (N_6335,N_6015,N_6109);
or U6336 (N_6336,N_6092,N_6004);
nand U6337 (N_6337,N_6094,N_6074);
nand U6338 (N_6338,N_6075,N_6006);
and U6339 (N_6339,N_6199,N_6233);
and U6340 (N_6340,N_6035,N_6125);
nor U6341 (N_6341,N_6130,N_6179);
nor U6342 (N_6342,N_6039,N_6139);
nand U6343 (N_6343,N_6153,N_6103);
nand U6344 (N_6344,N_6065,N_6076);
xnor U6345 (N_6345,N_6100,N_6208);
and U6346 (N_6346,N_6227,N_6107);
or U6347 (N_6347,N_6079,N_6214);
xor U6348 (N_6348,N_6108,N_6137);
or U6349 (N_6349,N_6170,N_6072);
and U6350 (N_6350,N_6198,N_6042);
and U6351 (N_6351,N_6236,N_6019);
or U6352 (N_6352,N_6201,N_6148);
xnor U6353 (N_6353,N_6034,N_6203);
or U6354 (N_6354,N_6010,N_6024);
or U6355 (N_6355,N_6191,N_6123);
xor U6356 (N_6356,N_6008,N_6230);
or U6357 (N_6357,N_6202,N_6249);
or U6358 (N_6358,N_6223,N_6055);
and U6359 (N_6359,N_6048,N_6200);
or U6360 (N_6360,N_6120,N_6156);
nor U6361 (N_6361,N_6051,N_6111);
nand U6362 (N_6362,N_6080,N_6119);
and U6363 (N_6363,N_6141,N_6098);
or U6364 (N_6364,N_6159,N_6147);
and U6365 (N_6365,N_6224,N_6217);
and U6366 (N_6366,N_6104,N_6218);
nor U6367 (N_6367,N_6028,N_6231);
xnor U6368 (N_6368,N_6009,N_6013);
or U6369 (N_6369,N_6127,N_6031);
or U6370 (N_6370,N_6215,N_6096);
or U6371 (N_6371,N_6041,N_6118);
or U6372 (N_6372,N_6116,N_6144);
nand U6373 (N_6373,N_6131,N_6090);
nand U6374 (N_6374,N_6000,N_6194);
xnor U6375 (N_6375,N_6245,N_6240);
and U6376 (N_6376,N_6031,N_6065);
or U6377 (N_6377,N_6185,N_6082);
or U6378 (N_6378,N_6233,N_6052);
or U6379 (N_6379,N_6105,N_6191);
nor U6380 (N_6380,N_6127,N_6107);
nor U6381 (N_6381,N_6227,N_6068);
nor U6382 (N_6382,N_6233,N_6085);
xnor U6383 (N_6383,N_6241,N_6172);
xnor U6384 (N_6384,N_6002,N_6230);
nor U6385 (N_6385,N_6006,N_6112);
xnor U6386 (N_6386,N_6000,N_6123);
and U6387 (N_6387,N_6209,N_6108);
nand U6388 (N_6388,N_6184,N_6241);
nor U6389 (N_6389,N_6022,N_6213);
or U6390 (N_6390,N_6195,N_6093);
and U6391 (N_6391,N_6025,N_6061);
nand U6392 (N_6392,N_6210,N_6134);
nor U6393 (N_6393,N_6015,N_6158);
or U6394 (N_6394,N_6157,N_6021);
nand U6395 (N_6395,N_6231,N_6185);
xor U6396 (N_6396,N_6230,N_6153);
nand U6397 (N_6397,N_6233,N_6081);
xor U6398 (N_6398,N_6168,N_6230);
and U6399 (N_6399,N_6125,N_6208);
or U6400 (N_6400,N_6059,N_6212);
xnor U6401 (N_6401,N_6153,N_6151);
and U6402 (N_6402,N_6002,N_6130);
nand U6403 (N_6403,N_6073,N_6095);
nor U6404 (N_6404,N_6056,N_6033);
and U6405 (N_6405,N_6079,N_6072);
nor U6406 (N_6406,N_6073,N_6084);
nor U6407 (N_6407,N_6185,N_6049);
xnor U6408 (N_6408,N_6056,N_6180);
nand U6409 (N_6409,N_6096,N_6247);
nor U6410 (N_6410,N_6092,N_6174);
and U6411 (N_6411,N_6166,N_6105);
and U6412 (N_6412,N_6097,N_6167);
or U6413 (N_6413,N_6198,N_6111);
nor U6414 (N_6414,N_6144,N_6149);
and U6415 (N_6415,N_6080,N_6059);
xnor U6416 (N_6416,N_6015,N_6132);
nor U6417 (N_6417,N_6088,N_6103);
nor U6418 (N_6418,N_6031,N_6207);
nand U6419 (N_6419,N_6162,N_6167);
nor U6420 (N_6420,N_6173,N_6044);
or U6421 (N_6421,N_6190,N_6143);
xnor U6422 (N_6422,N_6141,N_6033);
nand U6423 (N_6423,N_6156,N_6044);
and U6424 (N_6424,N_6062,N_6156);
or U6425 (N_6425,N_6222,N_6141);
or U6426 (N_6426,N_6134,N_6094);
or U6427 (N_6427,N_6208,N_6221);
xor U6428 (N_6428,N_6081,N_6185);
nor U6429 (N_6429,N_6135,N_6032);
or U6430 (N_6430,N_6010,N_6033);
or U6431 (N_6431,N_6173,N_6009);
nor U6432 (N_6432,N_6175,N_6208);
xnor U6433 (N_6433,N_6031,N_6074);
and U6434 (N_6434,N_6130,N_6135);
and U6435 (N_6435,N_6199,N_6181);
xnor U6436 (N_6436,N_6160,N_6060);
nand U6437 (N_6437,N_6081,N_6193);
nand U6438 (N_6438,N_6085,N_6232);
nor U6439 (N_6439,N_6211,N_6044);
or U6440 (N_6440,N_6234,N_6195);
or U6441 (N_6441,N_6203,N_6225);
nor U6442 (N_6442,N_6178,N_6180);
nor U6443 (N_6443,N_6206,N_6015);
nand U6444 (N_6444,N_6171,N_6156);
and U6445 (N_6445,N_6052,N_6150);
or U6446 (N_6446,N_6148,N_6184);
nor U6447 (N_6447,N_6048,N_6129);
or U6448 (N_6448,N_6128,N_6101);
and U6449 (N_6449,N_6189,N_6120);
or U6450 (N_6450,N_6044,N_6206);
and U6451 (N_6451,N_6052,N_6116);
nand U6452 (N_6452,N_6071,N_6248);
nand U6453 (N_6453,N_6227,N_6018);
nor U6454 (N_6454,N_6034,N_6145);
or U6455 (N_6455,N_6162,N_6211);
nand U6456 (N_6456,N_6133,N_6058);
or U6457 (N_6457,N_6062,N_6046);
and U6458 (N_6458,N_6125,N_6199);
and U6459 (N_6459,N_6123,N_6243);
and U6460 (N_6460,N_6014,N_6135);
xor U6461 (N_6461,N_6171,N_6177);
xor U6462 (N_6462,N_6195,N_6235);
and U6463 (N_6463,N_6008,N_6171);
and U6464 (N_6464,N_6128,N_6239);
xnor U6465 (N_6465,N_6097,N_6037);
nand U6466 (N_6466,N_6212,N_6095);
nor U6467 (N_6467,N_6139,N_6161);
nor U6468 (N_6468,N_6182,N_6079);
and U6469 (N_6469,N_6049,N_6159);
nand U6470 (N_6470,N_6135,N_6249);
nand U6471 (N_6471,N_6181,N_6016);
xnor U6472 (N_6472,N_6120,N_6058);
or U6473 (N_6473,N_6192,N_6084);
nand U6474 (N_6474,N_6006,N_6073);
nand U6475 (N_6475,N_6073,N_6225);
and U6476 (N_6476,N_6115,N_6204);
nor U6477 (N_6477,N_6103,N_6112);
nand U6478 (N_6478,N_6174,N_6171);
nand U6479 (N_6479,N_6153,N_6055);
or U6480 (N_6480,N_6075,N_6079);
nand U6481 (N_6481,N_6088,N_6129);
and U6482 (N_6482,N_6205,N_6222);
or U6483 (N_6483,N_6174,N_6120);
nor U6484 (N_6484,N_6211,N_6134);
and U6485 (N_6485,N_6166,N_6019);
nor U6486 (N_6486,N_6103,N_6119);
or U6487 (N_6487,N_6134,N_6006);
nand U6488 (N_6488,N_6156,N_6175);
xor U6489 (N_6489,N_6021,N_6126);
or U6490 (N_6490,N_6195,N_6064);
nand U6491 (N_6491,N_6003,N_6168);
nand U6492 (N_6492,N_6153,N_6122);
and U6493 (N_6493,N_6083,N_6220);
nand U6494 (N_6494,N_6083,N_6016);
nor U6495 (N_6495,N_6055,N_6133);
xor U6496 (N_6496,N_6140,N_6172);
nand U6497 (N_6497,N_6218,N_6171);
and U6498 (N_6498,N_6185,N_6184);
nor U6499 (N_6499,N_6112,N_6003);
xor U6500 (N_6500,N_6493,N_6483);
or U6501 (N_6501,N_6388,N_6251);
and U6502 (N_6502,N_6426,N_6357);
xor U6503 (N_6503,N_6329,N_6273);
nor U6504 (N_6504,N_6438,N_6334);
or U6505 (N_6505,N_6416,N_6284);
or U6506 (N_6506,N_6371,N_6456);
nand U6507 (N_6507,N_6451,N_6318);
or U6508 (N_6508,N_6420,N_6260);
nor U6509 (N_6509,N_6399,N_6335);
or U6510 (N_6510,N_6321,N_6323);
nand U6511 (N_6511,N_6348,N_6269);
or U6512 (N_6512,N_6376,N_6356);
or U6513 (N_6513,N_6315,N_6464);
xnor U6514 (N_6514,N_6276,N_6496);
and U6515 (N_6515,N_6250,N_6398);
xnor U6516 (N_6516,N_6463,N_6444);
and U6517 (N_6517,N_6450,N_6333);
xor U6518 (N_6518,N_6401,N_6274);
nor U6519 (N_6519,N_6270,N_6395);
and U6520 (N_6520,N_6405,N_6308);
nand U6521 (N_6521,N_6253,N_6382);
nor U6522 (N_6522,N_6298,N_6462);
xor U6523 (N_6523,N_6494,N_6380);
nor U6524 (N_6524,N_6268,N_6312);
and U6525 (N_6525,N_6411,N_6425);
or U6526 (N_6526,N_6294,N_6375);
xnor U6527 (N_6527,N_6275,N_6351);
and U6528 (N_6528,N_6455,N_6467);
xnor U6529 (N_6529,N_6349,N_6396);
nand U6530 (N_6530,N_6277,N_6385);
nor U6531 (N_6531,N_6272,N_6449);
nor U6532 (N_6532,N_6364,N_6341);
xor U6533 (N_6533,N_6254,N_6390);
and U6534 (N_6534,N_6470,N_6338);
nand U6535 (N_6535,N_6422,N_6305);
nor U6536 (N_6536,N_6384,N_6337);
nand U6537 (N_6537,N_6471,N_6497);
or U6538 (N_6538,N_6423,N_6287);
and U6539 (N_6539,N_6336,N_6289);
nor U6540 (N_6540,N_6307,N_6407);
nand U6541 (N_6541,N_6309,N_6292);
or U6542 (N_6542,N_6419,N_6295);
nor U6543 (N_6543,N_6358,N_6263);
nand U6544 (N_6544,N_6331,N_6316);
nor U6545 (N_6545,N_6352,N_6415);
nand U6546 (N_6546,N_6327,N_6387);
nor U6547 (N_6547,N_6368,N_6320);
nand U6548 (N_6548,N_6354,N_6491);
nor U6549 (N_6549,N_6343,N_6266);
nor U6550 (N_6550,N_6432,N_6412);
or U6551 (N_6551,N_6381,N_6466);
nor U6552 (N_6552,N_6428,N_6252);
nor U6553 (N_6553,N_6486,N_6404);
and U6554 (N_6554,N_6392,N_6296);
nor U6555 (N_6555,N_6319,N_6402);
and U6556 (N_6556,N_6437,N_6469);
xor U6557 (N_6557,N_6445,N_6436);
nand U6558 (N_6558,N_6383,N_6324);
nand U6559 (N_6559,N_6300,N_6353);
nor U6560 (N_6560,N_6408,N_6282);
nor U6561 (N_6561,N_6286,N_6468);
xor U6562 (N_6562,N_6424,N_6281);
nand U6563 (N_6563,N_6421,N_6325);
nand U6564 (N_6564,N_6367,N_6256);
and U6565 (N_6565,N_6394,N_6498);
nand U6566 (N_6566,N_6413,N_6257);
nor U6567 (N_6567,N_6359,N_6283);
or U6568 (N_6568,N_6365,N_6389);
nor U6569 (N_6569,N_6363,N_6397);
nor U6570 (N_6570,N_6410,N_6439);
and U6571 (N_6571,N_6303,N_6453);
nand U6572 (N_6572,N_6480,N_6313);
nor U6573 (N_6573,N_6372,N_6434);
nand U6574 (N_6574,N_6442,N_6339);
xnor U6575 (N_6575,N_6291,N_6360);
nand U6576 (N_6576,N_6386,N_6379);
xor U6577 (N_6577,N_6447,N_6278);
and U6578 (N_6578,N_6374,N_6265);
and U6579 (N_6579,N_6409,N_6490);
or U6580 (N_6580,N_6403,N_6479);
nand U6581 (N_6581,N_6328,N_6264);
nor U6582 (N_6582,N_6350,N_6433);
nor U6583 (N_6583,N_6435,N_6458);
or U6584 (N_6584,N_6267,N_6474);
nor U6585 (N_6585,N_6346,N_6452);
nand U6586 (N_6586,N_6487,N_6448);
nor U6587 (N_6587,N_6484,N_6393);
or U6588 (N_6588,N_6285,N_6400);
nand U6589 (N_6589,N_6262,N_6340);
or U6590 (N_6590,N_6472,N_6482);
nor U6591 (N_6591,N_6417,N_6418);
nand U6592 (N_6592,N_6299,N_6304);
xor U6593 (N_6593,N_6377,N_6332);
nand U6594 (N_6594,N_6306,N_6443);
and U6595 (N_6595,N_6475,N_6427);
or U6596 (N_6596,N_6414,N_6440);
or U6597 (N_6597,N_6344,N_6481);
and U6598 (N_6598,N_6342,N_6280);
xnor U6599 (N_6599,N_6326,N_6355);
nand U6600 (N_6600,N_6255,N_6293);
xnor U6601 (N_6601,N_6391,N_6288);
nor U6602 (N_6602,N_6477,N_6362);
nor U6603 (N_6603,N_6495,N_6366);
and U6604 (N_6604,N_6431,N_6489);
xnor U6605 (N_6605,N_6406,N_6485);
and U6606 (N_6606,N_6492,N_6441);
nor U6607 (N_6607,N_6311,N_6258);
xnor U6608 (N_6608,N_6459,N_6369);
and U6609 (N_6609,N_6290,N_6301);
xnor U6610 (N_6610,N_6461,N_6454);
or U6611 (N_6611,N_6361,N_6271);
xnor U6612 (N_6612,N_6279,N_6370);
and U6613 (N_6613,N_6345,N_6499);
or U6614 (N_6614,N_6457,N_6460);
and U6615 (N_6615,N_6322,N_6330);
nor U6616 (N_6616,N_6261,N_6378);
and U6617 (N_6617,N_6465,N_6429);
and U6618 (N_6618,N_6488,N_6430);
and U6619 (N_6619,N_6259,N_6473);
or U6620 (N_6620,N_6446,N_6302);
and U6621 (N_6621,N_6310,N_6317);
and U6622 (N_6622,N_6347,N_6297);
and U6623 (N_6623,N_6476,N_6478);
xnor U6624 (N_6624,N_6314,N_6373);
nor U6625 (N_6625,N_6271,N_6487);
nor U6626 (N_6626,N_6341,N_6312);
nand U6627 (N_6627,N_6351,N_6288);
nor U6628 (N_6628,N_6399,N_6355);
and U6629 (N_6629,N_6438,N_6403);
xnor U6630 (N_6630,N_6453,N_6454);
and U6631 (N_6631,N_6375,N_6442);
nor U6632 (N_6632,N_6325,N_6439);
or U6633 (N_6633,N_6272,N_6393);
nor U6634 (N_6634,N_6252,N_6274);
and U6635 (N_6635,N_6384,N_6250);
nor U6636 (N_6636,N_6405,N_6297);
xor U6637 (N_6637,N_6271,N_6404);
and U6638 (N_6638,N_6343,N_6384);
nand U6639 (N_6639,N_6260,N_6465);
nand U6640 (N_6640,N_6266,N_6420);
and U6641 (N_6641,N_6483,N_6280);
xor U6642 (N_6642,N_6478,N_6276);
or U6643 (N_6643,N_6453,N_6355);
or U6644 (N_6644,N_6436,N_6390);
xnor U6645 (N_6645,N_6293,N_6313);
nand U6646 (N_6646,N_6281,N_6343);
nor U6647 (N_6647,N_6338,N_6297);
nand U6648 (N_6648,N_6285,N_6421);
xnor U6649 (N_6649,N_6332,N_6366);
nor U6650 (N_6650,N_6317,N_6270);
or U6651 (N_6651,N_6349,N_6392);
xor U6652 (N_6652,N_6377,N_6382);
nor U6653 (N_6653,N_6470,N_6250);
nand U6654 (N_6654,N_6404,N_6327);
xor U6655 (N_6655,N_6282,N_6285);
xor U6656 (N_6656,N_6348,N_6437);
nand U6657 (N_6657,N_6256,N_6302);
nor U6658 (N_6658,N_6365,N_6252);
xnor U6659 (N_6659,N_6460,N_6477);
xor U6660 (N_6660,N_6261,N_6298);
nand U6661 (N_6661,N_6478,N_6439);
and U6662 (N_6662,N_6351,N_6274);
nor U6663 (N_6663,N_6397,N_6482);
nand U6664 (N_6664,N_6424,N_6291);
or U6665 (N_6665,N_6445,N_6373);
and U6666 (N_6666,N_6343,N_6328);
xnor U6667 (N_6667,N_6377,N_6277);
nor U6668 (N_6668,N_6404,N_6287);
and U6669 (N_6669,N_6472,N_6414);
and U6670 (N_6670,N_6444,N_6283);
nand U6671 (N_6671,N_6339,N_6421);
nand U6672 (N_6672,N_6350,N_6377);
nor U6673 (N_6673,N_6281,N_6336);
nand U6674 (N_6674,N_6390,N_6400);
nor U6675 (N_6675,N_6392,N_6391);
or U6676 (N_6676,N_6474,N_6439);
and U6677 (N_6677,N_6415,N_6333);
or U6678 (N_6678,N_6269,N_6414);
and U6679 (N_6679,N_6346,N_6371);
xnor U6680 (N_6680,N_6334,N_6324);
and U6681 (N_6681,N_6491,N_6429);
nand U6682 (N_6682,N_6349,N_6256);
xnor U6683 (N_6683,N_6280,N_6348);
and U6684 (N_6684,N_6495,N_6250);
or U6685 (N_6685,N_6496,N_6360);
xnor U6686 (N_6686,N_6379,N_6275);
or U6687 (N_6687,N_6426,N_6279);
or U6688 (N_6688,N_6416,N_6358);
nor U6689 (N_6689,N_6486,N_6252);
xnor U6690 (N_6690,N_6396,N_6375);
xnor U6691 (N_6691,N_6412,N_6262);
nor U6692 (N_6692,N_6408,N_6385);
or U6693 (N_6693,N_6427,N_6496);
nand U6694 (N_6694,N_6378,N_6373);
nand U6695 (N_6695,N_6278,N_6431);
or U6696 (N_6696,N_6432,N_6274);
and U6697 (N_6697,N_6257,N_6412);
and U6698 (N_6698,N_6489,N_6262);
and U6699 (N_6699,N_6397,N_6359);
and U6700 (N_6700,N_6385,N_6276);
nand U6701 (N_6701,N_6312,N_6253);
xor U6702 (N_6702,N_6344,N_6493);
xnor U6703 (N_6703,N_6390,N_6395);
or U6704 (N_6704,N_6381,N_6445);
nor U6705 (N_6705,N_6303,N_6407);
nor U6706 (N_6706,N_6275,N_6454);
xor U6707 (N_6707,N_6327,N_6496);
or U6708 (N_6708,N_6304,N_6381);
xnor U6709 (N_6709,N_6406,N_6408);
and U6710 (N_6710,N_6370,N_6451);
xor U6711 (N_6711,N_6349,N_6328);
and U6712 (N_6712,N_6486,N_6344);
nor U6713 (N_6713,N_6482,N_6403);
xor U6714 (N_6714,N_6433,N_6376);
xnor U6715 (N_6715,N_6414,N_6451);
nand U6716 (N_6716,N_6342,N_6287);
nand U6717 (N_6717,N_6483,N_6308);
nand U6718 (N_6718,N_6420,N_6348);
nand U6719 (N_6719,N_6270,N_6288);
nor U6720 (N_6720,N_6371,N_6417);
xor U6721 (N_6721,N_6432,N_6442);
nor U6722 (N_6722,N_6324,N_6270);
and U6723 (N_6723,N_6327,N_6350);
xnor U6724 (N_6724,N_6473,N_6470);
or U6725 (N_6725,N_6347,N_6479);
nand U6726 (N_6726,N_6332,N_6326);
nor U6727 (N_6727,N_6304,N_6398);
nand U6728 (N_6728,N_6461,N_6269);
xnor U6729 (N_6729,N_6449,N_6390);
or U6730 (N_6730,N_6309,N_6362);
nor U6731 (N_6731,N_6256,N_6310);
and U6732 (N_6732,N_6473,N_6328);
xnor U6733 (N_6733,N_6346,N_6310);
or U6734 (N_6734,N_6274,N_6377);
nor U6735 (N_6735,N_6457,N_6364);
or U6736 (N_6736,N_6420,N_6352);
and U6737 (N_6737,N_6311,N_6254);
nor U6738 (N_6738,N_6494,N_6441);
nor U6739 (N_6739,N_6325,N_6365);
nand U6740 (N_6740,N_6277,N_6300);
and U6741 (N_6741,N_6423,N_6456);
nor U6742 (N_6742,N_6357,N_6279);
nand U6743 (N_6743,N_6297,N_6429);
and U6744 (N_6744,N_6342,N_6292);
or U6745 (N_6745,N_6304,N_6393);
nand U6746 (N_6746,N_6341,N_6338);
xnor U6747 (N_6747,N_6347,N_6408);
xor U6748 (N_6748,N_6415,N_6304);
xnor U6749 (N_6749,N_6479,N_6396);
nor U6750 (N_6750,N_6658,N_6674);
or U6751 (N_6751,N_6609,N_6745);
or U6752 (N_6752,N_6613,N_6727);
or U6753 (N_6753,N_6662,N_6749);
nand U6754 (N_6754,N_6567,N_6734);
or U6755 (N_6755,N_6502,N_6612);
and U6756 (N_6756,N_6530,N_6523);
nand U6757 (N_6757,N_6591,N_6542);
or U6758 (N_6758,N_6512,N_6554);
xor U6759 (N_6759,N_6677,N_6563);
and U6760 (N_6760,N_6635,N_6521);
or U6761 (N_6761,N_6735,N_6743);
xnor U6762 (N_6762,N_6684,N_6701);
xor U6763 (N_6763,N_6644,N_6723);
nand U6764 (N_6764,N_6673,N_6524);
xnor U6765 (N_6765,N_6671,N_6592);
nor U6766 (N_6766,N_6503,N_6648);
nand U6767 (N_6767,N_6670,N_6652);
nand U6768 (N_6768,N_6509,N_6620);
nor U6769 (N_6769,N_6600,N_6666);
nor U6770 (N_6770,N_6585,N_6514);
and U6771 (N_6771,N_6656,N_6541);
xor U6772 (N_6772,N_6570,N_6551);
and U6773 (N_6773,N_6692,N_6624);
or U6774 (N_6774,N_6716,N_6707);
xor U6775 (N_6775,N_6578,N_6690);
nor U6776 (N_6776,N_6534,N_6619);
or U6777 (N_6777,N_6614,N_6737);
nand U6778 (N_6778,N_6519,N_6650);
nor U6779 (N_6779,N_6621,N_6558);
and U6780 (N_6780,N_6522,N_6576);
xor U6781 (N_6781,N_6729,N_6746);
nand U6782 (N_6782,N_6642,N_6575);
nand U6783 (N_6783,N_6733,N_6546);
and U6784 (N_6784,N_6748,N_6640);
xor U6785 (N_6785,N_6557,N_6504);
and U6786 (N_6786,N_6643,N_6685);
nor U6787 (N_6787,N_6728,N_6708);
nand U6788 (N_6788,N_6604,N_6527);
and U6789 (N_6789,N_6518,N_6550);
or U6790 (N_6790,N_6501,N_6583);
or U6791 (N_6791,N_6726,N_6584);
and U6792 (N_6792,N_6549,N_6725);
xnor U6793 (N_6793,N_6711,N_6694);
nand U6794 (N_6794,N_6632,N_6535);
or U6795 (N_6795,N_6599,N_6507);
or U6796 (N_6796,N_6704,N_6722);
and U6797 (N_6797,N_6532,N_6589);
nand U6798 (N_6798,N_6568,N_6742);
or U6799 (N_6799,N_6700,N_6696);
xor U6800 (N_6800,N_6681,N_6705);
nand U6801 (N_6801,N_6718,N_6610);
nor U6802 (N_6802,N_6622,N_6676);
nand U6803 (N_6803,N_6608,N_6672);
xnor U6804 (N_6804,N_6714,N_6616);
nand U6805 (N_6805,N_6679,N_6543);
nor U6806 (N_6806,N_6528,N_6577);
and U6807 (N_6807,N_6628,N_6669);
nor U6808 (N_6808,N_6697,N_6544);
nand U6809 (N_6809,N_6686,N_6590);
nor U6810 (N_6810,N_6598,N_6715);
or U6811 (N_6811,N_6653,N_6562);
nand U6812 (N_6812,N_6515,N_6525);
nand U6813 (N_6813,N_6517,N_6680);
nand U6814 (N_6814,N_6626,N_6637);
and U6815 (N_6815,N_6538,N_6654);
nor U6816 (N_6816,N_6691,N_6675);
or U6817 (N_6817,N_6688,N_6655);
and U6818 (N_6818,N_6537,N_6645);
nor U6819 (N_6819,N_6573,N_6665);
nand U6820 (N_6820,N_6566,N_6601);
nor U6821 (N_6821,N_6533,N_6529);
xnor U6822 (N_6822,N_6661,N_6500);
nor U6823 (N_6823,N_6564,N_6699);
xnor U6824 (N_6824,N_6739,N_6617);
and U6825 (N_6825,N_6709,N_6513);
or U6826 (N_6826,N_6683,N_6582);
xor U6827 (N_6827,N_6702,N_6615);
and U6828 (N_6828,N_6607,N_6630);
and U6829 (N_6829,N_6717,N_6510);
or U6830 (N_6830,N_6603,N_6580);
nand U6831 (N_6831,N_6657,N_6703);
and U6832 (N_6832,N_6724,N_6596);
xnor U6833 (N_6833,N_6730,N_6663);
and U6834 (N_6834,N_6627,N_6553);
nand U6835 (N_6835,N_6719,N_6581);
xnor U6836 (N_6836,N_6594,N_6526);
nor U6837 (N_6837,N_6516,N_6511);
nand U6838 (N_6838,N_6682,N_6741);
nor U6839 (N_6839,N_6559,N_6588);
nand U6840 (N_6840,N_6713,N_6740);
nand U6841 (N_6841,N_6540,N_6605);
nor U6842 (N_6842,N_6625,N_6721);
and U6843 (N_6843,N_6660,N_6667);
nand U6844 (N_6844,N_6695,N_6579);
nand U6845 (N_6845,N_6687,N_6539);
and U6846 (N_6846,N_6641,N_6506);
nand U6847 (N_6847,N_6561,N_6611);
or U6848 (N_6848,N_6651,N_6569);
xor U6849 (N_6849,N_6623,N_6548);
xor U6850 (N_6850,N_6706,N_6629);
nand U6851 (N_6851,N_6587,N_6636);
and U6852 (N_6852,N_6536,N_6634);
xor U6853 (N_6853,N_6572,N_6593);
or U6854 (N_6854,N_6602,N_6678);
nand U6855 (N_6855,N_6712,N_6520);
and U6856 (N_6856,N_6571,N_6606);
xor U6857 (N_6857,N_6552,N_6586);
and U6858 (N_6858,N_6545,N_6647);
nor U6859 (N_6859,N_6618,N_6597);
or U6860 (N_6860,N_6595,N_6531);
or U6861 (N_6861,N_6574,N_6633);
nor U6862 (N_6862,N_6555,N_6639);
and U6863 (N_6863,N_6732,N_6547);
nand U6864 (N_6864,N_6565,N_6668);
xor U6865 (N_6865,N_6556,N_6560);
and U6866 (N_6866,N_6738,N_6744);
or U6867 (N_6867,N_6720,N_6508);
and U6868 (N_6868,N_6736,N_6731);
and U6869 (N_6869,N_6710,N_6646);
and U6870 (N_6870,N_6631,N_6698);
or U6871 (N_6871,N_6664,N_6649);
and U6872 (N_6872,N_6659,N_6693);
or U6873 (N_6873,N_6747,N_6505);
and U6874 (N_6874,N_6689,N_6638);
and U6875 (N_6875,N_6749,N_6591);
nor U6876 (N_6876,N_6695,N_6742);
or U6877 (N_6877,N_6668,N_6655);
nor U6878 (N_6878,N_6682,N_6513);
and U6879 (N_6879,N_6639,N_6729);
nand U6880 (N_6880,N_6628,N_6551);
nand U6881 (N_6881,N_6557,N_6606);
and U6882 (N_6882,N_6669,N_6661);
or U6883 (N_6883,N_6511,N_6717);
or U6884 (N_6884,N_6645,N_6717);
or U6885 (N_6885,N_6580,N_6723);
xnor U6886 (N_6886,N_6712,N_6562);
xor U6887 (N_6887,N_6578,N_6675);
xnor U6888 (N_6888,N_6532,N_6549);
xor U6889 (N_6889,N_6586,N_6696);
nand U6890 (N_6890,N_6588,N_6540);
nor U6891 (N_6891,N_6602,N_6605);
or U6892 (N_6892,N_6605,N_6519);
xnor U6893 (N_6893,N_6507,N_6500);
nor U6894 (N_6894,N_6522,N_6692);
nor U6895 (N_6895,N_6542,N_6553);
and U6896 (N_6896,N_6616,N_6617);
nand U6897 (N_6897,N_6536,N_6635);
nor U6898 (N_6898,N_6720,N_6684);
nor U6899 (N_6899,N_6531,N_6666);
or U6900 (N_6900,N_6716,N_6531);
and U6901 (N_6901,N_6569,N_6585);
nor U6902 (N_6902,N_6590,N_6613);
nor U6903 (N_6903,N_6576,N_6615);
nand U6904 (N_6904,N_6556,N_6539);
and U6905 (N_6905,N_6674,N_6664);
nor U6906 (N_6906,N_6697,N_6721);
xnor U6907 (N_6907,N_6741,N_6748);
or U6908 (N_6908,N_6554,N_6520);
and U6909 (N_6909,N_6573,N_6717);
nand U6910 (N_6910,N_6640,N_6535);
nand U6911 (N_6911,N_6613,N_6577);
nand U6912 (N_6912,N_6516,N_6602);
and U6913 (N_6913,N_6577,N_6605);
and U6914 (N_6914,N_6664,N_6519);
and U6915 (N_6915,N_6567,N_6548);
or U6916 (N_6916,N_6649,N_6744);
xor U6917 (N_6917,N_6576,N_6619);
nand U6918 (N_6918,N_6657,N_6511);
and U6919 (N_6919,N_6582,N_6744);
xnor U6920 (N_6920,N_6723,N_6542);
nor U6921 (N_6921,N_6516,N_6650);
nand U6922 (N_6922,N_6502,N_6736);
and U6923 (N_6923,N_6731,N_6522);
nand U6924 (N_6924,N_6670,N_6575);
and U6925 (N_6925,N_6710,N_6588);
and U6926 (N_6926,N_6734,N_6526);
or U6927 (N_6927,N_6583,N_6513);
nand U6928 (N_6928,N_6637,N_6733);
and U6929 (N_6929,N_6538,N_6603);
xnor U6930 (N_6930,N_6670,N_6503);
xnor U6931 (N_6931,N_6643,N_6555);
nand U6932 (N_6932,N_6593,N_6667);
xor U6933 (N_6933,N_6651,N_6686);
nand U6934 (N_6934,N_6640,N_6508);
nand U6935 (N_6935,N_6529,N_6560);
nor U6936 (N_6936,N_6595,N_6681);
nor U6937 (N_6937,N_6611,N_6726);
or U6938 (N_6938,N_6643,N_6566);
nand U6939 (N_6939,N_6633,N_6590);
and U6940 (N_6940,N_6548,N_6511);
nand U6941 (N_6941,N_6624,N_6701);
nand U6942 (N_6942,N_6524,N_6582);
xor U6943 (N_6943,N_6553,N_6576);
nor U6944 (N_6944,N_6642,N_6532);
nand U6945 (N_6945,N_6591,N_6702);
or U6946 (N_6946,N_6501,N_6670);
and U6947 (N_6947,N_6703,N_6550);
nand U6948 (N_6948,N_6598,N_6507);
nor U6949 (N_6949,N_6655,N_6600);
and U6950 (N_6950,N_6720,N_6687);
nand U6951 (N_6951,N_6689,N_6593);
and U6952 (N_6952,N_6590,N_6648);
nor U6953 (N_6953,N_6618,N_6552);
nor U6954 (N_6954,N_6540,N_6539);
xnor U6955 (N_6955,N_6625,N_6666);
xor U6956 (N_6956,N_6697,N_6560);
nor U6957 (N_6957,N_6623,N_6516);
nor U6958 (N_6958,N_6558,N_6664);
or U6959 (N_6959,N_6639,N_6690);
nand U6960 (N_6960,N_6664,N_6556);
xnor U6961 (N_6961,N_6510,N_6728);
and U6962 (N_6962,N_6609,N_6545);
and U6963 (N_6963,N_6707,N_6501);
or U6964 (N_6964,N_6668,N_6626);
or U6965 (N_6965,N_6582,N_6547);
or U6966 (N_6966,N_6619,N_6592);
or U6967 (N_6967,N_6608,N_6563);
or U6968 (N_6968,N_6558,N_6652);
nand U6969 (N_6969,N_6657,N_6595);
xor U6970 (N_6970,N_6525,N_6696);
nor U6971 (N_6971,N_6659,N_6643);
nor U6972 (N_6972,N_6713,N_6655);
and U6973 (N_6973,N_6694,N_6736);
and U6974 (N_6974,N_6543,N_6748);
or U6975 (N_6975,N_6614,N_6588);
nor U6976 (N_6976,N_6640,N_6679);
or U6977 (N_6977,N_6710,N_6644);
and U6978 (N_6978,N_6693,N_6573);
nor U6979 (N_6979,N_6741,N_6631);
nand U6980 (N_6980,N_6511,N_6566);
or U6981 (N_6981,N_6546,N_6716);
nand U6982 (N_6982,N_6571,N_6566);
nand U6983 (N_6983,N_6567,N_6630);
and U6984 (N_6984,N_6540,N_6644);
nand U6985 (N_6985,N_6547,N_6575);
and U6986 (N_6986,N_6537,N_6591);
nor U6987 (N_6987,N_6687,N_6620);
nor U6988 (N_6988,N_6649,N_6647);
nand U6989 (N_6989,N_6658,N_6618);
xor U6990 (N_6990,N_6634,N_6732);
xnor U6991 (N_6991,N_6593,N_6598);
or U6992 (N_6992,N_6540,N_6630);
and U6993 (N_6993,N_6717,N_6589);
nor U6994 (N_6994,N_6728,N_6744);
nor U6995 (N_6995,N_6611,N_6524);
or U6996 (N_6996,N_6622,N_6719);
or U6997 (N_6997,N_6739,N_6712);
or U6998 (N_6998,N_6741,N_6671);
and U6999 (N_6999,N_6709,N_6622);
nor U7000 (N_7000,N_6798,N_6785);
nand U7001 (N_7001,N_6793,N_6811);
xor U7002 (N_7002,N_6834,N_6910);
and U7003 (N_7003,N_6919,N_6759);
or U7004 (N_7004,N_6998,N_6977);
nand U7005 (N_7005,N_6787,N_6974);
xnor U7006 (N_7006,N_6973,N_6937);
nor U7007 (N_7007,N_6800,N_6965);
xor U7008 (N_7008,N_6862,N_6967);
xnor U7009 (N_7009,N_6752,N_6870);
or U7010 (N_7010,N_6874,N_6959);
nand U7011 (N_7011,N_6762,N_6783);
and U7012 (N_7012,N_6864,N_6810);
nor U7013 (N_7013,N_6952,N_6823);
xnor U7014 (N_7014,N_6946,N_6838);
nor U7015 (N_7015,N_6782,N_6917);
nand U7016 (N_7016,N_6799,N_6992);
and U7017 (N_7017,N_6833,N_6776);
and U7018 (N_7018,N_6927,N_6893);
and U7019 (N_7019,N_6915,N_6871);
nor U7020 (N_7020,N_6891,N_6849);
nor U7021 (N_7021,N_6987,N_6896);
and U7022 (N_7022,N_6822,N_6832);
nand U7023 (N_7023,N_6755,N_6808);
or U7024 (N_7024,N_6953,N_6771);
xnor U7025 (N_7025,N_6904,N_6983);
and U7026 (N_7026,N_6886,N_6957);
nand U7027 (N_7027,N_6895,N_6958);
xnor U7028 (N_7028,N_6906,N_6754);
nand U7029 (N_7029,N_6770,N_6774);
xnor U7030 (N_7030,N_6994,N_6913);
and U7031 (N_7031,N_6932,N_6963);
nand U7032 (N_7032,N_6750,N_6941);
xnor U7033 (N_7033,N_6772,N_6855);
and U7034 (N_7034,N_6969,N_6824);
xnor U7035 (N_7035,N_6831,N_6942);
nand U7036 (N_7036,N_6817,N_6916);
or U7037 (N_7037,N_6989,N_6873);
xor U7038 (N_7038,N_6841,N_6812);
xnor U7039 (N_7039,N_6966,N_6769);
nand U7040 (N_7040,N_6997,N_6802);
and U7041 (N_7041,N_6968,N_6827);
xor U7042 (N_7042,N_6843,N_6935);
nor U7043 (N_7043,N_6788,N_6988);
nand U7044 (N_7044,N_6890,N_6933);
nor U7045 (N_7045,N_6764,N_6775);
or U7046 (N_7046,N_6840,N_6999);
or U7047 (N_7047,N_6819,N_6846);
xnor U7048 (N_7048,N_6894,N_6865);
and U7049 (N_7049,N_6818,N_6951);
and U7050 (N_7050,N_6851,N_6956);
and U7051 (N_7051,N_6837,N_6961);
or U7052 (N_7052,N_6878,N_6760);
or U7053 (N_7053,N_6863,N_6792);
or U7054 (N_7054,N_6887,N_6938);
nand U7055 (N_7055,N_6784,N_6820);
or U7056 (N_7056,N_6850,N_6786);
or U7057 (N_7057,N_6909,N_6885);
nand U7058 (N_7058,N_6908,N_6881);
nor U7059 (N_7059,N_6939,N_6758);
xor U7060 (N_7060,N_6828,N_6847);
and U7061 (N_7061,N_6955,N_6753);
nand U7062 (N_7062,N_6912,N_6761);
xor U7063 (N_7063,N_6867,N_6765);
or U7064 (N_7064,N_6940,N_6995);
nor U7065 (N_7065,N_6781,N_6945);
nor U7066 (N_7066,N_6982,N_6829);
nand U7067 (N_7067,N_6853,N_6970);
and U7068 (N_7068,N_6803,N_6950);
and U7069 (N_7069,N_6805,N_6930);
or U7070 (N_7070,N_6990,N_6844);
nand U7071 (N_7071,N_6858,N_6901);
nor U7072 (N_7072,N_6980,N_6981);
and U7073 (N_7073,N_6763,N_6790);
and U7074 (N_7074,N_6804,N_6825);
nor U7075 (N_7075,N_6869,N_6861);
or U7076 (N_7076,N_6766,N_6920);
xnor U7077 (N_7077,N_6877,N_6815);
and U7078 (N_7078,N_6875,N_6964);
and U7079 (N_7079,N_6925,N_6836);
xor U7080 (N_7080,N_6852,N_6922);
nor U7081 (N_7081,N_6860,N_6902);
or U7082 (N_7082,N_6924,N_6979);
and U7083 (N_7083,N_6975,N_6821);
or U7084 (N_7084,N_6777,N_6848);
nand U7085 (N_7085,N_6801,N_6918);
and U7086 (N_7086,N_6996,N_6991);
nor U7087 (N_7087,N_6944,N_6962);
nor U7088 (N_7088,N_6789,N_6830);
and U7089 (N_7089,N_6797,N_6931);
nand U7090 (N_7090,N_6814,N_6883);
xnor U7091 (N_7091,N_6985,N_6899);
xnor U7092 (N_7092,N_6854,N_6795);
nand U7093 (N_7093,N_6882,N_6948);
or U7094 (N_7094,N_6807,N_6778);
xor U7095 (N_7095,N_6971,N_6780);
nor U7096 (N_7096,N_6856,N_6984);
nand U7097 (N_7097,N_6897,N_6905);
xor U7098 (N_7098,N_6900,N_6757);
nand U7099 (N_7099,N_6751,N_6923);
nor U7100 (N_7100,N_6791,N_6773);
xnor U7101 (N_7101,N_6960,N_6872);
and U7102 (N_7102,N_6884,N_6929);
and U7103 (N_7103,N_6978,N_6857);
or U7104 (N_7104,N_6845,N_6903);
or U7105 (N_7105,N_6986,N_6976);
nor U7106 (N_7106,N_6947,N_6892);
and U7107 (N_7107,N_6767,N_6839);
xor U7108 (N_7108,N_6928,N_6914);
and U7109 (N_7109,N_6826,N_6954);
nor U7110 (N_7110,N_6779,N_6768);
and U7111 (N_7111,N_6866,N_6926);
xnor U7112 (N_7112,N_6943,N_6835);
or U7113 (N_7113,N_6756,N_6880);
or U7114 (N_7114,N_6816,N_6806);
xor U7115 (N_7115,N_6876,N_6842);
nand U7116 (N_7116,N_6796,N_6794);
or U7117 (N_7117,N_6868,N_6911);
xor U7118 (N_7118,N_6949,N_6879);
nand U7119 (N_7119,N_6859,N_6888);
nand U7120 (N_7120,N_6972,N_6921);
nor U7121 (N_7121,N_6934,N_6889);
nor U7122 (N_7122,N_6907,N_6809);
nor U7123 (N_7123,N_6898,N_6813);
or U7124 (N_7124,N_6936,N_6993);
nand U7125 (N_7125,N_6833,N_6921);
nand U7126 (N_7126,N_6796,N_6801);
xor U7127 (N_7127,N_6952,N_6967);
nor U7128 (N_7128,N_6765,N_6800);
and U7129 (N_7129,N_6764,N_6789);
nand U7130 (N_7130,N_6936,N_6986);
xnor U7131 (N_7131,N_6943,N_6803);
nand U7132 (N_7132,N_6838,N_6752);
nand U7133 (N_7133,N_6902,N_6825);
nand U7134 (N_7134,N_6985,N_6862);
and U7135 (N_7135,N_6796,N_6770);
and U7136 (N_7136,N_6912,N_6791);
or U7137 (N_7137,N_6818,N_6829);
or U7138 (N_7138,N_6927,N_6912);
and U7139 (N_7139,N_6835,N_6755);
xnor U7140 (N_7140,N_6772,N_6796);
nor U7141 (N_7141,N_6936,N_6945);
nor U7142 (N_7142,N_6851,N_6764);
nand U7143 (N_7143,N_6857,N_6961);
nor U7144 (N_7144,N_6891,N_6939);
nor U7145 (N_7145,N_6930,N_6876);
xnor U7146 (N_7146,N_6931,N_6832);
xor U7147 (N_7147,N_6958,N_6828);
nand U7148 (N_7148,N_6940,N_6972);
and U7149 (N_7149,N_6756,N_6933);
nand U7150 (N_7150,N_6951,N_6829);
or U7151 (N_7151,N_6820,N_6823);
nor U7152 (N_7152,N_6781,N_6776);
or U7153 (N_7153,N_6803,N_6968);
xnor U7154 (N_7154,N_6954,N_6789);
nor U7155 (N_7155,N_6977,N_6755);
xor U7156 (N_7156,N_6844,N_6888);
xor U7157 (N_7157,N_6941,N_6946);
xor U7158 (N_7158,N_6856,N_6764);
xnor U7159 (N_7159,N_6949,N_6995);
nand U7160 (N_7160,N_6996,N_6755);
xnor U7161 (N_7161,N_6808,N_6996);
and U7162 (N_7162,N_6918,N_6903);
and U7163 (N_7163,N_6937,N_6761);
and U7164 (N_7164,N_6834,N_6931);
or U7165 (N_7165,N_6838,N_6982);
nand U7166 (N_7166,N_6821,N_6872);
nor U7167 (N_7167,N_6989,N_6897);
nand U7168 (N_7168,N_6947,N_6895);
or U7169 (N_7169,N_6753,N_6996);
or U7170 (N_7170,N_6781,N_6923);
and U7171 (N_7171,N_6909,N_6791);
and U7172 (N_7172,N_6774,N_6777);
nand U7173 (N_7173,N_6838,N_6793);
xor U7174 (N_7174,N_6781,N_6805);
xor U7175 (N_7175,N_6811,N_6910);
nand U7176 (N_7176,N_6776,N_6839);
and U7177 (N_7177,N_6813,N_6848);
or U7178 (N_7178,N_6786,N_6817);
nor U7179 (N_7179,N_6842,N_6867);
or U7180 (N_7180,N_6809,N_6914);
and U7181 (N_7181,N_6963,N_6887);
nor U7182 (N_7182,N_6813,N_6792);
nor U7183 (N_7183,N_6895,N_6876);
xnor U7184 (N_7184,N_6823,N_6872);
nand U7185 (N_7185,N_6965,N_6898);
xor U7186 (N_7186,N_6799,N_6791);
nand U7187 (N_7187,N_6933,N_6951);
nor U7188 (N_7188,N_6917,N_6915);
xnor U7189 (N_7189,N_6903,N_6981);
and U7190 (N_7190,N_6787,N_6811);
and U7191 (N_7191,N_6820,N_6816);
or U7192 (N_7192,N_6905,N_6796);
nand U7193 (N_7193,N_6959,N_6808);
and U7194 (N_7194,N_6964,N_6894);
nand U7195 (N_7195,N_6943,N_6925);
nor U7196 (N_7196,N_6763,N_6929);
nor U7197 (N_7197,N_6969,N_6798);
nand U7198 (N_7198,N_6760,N_6766);
and U7199 (N_7199,N_6946,N_6882);
nor U7200 (N_7200,N_6988,N_6875);
nor U7201 (N_7201,N_6857,N_6885);
nand U7202 (N_7202,N_6989,N_6938);
nor U7203 (N_7203,N_6798,N_6800);
and U7204 (N_7204,N_6885,N_6908);
xor U7205 (N_7205,N_6986,N_6792);
nand U7206 (N_7206,N_6950,N_6771);
xor U7207 (N_7207,N_6958,N_6944);
and U7208 (N_7208,N_6838,N_6863);
and U7209 (N_7209,N_6869,N_6786);
nor U7210 (N_7210,N_6783,N_6776);
or U7211 (N_7211,N_6852,N_6870);
nor U7212 (N_7212,N_6832,N_6755);
nand U7213 (N_7213,N_6932,N_6957);
nand U7214 (N_7214,N_6862,N_6768);
nand U7215 (N_7215,N_6827,N_6971);
and U7216 (N_7216,N_6944,N_6852);
xor U7217 (N_7217,N_6764,N_6767);
nand U7218 (N_7218,N_6800,N_6923);
nand U7219 (N_7219,N_6767,N_6829);
nor U7220 (N_7220,N_6797,N_6990);
nand U7221 (N_7221,N_6769,N_6816);
and U7222 (N_7222,N_6794,N_6925);
nand U7223 (N_7223,N_6804,N_6957);
nand U7224 (N_7224,N_6794,N_6904);
nand U7225 (N_7225,N_6842,N_6868);
nor U7226 (N_7226,N_6835,N_6904);
xor U7227 (N_7227,N_6887,N_6949);
xnor U7228 (N_7228,N_6939,N_6999);
or U7229 (N_7229,N_6940,N_6777);
nand U7230 (N_7230,N_6764,N_6945);
xor U7231 (N_7231,N_6751,N_6881);
or U7232 (N_7232,N_6921,N_6938);
or U7233 (N_7233,N_6844,N_6996);
xor U7234 (N_7234,N_6982,N_6760);
nand U7235 (N_7235,N_6772,N_6840);
nand U7236 (N_7236,N_6945,N_6891);
and U7237 (N_7237,N_6870,N_6765);
nand U7238 (N_7238,N_6981,N_6953);
and U7239 (N_7239,N_6821,N_6990);
or U7240 (N_7240,N_6805,N_6931);
or U7241 (N_7241,N_6920,N_6971);
nand U7242 (N_7242,N_6979,N_6897);
nand U7243 (N_7243,N_6788,N_6785);
and U7244 (N_7244,N_6789,N_6965);
nor U7245 (N_7245,N_6984,N_6945);
xor U7246 (N_7246,N_6791,N_6948);
and U7247 (N_7247,N_6977,N_6831);
nor U7248 (N_7248,N_6784,N_6928);
nor U7249 (N_7249,N_6945,N_6802);
or U7250 (N_7250,N_7206,N_7201);
and U7251 (N_7251,N_7231,N_7059);
and U7252 (N_7252,N_7116,N_7240);
nor U7253 (N_7253,N_7121,N_7029);
or U7254 (N_7254,N_7131,N_7171);
xnor U7255 (N_7255,N_7101,N_7045);
xor U7256 (N_7256,N_7165,N_7153);
nor U7257 (N_7257,N_7112,N_7071);
and U7258 (N_7258,N_7233,N_7085);
nand U7259 (N_7259,N_7221,N_7056);
xor U7260 (N_7260,N_7097,N_7098);
nor U7261 (N_7261,N_7009,N_7193);
xor U7262 (N_7262,N_7030,N_7140);
nand U7263 (N_7263,N_7016,N_7039);
and U7264 (N_7264,N_7027,N_7086);
xor U7265 (N_7265,N_7161,N_7008);
nand U7266 (N_7266,N_7237,N_7049);
nor U7267 (N_7267,N_7179,N_7002);
or U7268 (N_7268,N_7119,N_7105);
or U7269 (N_7269,N_7132,N_7155);
or U7270 (N_7270,N_7176,N_7099);
nor U7271 (N_7271,N_7134,N_7074);
xor U7272 (N_7272,N_7218,N_7149);
or U7273 (N_7273,N_7157,N_7189);
xor U7274 (N_7274,N_7247,N_7235);
nor U7275 (N_7275,N_7248,N_7023);
and U7276 (N_7276,N_7079,N_7232);
or U7277 (N_7277,N_7075,N_7128);
and U7278 (N_7278,N_7117,N_7143);
xnor U7279 (N_7279,N_7230,N_7152);
nor U7280 (N_7280,N_7151,N_7104);
nor U7281 (N_7281,N_7126,N_7110);
nor U7282 (N_7282,N_7042,N_7166);
and U7283 (N_7283,N_7224,N_7181);
xnor U7284 (N_7284,N_7052,N_7107);
and U7285 (N_7285,N_7216,N_7139);
or U7286 (N_7286,N_7219,N_7154);
or U7287 (N_7287,N_7167,N_7138);
nor U7288 (N_7288,N_7146,N_7072);
or U7289 (N_7289,N_7196,N_7156);
nor U7290 (N_7290,N_7177,N_7094);
nor U7291 (N_7291,N_7239,N_7184);
and U7292 (N_7292,N_7066,N_7035);
and U7293 (N_7293,N_7013,N_7018);
xnor U7294 (N_7294,N_7062,N_7080);
nor U7295 (N_7295,N_7111,N_7185);
xnor U7296 (N_7296,N_7047,N_7217);
nand U7297 (N_7297,N_7067,N_7000);
nor U7298 (N_7298,N_7103,N_7077);
and U7299 (N_7299,N_7054,N_7198);
nor U7300 (N_7300,N_7043,N_7236);
nand U7301 (N_7301,N_7125,N_7144);
nor U7302 (N_7302,N_7174,N_7160);
and U7303 (N_7303,N_7038,N_7243);
xor U7304 (N_7304,N_7053,N_7017);
nor U7305 (N_7305,N_7192,N_7246);
nand U7306 (N_7306,N_7106,N_7057);
nand U7307 (N_7307,N_7084,N_7203);
xor U7308 (N_7308,N_7007,N_7006);
nand U7309 (N_7309,N_7076,N_7142);
and U7310 (N_7310,N_7183,N_7050);
and U7311 (N_7311,N_7197,N_7005);
nor U7312 (N_7312,N_7202,N_7058);
xnor U7313 (N_7313,N_7032,N_7170);
xnor U7314 (N_7314,N_7133,N_7069);
and U7315 (N_7315,N_7015,N_7044);
xnor U7316 (N_7316,N_7083,N_7172);
xnor U7317 (N_7317,N_7122,N_7242);
or U7318 (N_7318,N_7180,N_7031);
nand U7319 (N_7319,N_7208,N_7003);
or U7320 (N_7320,N_7115,N_7065);
xnor U7321 (N_7321,N_7088,N_7063);
or U7322 (N_7322,N_7178,N_7014);
xor U7323 (N_7323,N_7034,N_7129);
nand U7324 (N_7324,N_7162,N_7093);
xnor U7325 (N_7325,N_7175,N_7227);
nor U7326 (N_7326,N_7092,N_7026);
nand U7327 (N_7327,N_7186,N_7187);
nand U7328 (N_7328,N_7225,N_7070);
xor U7329 (N_7329,N_7148,N_7114);
or U7330 (N_7330,N_7001,N_7012);
or U7331 (N_7331,N_7222,N_7048);
nor U7332 (N_7332,N_7147,N_7082);
xnor U7333 (N_7333,N_7159,N_7037);
or U7334 (N_7334,N_7212,N_7090);
nor U7335 (N_7335,N_7204,N_7164);
or U7336 (N_7336,N_7213,N_7078);
or U7337 (N_7337,N_7011,N_7073);
or U7338 (N_7338,N_7214,N_7091);
nor U7339 (N_7339,N_7124,N_7209);
xnor U7340 (N_7340,N_7130,N_7169);
xor U7341 (N_7341,N_7108,N_7089);
or U7342 (N_7342,N_7141,N_7120);
or U7343 (N_7343,N_7191,N_7137);
xnor U7344 (N_7344,N_7234,N_7223);
xor U7345 (N_7345,N_7033,N_7158);
xnor U7346 (N_7346,N_7040,N_7060);
or U7347 (N_7347,N_7022,N_7194);
xor U7348 (N_7348,N_7064,N_7188);
or U7349 (N_7349,N_7199,N_7182);
or U7350 (N_7350,N_7226,N_7228);
nor U7351 (N_7351,N_7020,N_7036);
nor U7352 (N_7352,N_7207,N_7195);
xnor U7353 (N_7353,N_7210,N_7081);
and U7354 (N_7354,N_7123,N_7025);
xnor U7355 (N_7355,N_7249,N_7211);
and U7356 (N_7356,N_7229,N_7028);
nand U7357 (N_7357,N_7200,N_7095);
nor U7358 (N_7358,N_7100,N_7087);
or U7359 (N_7359,N_7046,N_7068);
nand U7360 (N_7360,N_7205,N_7244);
nor U7361 (N_7361,N_7190,N_7113);
or U7362 (N_7362,N_7109,N_7245);
or U7363 (N_7363,N_7136,N_7004);
nor U7364 (N_7364,N_7127,N_7051);
xnor U7365 (N_7365,N_7118,N_7096);
and U7366 (N_7366,N_7010,N_7173);
or U7367 (N_7367,N_7215,N_7163);
nand U7368 (N_7368,N_7061,N_7135);
xor U7369 (N_7369,N_7238,N_7150);
and U7370 (N_7370,N_7024,N_7220);
xor U7371 (N_7371,N_7241,N_7168);
nand U7372 (N_7372,N_7021,N_7145);
xnor U7373 (N_7373,N_7041,N_7055);
xor U7374 (N_7374,N_7102,N_7019);
or U7375 (N_7375,N_7132,N_7196);
and U7376 (N_7376,N_7111,N_7161);
nor U7377 (N_7377,N_7085,N_7106);
nand U7378 (N_7378,N_7089,N_7126);
nand U7379 (N_7379,N_7191,N_7187);
nor U7380 (N_7380,N_7138,N_7060);
xnor U7381 (N_7381,N_7149,N_7066);
or U7382 (N_7382,N_7241,N_7104);
nor U7383 (N_7383,N_7210,N_7087);
nand U7384 (N_7384,N_7015,N_7180);
xnor U7385 (N_7385,N_7003,N_7156);
nand U7386 (N_7386,N_7105,N_7071);
xnor U7387 (N_7387,N_7196,N_7198);
xor U7388 (N_7388,N_7024,N_7081);
xnor U7389 (N_7389,N_7199,N_7223);
xor U7390 (N_7390,N_7110,N_7081);
and U7391 (N_7391,N_7086,N_7163);
xnor U7392 (N_7392,N_7234,N_7198);
or U7393 (N_7393,N_7221,N_7218);
and U7394 (N_7394,N_7236,N_7128);
nor U7395 (N_7395,N_7202,N_7080);
or U7396 (N_7396,N_7032,N_7181);
xnor U7397 (N_7397,N_7146,N_7165);
nand U7398 (N_7398,N_7130,N_7181);
nand U7399 (N_7399,N_7037,N_7069);
xor U7400 (N_7400,N_7091,N_7236);
xor U7401 (N_7401,N_7192,N_7225);
and U7402 (N_7402,N_7182,N_7108);
and U7403 (N_7403,N_7147,N_7172);
or U7404 (N_7404,N_7052,N_7046);
nand U7405 (N_7405,N_7152,N_7167);
and U7406 (N_7406,N_7241,N_7179);
nand U7407 (N_7407,N_7000,N_7171);
or U7408 (N_7408,N_7027,N_7060);
or U7409 (N_7409,N_7244,N_7005);
or U7410 (N_7410,N_7073,N_7159);
and U7411 (N_7411,N_7138,N_7136);
nand U7412 (N_7412,N_7195,N_7059);
xnor U7413 (N_7413,N_7133,N_7155);
nand U7414 (N_7414,N_7141,N_7213);
or U7415 (N_7415,N_7234,N_7018);
nand U7416 (N_7416,N_7008,N_7003);
xor U7417 (N_7417,N_7234,N_7144);
or U7418 (N_7418,N_7239,N_7016);
nor U7419 (N_7419,N_7230,N_7213);
or U7420 (N_7420,N_7125,N_7135);
xnor U7421 (N_7421,N_7209,N_7036);
xor U7422 (N_7422,N_7116,N_7198);
nand U7423 (N_7423,N_7116,N_7231);
nand U7424 (N_7424,N_7055,N_7047);
nor U7425 (N_7425,N_7110,N_7244);
nor U7426 (N_7426,N_7107,N_7169);
and U7427 (N_7427,N_7098,N_7046);
and U7428 (N_7428,N_7215,N_7248);
or U7429 (N_7429,N_7118,N_7041);
and U7430 (N_7430,N_7168,N_7025);
xnor U7431 (N_7431,N_7194,N_7247);
xor U7432 (N_7432,N_7018,N_7069);
xnor U7433 (N_7433,N_7070,N_7176);
and U7434 (N_7434,N_7123,N_7053);
or U7435 (N_7435,N_7123,N_7093);
nor U7436 (N_7436,N_7168,N_7027);
nand U7437 (N_7437,N_7116,N_7009);
or U7438 (N_7438,N_7109,N_7050);
or U7439 (N_7439,N_7085,N_7073);
nor U7440 (N_7440,N_7101,N_7134);
xnor U7441 (N_7441,N_7056,N_7199);
and U7442 (N_7442,N_7195,N_7016);
nand U7443 (N_7443,N_7012,N_7047);
or U7444 (N_7444,N_7223,N_7170);
nor U7445 (N_7445,N_7144,N_7030);
or U7446 (N_7446,N_7154,N_7087);
nor U7447 (N_7447,N_7178,N_7036);
nand U7448 (N_7448,N_7144,N_7021);
or U7449 (N_7449,N_7177,N_7070);
nand U7450 (N_7450,N_7137,N_7016);
and U7451 (N_7451,N_7043,N_7095);
xnor U7452 (N_7452,N_7026,N_7187);
and U7453 (N_7453,N_7101,N_7089);
xor U7454 (N_7454,N_7127,N_7122);
nand U7455 (N_7455,N_7163,N_7172);
xor U7456 (N_7456,N_7044,N_7240);
and U7457 (N_7457,N_7085,N_7100);
nand U7458 (N_7458,N_7041,N_7149);
and U7459 (N_7459,N_7226,N_7047);
nand U7460 (N_7460,N_7065,N_7129);
nor U7461 (N_7461,N_7005,N_7059);
and U7462 (N_7462,N_7036,N_7093);
xor U7463 (N_7463,N_7125,N_7086);
or U7464 (N_7464,N_7132,N_7220);
and U7465 (N_7465,N_7144,N_7128);
and U7466 (N_7466,N_7055,N_7044);
nor U7467 (N_7467,N_7143,N_7074);
xor U7468 (N_7468,N_7014,N_7246);
and U7469 (N_7469,N_7103,N_7040);
and U7470 (N_7470,N_7203,N_7078);
or U7471 (N_7471,N_7053,N_7082);
xnor U7472 (N_7472,N_7140,N_7012);
nor U7473 (N_7473,N_7053,N_7246);
and U7474 (N_7474,N_7003,N_7149);
and U7475 (N_7475,N_7073,N_7061);
nor U7476 (N_7476,N_7146,N_7109);
nand U7477 (N_7477,N_7234,N_7102);
or U7478 (N_7478,N_7122,N_7128);
or U7479 (N_7479,N_7101,N_7241);
xnor U7480 (N_7480,N_7068,N_7081);
and U7481 (N_7481,N_7034,N_7234);
and U7482 (N_7482,N_7105,N_7082);
nor U7483 (N_7483,N_7248,N_7106);
nand U7484 (N_7484,N_7020,N_7157);
nand U7485 (N_7485,N_7200,N_7153);
and U7486 (N_7486,N_7238,N_7209);
and U7487 (N_7487,N_7080,N_7011);
nand U7488 (N_7488,N_7145,N_7193);
xor U7489 (N_7489,N_7057,N_7164);
or U7490 (N_7490,N_7104,N_7027);
nor U7491 (N_7491,N_7082,N_7055);
or U7492 (N_7492,N_7127,N_7000);
nand U7493 (N_7493,N_7204,N_7007);
xnor U7494 (N_7494,N_7003,N_7152);
or U7495 (N_7495,N_7099,N_7132);
nand U7496 (N_7496,N_7076,N_7228);
nor U7497 (N_7497,N_7119,N_7143);
or U7498 (N_7498,N_7203,N_7036);
nand U7499 (N_7499,N_7185,N_7219);
or U7500 (N_7500,N_7327,N_7459);
nor U7501 (N_7501,N_7364,N_7392);
or U7502 (N_7502,N_7448,N_7413);
or U7503 (N_7503,N_7368,N_7325);
xnor U7504 (N_7504,N_7428,N_7363);
and U7505 (N_7505,N_7354,N_7317);
or U7506 (N_7506,N_7328,N_7398);
xnor U7507 (N_7507,N_7485,N_7443);
nand U7508 (N_7508,N_7261,N_7296);
xnor U7509 (N_7509,N_7336,N_7492);
nor U7510 (N_7510,N_7400,N_7391);
or U7511 (N_7511,N_7268,N_7463);
or U7512 (N_7512,N_7300,N_7343);
or U7513 (N_7513,N_7381,N_7265);
or U7514 (N_7514,N_7480,N_7431);
nor U7515 (N_7515,N_7433,N_7313);
xor U7516 (N_7516,N_7326,N_7435);
nand U7517 (N_7517,N_7407,N_7284);
or U7518 (N_7518,N_7434,N_7259);
and U7519 (N_7519,N_7461,N_7399);
nor U7520 (N_7520,N_7274,N_7387);
nor U7521 (N_7521,N_7348,N_7453);
or U7522 (N_7522,N_7419,N_7331);
nor U7523 (N_7523,N_7333,N_7360);
nor U7524 (N_7524,N_7370,N_7417);
nor U7525 (N_7525,N_7385,N_7332);
nand U7526 (N_7526,N_7340,N_7257);
or U7527 (N_7527,N_7457,N_7452);
nand U7528 (N_7528,N_7386,N_7302);
and U7529 (N_7529,N_7335,N_7478);
or U7530 (N_7530,N_7491,N_7495);
or U7531 (N_7531,N_7319,N_7402);
and U7532 (N_7532,N_7476,N_7321);
nor U7533 (N_7533,N_7358,N_7487);
and U7534 (N_7534,N_7490,N_7393);
and U7535 (N_7535,N_7432,N_7384);
nor U7536 (N_7536,N_7493,N_7305);
nand U7537 (N_7537,N_7494,N_7424);
nor U7538 (N_7538,N_7499,N_7451);
or U7539 (N_7539,N_7349,N_7395);
xor U7540 (N_7540,N_7446,N_7460);
and U7541 (N_7541,N_7263,N_7405);
nand U7542 (N_7542,N_7447,N_7465);
nor U7543 (N_7543,N_7345,N_7477);
nand U7544 (N_7544,N_7322,N_7430);
nand U7545 (N_7545,N_7362,N_7301);
and U7546 (N_7546,N_7308,N_7323);
nor U7547 (N_7547,N_7454,N_7421);
xnor U7548 (N_7548,N_7472,N_7359);
nor U7549 (N_7549,N_7464,N_7283);
xnor U7550 (N_7550,N_7266,N_7254);
nand U7551 (N_7551,N_7339,N_7286);
nor U7552 (N_7552,N_7437,N_7466);
nor U7553 (N_7553,N_7404,N_7275);
nand U7554 (N_7554,N_7473,N_7438);
nand U7555 (N_7555,N_7397,N_7252);
nand U7556 (N_7556,N_7316,N_7422);
nor U7557 (N_7557,N_7379,N_7350);
nor U7558 (N_7558,N_7444,N_7450);
or U7559 (N_7559,N_7279,N_7479);
xor U7560 (N_7560,N_7481,N_7310);
and U7561 (N_7561,N_7426,N_7408);
or U7562 (N_7562,N_7436,N_7489);
nand U7563 (N_7563,N_7415,N_7267);
and U7564 (N_7564,N_7356,N_7341);
nand U7565 (N_7565,N_7324,N_7378);
nor U7566 (N_7566,N_7344,N_7250);
and U7567 (N_7567,N_7297,N_7309);
and U7568 (N_7568,N_7409,N_7445);
nand U7569 (N_7569,N_7277,N_7449);
xor U7570 (N_7570,N_7292,N_7410);
nor U7571 (N_7571,N_7291,N_7272);
nand U7572 (N_7572,N_7373,N_7488);
xor U7573 (N_7573,N_7470,N_7375);
or U7574 (N_7574,N_7251,N_7423);
and U7575 (N_7575,N_7312,N_7276);
nand U7576 (N_7576,N_7353,N_7256);
and U7577 (N_7577,N_7469,N_7440);
xnor U7578 (N_7578,N_7486,N_7416);
or U7579 (N_7579,N_7427,N_7498);
xnor U7580 (N_7580,N_7337,N_7377);
nand U7581 (N_7581,N_7285,N_7273);
or U7582 (N_7582,N_7346,N_7329);
xor U7583 (N_7583,N_7269,N_7456);
xor U7584 (N_7584,N_7411,N_7347);
or U7585 (N_7585,N_7303,N_7278);
nor U7586 (N_7586,N_7280,N_7382);
nand U7587 (N_7587,N_7320,N_7371);
nor U7588 (N_7588,N_7388,N_7420);
nor U7589 (N_7589,N_7304,N_7366);
nand U7590 (N_7590,N_7264,N_7475);
xor U7591 (N_7591,N_7293,N_7258);
xor U7592 (N_7592,N_7455,N_7338);
nor U7593 (N_7593,N_7401,N_7414);
nor U7594 (N_7594,N_7474,N_7351);
xnor U7595 (N_7595,N_7497,N_7429);
and U7596 (N_7596,N_7471,N_7482);
xnor U7597 (N_7597,N_7255,N_7403);
or U7598 (N_7598,N_7334,N_7390);
nor U7599 (N_7599,N_7496,N_7367);
nor U7600 (N_7600,N_7287,N_7298);
nor U7601 (N_7601,N_7294,N_7361);
or U7602 (N_7602,N_7270,N_7374);
nand U7603 (N_7603,N_7468,N_7484);
nor U7604 (N_7604,N_7372,N_7383);
nand U7605 (N_7605,N_7467,N_7299);
and U7606 (N_7606,N_7342,N_7271);
or U7607 (N_7607,N_7357,N_7365);
xnor U7608 (N_7608,N_7483,N_7442);
nand U7609 (N_7609,N_7406,N_7441);
nor U7610 (N_7610,N_7389,N_7462);
nor U7611 (N_7611,N_7282,N_7355);
nor U7612 (N_7612,N_7289,N_7412);
or U7613 (N_7613,N_7330,N_7394);
and U7614 (N_7614,N_7307,N_7306);
or U7615 (N_7615,N_7288,N_7380);
nand U7616 (N_7616,N_7396,N_7352);
and U7617 (N_7617,N_7418,N_7295);
nand U7618 (N_7618,N_7369,N_7314);
and U7619 (N_7619,N_7262,N_7439);
and U7620 (N_7620,N_7315,N_7281);
nand U7621 (N_7621,N_7290,N_7425);
xor U7622 (N_7622,N_7318,N_7260);
or U7623 (N_7623,N_7458,N_7376);
nand U7624 (N_7624,N_7253,N_7311);
or U7625 (N_7625,N_7315,N_7286);
or U7626 (N_7626,N_7452,N_7475);
nand U7627 (N_7627,N_7262,N_7254);
or U7628 (N_7628,N_7362,N_7294);
or U7629 (N_7629,N_7250,N_7320);
nor U7630 (N_7630,N_7495,N_7270);
or U7631 (N_7631,N_7315,N_7464);
nor U7632 (N_7632,N_7417,N_7357);
and U7633 (N_7633,N_7267,N_7412);
and U7634 (N_7634,N_7475,N_7253);
xnor U7635 (N_7635,N_7328,N_7429);
nor U7636 (N_7636,N_7338,N_7384);
nor U7637 (N_7637,N_7473,N_7300);
nand U7638 (N_7638,N_7493,N_7428);
nand U7639 (N_7639,N_7290,N_7402);
and U7640 (N_7640,N_7428,N_7377);
nand U7641 (N_7641,N_7407,N_7497);
or U7642 (N_7642,N_7462,N_7347);
or U7643 (N_7643,N_7318,N_7458);
and U7644 (N_7644,N_7255,N_7283);
nor U7645 (N_7645,N_7331,N_7410);
nor U7646 (N_7646,N_7480,N_7271);
nand U7647 (N_7647,N_7284,N_7362);
and U7648 (N_7648,N_7401,N_7422);
nand U7649 (N_7649,N_7366,N_7488);
or U7650 (N_7650,N_7313,N_7386);
and U7651 (N_7651,N_7377,N_7497);
or U7652 (N_7652,N_7395,N_7398);
and U7653 (N_7653,N_7367,N_7292);
nor U7654 (N_7654,N_7383,N_7429);
nor U7655 (N_7655,N_7431,N_7319);
nor U7656 (N_7656,N_7372,N_7303);
xor U7657 (N_7657,N_7327,N_7446);
nor U7658 (N_7658,N_7451,N_7261);
nand U7659 (N_7659,N_7420,N_7301);
nor U7660 (N_7660,N_7287,N_7297);
nand U7661 (N_7661,N_7252,N_7365);
xnor U7662 (N_7662,N_7449,N_7265);
or U7663 (N_7663,N_7383,N_7403);
nor U7664 (N_7664,N_7398,N_7410);
and U7665 (N_7665,N_7280,N_7391);
and U7666 (N_7666,N_7367,N_7360);
xnor U7667 (N_7667,N_7417,N_7424);
xor U7668 (N_7668,N_7470,N_7335);
and U7669 (N_7669,N_7275,N_7345);
xnor U7670 (N_7670,N_7493,N_7444);
nand U7671 (N_7671,N_7355,N_7299);
nor U7672 (N_7672,N_7410,N_7425);
or U7673 (N_7673,N_7319,N_7305);
or U7674 (N_7674,N_7305,N_7448);
or U7675 (N_7675,N_7298,N_7449);
and U7676 (N_7676,N_7320,N_7313);
xor U7677 (N_7677,N_7447,N_7369);
nand U7678 (N_7678,N_7499,N_7476);
or U7679 (N_7679,N_7390,N_7460);
xnor U7680 (N_7680,N_7476,N_7484);
and U7681 (N_7681,N_7264,N_7423);
nand U7682 (N_7682,N_7411,N_7339);
nand U7683 (N_7683,N_7355,N_7496);
or U7684 (N_7684,N_7460,N_7419);
xor U7685 (N_7685,N_7321,N_7429);
nor U7686 (N_7686,N_7431,N_7476);
and U7687 (N_7687,N_7309,N_7266);
and U7688 (N_7688,N_7342,N_7435);
and U7689 (N_7689,N_7304,N_7473);
nor U7690 (N_7690,N_7320,N_7480);
nor U7691 (N_7691,N_7420,N_7460);
nand U7692 (N_7692,N_7423,N_7397);
xnor U7693 (N_7693,N_7306,N_7488);
and U7694 (N_7694,N_7401,N_7309);
or U7695 (N_7695,N_7471,N_7299);
and U7696 (N_7696,N_7400,N_7414);
nand U7697 (N_7697,N_7449,N_7398);
nand U7698 (N_7698,N_7423,N_7458);
nor U7699 (N_7699,N_7446,N_7468);
or U7700 (N_7700,N_7375,N_7303);
and U7701 (N_7701,N_7388,N_7425);
nand U7702 (N_7702,N_7396,N_7284);
and U7703 (N_7703,N_7267,N_7356);
or U7704 (N_7704,N_7453,N_7438);
xor U7705 (N_7705,N_7494,N_7317);
xnor U7706 (N_7706,N_7486,N_7299);
xor U7707 (N_7707,N_7359,N_7425);
xnor U7708 (N_7708,N_7427,N_7482);
and U7709 (N_7709,N_7426,N_7277);
or U7710 (N_7710,N_7295,N_7288);
xnor U7711 (N_7711,N_7418,N_7269);
nand U7712 (N_7712,N_7422,N_7388);
nand U7713 (N_7713,N_7402,N_7384);
or U7714 (N_7714,N_7313,N_7252);
and U7715 (N_7715,N_7472,N_7408);
or U7716 (N_7716,N_7277,N_7287);
and U7717 (N_7717,N_7310,N_7321);
or U7718 (N_7718,N_7309,N_7285);
and U7719 (N_7719,N_7361,N_7262);
nand U7720 (N_7720,N_7454,N_7268);
and U7721 (N_7721,N_7354,N_7474);
nor U7722 (N_7722,N_7478,N_7494);
nor U7723 (N_7723,N_7297,N_7407);
nand U7724 (N_7724,N_7330,N_7408);
xor U7725 (N_7725,N_7355,N_7398);
nor U7726 (N_7726,N_7433,N_7337);
nand U7727 (N_7727,N_7402,N_7491);
and U7728 (N_7728,N_7305,N_7416);
nand U7729 (N_7729,N_7382,N_7451);
or U7730 (N_7730,N_7419,N_7428);
xor U7731 (N_7731,N_7470,N_7405);
or U7732 (N_7732,N_7392,N_7461);
xor U7733 (N_7733,N_7482,N_7307);
nor U7734 (N_7734,N_7448,N_7278);
nor U7735 (N_7735,N_7270,N_7489);
xor U7736 (N_7736,N_7463,N_7302);
xnor U7737 (N_7737,N_7259,N_7325);
nor U7738 (N_7738,N_7391,N_7269);
xor U7739 (N_7739,N_7452,N_7358);
and U7740 (N_7740,N_7266,N_7304);
or U7741 (N_7741,N_7393,N_7347);
or U7742 (N_7742,N_7301,N_7273);
xnor U7743 (N_7743,N_7285,N_7409);
or U7744 (N_7744,N_7433,N_7426);
xnor U7745 (N_7745,N_7323,N_7466);
or U7746 (N_7746,N_7333,N_7361);
or U7747 (N_7747,N_7377,N_7328);
or U7748 (N_7748,N_7489,N_7396);
nand U7749 (N_7749,N_7455,N_7302);
xor U7750 (N_7750,N_7704,N_7587);
xor U7751 (N_7751,N_7666,N_7656);
or U7752 (N_7752,N_7739,N_7502);
and U7753 (N_7753,N_7642,N_7714);
nor U7754 (N_7754,N_7525,N_7690);
nor U7755 (N_7755,N_7667,N_7670);
nor U7756 (N_7756,N_7677,N_7685);
and U7757 (N_7757,N_7635,N_7725);
nor U7758 (N_7758,N_7747,N_7588);
xnor U7759 (N_7759,N_7535,N_7584);
nand U7760 (N_7760,N_7537,N_7689);
or U7761 (N_7761,N_7555,N_7679);
xor U7762 (N_7762,N_7683,N_7572);
nor U7763 (N_7763,N_7583,N_7665);
nor U7764 (N_7764,N_7591,N_7580);
xnor U7765 (N_7765,N_7669,N_7523);
or U7766 (N_7766,N_7516,N_7713);
nand U7767 (N_7767,N_7738,N_7595);
and U7768 (N_7768,N_7673,N_7547);
nor U7769 (N_7769,N_7614,N_7631);
or U7770 (N_7770,N_7606,N_7508);
xnor U7771 (N_7771,N_7564,N_7640);
nor U7772 (N_7772,N_7705,N_7624);
and U7773 (N_7773,N_7645,N_7539);
and U7774 (N_7774,N_7597,N_7611);
xnor U7775 (N_7775,N_7680,N_7695);
nand U7776 (N_7776,N_7744,N_7616);
xnor U7777 (N_7777,N_7742,N_7592);
nand U7778 (N_7778,N_7657,N_7626);
nor U7779 (N_7779,N_7603,N_7543);
nand U7780 (N_7780,N_7678,N_7732);
nor U7781 (N_7781,N_7629,N_7636);
nor U7782 (N_7782,N_7686,N_7723);
nand U7783 (N_7783,N_7688,N_7736);
nor U7784 (N_7784,N_7724,N_7722);
nor U7785 (N_7785,N_7522,N_7659);
and U7786 (N_7786,N_7549,N_7701);
nor U7787 (N_7787,N_7556,N_7548);
and U7788 (N_7788,N_7552,N_7733);
and U7789 (N_7789,N_7536,N_7530);
and U7790 (N_7790,N_7716,N_7506);
nor U7791 (N_7791,N_7565,N_7646);
or U7792 (N_7792,N_7540,N_7660);
xnor U7793 (N_7793,N_7692,N_7651);
nand U7794 (N_7794,N_7568,N_7641);
nor U7795 (N_7795,N_7623,N_7630);
nor U7796 (N_7796,N_7531,N_7517);
nor U7797 (N_7797,N_7503,N_7617);
nor U7798 (N_7798,N_7562,N_7600);
and U7799 (N_7799,N_7561,N_7699);
or U7800 (N_7800,N_7745,N_7697);
nand U7801 (N_7801,N_7727,N_7712);
or U7802 (N_7802,N_7598,N_7709);
nor U7803 (N_7803,N_7718,N_7663);
and U7804 (N_7804,N_7538,N_7649);
and U7805 (N_7805,N_7520,N_7620);
and U7806 (N_7806,N_7638,N_7578);
nor U7807 (N_7807,N_7515,N_7654);
and U7808 (N_7808,N_7563,N_7526);
and U7809 (N_7809,N_7596,N_7613);
nor U7810 (N_7810,N_7601,N_7507);
xor U7811 (N_7811,N_7687,N_7622);
or U7812 (N_7812,N_7544,N_7633);
or U7813 (N_7813,N_7741,N_7625);
nor U7814 (N_7814,N_7737,N_7571);
and U7815 (N_7815,N_7615,N_7675);
and U7816 (N_7816,N_7610,N_7557);
nor U7817 (N_7817,N_7546,N_7550);
and U7818 (N_7818,N_7585,N_7590);
nor U7819 (N_7819,N_7586,N_7662);
or U7820 (N_7820,N_7627,N_7570);
or U7821 (N_7821,N_7647,N_7719);
nand U7822 (N_7822,N_7740,N_7681);
nor U7823 (N_7823,N_7529,N_7589);
nand U7824 (N_7824,N_7505,N_7612);
xnor U7825 (N_7825,N_7749,N_7609);
nand U7826 (N_7826,N_7655,N_7728);
or U7827 (N_7827,N_7671,N_7527);
xor U7828 (N_7828,N_7608,N_7512);
nor U7829 (N_7829,N_7694,N_7545);
or U7830 (N_7830,N_7542,N_7519);
and U7831 (N_7831,N_7730,N_7729);
nor U7832 (N_7832,N_7533,N_7710);
nor U7833 (N_7833,N_7628,N_7599);
nor U7834 (N_7834,N_7717,N_7734);
or U7835 (N_7835,N_7501,N_7573);
nor U7836 (N_7836,N_7518,N_7637);
xnor U7837 (N_7837,N_7658,N_7668);
and U7838 (N_7838,N_7619,N_7743);
xor U7839 (N_7839,N_7510,N_7720);
or U7840 (N_7840,N_7602,N_7579);
or U7841 (N_7841,N_7721,N_7504);
xor U7842 (N_7842,N_7639,N_7711);
and U7843 (N_7843,N_7582,N_7511);
or U7844 (N_7844,N_7576,N_7652);
or U7845 (N_7845,N_7706,N_7551);
nand U7846 (N_7846,N_7702,N_7735);
nor U7847 (N_7847,N_7691,N_7684);
nand U7848 (N_7848,N_7634,N_7643);
nand U7849 (N_7849,N_7553,N_7513);
nand U7850 (N_7850,N_7541,N_7693);
nand U7851 (N_7851,N_7682,N_7708);
nand U7852 (N_7852,N_7567,N_7605);
nand U7853 (N_7853,N_7726,N_7560);
and U7854 (N_7854,N_7661,N_7746);
nor U7855 (N_7855,N_7593,N_7569);
nor U7856 (N_7856,N_7731,N_7648);
xnor U7857 (N_7857,N_7554,N_7575);
and U7858 (N_7858,N_7534,N_7532);
nor U7859 (N_7859,N_7700,N_7604);
and U7860 (N_7860,N_7632,N_7607);
xnor U7861 (N_7861,N_7574,N_7524);
xor U7862 (N_7862,N_7618,N_7594);
or U7863 (N_7863,N_7698,N_7528);
nor U7864 (N_7864,N_7514,N_7509);
nor U7865 (N_7865,N_7566,N_7559);
or U7866 (N_7866,N_7558,N_7664);
xnor U7867 (N_7867,N_7707,N_7644);
or U7868 (N_7868,N_7650,N_7577);
nor U7869 (N_7869,N_7674,N_7703);
nor U7870 (N_7870,N_7696,N_7500);
nor U7871 (N_7871,N_7672,N_7653);
nor U7872 (N_7872,N_7581,N_7748);
nor U7873 (N_7873,N_7521,N_7676);
or U7874 (N_7874,N_7715,N_7621);
and U7875 (N_7875,N_7508,N_7726);
and U7876 (N_7876,N_7512,N_7585);
nand U7877 (N_7877,N_7612,N_7655);
nor U7878 (N_7878,N_7641,N_7552);
xnor U7879 (N_7879,N_7738,N_7531);
nand U7880 (N_7880,N_7502,N_7514);
and U7881 (N_7881,N_7583,N_7746);
nor U7882 (N_7882,N_7720,N_7605);
and U7883 (N_7883,N_7647,N_7567);
or U7884 (N_7884,N_7550,N_7695);
nor U7885 (N_7885,N_7555,N_7579);
and U7886 (N_7886,N_7640,N_7595);
xor U7887 (N_7887,N_7675,N_7549);
nor U7888 (N_7888,N_7519,N_7626);
and U7889 (N_7889,N_7679,N_7612);
and U7890 (N_7890,N_7653,N_7657);
nand U7891 (N_7891,N_7542,N_7659);
xnor U7892 (N_7892,N_7587,N_7738);
xor U7893 (N_7893,N_7693,N_7682);
nor U7894 (N_7894,N_7616,N_7521);
xnor U7895 (N_7895,N_7637,N_7669);
xnor U7896 (N_7896,N_7697,N_7692);
and U7897 (N_7897,N_7619,N_7731);
or U7898 (N_7898,N_7502,N_7725);
nand U7899 (N_7899,N_7623,N_7684);
nand U7900 (N_7900,N_7739,N_7609);
xnor U7901 (N_7901,N_7502,N_7728);
and U7902 (N_7902,N_7519,N_7588);
xnor U7903 (N_7903,N_7504,N_7711);
xor U7904 (N_7904,N_7641,N_7660);
xnor U7905 (N_7905,N_7582,N_7657);
nand U7906 (N_7906,N_7660,N_7555);
xor U7907 (N_7907,N_7571,N_7511);
xor U7908 (N_7908,N_7520,N_7741);
xnor U7909 (N_7909,N_7503,N_7747);
xor U7910 (N_7910,N_7580,N_7677);
nand U7911 (N_7911,N_7707,N_7572);
nor U7912 (N_7912,N_7733,N_7585);
nand U7913 (N_7913,N_7650,N_7669);
and U7914 (N_7914,N_7644,N_7598);
and U7915 (N_7915,N_7671,N_7655);
or U7916 (N_7916,N_7603,N_7583);
nor U7917 (N_7917,N_7547,N_7548);
and U7918 (N_7918,N_7514,N_7566);
nor U7919 (N_7919,N_7699,N_7707);
nor U7920 (N_7920,N_7566,N_7667);
nand U7921 (N_7921,N_7533,N_7663);
nand U7922 (N_7922,N_7518,N_7685);
and U7923 (N_7923,N_7599,N_7631);
and U7924 (N_7924,N_7708,N_7540);
or U7925 (N_7925,N_7718,N_7595);
nor U7926 (N_7926,N_7602,N_7571);
and U7927 (N_7927,N_7565,N_7700);
xor U7928 (N_7928,N_7506,N_7555);
xor U7929 (N_7929,N_7657,N_7602);
nor U7930 (N_7930,N_7566,N_7596);
nor U7931 (N_7931,N_7572,N_7589);
nor U7932 (N_7932,N_7739,N_7715);
nor U7933 (N_7933,N_7640,N_7579);
or U7934 (N_7934,N_7643,N_7514);
or U7935 (N_7935,N_7600,N_7708);
or U7936 (N_7936,N_7719,N_7540);
xor U7937 (N_7937,N_7734,N_7507);
xnor U7938 (N_7938,N_7691,N_7526);
xnor U7939 (N_7939,N_7564,N_7605);
or U7940 (N_7940,N_7564,N_7514);
nor U7941 (N_7941,N_7658,N_7558);
nor U7942 (N_7942,N_7651,N_7502);
or U7943 (N_7943,N_7591,N_7635);
nor U7944 (N_7944,N_7710,N_7728);
or U7945 (N_7945,N_7506,N_7731);
nand U7946 (N_7946,N_7679,N_7564);
nor U7947 (N_7947,N_7639,N_7706);
nand U7948 (N_7948,N_7598,N_7717);
or U7949 (N_7949,N_7588,N_7667);
xor U7950 (N_7950,N_7708,N_7542);
and U7951 (N_7951,N_7622,N_7525);
nand U7952 (N_7952,N_7622,N_7519);
nor U7953 (N_7953,N_7540,N_7743);
xor U7954 (N_7954,N_7545,N_7522);
nand U7955 (N_7955,N_7562,N_7732);
xor U7956 (N_7956,N_7573,N_7597);
xor U7957 (N_7957,N_7734,N_7680);
or U7958 (N_7958,N_7559,N_7616);
nand U7959 (N_7959,N_7562,N_7684);
xnor U7960 (N_7960,N_7616,N_7589);
or U7961 (N_7961,N_7540,N_7606);
and U7962 (N_7962,N_7713,N_7748);
or U7963 (N_7963,N_7743,N_7740);
nand U7964 (N_7964,N_7644,N_7570);
nor U7965 (N_7965,N_7702,N_7568);
or U7966 (N_7966,N_7548,N_7694);
nor U7967 (N_7967,N_7535,N_7686);
and U7968 (N_7968,N_7628,N_7663);
nand U7969 (N_7969,N_7517,N_7616);
nand U7970 (N_7970,N_7627,N_7696);
xor U7971 (N_7971,N_7527,N_7748);
nor U7972 (N_7972,N_7565,N_7517);
or U7973 (N_7973,N_7552,N_7602);
or U7974 (N_7974,N_7684,N_7741);
or U7975 (N_7975,N_7532,N_7675);
and U7976 (N_7976,N_7725,N_7696);
nor U7977 (N_7977,N_7691,N_7666);
or U7978 (N_7978,N_7688,N_7563);
nand U7979 (N_7979,N_7670,N_7548);
nand U7980 (N_7980,N_7694,N_7689);
nor U7981 (N_7981,N_7653,N_7687);
and U7982 (N_7982,N_7605,N_7571);
and U7983 (N_7983,N_7713,N_7515);
nand U7984 (N_7984,N_7612,N_7538);
nand U7985 (N_7985,N_7709,N_7720);
xnor U7986 (N_7986,N_7691,N_7576);
or U7987 (N_7987,N_7608,N_7542);
nand U7988 (N_7988,N_7699,N_7683);
nor U7989 (N_7989,N_7746,N_7638);
nor U7990 (N_7990,N_7508,N_7641);
or U7991 (N_7991,N_7552,N_7595);
or U7992 (N_7992,N_7724,N_7660);
nor U7993 (N_7993,N_7702,N_7699);
xnor U7994 (N_7994,N_7696,N_7529);
nor U7995 (N_7995,N_7563,N_7565);
nand U7996 (N_7996,N_7650,N_7585);
or U7997 (N_7997,N_7707,N_7566);
and U7998 (N_7998,N_7726,N_7676);
and U7999 (N_7999,N_7551,N_7651);
xnor U8000 (N_8000,N_7958,N_7872);
or U8001 (N_8001,N_7992,N_7957);
nand U8002 (N_8002,N_7769,N_7883);
nor U8003 (N_8003,N_7761,N_7930);
nand U8004 (N_8004,N_7941,N_7829);
or U8005 (N_8005,N_7822,N_7905);
nor U8006 (N_8006,N_7867,N_7971);
xor U8007 (N_8007,N_7979,N_7871);
or U8008 (N_8008,N_7762,N_7760);
xnor U8009 (N_8009,N_7868,N_7942);
or U8010 (N_8010,N_7980,N_7965);
nor U8011 (N_8011,N_7983,N_7777);
or U8012 (N_8012,N_7766,N_7989);
xor U8013 (N_8013,N_7895,N_7811);
or U8014 (N_8014,N_7984,N_7994);
or U8015 (N_8015,N_7865,N_7850);
xnor U8016 (N_8016,N_7828,N_7785);
xor U8017 (N_8017,N_7801,N_7946);
nor U8018 (N_8018,N_7982,N_7898);
xor U8019 (N_8019,N_7904,N_7913);
nand U8020 (N_8020,N_7839,N_7917);
and U8021 (N_8021,N_7852,N_7998);
nand U8022 (N_8022,N_7914,N_7849);
nand U8023 (N_8023,N_7949,N_7756);
or U8024 (N_8024,N_7893,N_7987);
nor U8025 (N_8025,N_7919,N_7915);
and U8026 (N_8026,N_7906,N_7977);
nand U8027 (N_8027,N_7790,N_7869);
and U8028 (N_8028,N_7955,N_7800);
nor U8029 (N_8029,N_7853,N_7887);
nor U8030 (N_8030,N_7805,N_7773);
xnor U8031 (N_8031,N_7813,N_7962);
xnor U8032 (N_8032,N_7837,N_7826);
nor U8033 (N_8033,N_7951,N_7842);
or U8034 (N_8034,N_7873,N_7870);
or U8035 (N_8035,N_7818,N_7920);
xor U8036 (N_8036,N_7959,N_7978);
nor U8037 (N_8037,N_7990,N_7963);
nand U8038 (N_8038,N_7832,N_7967);
nand U8039 (N_8039,N_7831,N_7792);
nor U8040 (N_8040,N_7848,N_7975);
nor U8041 (N_8041,N_7931,N_7754);
nor U8042 (N_8042,N_7774,N_7786);
and U8043 (N_8043,N_7938,N_7835);
nor U8044 (N_8044,N_7945,N_7966);
xor U8045 (N_8045,N_7807,N_7784);
and U8046 (N_8046,N_7929,N_7934);
xor U8047 (N_8047,N_7874,N_7823);
nor U8048 (N_8048,N_7863,N_7882);
or U8049 (N_8049,N_7937,N_7976);
xor U8050 (N_8050,N_7846,N_7866);
or U8051 (N_8051,N_7940,N_7803);
or U8052 (N_8052,N_7986,N_7857);
and U8053 (N_8053,N_7770,N_7802);
nor U8054 (N_8054,N_7833,N_7772);
nor U8055 (N_8055,N_7763,N_7935);
xor U8056 (N_8056,N_7824,N_7890);
xnor U8057 (N_8057,N_7993,N_7859);
nand U8058 (N_8058,N_7969,N_7750);
nand U8059 (N_8059,N_7796,N_7776);
nor U8060 (N_8060,N_7759,N_7972);
and U8061 (N_8061,N_7845,N_7755);
xnor U8062 (N_8062,N_7765,N_7862);
and U8063 (N_8063,N_7816,N_7891);
nand U8064 (N_8064,N_7948,N_7821);
nand U8065 (N_8065,N_7751,N_7791);
nand U8066 (N_8066,N_7960,N_7794);
xor U8067 (N_8067,N_7954,N_7936);
or U8068 (N_8068,N_7795,N_7974);
and U8069 (N_8069,N_7787,N_7970);
and U8070 (N_8070,N_7806,N_7880);
or U8071 (N_8071,N_7926,N_7855);
or U8072 (N_8072,N_7961,N_7864);
xnor U8073 (N_8073,N_7899,N_7834);
or U8074 (N_8074,N_7921,N_7973);
nor U8075 (N_8075,N_7782,N_7999);
nor U8076 (N_8076,N_7985,N_7902);
or U8077 (N_8077,N_7922,N_7753);
xnor U8078 (N_8078,N_7783,N_7861);
nand U8079 (N_8079,N_7881,N_7780);
nand U8080 (N_8080,N_7988,N_7996);
or U8081 (N_8081,N_7793,N_7927);
nor U8082 (N_8082,N_7916,N_7885);
xnor U8083 (N_8083,N_7814,N_7876);
nor U8084 (N_8084,N_7968,N_7918);
nor U8085 (N_8085,N_7953,N_7854);
nor U8086 (N_8086,N_7847,N_7757);
nor U8087 (N_8087,N_7771,N_7911);
and U8088 (N_8088,N_7879,N_7815);
and U8089 (N_8089,N_7838,N_7925);
xor U8090 (N_8090,N_7819,N_7896);
nor U8091 (N_8091,N_7924,N_7798);
or U8092 (N_8092,N_7843,N_7884);
xor U8093 (N_8093,N_7860,N_7836);
and U8094 (N_8094,N_7900,N_7878);
nand U8095 (N_8095,N_7775,N_7825);
nand U8096 (N_8096,N_7817,N_7907);
or U8097 (N_8097,N_7932,N_7768);
and U8098 (N_8098,N_7797,N_7892);
nor U8099 (N_8099,N_7809,N_7995);
and U8100 (N_8100,N_7840,N_7928);
xor U8101 (N_8101,N_7778,N_7897);
and U8102 (N_8102,N_7830,N_7767);
nor U8103 (N_8103,N_7804,N_7910);
or U8104 (N_8104,N_7875,N_7851);
or U8105 (N_8105,N_7894,N_7877);
nand U8106 (N_8106,N_7781,N_7964);
and U8107 (N_8107,N_7788,N_7956);
and U8108 (N_8108,N_7908,N_7844);
nand U8109 (N_8109,N_7810,N_7943);
nand U8110 (N_8110,N_7944,N_7888);
and U8111 (N_8111,N_7886,N_7939);
nor U8112 (N_8112,N_7779,N_7923);
or U8113 (N_8113,N_7752,N_7799);
nor U8114 (N_8114,N_7947,N_7912);
and U8115 (N_8115,N_7858,N_7764);
nor U8116 (N_8116,N_7909,N_7981);
xor U8117 (N_8117,N_7903,N_7812);
and U8118 (N_8118,N_7991,N_7820);
and U8119 (N_8119,N_7901,N_7997);
and U8120 (N_8120,N_7952,N_7950);
xnor U8121 (N_8121,N_7758,N_7789);
xnor U8122 (N_8122,N_7933,N_7808);
xnor U8123 (N_8123,N_7827,N_7889);
or U8124 (N_8124,N_7856,N_7841);
or U8125 (N_8125,N_7831,N_7939);
and U8126 (N_8126,N_7811,N_7823);
and U8127 (N_8127,N_7760,N_7996);
nand U8128 (N_8128,N_7811,N_7838);
and U8129 (N_8129,N_7970,N_7798);
nor U8130 (N_8130,N_7758,N_7944);
or U8131 (N_8131,N_7985,N_7836);
and U8132 (N_8132,N_7942,N_7993);
xnor U8133 (N_8133,N_7978,N_7948);
xnor U8134 (N_8134,N_7845,N_7981);
nor U8135 (N_8135,N_7753,N_7946);
and U8136 (N_8136,N_7833,N_7973);
xor U8137 (N_8137,N_7828,N_7777);
nand U8138 (N_8138,N_7848,N_7765);
nor U8139 (N_8139,N_7788,N_7761);
xor U8140 (N_8140,N_7835,N_7817);
xor U8141 (N_8141,N_7943,N_7978);
xnor U8142 (N_8142,N_7894,N_7847);
and U8143 (N_8143,N_7946,N_7759);
and U8144 (N_8144,N_7858,N_7905);
nand U8145 (N_8145,N_7817,N_7781);
and U8146 (N_8146,N_7932,N_7848);
xor U8147 (N_8147,N_7893,N_7834);
nand U8148 (N_8148,N_7890,N_7787);
and U8149 (N_8149,N_7988,N_7837);
or U8150 (N_8150,N_7756,N_7932);
nand U8151 (N_8151,N_7896,N_7792);
and U8152 (N_8152,N_7971,N_7904);
nand U8153 (N_8153,N_7957,N_7874);
and U8154 (N_8154,N_7775,N_7996);
and U8155 (N_8155,N_7949,N_7817);
nor U8156 (N_8156,N_7961,N_7825);
or U8157 (N_8157,N_7756,N_7953);
or U8158 (N_8158,N_7770,N_7896);
xor U8159 (N_8159,N_7751,N_7963);
and U8160 (N_8160,N_7753,N_7927);
and U8161 (N_8161,N_7767,N_7815);
xnor U8162 (N_8162,N_7979,N_7893);
nor U8163 (N_8163,N_7787,N_7834);
xor U8164 (N_8164,N_7915,N_7765);
xnor U8165 (N_8165,N_7826,N_7982);
or U8166 (N_8166,N_7788,N_7851);
nand U8167 (N_8167,N_7806,N_7809);
nand U8168 (N_8168,N_7865,N_7956);
nand U8169 (N_8169,N_7878,N_7905);
and U8170 (N_8170,N_7785,N_7794);
nor U8171 (N_8171,N_7906,N_7843);
or U8172 (N_8172,N_7993,N_7939);
nor U8173 (N_8173,N_7873,N_7981);
nand U8174 (N_8174,N_7971,N_7925);
xor U8175 (N_8175,N_7888,N_7852);
nor U8176 (N_8176,N_7826,N_7798);
nor U8177 (N_8177,N_7805,N_7989);
and U8178 (N_8178,N_7862,N_7915);
nand U8179 (N_8179,N_7791,N_7767);
and U8180 (N_8180,N_7781,N_7895);
xnor U8181 (N_8181,N_7927,N_7923);
nor U8182 (N_8182,N_7999,N_7754);
and U8183 (N_8183,N_7870,N_7894);
and U8184 (N_8184,N_7869,N_7927);
and U8185 (N_8185,N_7900,N_7846);
nand U8186 (N_8186,N_7847,N_7927);
nand U8187 (N_8187,N_7777,N_7949);
or U8188 (N_8188,N_7838,N_7994);
nor U8189 (N_8189,N_7772,N_7928);
xnor U8190 (N_8190,N_7751,N_7935);
nand U8191 (N_8191,N_7768,N_7981);
xnor U8192 (N_8192,N_7920,N_7911);
xor U8193 (N_8193,N_7984,N_7908);
nor U8194 (N_8194,N_7751,N_7973);
nor U8195 (N_8195,N_7870,N_7807);
xnor U8196 (N_8196,N_7781,N_7976);
and U8197 (N_8197,N_7751,N_7913);
and U8198 (N_8198,N_7769,N_7910);
or U8199 (N_8199,N_7953,N_7960);
or U8200 (N_8200,N_7962,N_7937);
nor U8201 (N_8201,N_7970,N_7891);
xor U8202 (N_8202,N_7799,N_7854);
or U8203 (N_8203,N_7864,N_7837);
and U8204 (N_8204,N_7807,N_7952);
or U8205 (N_8205,N_7892,N_7804);
nand U8206 (N_8206,N_7987,N_7796);
and U8207 (N_8207,N_7969,N_7898);
or U8208 (N_8208,N_7754,N_7886);
or U8209 (N_8209,N_7922,N_7940);
or U8210 (N_8210,N_7857,N_7991);
nand U8211 (N_8211,N_7886,N_7872);
xnor U8212 (N_8212,N_7984,N_7791);
or U8213 (N_8213,N_7861,N_7882);
nor U8214 (N_8214,N_7927,N_7766);
nand U8215 (N_8215,N_7995,N_7889);
nand U8216 (N_8216,N_7992,N_7921);
nand U8217 (N_8217,N_7995,N_7946);
xnor U8218 (N_8218,N_7949,N_7883);
xor U8219 (N_8219,N_7877,N_7916);
or U8220 (N_8220,N_7986,N_7910);
and U8221 (N_8221,N_7934,N_7780);
or U8222 (N_8222,N_7995,N_7773);
nand U8223 (N_8223,N_7904,N_7832);
nand U8224 (N_8224,N_7839,N_7933);
nor U8225 (N_8225,N_7832,N_7757);
nor U8226 (N_8226,N_7751,N_7801);
and U8227 (N_8227,N_7838,N_7885);
nor U8228 (N_8228,N_7799,N_7771);
and U8229 (N_8229,N_7843,N_7930);
or U8230 (N_8230,N_7796,N_7846);
nor U8231 (N_8231,N_7896,N_7979);
nand U8232 (N_8232,N_7908,N_7761);
and U8233 (N_8233,N_7810,N_7790);
xnor U8234 (N_8234,N_7901,N_7785);
xnor U8235 (N_8235,N_7963,N_7846);
and U8236 (N_8236,N_7936,N_7943);
or U8237 (N_8237,N_7753,N_7958);
xor U8238 (N_8238,N_7970,N_7799);
xor U8239 (N_8239,N_7833,N_7797);
and U8240 (N_8240,N_7851,N_7915);
or U8241 (N_8241,N_7947,N_7827);
nand U8242 (N_8242,N_7864,N_7890);
nor U8243 (N_8243,N_7997,N_7891);
or U8244 (N_8244,N_7872,N_7901);
nor U8245 (N_8245,N_7868,N_7904);
xnor U8246 (N_8246,N_7847,N_7834);
nor U8247 (N_8247,N_7794,N_7923);
nand U8248 (N_8248,N_7859,N_7969);
nor U8249 (N_8249,N_7838,N_7959);
nand U8250 (N_8250,N_8156,N_8196);
or U8251 (N_8251,N_8108,N_8098);
and U8252 (N_8252,N_8002,N_8168);
nand U8253 (N_8253,N_8165,N_8059);
or U8254 (N_8254,N_8241,N_8082);
xor U8255 (N_8255,N_8167,N_8062);
or U8256 (N_8256,N_8133,N_8183);
and U8257 (N_8257,N_8200,N_8112);
nand U8258 (N_8258,N_8026,N_8130);
xnor U8259 (N_8259,N_8153,N_8094);
and U8260 (N_8260,N_8069,N_8243);
nand U8261 (N_8261,N_8047,N_8131);
nor U8262 (N_8262,N_8093,N_8074);
or U8263 (N_8263,N_8143,N_8119);
and U8264 (N_8264,N_8234,N_8135);
xor U8265 (N_8265,N_8237,N_8212);
and U8266 (N_8266,N_8001,N_8027);
nand U8267 (N_8267,N_8189,N_8058);
nand U8268 (N_8268,N_8201,N_8091);
nand U8269 (N_8269,N_8157,N_8014);
xnor U8270 (N_8270,N_8194,N_8247);
xnor U8271 (N_8271,N_8046,N_8086);
nor U8272 (N_8272,N_8159,N_8177);
or U8273 (N_8273,N_8240,N_8096);
nor U8274 (N_8274,N_8104,N_8100);
nor U8275 (N_8275,N_8097,N_8042);
nand U8276 (N_8276,N_8012,N_8205);
nor U8277 (N_8277,N_8066,N_8206);
nand U8278 (N_8278,N_8077,N_8050);
or U8279 (N_8279,N_8102,N_8071);
xor U8280 (N_8280,N_8150,N_8184);
and U8281 (N_8281,N_8145,N_8182);
nand U8282 (N_8282,N_8217,N_8080);
nor U8283 (N_8283,N_8181,N_8161);
nor U8284 (N_8284,N_8016,N_8210);
nand U8285 (N_8285,N_8029,N_8079);
or U8286 (N_8286,N_8083,N_8054);
or U8287 (N_8287,N_8146,N_8129);
nand U8288 (N_8288,N_8176,N_8236);
or U8289 (N_8289,N_8211,N_8220);
nor U8290 (N_8290,N_8018,N_8073);
nand U8291 (N_8291,N_8137,N_8152);
and U8292 (N_8292,N_8036,N_8118);
or U8293 (N_8293,N_8034,N_8140);
or U8294 (N_8294,N_8171,N_8117);
nand U8295 (N_8295,N_8044,N_8224);
nand U8296 (N_8296,N_8185,N_8116);
and U8297 (N_8297,N_8215,N_8227);
xnor U8298 (N_8298,N_8110,N_8028);
nor U8299 (N_8299,N_8198,N_8221);
nor U8300 (N_8300,N_8040,N_8125);
or U8301 (N_8301,N_8008,N_8010);
nand U8302 (N_8302,N_8123,N_8070);
and U8303 (N_8303,N_8122,N_8005);
nor U8304 (N_8304,N_8192,N_8193);
nand U8305 (N_8305,N_8172,N_8126);
nand U8306 (N_8306,N_8090,N_8249);
nand U8307 (N_8307,N_8033,N_8208);
nand U8308 (N_8308,N_8158,N_8141);
nor U8309 (N_8309,N_8154,N_8056);
or U8310 (N_8310,N_8162,N_8085);
xnor U8311 (N_8311,N_8160,N_8178);
nor U8312 (N_8312,N_8191,N_8048);
nor U8313 (N_8313,N_8173,N_8007);
nor U8314 (N_8314,N_8095,N_8197);
xor U8315 (N_8315,N_8190,N_8127);
and U8316 (N_8316,N_8164,N_8052);
nand U8317 (N_8317,N_8246,N_8015);
nand U8318 (N_8318,N_8213,N_8017);
nor U8319 (N_8319,N_8128,N_8019);
and U8320 (N_8320,N_8120,N_8186);
nand U8321 (N_8321,N_8009,N_8105);
nand U8322 (N_8322,N_8216,N_8204);
nor U8323 (N_8323,N_8202,N_8113);
xnor U8324 (N_8324,N_8223,N_8004);
nand U8325 (N_8325,N_8031,N_8132);
xnor U8326 (N_8326,N_8057,N_8101);
nor U8327 (N_8327,N_8078,N_8068);
nor U8328 (N_8328,N_8169,N_8195);
nand U8329 (N_8329,N_8041,N_8013);
or U8330 (N_8330,N_8025,N_8021);
nor U8331 (N_8331,N_8003,N_8089);
nor U8332 (N_8332,N_8024,N_8148);
nand U8333 (N_8333,N_8239,N_8231);
nor U8334 (N_8334,N_8061,N_8238);
and U8335 (N_8335,N_8055,N_8006);
xor U8336 (N_8336,N_8228,N_8000);
nor U8337 (N_8337,N_8147,N_8179);
and U8338 (N_8338,N_8072,N_8138);
or U8339 (N_8339,N_8087,N_8106);
nor U8340 (N_8340,N_8244,N_8045);
and U8341 (N_8341,N_8115,N_8180);
or U8342 (N_8342,N_8235,N_8134);
and U8343 (N_8343,N_8114,N_8209);
nor U8344 (N_8344,N_8065,N_8092);
nand U8345 (N_8345,N_8030,N_8187);
nor U8346 (N_8346,N_8088,N_8219);
nand U8347 (N_8347,N_8060,N_8035);
nor U8348 (N_8348,N_8174,N_8037);
and U8349 (N_8349,N_8136,N_8099);
or U8350 (N_8350,N_8222,N_8225);
xnor U8351 (N_8351,N_8109,N_8032);
and U8352 (N_8352,N_8038,N_8107);
or U8353 (N_8353,N_8023,N_8230);
nand U8354 (N_8354,N_8170,N_8051);
nor U8355 (N_8355,N_8175,N_8139);
xnor U8356 (N_8356,N_8111,N_8242);
xnor U8357 (N_8357,N_8081,N_8075);
nand U8358 (N_8358,N_8039,N_8232);
nor U8359 (N_8359,N_8188,N_8218);
and U8360 (N_8360,N_8049,N_8064);
or U8361 (N_8361,N_8053,N_8199);
or U8362 (N_8362,N_8142,N_8020);
or U8363 (N_8363,N_8151,N_8245);
nor U8364 (N_8364,N_8063,N_8067);
nor U8365 (N_8365,N_8084,N_8226);
nand U8366 (N_8366,N_8043,N_8166);
nor U8367 (N_8367,N_8233,N_8011);
or U8368 (N_8368,N_8121,N_8203);
nor U8369 (N_8369,N_8163,N_8155);
xor U8370 (N_8370,N_8076,N_8229);
nor U8371 (N_8371,N_8144,N_8248);
and U8372 (N_8372,N_8103,N_8207);
nand U8373 (N_8373,N_8214,N_8124);
nor U8374 (N_8374,N_8149,N_8022);
nand U8375 (N_8375,N_8078,N_8053);
and U8376 (N_8376,N_8108,N_8142);
xor U8377 (N_8377,N_8080,N_8018);
nand U8378 (N_8378,N_8155,N_8012);
nand U8379 (N_8379,N_8051,N_8052);
xor U8380 (N_8380,N_8156,N_8189);
nor U8381 (N_8381,N_8144,N_8006);
nor U8382 (N_8382,N_8191,N_8136);
and U8383 (N_8383,N_8184,N_8022);
nand U8384 (N_8384,N_8242,N_8011);
and U8385 (N_8385,N_8059,N_8139);
or U8386 (N_8386,N_8055,N_8177);
nor U8387 (N_8387,N_8015,N_8046);
xor U8388 (N_8388,N_8247,N_8235);
nor U8389 (N_8389,N_8074,N_8222);
nor U8390 (N_8390,N_8138,N_8065);
nor U8391 (N_8391,N_8144,N_8043);
xor U8392 (N_8392,N_8121,N_8048);
nor U8393 (N_8393,N_8000,N_8184);
or U8394 (N_8394,N_8198,N_8201);
or U8395 (N_8395,N_8078,N_8127);
and U8396 (N_8396,N_8076,N_8174);
nand U8397 (N_8397,N_8212,N_8029);
nand U8398 (N_8398,N_8004,N_8088);
or U8399 (N_8399,N_8014,N_8100);
xor U8400 (N_8400,N_8072,N_8005);
nor U8401 (N_8401,N_8096,N_8065);
nand U8402 (N_8402,N_8043,N_8225);
xnor U8403 (N_8403,N_8197,N_8134);
nand U8404 (N_8404,N_8069,N_8079);
or U8405 (N_8405,N_8099,N_8025);
nor U8406 (N_8406,N_8205,N_8127);
nand U8407 (N_8407,N_8168,N_8232);
xnor U8408 (N_8408,N_8060,N_8069);
nor U8409 (N_8409,N_8204,N_8122);
xnor U8410 (N_8410,N_8202,N_8117);
xnor U8411 (N_8411,N_8138,N_8146);
nor U8412 (N_8412,N_8165,N_8128);
or U8413 (N_8413,N_8114,N_8073);
nor U8414 (N_8414,N_8050,N_8194);
xnor U8415 (N_8415,N_8049,N_8081);
nand U8416 (N_8416,N_8126,N_8093);
or U8417 (N_8417,N_8071,N_8059);
nor U8418 (N_8418,N_8220,N_8169);
nand U8419 (N_8419,N_8025,N_8126);
xor U8420 (N_8420,N_8247,N_8160);
xnor U8421 (N_8421,N_8205,N_8178);
and U8422 (N_8422,N_8173,N_8146);
or U8423 (N_8423,N_8155,N_8018);
nand U8424 (N_8424,N_8049,N_8135);
xor U8425 (N_8425,N_8150,N_8103);
and U8426 (N_8426,N_8137,N_8059);
and U8427 (N_8427,N_8017,N_8196);
and U8428 (N_8428,N_8117,N_8125);
xnor U8429 (N_8429,N_8147,N_8053);
or U8430 (N_8430,N_8152,N_8040);
or U8431 (N_8431,N_8004,N_8061);
nand U8432 (N_8432,N_8106,N_8248);
or U8433 (N_8433,N_8166,N_8238);
nand U8434 (N_8434,N_8141,N_8122);
and U8435 (N_8435,N_8105,N_8036);
or U8436 (N_8436,N_8114,N_8160);
xnor U8437 (N_8437,N_8226,N_8172);
and U8438 (N_8438,N_8076,N_8206);
nand U8439 (N_8439,N_8012,N_8020);
nand U8440 (N_8440,N_8016,N_8047);
nor U8441 (N_8441,N_8149,N_8154);
xnor U8442 (N_8442,N_8174,N_8241);
xnor U8443 (N_8443,N_8034,N_8151);
xor U8444 (N_8444,N_8237,N_8058);
nand U8445 (N_8445,N_8159,N_8019);
and U8446 (N_8446,N_8159,N_8188);
or U8447 (N_8447,N_8101,N_8073);
nor U8448 (N_8448,N_8152,N_8087);
xor U8449 (N_8449,N_8202,N_8111);
and U8450 (N_8450,N_8051,N_8102);
xor U8451 (N_8451,N_8240,N_8014);
or U8452 (N_8452,N_8140,N_8061);
nor U8453 (N_8453,N_8139,N_8174);
xnor U8454 (N_8454,N_8174,N_8213);
xor U8455 (N_8455,N_8024,N_8111);
nor U8456 (N_8456,N_8127,N_8097);
and U8457 (N_8457,N_8169,N_8056);
nor U8458 (N_8458,N_8050,N_8216);
nand U8459 (N_8459,N_8133,N_8161);
or U8460 (N_8460,N_8123,N_8117);
and U8461 (N_8461,N_8054,N_8174);
and U8462 (N_8462,N_8061,N_8001);
xnor U8463 (N_8463,N_8132,N_8152);
nand U8464 (N_8464,N_8192,N_8009);
and U8465 (N_8465,N_8110,N_8032);
nor U8466 (N_8466,N_8214,N_8023);
or U8467 (N_8467,N_8238,N_8062);
nor U8468 (N_8468,N_8143,N_8089);
nand U8469 (N_8469,N_8035,N_8014);
or U8470 (N_8470,N_8030,N_8221);
or U8471 (N_8471,N_8193,N_8160);
nor U8472 (N_8472,N_8134,N_8246);
or U8473 (N_8473,N_8054,N_8031);
and U8474 (N_8474,N_8041,N_8185);
xor U8475 (N_8475,N_8194,N_8161);
nor U8476 (N_8476,N_8222,N_8082);
nand U8477 (N_8477,N_8214,N_8248);
nor U8478 (N_8478,N_8070,N_8014);
xor U8479 (N_8479,N_8201,N_8062);
or U8480 (N_8480,N_8147,N_8155);
nor U8481 (N_8481,N_8125,N_8058);
nand U8482 (N_8482,N_8033,N_8201);
nand U8483 (N_8483,N_8093,N_8220);
and U8484 (N_8484,N_8237,N_8150);
nor U8485 (N_8485,N_8165,N_8108);
or U8486 (N_8486,N_8177,N_8013);
or U8487 (N_8487,N_8011,N_8179);
and U8488 (N_8488,N_8065,N_8174);
or U8489 (N_8489,N_8058,N_8230);
xor U8490 (N_8490,N_8243,N_8035);
xor U8491 (N_8491,N_8056,N_8170);
nor U8492 (N_8492,N_8056,N_8104);
or U8493 (N_8493,N_8155,N_8159);
and U8494 (N_8494,N_8083,N_8178);
nor U8495 (N_8495,N_8071,N_8007);
or U8496 (N_8496,N_8184,N_8193);
nor U8497 (N_8497,N_8194,N_8127);
nor U8498 (N_8498,N_8175,N_8167);
or U8499 (N_8499,N_8019,N_8142);
nor U8500 (N_8500,N_8468,N_8335);
xnor U8501 (N_8501,N_8277,N_8326);
xnor U8502 (N_8502,N_8453,N_8374);
or U8503 (N_8503,N_8255,N_8430);
and U8504 (N_8504,N_8319,N_8438);
nand U8505 (N_8505,N_8352,N_8300);
xnor U8506 (N_8506,N_8369,N_8309);
or U8507 (N_8507,N_8336,N_8279);
xnor U8508 (N_8508,N_8350,N_8486);
nor U8509 (N_8509,N_8351,N_8473);
nor U8510 (N_8510,N_8261,N_8358);
nor U8511 (N_8511,N_8435,N_8334);
or U8512 (N_8512,N_8410,N_8490);
nor U8513 (N_8513,N_8362,N_8411);
and U8514 (N_8514,N_8429,N_8360);
or U8515 (N_8515,N_8479,N_8390);
and U8516 (N_8516,N_8316,N_8339);
nand U8517 (N_8517,N_8408,N_8443);
nand U8518 (N_8518,N_8270,N_8424);
and U8519 (N_8519,N_8320,N_8493);
and U8520 (N_8520,N_8262,N_8268);
nand U8521 (N_8521,N_8302,N_8396);
nand U8522 (N_8522,N_8449,N_8275);
nand U8523 (N_8523,N_8381,N_8426);
and U8524 (N_8524,N_8285,N_8394);
nand U8525 (N_8525,N_8422,N_8367);
nand U8526 (N_8526,N_8370,N_8444);
and U8527 (N_8527,N_8323,N_8273);
and U8528 (N_8528,N_8330,N_8264);
xnor U8529 (N_8529,N_8256,N_8445);
xor U8530 (N_8530,N_8483,N_8318);
and U8531 (N_8531,N_8492,N_8417);
nand U8532 (N_8532,N_8267,N_8494);
xnor U8533 (N_8533,N_8375,N_8291);
nor U8534 (N_8534,N_8254,N_8398);
and U8535 (N_8535,N_8299,N_8383);
xnor U8536 (N_8536,N_8402,N_8372);
or U8537 (N_8537,N_8481,N_8466);
nor U8538 (N_8538,N_8377,N_8333);
nor U8539 (N_8539,N_8469,N_8345);
nand U8540 (N_8540,N_8293,N_8471);
or U8541 (N_8541,N_8423,N_8365);
xnor U8542 (N_8542,N_8271,N_8458);
xor U8543 (N_8543,N_8400,N_8265);
xor U8544 (N_8544,N_8373,N_8361);
nand U8545 (N_8545,N_8322,N_8329);
nor U8546 (N_8546,N_8354,N_8464);
or U8547 (N_8547,N_8437,N_8306);
or U8548 (N_8548,N_8287,N_8407);
nor U8549 (N_8549,N_8272,N_8263);
nor U8550 (N_8550,N_8276,N_8484);
xnor U8551 (N_8551,N_8455,N_8491);
xnor U8552 (N_8552,N_8399,N_8462);
xor U8553 (N_8553,N_8310,N_8414);
nor U8554 (N_8554,N_8363,N_8477);
nor U8555 (N_8555,N_8295,N_8465);
nand U8556 (N_8556,N_8496,N_8340);
xnor U8557 (N_8557,N_8253,N_8406);
and U8558 (N_8558,N_8397,N_8257);
nor U8559 (N_8559,N_8405,N_8446);
xor U8560 (N_8560,N_8391,N_8431);
nand U8561 (N_8561,N_8298,N_8342);
xnor U8562 (N_8562,N_8301,N_8482);
xor U8563 (N_8563,N_8280,N_8393);
xor U8564 (N_8564,N_8454,N_8448);
and U8565 (N_8565,N_8376,N_8344);
xor U8566 (N_8566,N_8284,N_8353);
nand U8567 (N_8567,N_8480,N_8368);
or U8568 (N_8568,N_8495,N_8337);
or U8569 (N_8569,N_8409,N_8389);
nand U8570 (N_8570,N_8380,N_8425);
or U8571 (N_8571,N_8436,N_8307);
and U8572 (N_8572,N_8379,N_8382);
nor U8573 (N_8573,N_8488,N_8331);
nand U8574 (N_8574,N_8341,N_8364);
xnor U8575 (N_8575,N_8392,N_8413);
nor U8576 (N_8576,N_8324,N_8415);
xor U8577 (N_8577,N_8290,N_8489);
and U8578 (N_8578,N_8314,N_8266);
nor U8579 (N_8579,N_8269,N_8348);
xor U8580 (N_8580,N_8434,N_8321);
nor U8581 (N_8581,N_8499,N_8378);
nand U8582 (N_8582,N_8470,N_8259);
nand U8583 (N_8583,N_8292,N_8359);
and U8584 (N_8584,N_8476,N_8343);
and U8585 (N_8585,N_8250,N_8467);
xor U8586 (N_8586,N_8311,N_8487);
nand U8587 (N_8587,N_8432,N_8404);
or U8588 (N_8588,N_8451,N_8447);
xor U8589 (N_8589,N_8427,N_8441);
nand U8590 (N_8590,N_8297,N_8459);
nand U8591 (N_8591,N_8303,N_8385);
nand U8592 (N_8592,N_8286,N_8401);
xor U8593 (N_8593,N_8428,N_8356);
and U8594 (N_8594,N_8288,N_8327);
and U8595 (N_8595,N_8463,N_8283);
or U8596 (N_8596,N_8420,N_8371);
nor U8597 (N_8597,N_8384,N_8472);
nand U8598 (N_8598,N_8366,N_8421);
or U8599 (N_8599,N_8251,N_8294);
nor U8600 (N_8600,N_8403,N_8386);
nand U8601 (N_8601,N_8328,N_8418);
and U8602 (N_8602,N_8289,N_8274);
nand U8603 (N_8603,N_8497,N_8474);
or U8604 (N_8604,N_8457,N_8498);
or U8605 (N_8605,N_8315,N_8304);
nand U8606 (N_8606,N_8452,N_8349);
nor U8607 (N_8607,N_8433,N_8419);
or U8608 (N_8608,N_8347,N_8282);
nor U8609 (N_8609,N_8258,N_8317);
and U8610 (N_8610,N_8260,N_8325);
xor U8611 (N_8611,N_8450,N_8355);
or U8612 (N_8612,N_8305,N_8461);
xnor U8613 (N_8613,N_8460,N_8478);
or U8614 (N_8614,N_8395,N_8412);
nand U8615 (N_8615,N_8485,N_8442);
nor U8616 (N_8616,N_8456,N_8281);
and U8617 (N_8617,N_8357,N_8346);
nand U8618 (N_8618,N_8475,N_8416);
xnor U8619 (N_8619,N_8439,N_8252);
or U8620 (N_8620,N_8332,N_8387);
nand U8621 (N_8621,N_8308,N_8312);
or U8622 (N_8622,N_8313,N_8388);
or U8623 (N_8623,N_8278,N_8338);
nand U8624 (N_8624,N_8440,N_8296);
or U8625 (N_8625,N_8283,N_8304);
nand U8626 (N_8626,N_8481,N_8396);
nand U8627 (N_8627,N_8255,N_8330);
or U8628 (N_8628,N_8348,N_8295);
or U8629 (N_8629,N_8250,N_8476);
nor U8630 (N_8630,N_8296,N_8458);
xnor U8631 (N_8631,N_8436,N_8315);
nor U8632 (N_8632,N_8462,N_8366);
nor U8633 (N_8633,N_8440,N_8338);
xor U8634 (N_8634,N_8380,N_8486);
nand U8635 (N_8635,N_8393,N_8257);
nand U8636 (N_8636,N_8464,N_8431);
or U8637 (N_8637,N_8278,N_8481);
and U8638 (N_8638,N_8262,N_8461);
and U8639 (N_8639,N_8334,N_8439);
nand U8640 (N_8640,N_8490,N_8251);
and U8641 (N_8641,N_8373,N_8318);
and U8642 (N_8642,N_8328,N_8364);
or U8643 (N_8643,N_8389,N_8366);
xor U8644 (N_8644,N_8413,N_8473);
and U8645 (N_8645,N_8254,N_8488);
nand U8646 (N_8646,N_8467,N_8327);
or U8647 (N_8647,N_8459,N_8478);
nor U8648 (N_8648,N_8424,N_8354);
and U8649 (N_8649,N_8471,N_8466);
and U8650 (N_8650,N_8328,N_8412);
nor U8651 (N_8651,N_8276,N_8415);
and U8652 (N_8652,N_8427,N_8489);
or U8653 (N_8653,N_8464,N_8383);
or U8654 (N_8654,N_8466,N_8413);
nor U8655 (N_8655,N_8385,N_8410);
xor U8656 (N_8656,N_8290,N_8413);
xor U8657 (N_8657,N_8413,N_8332);
and U8658 (N_8658,N_8280,N_8296);
and U8659 (N_8659,N_8268,N_8378);
nand U8660 (N_8660,N_8388,N_8464);
and U8661 (N_8661,N_8303,N_8314);
or U8662 (N_8662,N_8270,N_8287);
nand U8663 (N_8663,N_8418,N_8452);
nor U8664 (N_8664,N_8431,N_8253);
xnor U8665 (N_8665,N_8287,N_8333);
and U8666 (N_8666,N_8362,N_8398);
xnor U8667 (N_8667,N_8465,N_8466);
or U8668 (N_8668,N_8407,N_8305);
or U8669 (N_8669,N_8279,N_8304);
nor U8670 (N_8670,N_8287,N_8362);
nand U8671 (N_8671,N_8478,N_8291);
and U8672 (N_8672,N_8253,N_8342);
or U8673 (N_8673,N_8353,N_8444);
and U8674 (N_8674,N_8399,N_8389);
nand U8675 (N_8675,N_8365,N_8396);
or U8676 (N_8676,N_8391,N_8274);
or U8677 (N_8677,N_8388,N_8448);
nor U8678 (N_8678,N_8342,N_8410);
nor U8679 (N_8679,N_8333,N_8283);
or U8680 (N_8680,N_8257,N_8459);
or U8681 (N_8681,N_8375,N_8334);
xor U8682 (N_8682,N_8283,N_8445);
nand U8683 (N_8683,N_8428,N_8277);
or U8684 (N_8684,N_8387,N_8306);
and U8685 (N_8685,N_8257,N_8479);
nand U8686 (N_8686,N_8358,N_8305);
and U8687 (N_8687,N_8433,N_8266);
nor U8688 (N_8688,N_8462,N_8406);
nor U8689 (N_8689,N_8478,N_8334);
or U8690 (N_8690,N_8498,N_8410);
and U8691 (N_8691,N_8480,N_8417);
nand U8692 (N_8692,N_8303,N_8459);
nor U8693 (N_8693,N_8347,N_8396);
and U8694 (N_8694,N_8384,N_8279);
xor U8695 (N_8695,N_8418,N_8274);
nor U8696 (N_8696,N_8406,N_8414);
nor U8697 (N_8697,N_8379,N_8489);
and U8698 (N_8698,N_8381,N_8484);
and U8699 (N_8699,N_8260,N_8344);
nor U8700 (N_8700,N_8396,N_8288);
nor U8701 (N_8701,N_8431,N_8429);
nor U8702 (N_8702,N_8340,N_8365);
xnor U8703 (N_8703,N_8395,N_8424);
xor U8704 (N_8704,N_8456,N_8446);
nor U8705 (N_8705,N_8304,N_8324);
and U8706 (N_8706,N_8465,N_8417);
nand U8707 (N_8707,N_8274,N_8310);
nor U8708 (N_8708,N_8263,N_8356);
xor U8709 (N_8709,N_8339,N_8276);
xor U8710 (N_8710,N_8340,N_8329);
or U8711 (N_8711,N_8376,N_8411);
xor U8712 (N_8712,N_8399,N_8337);
nor U8713 (N_8713,N_8436,N_8250);
and U8714 (N_8714,N_8363,N_8303);
nand U8715 (N_8715,N_8300,N_8375);
nand U8716 (N_8716,N_8396,N_8269);
nand U8717 (N_8717,N_8397,N_8461);
or U8718 (N_8718,N_8482,N_8256);
and U8719 (N_8719,N_8320,N_8362);
and U8720 (N_8720,N_8413,N_8388);
nand U8721 (N_8721,N_8354,N_8285);
nand U8722 (N_8722,N_8497,N_8338);
nor U8723 (N_8723,N_8485,N_8462);
xnor U8724 (N_8724,N_8441,N_8467);
nand U8725 (N_8725,N_8472,N_8357);
or U8726 (N_8726,N_8279,N_8460);
xnor U8727 (N_8727,N_8346,N_8364);
or U8728 (N_8728,N_8357,N_8395);
nor U8729 (N_8729,N_8417,N_8330);
and U8730 (N_8730,N_8419,N_8453);
xnor U8731 (N_8731,N_8476,N_8298);
or U8732 (N_8732,N_8435,N_8372);
and U8733 (N_8733,N_8272,N_8407);
and U8734 (N_8734,N_8299,N_8496);
nor U8735 (N_8735,N_8464,N_8401);
or U8736 (N_8736,N_8255,N_8272);
and U8737 (N_8737,N_8382,N_8281);
xor U8738 (N_8738,N_8263,N_8412);
nand U8739 (N_8739,N_8372,N_8468);
nor U8740 (N_8740,N_8463,N_8394);
nor U8741 (N_8741,N_8438,N_8299);
xor U8742 (N_8742,N_8338,N_8384);
and U8743 (N_8743,N_8291,N_8292);
xor U8744 (N_8744,N_8336,N_8499);
nand U8745 (N_8745,N_8386,N_8494);
nor U8746 (N_8746,N_8277,N_8292);
xnor U8747 (N_8747,N_8414,N_8334);
and U8748 (N_8748,N_8259,N_8320);
nand U8749 (N_8749,N_8436,N_8440);
and U8750 (N_8750,N_8524,N_8554);
or U8751 (N_8751,N_8690,N_8523);
or U8752 (N_8752,N_8666,N_8585);
and U8753 (N_8753,N_8742,N_8673);
nand U8754 (N_8754,N_8706,N_8534);
nor U8755 (N_8755,N_8711,N_8612);
and U8756 (N_8756,N_8705,N_8682);
and U8757 (N_8757,N_8719,N_8670);
nor U8758 (N_8758,N_8683,N_8736);
and U8759 (N_8759,N_8729,N_8631);
nand U8760 (N_8760,N_8727,N_8720);
and U8761 (N_8761,N_8616,N_8560);
nand U8762 (N_8762,N_8639,N_8595);
and U8763 (N_8763,N_8568,N_8532);
or U8764 (N_8764,N_8671,N_8714);
nor U8765 (N_8765,N_8618,N_8624);
nor U8766 (N_8766,N_8702,N_8712);
xor U8767 (N_8767,N_8621,N_8557);
nand U8768 (N_8768,N_8668,N_8544);
or U8769 (N_8769,N_8569,N_8541);
xnor U8770 (N_8770,N_8687,N_8520);
and U8771 (N_8771,N_8748,N_8698);
xnor U8772 (N_8772,N_8678,N_8741);
nand U8773 (N_8773,N_8578,N_8556);
nand U8774 (N_8774,N_8550,N_8649);
or U8775 (N_8775,N_8635,N_8661);
and U8776 (N_8776,N_8732,N_8601);
nor U8777 (N_8777,N_8504,N_8725);
nand U8778 (N_8778,N_8521,N_8609);
nand U8779 (N_8779,N_8611,N_8610);
or U8780 (N_8780,N_8553,N_8630);
or U8781 (N_8781,N_8623,N_8652);
xnor U8782 (N_8782,N_8603,N_8708);
xnor U8783 (N_8783,N_8648,N_8703);
nand U8784 (N_8784,N_8655,N_8566);
nor U8785 (N_8785,N_8584,N_8679);
nor U8786 (N_8786,N_8562,N_8614);
and U8787 (N_8787,N_8509,N_8582);
and U8788 (N_8788,N_8604,N_8570);
nor U8789 (N_8789,N_8647,N_8626);
nor U8790 (N_8790,N_8519,N_8685);
xor U8791 (N_8791,N_8539,N_8564);
nor U8792 (N_8792,N_8575,N_8654);
xnor U8793 (N_8793,N_8695,N_8512);
and U8794 (N_8794,N_8625,N_8650);
or U8795 (N_8795,N_8726,N_8728);
xor U8796 (N_8796,N_8627,N_8571);
nand U8797 (N_8797,N_8583,N_8660);
xnor U8798 (N_8798,N_8597,N_8658);
nor U8799 (N_8799,N_8542,N_8596);
and U8800 (N_8800,N_8722,N_8589);
and U8801 (N_8801,N_8716,N_8530);
nand U8802 (N_8802,N_8573,N_8694);
nor U8803 (N_8803,N_8653,N_8528);
and U8804 (N_8804,N_8598,N_8591);
nand U8805 (N_8805,N_8500,N_8533);
nand U8806 (N_8806,N_8662,N_8574);
or U8807 (N_8807,N_8622,N_8738);
xor U8808 (N_8808,N_8517,N_8643);
nand U8809 (N_8809,N_8644,N_8718);
nor U8810 (N_8810,N_8681,N_8731);
nand U8811 (N_8811,N_8745,N_8592);
nand U8812 (N_8812,N_8527,N_8645);
nand U8813 (N_8813,N_8740,N_8669);
xnor U8814 (N_8814,N_8677,N_8563);
nand U8815 (N_8815,N_8508,N_8646);
nor U8816 (N_8816,N_8713,N_8619);
and U8817 (N_8817,N_8518,N_8700);
and U8818 (N_8818,N_8515,N_8565);
xnor U8819 (N_8819,N_8696,N_8540);
and U8820 (N_8820,N_8680,N_8739);
nand U8821 (N_8821,N_8674,N_8615);
nor U8822 (N_8822,N_8605,N_8513);
and U8823 (N_8823,N_8721,N_8663);
and U8824 (N_8824,N_8636,N_8723);
xnor U8825 (N_8825,N_8628,N_8510);
and U8826 (N_8826,N_8638,N_8665);
nand U8827 (N_8827,N_8581,N_8693);
or U8828 (N_8828,N_8737,N_8535);
or U8829 (N_8829,N_8749,N_8559);
and U8830 (N_8830,N_8522,N_8561);
nand U8831 (N_8831,N_8642,N_8529);
or U8832 (N_8832,N_8593,N_8686);
nor U8833 (N_8833,N_8548,N_8735);
nor U8834 (N_8834,N_8617,N_8600);
nor U8835 (N_8835,N_8697,N_8538);
and U8836 (N_8836,N_8699,N_8608);
and U8837 (N_8837,N_8733,N_8709);
nand U8838 (N_8838,N_8701,N_8545);
and U8839 (N_8839,N_8606,N_8715);
nor U8840 (N_8840,N_8667,N_8594);
nor U8841 (N_8841,N_8501,N_8507);
or U8842 (N_8842,N_8546,N_8531);
nand U8843 (N_8843,N_8558,N_8576);
nor U8844 (N_8844,N_8551,N_8730);
nand U8845 (N_8845,N_8525,N_8704);
nand U8846 (N_8846,N_8580,N_8641);
xnor U8847 (N_8847,N_8613,N_8511);
nand U8848 (N_8848,N_8744,N_8637);
nand U8849 (N_8849,N_8657,N_8526);
xor U8850 (N_8850,N_8692,N_8688);
nor U8851 (N_8851,N_8675,N_8676);
nor U8852 (N_8852,N_8514,N_8572);
nand U8853 (N_8853,N_8746,N_8710);
nor U8854 (N_8854,N_8633,N_8691);
xnor U8855 (N_8855,N_8543,N_8640);
and U8856 (N_8856,N_8689,N_8634);
xnor U8857 (N_8857,N_8724,N_8664);
nand U8858 (N_8858,N_8629,N_8549);
and U8859 (N_8859,N_8586,N_8579);
nand U8860 (N_8860,N_8684,N_8602);
nand U8861 (N_8861,N_8672,N_8743);
nand U8862 (N_8862,N_8656,N_8567);
nand U8863 (N_8863,N_8659,N_8632);
nor U8864 (N_8864,N_8620,N_8651);
and U8865 (N_8865,N_8536,N_8607);
and U8866 (N_8866,N_8587,N_8503);
nor U8867 (N_8867,N_8506,N_8537);
and U8868 (N_8868,N_8590,N_8577);
nor U8869 (N_8869,N_8547,N_8734);
xnor U8870 (N_8870,N_8555,N_8505);
xor U8871 (N_8871,N_8747,N_8707);
nor U8872 (N_8872,N_8552,N_8717);
nand U8873 (N_8873,N_8516,N_8588);
or U8874 (N_8874,N_8599,N_8502);
xnor U8875 (N_8875,N_8749,N_8659);
nor U8876 (N_8876,N_8669,N_8714);
or U8877 (N_8877,N_8665,N_8539);
xnor U8878 (N_8878,N_8676,N_8661);
and U8879 (N_8879,N_8557,N_8591);
nor U8880 (N_8880,N_8541,N_8640);
and U8881 (N_8881,N_8590,N_8632);
nand U8882 (N_8882,N_8592,N_8590);
nor U8883 (N_8883,N_8501,N_8565);
nand U8884 (N_8884,N_8540,N_8691);
xor U8885 (N_8885,N_8669,N_8736);
nand U8886 (N_8886,N_8524,N_8629);
and U8887 (N_8887,N_8532,N_8689);
or U8888 (N_8888,N_8528,N_8708);
nand U8889 (N_8889,N_8680,N_8595);
nand U8890 (N_8890,N_8545,N_8716);
or U8891 (N_8891,N_8511,N_8558);
nand U8892 (N_8892,N_8616,N_8732);
and U8893 (N_8893,N_8641,N_8737);
and U8894 (N_8894,N_8557,N_8665);
nand U8895 (N_8895,N_8673,N_8502);
xor U8896 (N_8896,N_8670,N_8612);
and U8897 (N_8897,N_8579,N_8679);
xnor U8898 (N_8898,N_8693,N_8587);
and U8899 (N_8899,N_8566,N_8596);
and U8900 (N_8900,N_8503,N_8703);
nand U8901 (N_8901,N_8702,N_8701);
xor U8902 (N_8902,N_8511,N_8749);
and U8903 (N_8903,N_8644,N_8633);
xor U8904 (N_8904,N_8654,N_8510);
nor U8905 (N_8905,N_8696,N_8662);
nand U8906 (N_8906,N_8746,N_8588);
xor U8907 (N_8907,N_8572,N_8707);
and U8908 (N_8908,N_8639,N_8622);
nor U8909 (N_8909,N_8569,N_8518);
nand U8910 (N_8910,N_8567,N_8678);
and U8911 (N_8911,N_8500,N_8589);
nor U8912 (N_8912,N_8532,N_8615);
or U8913 (N_8913,N_8732,N_8525);
and U8914 (N_8914,N_8540,N_8653);
nand U8915 (N_8915,N_8737,N_8541);
or U8916 (N_8916,N_8516,N_8697);
or U8917 (N_8917,N_8692,N_8611);
nor U8918 (N_8918,N_8625,N_8687);
or U8919 (N_8919,N_8711,N_8501);
and U8920 (N_8920,N_8513,N_8724);
or U8921 (N_8921,N_8639,N_8556);
xor U8922 (N_8922,N_8688,N_8563);
and U8923 (N_8923,N_8701,N_8732);
xor U8924 (N_8924,N_8607,N_8608);
xnor U8925 (N_8925,N_8551,N_8606);
and U8926 (N_8926,N_8666,N_8677);
nor U8927 (N_8927,N_8665,N_8719);
nor U8928 (N_8928,N_8513,N_8690);
nand U8929 (N_8929,N_8555,N_8531);
nor U8930 (N_8930,N_8609,N_8522);
or U8931 (N_8931,N_8629,N_8574);
and U8932 (N_8932,N_8635,N_8550);
nand U8933 (N_8933,N_8516,N_8565);
xnor U8934 (N_8934,N_8680,N_8584);
nand U8935 (N_8935,N_8742,N_8729);
or U8936 (N_8936,N_8516,N_8515);
nand U8937 (N_8937,N_8643,N_8627);
or U8938 (N_8938,N_8706,N_8626);
xor U8939 (N_8939,N_8577,N_8670);
nand U8940 (N_8940,N_8708,N_8740);
nor U8941 (N_8941,N_8669,N_8630);
and U8942 (N_8942,N_8695,N_8555);
nand U8943 (N_8943,N_8707,N_8602);
nor U8944 (N_8944,N_8744,N_8574);
nand U8945 (N_8945,N_8731,N_8615);
nor U8946 (N_8946,N_8613,N_8652);
or U8947 (N_8947,N_8656,N_8632);
and U8948 (N_8948,N_8609,N_8667);
nor U8949 (N_8949,N_8742,N_8619);
or U8950 (N_8950,N_8738,N_8540);
xnor U8951 (N_8951,N_8621,N_8538);
nand U8952 (N_8952,N_8627,N_8650);
and U8953 (N_8953,N_8686,N_8708);
nor U8954 (N_8954,N_8650,N_8702);
and U8955 (N_8955,N_8614,N_8609);
nand U8956 (N_8956,N_8572,N_8622);
or U8957 (N_8957,N_8524,N_8666);
and U8958 (N_8958,N_8558,N_8521);
nor U8959 (N_8959,N_8667,N_8683);
and U8960 (N_8960,N_8574,N_8522);
xnor U8961 (N_8961,N_8563,N_8587);
nand U8962 (N_8962,N_8697,N_8650);
and U8963 (N_8963,N_8613,N_8506);
nand U8964 (N_8964,N_8695,N_8640);
nor U8965 (N_8965,N_8731,N_8551);
and U8966 (N_8966,N_8723,N_8654);
xor U8967 (N_8967,N_8683,N_8706);
nor U8968 (N_8968,N_8534,N_8616);
nand U8969 (N_8969,N_8557,N_8683);
and U8970 (N_8970,N_8697,N_8659);
nand U8971 (N_8971,N_8616,N_8531);
nor U8972 (N_8972,N_8727,N_8568);
nand U8973 (N_8973,N_8651,N_8528);
xnor U8974 (N_8974,N_8738,N_8532);
and U8975 (N_8975,N_8585,N_8517);
nand U8976 (N_8976,N_8740,N_8714);
nand U8977 (N_8977,N_8526,N_8622);
or U8978 (N_8978,N_8557,N_8708);
nor U8979 (N_8979,N_8694,N_8662);
nand U8980 (N_8980,N_8719,N_8724);
and U8981 (N_8981,N_8601,N_8506);
nor U8982 (N_8982,N_8703,N_8686);
or U8983 (N_8983,N_8680,N_8555);
nor U8984 (N_8984,N_8503,N_8737);
nor U8985 (N_8985,N_8534,N_8700);
nor U8986 (N_8986,N_8617,N_8550);
nor U8987 (N_8987,N_8715,N_8680);
and U8988 (N_8988,N_8651,N_8677);
and U8989 (N_8989,N_8681,N_8629);
or U8990 (N_8990,N_8624,N_8530);
nor U8991 (N_8991,N_8632,N_8554);
or U8992 (N_8992,N_8748,N_8575);
nand U8993 (N_8993,N_8677,N_8616);
and U8994 (N_8994,N_8609,N_8633);
and U8995 (N_8995,N_8582,N_8661);
nand U8996 (N_8996,N_8526,N_8740);
xnor U8997 (N_8997,N_8576,N_8728);
nand U8998 (N_8998,N_8745,N_8590);
or U8999 (N_8999,N_8682,N_8645);
nand U9000 (N_9000,N_8789,N_8858);
xor U9001 (N_9001,N_8765,N_8953);
or U9002 (N_9002,N_8818,N_8831);
nor U9003 (N_9003,N_8905,N_8879);
xor U9004 (N_9004,N_8780,N_8988);
or U9005 (N_9005,N_8984,N_8929);
nand U9006 (N_9006,N_8906,N_8894);
and U9007 (N_9007,N_8882,N_8811);
and U9008 (N_9008,N_8951,N_8838);
and U9009 (N_9009,N_8813,N_8790);
nand U9010 (N_9010,N_8852,N_8792);
xnor U9011 (N_9011,N_8812,N_8981);
nand U9012 (N_9012,N_8952,N_8799);
nand U9013 (N_9013,N_8753,N_8870);
or U9014 (N_9014,N_8846,N_8786);
or U9015 (N_9015,N_8986,N_8793);
xnor U9016 (N_9016,N_8758,N_8903);
nand U9017 (N_9017,N_8755,N_8943);
and U9018 (N_9018,N_8805,N_8817);
and U9019 (N_9019,N_8841,N_8955);
and U9020 (N_9020,N_8759,N_8830);
xnor U9021 (N_9021,N_8959,N_8787);
or U9022 (N_9022,N_8828,N_8993);
or U9023 (N_9023,N_8960,N_8990);
xor U9024 (N_9024,N_8938,N_8750);
or U9025 (N_9025,N_8992,N_8770);
nand U9026 (N_9026,N_8756,N_8874);
nor U9027 (N_9027,N_8883,N_8875);
or U9028 (N_9028,N_8829,N_8801);
and U9029 (N_9029,N_8784,N_8900);
xnor U9030 (N_9030,N_8816,N_8810);
xnor U9031 (N_9031,N_8800,N_8954);
xor U9032 (N_9032,N_8980,N_8978);
or U9033 (N_9033,N_8845,N_8933);
xnor U9034 (N_9034,N_8809,N_8989);
nor U9035 (N_9035,N_8766,N_8934);
nor U9036 (N_9036,N_8824,N_8998);
nand U9037 (N_9037,N_8917,N_8876);
or U9038 (N_9038,N_8827,N_8968);
and U9039 (N_9039,N_8888,N_8956);
nor U9040 (N_9040,N_8898,N_8864);
xnor U9041 (N_9041,N_8791,N_8921);
nor U9042 (N_9042,N_8947,N_8842);
xor U9043 (N_9043,N_8868,N_8839);
nand U9044 (N_9044,N_8871,N_8856);
nand U9045 (N_9045,N_8872,N_8859);
xnor U9046 (N_9046,N_8946,N_8886);
nor U9047 (N_9047,N_8971,N_8918);
or U9048 (N_9048,N_8797,N_8863);
xnor U9049 (N_9049,N_8969,N_8957);
nor U9050 (N_9050,N_8849,N_8939);
nor U9051 (N_9051,N_8979,N_8944);
nand U9052 (N_9052,N_8865,N_8774);
and U9053 (N_9053,N_8924,N_8814);
and U9054 (N_9054,N_8950,N_8991);
or U9055 (N_9055,N_8823,N_8773);
nor U9056 (N_9056,N_8772,N_8974);
nand U9057 (N_9057,N_8945,N_8867);
xnor U9058 (N_9058,N_8808,N_8821);
and U9059 (N_9059,N_8776,N_8825);
nor U9060 (N_9060,N_8881,N_8923);
and U9061 (N_9061,N_8781,N_8912);
xor U9062 (N_9062,N_8994,N_8806);
or U9063 (N_9063,N_8893,N_8916);
nor U9064 (N_9064,N_8965,N_8822);
xor U9065 (N_9065,N_8930,N_8796);
or U9066 (N_9066,N_8885,N_8771);
and U9067 (N_9067,N_8832,N_8803);
nor U9068 (N_9068,N_8948,N_8995);
nor U9069 (N_9069,N_8795,N_8877);
or U9070 (N_9070,N_8804,N_8857);
or U9071 (N_9071,N_8985,N_8890);
and U9072 (N_9072,N_8764,N_8835);
and U9073 (N_9073,N_8785,N_8932);
and U9074 (N_9074,N_8925,N_8850);
and U9075 (N_9075,N_8937,N_8901);
and U9076 (N_9076,N_8826,N_8851);
nor U9077 (N_9077,N_8936,N_8982);
nand U9078 (N_9078,N_8909,N_8975);
nand U9079 (N_9079,N_8908,N_8961);
or U9080 (N_9080,N_8973,N_8884);
xnor U9081 (N_9081,N_8941,N_8895);
xnor U9082 (N_9082,N_8779,N_8862);
and U9083 (N_9083,N_8899,N_8880);
xnor U9084 (N_9084,N_8966,N_8997);
or U9085 (N_9085,N_8972,N_8802);
nand U9086 (N_9086,N_8942,N_8999);
xnor U9087 (N_9087,N_8920,N_8794);
and U9088 (N_9088,N_8949,N_8855);
nand U9089 (N_9089,N_8889,N_8887);
nor U9090 (N_9090,N_8757,N_8987);
and U9091 (N_9091,N_8977,N_8854);
nor U9092 (N_9092,N_8815,N_8983);
or U9093 (N_9093,N_8844,N_8913);
nor U9094 (N_9094,N_8807,N_8861);
nor U9095 (N_9095,N_8798,N_8964);
and U9096 (N_9096,N_8919,N_8904);
xor U9097 (N_9097,N_8928,N_8860);
or U9098 (N_9098,N_8922,N_8970);
nor U9099 (N_9099,N_8902,N_8848);
nor U9100 (N_9100,N_8878,N_8763);
or U9101 (N_9101,N_8834,N_8783);
xnor U9102 (N_9102,N_8915,N_8940);
nand U9103 (N_9103,N_8896,N_8976);
or U9104 (N_9104,N_8927,N_8958);
nand U9105 (N_9105,N_8847,N_8931);
xor U9106 (N_9106,N_8996,N_8840);
nor U9107 (N_9107,N_8820,N_8962);
and U9108 (N_9108,N_8914,N_8926);
xor U9109 (N_9109,N_8754,N_8775);
nand U9110 (N_9110,N_8767,N_8760);
nor U9111 (N_9111,N_8761,N_8911);
nor U9112 (N_9112,N_8836,N_8910);
or U9113 (N_9113,N_8778,N_8897);
or U9114 (N_9114,N_8843,N_8782);
or U9115 (N_9115,N_8752,N_8768);
and U9116 (N_9116,N_8869,N_8891);
and U9117 (N_9117,N_8892,N_8769);
or U9118 (N_9118,N_8853,N_8935);
xor U9119 (N_9119,N_8837,N_8866);
nand U9120 (N_9120,N_8762,N_8751);
and U9121 (N_9121,N_8777,N_8788);
nor U9122 (N_9122,N_8907,N_8963);
nand U9123 (N_9123,N_8819,N_8873);
and U9124 (N_9124,N_8967,N_8833);
xor U9125 (N_9125,N_8983,N_8899);
xnor U9126 (N_9126,N_8921,N_8959);
nand U9127 (N_9127,N_8806,N_8909);
xor U9128 (N_9128,N_8878,N_8967);
xor U9129 (N_9129,N_8856,N_8801);
and U9130 (N_9130,N_8928,N_8786);
xor U9131 (N_9131,N_8890,N_8877);
nand U9132 (N_9132,N_8768,N_8968);
nor U9133 (N_9133,N_8904,N_8750);
nand U9134 (N_9134,N_8760,N_8809);
or U9135 (N_9135,N_8916,N_8945);
nand U9136 (N_9136,N_8859,N_8919);
nand U9137 (N_9137,N_8915,N_8888);
and U9138 (N_9138,N_8907,N_8939);
nand U9139 (N_9139,N_8991,N_8887);
nor U9140 (N_9140,N_8879,N_8916);
or U9141 (N_9141,N_8869,N_8934);
xnor U9142 (N_9142,N_8752,N_8756);
nand U9143 (N_9143,N_8898,N_8781);
nor U9144 (N_9144,N_8974,N_8877);
and U9145 (N_9145,N_8768,N_8844);
nor U9146 (N_9146,N_8856,N_8788);
xor U9147 (N_9147,N_8835,N_8892);
nor U9148 (N_9148,N_8972,N_8858);
nor U9149 (N_9149,N_8761,N_8803);
xor U9150 (N_9150,N_8800,N_8794);
nor U9151 (N_9151,N_8883,N_8960);
xnor U9152 (N_9152,N_8931,N_8890);
and U9153 (N_9153,N_8903,N_8933);
and U9154 (N_9154,N_8980,N_8765);
nor U9155 (N_9155,N_8823,N_8788);
or U9156 (N_9156,N_8859,N_8971);
and U9157 (N_9157,N_8910,N_8774);
and U9158 (N_9158,N_8794,N_8762);
nand U9159 (N_9159,N_8868,N_8934);
nand U9160 (N_9160,N_8865,N_8825);
nand U9161 (N_9161,N_8871,N_8837);
nor U9162 (N_9162,N_8920,N_8771);
and U9163 (N_9163,N_8914,N_8889);
xor U9164 (N_9164,N_8891,N_8793);
and U9165 (N_9165,N_8882,N_8832);
and U9166 (N_9166,N_8939,N_8988);
or U9167 (N_9167,N_8863,N_8771);
nand U9168 (N_9168,N_8981,N_8821);
and U9169 (N_9169,N_8884,N_8879);
and U9170 (N_9170,N_8998,N_8872);
and U9171 (N_9171,N_8771,N_8968);
nand U9172 (N_9172,N_8844,N_8775);
and U9173 (N_9173,N_8978,N_8783);
nor U9174 (N_9174,N_8919,N_8868);
nor U9175 (N_9175,N_8842,N_8984);
nor U9176 (N_9176,N_8985,N_8913);
nand U9177 (N_9177,N_8996,N_8925);
nand U9178 (N_9178,N_8850,N_8917);
or U9179 (N_9179,N_8903,N_8981);
xor U9180 (N_9180,N_8848,N_8910);
or U9181 (N_9181,N_8880,N_8828);
nor U9182 (N_9182,N_8831,N_8962);
nor U9183 (N_9183,N_8948,N_8951);
or U9184 (N_9184,N_8812,N_8896);
nand U9185 (N_9185,N_8811,N_8946);
and U9186 (N_9186,N_8964,N_8813);
nand U9187 (N_9187,N_8942,N_8815);
xnor U9188 (N_9188,N_8958,N_8905);
nor U9189 (N_9189,N_8812,N_8822);
nand U9190 (N_9190,N_8983,N_8763);
nor U9191 (N_9191,N_8820,N_8832);
nand U9192 (N_9192,N_8931,N_8864);
and U9193 (N_9193,N_8853,N_8922);
nor U9194 (N_9194,N_8781,N_8803);
nand U9195 (N_9195,N_8776,N_8909);
nand U9196 (N_9196,N_8764,N_8843);
and U9197 (N_9197,N_8836,N_8973);
xor U9198 (N_9198,N_8868,N_8806);
and U9199 (N_9199,N_8886,N_8783);
xor U9200 (N_9200,N_8778,N_8943);
nand U9201 (N_9201,N_8836,N_8832);
or U9202 (N_9202,N_8870,N_8834);
and U9203 (N_9203,N_8790,N_8751);
and U9204 (N_9204,N_8907,N_8834);
nor U9205 (N_9205,N_8983,N_8951);
and U9206 (N_9206,N_8989,N_8929);
nand U9207 (N_9207,N_8808,N_8917);
or U9208 (N_9208,N_8908,N_8860);
and U9209 (N_9209,N_8765,N_8824);
or U9210 (N_9210,N_8854,N_8816);
nor U9211 (N_9211,N_8935,N_8840);
nor U9212 (N_9212,N_8855,N_8819);
and U9213 (N_9213,N_8903,N_8901);
nor U9214 (N_9214,N_8812,N_8838);
and U9215 (N_9215,N_8930,N_8759);
xor U9216 (N_9216,N_8985,N_8929);
xnor U9217 (N_9217,N_8959,N_8914);
nand U9218 (N_9218,N_8992,N_8752);
nand U9219 (N_9219,N_8791,N_8824);
and U9220 (N_9220,N_8842,N_8750);
xnor U9221 (N_9221,N_8840,N_8790);
nor U9222 (N_9222,N_8843,N_8935);
nor U9223 (N_9223,N_8931,N_8915);
xnor U9224 (N_9224,N_8812,N_8839);
nand U9225 (N_9225,N_8818,N_8801);
xnor U9226 (N_9226,N_8902,N_8763);
xor U9227 (N_9227,N_8879,N_8966);
and U9228 (N_9228,N_8975,N_8971);
or U9229 (N_9229,N_8954,N_8826);
and U9230 (N_9230,N_8927,N_8852);
and U9231 (N_9231,N_8963,N_8784);
and U9232 (N_9232,N_8776,N_8948);
xnor U9233 (N_9233,N_8943,N_8873);
or U9234 (N_9234,N_8895,N_8930);
nor U9235 (N_9235,N_8785,N_8897);
or U9236 (N_9236,N_8966,N_8919);
and U9237 (N_9237,N_8786,N_8861);
nor U9238 (N_9238,N_8877,N_8827);
nor U9239 (N_9239,N_8992,N_8847);
or U9240 (N_9240,N_8847,N_8989);
or U9241 (N_9241,N_8908,N_8799);
nand U9242 (N_9242,N_8846,N_8999);
and U9243 (N_9243,N_8844,N_8900);
or U9244 (N_9244,N_8972,N_8867);
xnor U9245 (N_9245,N_8843,N_8797);
and U9246 (N_9246,N_8820,N_8758);
or U9247 (N_9247,N_8887,N_8867);
nand U9248 (N_9248,N_8966,N_8781);
or U9249 (N_9249,N_8843,N_8864);
xor U9250 (N_9250,N_9111,N_9049);
or U9251 (N_9251,N_9102,N_9236);
nand U9252 (N_9252,N_9197,N_9124);
xnor U9253 (N_9253,N_9087,N_9159);
nand U9254 (N_9254,N_9069,N_9225);
or U9255 (N_9255,N_9040,N_9072);
or U9256 (N_9256,N_9136,N_9028);
and U9257 (N_9257,N_9218,N_9242);
xor U9258 (N_9258,N_9209,N_9041);
nor U9259 (N_9259,N_9164,N_9039);
xor U9260 (N_9260,N_9065,N_9141);
or U9261 (N_9261,N_9025,N_9214);
or U9262 (N_9262,N_9162,N_9057);
and U9263 (N_9263,N_9085,N_9077);
nor U9264 (N_9264,N_9175,N_9148);
nor U9265 (N_9265,N_9132,N_9027);
nand U9266 (N_9266,N_9064,N_9152);
xnor U9267 (N_9267,N_9226,N_9245);
nor U9268 (N_9268,N_9232,N_9120);
or U9269 (N_9269,N_9058,N_9217);
or U9270 (N_9270,N_9056,N_9103);
nor U9271 (N_9271,N_9042,N_9061);
or U9272 (N_9272,N_9083,N_9023);
nand U9273 (N_9273,N_9091,N_9168);
nand U9274 (N_9274,N_9150,N_9208);
nor U9275 (N_9275,N_9167,N_9095);
and U9276 (N_9276,N_9114,N_9107);
and U9277 (N_9277,N_9060,N_9047);
xor U9278 (N_9278,N_9076,N_9090);
xor U9279 (N_9279,N_9068,N_9231);
nor U9280 (N_9280,N_9219,N_9220);
or U9281 (N_9281,N_9235,N_9003);
nand U9282 (N_9282,N_9133,N_9238);
nand U9283 (N_9283,N_9081,N_9037);
xor U9284 (N_9284,N_9204,N_9130);
and U9285 (N_9285,N_9066,N_9192);
nor U9286 (N_9286,N_9012,N_9035);
and U9287 (N_9287,N_9029,N_9019);
xnor U9288 (N_9288,N_9045,N_9013);
xnor U9289 (N_9289,N_9198,N_9194);
and U9290 (N_9290,N_9154,N_9105);
nand U9291 (N_9291,N_9059,N_9005);
or U9292 (N_9292,N_9119,N_9067);
and U9293 (N_9293,N_9074,N_9014);
nor U9294 (N_9294,N_9094,N_9241);
or U9295 (N_9295,N_9015,N_9070);
nor U9296 (N_9296,N_9142,N_9149);
nor U9297 (N_9297,N_9145,N_9223);
nor U9298 (N_9298,N_9129,N_9031);
or U9299 (N_9299,N_9186,N_9008);
or U9300 (N_9300,N_9201,N_9088);
and U9301 (N_9301,N_9213,N_9187);
nand U9302 (N_9302,N_9207,N_9093);
nor U9303 (N_9303,N_9155,N_9044);
and U9304 (N_9304,N_9140,N_9082);
nand U9305 (N_9305,N_9123,N_9211);
xnor U9306 (N_9306,N_9215,N_9224);
and U9307 (N_9307,N_9050,N_9156);
nor U9308 (N_9308,N_9180,N_9196);
nand U9309 (N_9309,N_9054,N_9062);
nand U9310 (N_9310,N_9110,N_9170);
and U9311 (N_9311,N_9032,N_9115);
or U9312 (N_9312,N_9210,N_9135);
nand U9313 (N_9313,N_9248,N_9010);
nand U9314 (N_9314,N_9146,N_9227);
and U9315 (N_9315,N_9171,N_9092);
nor U9316 (N_9316,N_9228,N_9221);
and U9317 (N_9317,N_9143,N_9244);
or U9318 (N_9318,N_9021,N_9078);
xnor U9319 (N_9319,N_9202,N_9176);
nor U9320 (N_9320,N_9195,N_9009);
or U9321 (N_9321,N_9063,N_9104);
and U9322 (N_9322,N_9125,N_9178);
or U9323 (N_9323,N_9199,N_9165);
or U9324 (N_9324,N_9126,N_9075);
nand U9325 (N_9325,N_9188,N_9160);
nor U9326 (N_9326,N_9079,N_9158);
and U9327 (N_9327,N_9139,N_9134);
nand U9328 (N_9328,N_9203,N_9038);
or U9329 (N_9329,N_9173,N_9097);
nor U9330 (N_9330,N_9000,N_9022);
nor U9331 (N_9331,N_9099,N_9108);
nor U9332 (N_9332,N_9184,N_9080);
nand U9333 (N_9333,N_9098,N_9055);
or U9334 (N_9334,N_9051,N_9153);
and U9335 (N_9335,N_9166,N_9117);
xnor U9336 (N_9336,N_9084,N_9007);
or U9337 (N_9337,N_9185,N_9239);
xor U9338 (N_9338,N_9234,N_9200);
xor U9339 (N_9339,N_9016,N_9172);
nand U9340 (N_9340,N_9034,N_9237);
nor U9341 (N_9341,N_9205,N_9174);
xnor U9342 (N_9342,N_9177,N_9053);
xor U9343 (N_9343,N_9043,N_9183);
nand U9344 (N_9344,N_9036,N_9179);
nand U9345 (N_9345,N_9131,N_9046);
xnor U9346 (N_9346,N_9033,N_9144);
or U9347 (N_9347,N_9122,N_9018);
nor U9348 (N_9348,N_9233,N_9030);
nor U9349 (N_9349,N_9024,N_9112);
and U9350 (N_9350,N_9128,N_9089);
xor U9351 (N_9351,N_9086,N_9181);
xnor U9352 (N_9352,N_9118,N_9229);
xor U9353 (N_9353,N_9017,N_9246);
nand U9354 (N_9354,N_9071,N_9113);
and U9355 (N_9355,N_9137,N_9230);
nor U9356 (N_9356,N_9240,N_9006);
and U9357 (N_9357,N_9189,N_9002);
xor U9358 (N_9358,N_9020,N_9222);
and U9359 (N_9359,N_9163,N_9109);
nand U9360 (N_9360,N_9106,N_9190);
xor U9361 (N_9361,N_9243,N_9011);
and U9362 (N_9362,N_9052,N_9001);
nor U9363 (N_9363,N_9096,N_9147);
xor U9364 (N_9364,N_9193,N_9191);
nand U9365 (N_9365,N_9157,N_9247);
nor U9366 (N_9366,N_9116,N_9249);
and U9367 (N_9367,N_9169,N_9048);
and U9368 (N_9368,N_9206,N_9212);
or U9369 (N_9369,N_9101,N_9182);
and U9370 (N_9370,N_9073,N_9004);
nor U9371 (N_9371,N_9161,N_9121);
or U9372 (N_9372,N_9216,N_9127);
nor U9373 (N_9373,N_9151,N_9138);
xor U9374 (N_9374,N_9100,N_9026);
xnor U9375 (N_9375,N_9240,N_9158);
xor U9376 (N_9376,N_9087,N_9117);
or U9377 (N_9377,N_9055,N_9151);
and U9378 (N_9378,N_9023,N_9227);
nand U9379 (N_9379,N_9247,N_9215);
or U9380 (N_9380,N_9211,N_9100);
and U9381 (N_9381,N_9130,N_9236);
and U9382 (N_9382,N_9060,N_9082);
nor U9383 (N_9383,N_9043,N_9037);
xor U9384 (N_9384,N_9192,N_9059);
xnor U9385 (N_9385,N_9028,N_9009);
nor U9386 (N_9386,N_9208,N_9046);
xnor U9387 (N_9387,N_9167,N_9054);
and U9388 (N_9388,N_9053,N_9072);
nor U9389 (N_9389,N_9012,N_9054);
nor U9390 (N_9390,N_9050,N_9077);
xor U9391 (N_9391,N_9112,N_9084);
and U9392 (N_9392,N_9129,N_9045);
and U9393 (N_9393,N_9173,N_9142);
xnor U9394 (N_9394,N_9130,N_9002);
nor U9395 (N_9395,N_9227,N_9200);
nor U9396 (N_9396,N_9071,N_9238);
and U9397 (N_9397,N_9117,N_9054);
nor U9398 (N_9398,N_9177,N_9042);
and U9399 (N_9399,N_9197,N_9006);
and U9400 (N_9400,N_9059,N_9118);
nor U9401 (N_9401,N_9199,N_9155);
and U9402 (N_9402,N_9100,N_9081);
xor U9403 (N_9403,N_9160,N_9220);
nor U9404 (N_9404,N_9201,N_9146);
nor U9405 (N_9405,N_9110,N_9171);
nand U9406 (N_9406,N_9137,N_9051);
or U9407 (N_9407,N_9113,N_9179);
nand U9408 (N_9408,N_9115,N_9011);
and U9409 (N_9409,N_9189,N_9147);
xor U9410 (N_9410,N_9082,N_9139);
nor U9411 (N_9411,N_9141,N_9078);
nor U9412 (N_9412,N_9188,N_9029);
or U9413 (N_9413,N_9049,N_9038);
nor U9414 (N_9414,N_9206,N_9079);
and U9415 (N_9415,N_9093,N_9164);
nand U9416 (N_9416,N_9029,N_9245);
nand U9417 (N_9417,N_9040,N_9060);
and U9418 (N_9418,N_9092,N_9214);
nor U9419 (N_9419,N_9185,N_9223);
nor U9420 (N_9420,N_9029,N_9017);
or U9421 (N_9421,N_9056,N_9014);
nand U9422 (N_9422,N_9248,N_9214);
and U9423 (N_9423,N_9116,N_9147);
nor U9424 (N_9424,N_9073,N_9242);
xor U9425 (N_9425,N_9090,N_9192);
xor U9426 (N_9426,N_9099,N_9182);
nor U9427 (N_9427,N_9145,N_9169);
and U9428 (N_9428,N_9236,N_9005);
or U9429 (N_9429,N_9007,N_9079);
or U9430 (N_9430,N_9149,N_9025);
and U9431 (N_9431,N_9212,N_9162);
nand U9432 (N_9432,N_9154,N_9163);
or U9433 (N_9433,N_9074,N_9061);
and U9434 (N_9434,N_9127,N_9129);
nor U9435 (N_9435,N_9077,N_9130);
or U9436 (N_9436,N_9106,N_9069);
nand U9437 (N_9437,N_9172,N_9028);
nor U9438 (N_9438,N_9002,N_9133);
or U9439 (N_9439,N_9161,N_9162);
nor U9440 (N_9440,N_9194,N_9240);
and U9441 (N_9441,N_9199,N_9076);
xnor U9442 (N_9442,N_9216,N_9077);
xnor U9443 (N_9443,N_9182,N_9048);
xnor U9444 (N_9444,N_9011,N_9211);
nor U9445 (N_9445,N_9020,N_9189);
nand U9446 (N_9446,N_9142,N_9172);
nor U9447 (N_9447,N_9202,N_9063);
or U9448 (N_9448,N_9124,N_9143);
or U9449 (N_9449,N_9128,N_9177);
xnor U9450 (N_9450,N_9184,N_9161);
and U9451 (N_9451,N_9078,N_9080);
and U9452 (N_9452,N_9042,N_9015);
or U9453 (N_9453,N_9146,N_9021);
or U9454 (N_9454,N_9031,N_9072);
nand U9455 (N_9455,N_9032,N_9226);
xnor U9456 (N_9456,N_9055,N_9206);
xnor U9457 (N_9457,N_9047,N_9031);
and U9458 (N_9458,N_9183,N_9064);
and U9459 (N_9459,N_9172,N_9181);
and U9460 (N_9460,N_9075,N_9213);
xnor U9461 (N_9461,N_9115,N_9204);
or U9462 (N_9462,N_9210,N_9151);
and U9463 (N_9463,N_9037,N_9063);
nor U9464 (N_9464,N_9144,N_9176);
or U9465 (N_9465,N_9006,N_9142);
and U9466 (N_9466,N_9178,N_9038);
nor U9467 (N_9467,N_9077,N_9007);
nand U9468 (N_9468,N_9237,N_9185);
nor U9469 (N_9469,N_9117,N_9111);
or U9470 (N_9470,N_9098,N_9225);
or U9471 (N_9471,N_9022,N_9144);
or U9472 (N_9472,N_9013,N_9015);
nand U9473 (N_9473,N_9208,N_9115);
nand U9474 (N_9474,N_9157,N_9197);
or U9475 (N_9475,N_9092,N_9210);
nand U9476 (N_9476,N_9077,N_9147);
xor U9477 (N_9477,N_9090,N_9163);
xnor U9478 (N_9478,N_9202,N_9145);
xor U9479 (N_9479,N_9018,N_9038);
xor U9480 (N_9480,N_9163,N_9099);
xnor U9481 (N_9481,N_9121,N_9238);
nor U9482 (N_9482,N_9063,N_9022);
nor U9483 (N_9483,N_9009,N_9207);
xnor U9484 (N_9484,N_9043,N_9130);
xnor U9485 (N_9485,N_9142,N_9037);
xnor U9486 (N_9486,N_9074,N_9215);
nor U9487 (N_9487,N_9088,N_9211);
xor U9488 (N_9488,N_9017,N_9093);
and U9489 (N_9489,N_9098,N_9062);
nor U9490 (N_9490,N_9086,N_9107);
nor U9491 (N_9491,N_9168,N_9003);
nand U9492 (N_9492,N_9003,N_9139);
nand U9493 (N_9493,N_9059,N_9161);
nor U9494 (N_9494,N_9153,N_9162);
or U9495 (N_9495,N_9036,N_9185);
nor U9496 (N_9496,N_9066,N_9003);
nor U9497 (N_9497,N_9136,N_9169);
or U9498 (N_9498,N_9237,N_9055);
nand U9499 (N_9499,N_9089,N_9023);
nand U9500 (N_9500,N_9365,N_9289);
or U9501 (N_9501,N_9368,N_9388);
or U9502 (N_9502,N_9457,N_9349);
and U9503 (N_9503,N_9392,N_9411);
or U9504 (N_9504,N_9301,N_9353);
xnor U9505 (N_9505,N_9437,N_9434);
nor U9506 (N_9506,N_9407,N_9417);
nand U9507 (N_9507,N_9332,N_9258);
xnor U9508 (N_9508,N_9342,N_9408);
xnor U9509 (N_9509,N_9359,N_9478);
nand U9510 (N_9510,N_9309,N_9265);
or U9511 (N_9511,N_9259,N_9445);
nor U9512 (N_9512,N_9470,N_9340);
or U9513 (N_9513,N_9269,N_9410);
xnor U9514 (N_9514,N_9400,N_9383);
xnor U9515 (N_9515,N_9317,N_9472);
xnor U9516 (N_9516,N_9282,N_9352);
xor U9517 (N_9517,N_9311,N_9495);
xor U9518 (N_9518,N_9310,N_9394);
nor U9519 (N_9519,N_9380,N_9372);
xor U9520 (N_9520,N_9492,N_9313);
nand U9521 (N_9521,N_9389,N_9488);
or U9522 (N_9522,N_9412,N_9266);
nor U9523 (N_9523,N_9345,N_9497);
nor U9524 (N_9524,N_9415,N_9436);
and U9525 (N_9525,N_9275,N_9440);
nand U9526 (N_9526,N_9344,N_9491);
or U9527 (N_9527,N_9439,N_9336);
or U9528 (N_9528,N_9480,N_9490);
nand U9529 (N_9529,N_9350,N_9387);
or U9530 (N_9530,N_9493,N_9331);
and U9531 (N_9531,N_9355,N_9418);
or U9532 (N_9532,N_9446,N_9327);
nand U9533 (N_9533,N_9467,N_9348);
or U9534 (N_9534,N_9499,N_9376);
xor U9535 (N_9535,N_9402,N_9278);
nor U9536 (N_9536,N_9398,N_9391);
and U9537 (N_9537,N_9381,N_9333);
xor U9538 (N_9538,N_9338,N_9422);
and U9539 (N_9539,N_9430,N_9290);
and U9540 (N_9540,N_9298,N_9264);
and U9541 (N_9541,N_9471,N_9494);
xor U9542 (N_9542,N_9403,N_9452);
nor U9543 (N_9543,N_9496,N_9384);
and U9544 (N_9544,N_9320,N_9370);
xor U9545 (N_9545,N_9334,N_9465);
nand U9546 (N_9546,N_9432,N_9321);
xnor U9547 (N_9547,N_9339,N_9409);
nor U9548 (N_9548,N_9401,N_9267);
and U9549 (N_9549,N_9468,N_9285);
or U9550 (N_9550,N_9360,N_9295);
nand U9551 (N_9551,N_9405,N_9319);
or U9552 (N_9552,N_9296,N_9425);
nor U9553 (N_9553,N_9428,N_9252);
or U9554 (N_9554,N_9351,N_9438);
and U9555 (N_9555,N_9256,N_9335);
or U9556 (N_9556,N_9377,N_9451);
xnor U9557 (N_9557,N_9283,N_9460);
nor U9558 (N_9558,N_9420,N_9429);
and U9559 (N_9559,N_9291,N_9453);
and U9560 (N_9560,N_9444,N_9483);
xnor U9561 (N_9561,N_9250,N_9287);
xor U9562 (N_9562,N_9281,N_9469);
nand U9563 (N_9563,N_9450,N_9318);
nor U9564 (N_9564,N_9424,N_9274);
nand U9565 (N_9565,N_9343,N_9489);
xnor U9566 (N_9566,N_9463,N_9361);
nor U9567 (N_9567,N_9312,N_9431);
and U9568 (N_9568,N_9433,N_9399);
or U9569 (N_9569,N_9337,N_9328);
or U9570 (N_9570,N_9302,N_9262);
nand U9571 (N_9571,N_9456,N_9395);
nor U9572 (N_9572,N_9435,N_9260);
xor U9573 (N_9573,N_9253,N_9374);
nor U9574 (N_9574,N_9284,N_9406);
nor U9575 (N_9575,N_9263,N_9443);
xnor U9576 (N_9576,N_9357,N_9373);
or U9577 (N_9577,N_9427,N_9277);
nor U9578 (N_9578,N_9475,N_9461);
nand U9579 (N_9579,N_9390,N_9326);
nor U9580 (N_9580,N_9270,N_9276);
and U9581 (N_9581,N_9466,N_9257);
or U9582 (N_9582,N_9356,N_9485);
and U9583 (N_9583,N_9315,N_9288);
xor U9584 (N_9584,N_9305,N_9254);
nand U9585 (N_9585,N_9426,N_9323);
nand U9586 (N_9586,N_9308,N_9304);
nand U9587 (N_9587,N_9423,N_9441);
and U9588 (N_9588,N_9459,N_9366);
xor U9589 (N_9589,N_9413,N_9379);
nor U9590 (N_9590,N_9255,N_9481);
nor U9591 (N_9591,N_9375,N_9307);
nand U9592 (N_9592,N_9482,N_9448);
or U9593 (N_9593,N_9261,N_9325);
xnor U9594 (N_9594,N_9363,N_9280);
nand U9595 (N_9595,N_9386,N_9414);
nor U9596 (N_9596,N_9271,N_9322);
nor U9597 (N_9597,N_9454,N_9397);
or U9598 (N_9598,N_9479,N_9462);
or U9599 (N_9599,N_9484,N_9286);
nor U9600 (N_9600,N_9273,N_9416);
or U9601 (N_9601,N_9268,N_9455);
or U9602 (N_9602,N_9477,N_9300);
or U9603 (N_9603,N_9297,N_9324);
or U9604 (N_9604,N_9303,N_9293);
xor U9605 (N_9605,N_9292,N_9316);
nor U9606 (N_9606,N_9474,N_9447);
nand U9607 (N_9607,N_9371,N_9404);
nor U9608 (N_9608,N_9369,N_9419);
nor U9609 (N_9609,N_9476,N_9367);
xor U9610 (N_9610,N_9378,N_9364);
or U9611 (N_9611,N_9486,N_9498);
xor U9612 (N_9612,N_9294,N_9421);
nand U9613 (N_9613,N_9449,N_9341);
nor U9614 (N_9614,N_9346,N_9382);
xor U9615 (N_9615,N_9299,N_9396);
xor U9616 (N_9616,N_9306,N_9362);
and U9617 (N_9617,N_9354,N_9330);
and U9618 (N_9618,N_9458,N_9279);
or U9619 (N_9619,N_9358,N_9272);
and U9620 (N_9620,N_9442,N_9251);
and U9621 (N_9621,N_9329,N_9473);
nor U9622 (N_9622,N_9385,N_9464);
nand U9623 (N_9623,N_9487,N_9314);
nor U9624 (N_9624,N_9347,N_9393);
nand U9625 (N_9625,N_9270,N_9330);
and U9626 (N_9626,N_9465,N_9355);
or U9627 (N_9627,N_9377,N_9323);
and U9628 (N_9628,N_9411,N_9379);
nor U9629 (N_9629,N_9324,N_9465);
or U9630 (N_9630,N_9317,N_9437);
nor U9631 (N_9631,N_9251,N_9288);
nor U9632 (N_9632,N_9252,N_9282);
or U9633 (N_9633,N_9291,N_9393);
xor U9634 (N_9634,N_9485,N_9295);
and U9635 (N_9635,N_9283,N_9336);
xor U9636 (N_9636,N_9482,N_9486);
and U9637 (N_9637,N_9259,N_9256);
nor U9638 (N_9638,N_9353,N_9363);
and U9639 (N_9639,N_9470,N_9353);
or U9640 (N_9640,N_9341,N_9334);
xor U9641 (N_9641,N_9255,N_9399);
and U9642 (N_9642,N_9417,N_9422);
and U9643 (N_9643,N_9439,N_9310);
nand U9644 (N_9644,N_9344,N_9456);
or U9645 (N_9645,N_9349,N_9404);
nor U9646 (N_9646,N_9325,N_9316);
nand U9647 (N_9647,N_9357,N_9307);
nand U9648 (N_9648,N_9254,N_9465);
or U9649 (N_9649,N_9304,N_9383);
and U9650 (N_9650,N_9480,N_9407);
or U9651 (N_9651,N_9417,N_9476);
and U9652 (N_9652,N_9336,N_9313);
and U9653 (N_9653,N_9296,N_9437);
or U9654 (N_9654,N_9383,N_9470);
or U9655 (N_9655,N_9410,N_9336);
xor U9656 (N_9656,N_9474,N_9316);
and U9657 (N_9657,N_9484,N_9314);
nand U9658 (N_9658,N_9438,N_9254);
and U9659 (N_9659,N_9485,N_9315);
xnor U9660 (N_9660,N_9356,N_9395);
nand U9661 (N_9661,N_9264,N_9480);
and U9662 (N_9662,N_9495,N_9418);
and U9663 (N_9663,N_9359,N_9477);
nor U9664 (N_9664,N_9402,N_9393);
or U9665 (N_9665,N_9279,N_9396);
nand U9666 (N_9666,N_9334,N_9358);
xnor U9667 (N_9667,N_9253,N_9409);
nor U9668 (N_9668,N_9324,N_9287);
or U9669 (N_9669,N_9271,N_9346);
nand U9670 (N_9670,N_9330,N_9289);
xnor U9671 (N_9671,N_9410,N_9464);
nand U9672 (N_9672,N_9393,N_9254);
and U9673 (N_9673,N_9425,N_9310);
and U9674 (N_9674,N_9453,N_9391);
xor U9675 (N_9675,N_9441,N_9395);
or U9676 (N_9676,N_9363,N_9377);
or U9677 (N_9677,N_9423,N_9410);
nor U9678 (N_9678,N_9267,N_9490);
xnor U9679 (N_9679,N_9279,N_9283);
nand U9680 (N_9680,N_9407,N_9484);
and U9681 (N_9681,N_9499,N_9361);
or U9682 (N_9682,N_9400,N_9347);
and U9683 (N_9683,N_9309,N_9268);
nor U9684 (N_9684,N_9357,N_9311);
and U9685 (N_9685,N_9496,N_9465);
nand U9686 (N_9686,N_9286,N_9360);
or U9687 (N_9687,N_9490,N_9448);
and U9688 (N_9688,N_9266,N_9409);
or U9689 (N_9689,N_9391,N_9368);
nor U9690 (N_9690,N_9301,N_9414);
and U9691 (N_9691,N_9275,N_9253);
and U9692 (N_9692,N_9472,N_9498);
nor U9693 (N_9693,N_9295,N_9404);
nor U9694 (N_9694,N_9466,N_9352);
xnor U9695 (N_9695,N_9368,N_9374);
nor U9696 (N_9696,N_9480,N_9259);
and U9697 (N_9697,N_9406,N_9496);
xor U9698 (N_9698,N_9253,N_9490);
and U9699 (N_9699,N_9408,N_9277);
nor U9700 (N_9700,N_9343,N_9437);
xnor U9701 (N_9701,N_9352,N_9488);
nand U9702 (N_9702,N_9356,N_9305);
and U9703 (N_9703,N_9424,N_9278);
nand U9704 (N_9704,N_9271,N_9499);
and U9705 (N_9705,N_9297,N_9329);
or U9706 (N_9706,N_9422,N_9413);
nor U9707 (N_9707,N_9366,N_9282);
and U9708 (N_9708,N_9354,N_9435);
nor U9709 (N_9709,N_9454,N_9442);
and U9710 (N_9710,N_9279,N_9426);
and U9711 (N_9711,N_9497,N_9415);
xor U9712 (N_9712,N_9395,N_9262);
and U9713 (N_9713,N_9485,N_9346);
xor U9714 (N_9714,N_9444,N_9261);
nand U9715 (N_9715,N_9490,N_9287);
or U9716 (N_9716,N_9328,N_9374);
nor U9717 (N_9717,N_9319,N_9348);
nor U9718 (N_9718,N_9279,N_9316);
and U9719 (N_9719,N_9394,N_9289);
nand U9720 (N_9720,N_9495,N_9327);
and U9721 (N_9721,N_9323,N_9347);
or U9722 (N_9722,N_9341,N_9326);
and U9723 (N_9723,N_9328,N_9388);
and U9724 (N_9724,N_9271,N_9292);
or U9725 (N_9725,N_9463,N_9482);
and U9726 (N_9726,N_9310,N_9393);
or U9727 (N_9727,N_9365,N_9384);
xor U9728 (N_9728,N_9312,N_9299);
nor U9729 (N_9729,N_9289,N_9473);
xnor U9730 (N_9730,N_9316,N_9417);
nand U9731 (N_9731,N_9267,N_9375);
and U9732 (N_9732,N_9417,N_9374);
nor U9733 (N_9733,N_9369,N_9487);
nand U9734 (N_9734,N_9323,N_9340);
or U9735 (N_9735,N_9412,N_9482);
nor U9736 (N_9736,N_9325,N_9486);
nand U9737 (N_9737,N_9311,N_9392);
and U9738 (N_9738,N_9441,N_9377);
xor U9739 (N_9739,N_9386,N_9444);
nor U9740 (N_9740,N_9470,N_9256);
and U9741 (N_9741,N_9375,N_9412);
xnor U9742 (N_9742,N_9314,N_9427);
nand U9743 (N_9743,N_9465,N_9331);
xor U9744 (N_9744,N_9379,N_9424);
and U9745 (N_9745,N_9363,N_9452);
nand U9746 (N_9746,N_9338,N_9285);
nor U9747 (N_9747,N_9332,N_9309);
and U9748 (N_9748,N_9481,N_9386);
nor U9749 (N_9749,N_9335,N_9395);
and U9750 (N_9750,N_9742,N_9508);
nor U9751 (N_9751,N_9504,N_9618);
nor U9752 (N_9752,N_9575,N_9516);
nand U9753 (N_9753,N_9652,N_9670);
or U9754 (N_9754,N_9549,N_9706);
xor U9755 (N_9755,N_9714,N_9749);
nand U9756 (N_9756,N_9635,N_9564);
and U9757 (N_9757,N_9623,N_9722);
nor U9758 (N_9758,N_9580,N_9550);
nand U9759 (N_9759,N_9731,N_9691);
nand U9760 (N_9760,N_9638,N_9669);
nor U9761 (N_9761,N_9684,N_9736);
xor U9762 (N_9762,N_9645,N_9701);
nand U9763 (N_9763,N_9689,N_9692);
and U9764 (N_9764,N_9524,N_9636);
or U9765 (N_9765,N_9667,N_9723);
nor U9766 (N_9766,N_9582,N_9605);
or U9767 (N_9767,N_9690,N_9655);
xnor U9768 (N_9768,N_9513,N_9639);
or U9769 (N_9769,N_9525,N_9547);
nand U9770 (N_9770,N_9587,N_9576);
nand U9771 (N_9771,N_9558,N_9571);
and U9772 (N_9772,N_9688,N_9686);
and U9773 (N_9773,N_9588,N_9599);
nand U9774 (N_9774,N_9725,N_9730);
nand U9775 (N_9775,N_9642,N_9679);
xnor U9776 (N_9776,N_9519,N_9544);
nor U9777 (N_9777,N_9685,N_9552);
nand U9778 (N_9778,N_9712,N_9560);
nor U9779 (N_9779,N_9617,N_9649);
and U9780 (N_9780,N_9557,N_9718);
and U9781 (N_9781,N_9534,N_9633);
or U9782 (N_9782,N_9735,N_9680);
nor U9783 (N_9783,N_9563,N_9505);
xnor U9784 (N_9784,N_9514,N_9533);
xor U9785 (N_9785,N_9738,N_9711);
xor U9786 (N_9786,N_9693,N_9596);
nand U9787 (N_9787,N_9521,N_9610);
xnor U9788 (N_9788,N_9646,N_9607);
or U9789 (N_9789,N_9666,N_9594);
or U9790 (N_9790,N_9579,N_9578);
xnor U9791 (N_9791,N_9545,N_9637);
or U9792 (N_9792,N_9624,N_9553);
nor U9793 (N_9793,N_9506,N_9511);
or U9794 (N_9794,N_9627,N_9562);
and U9795 (N_9795,N_9682,N_9530);
xor U9796 (N_9796,N_9540,N_9674);
xor U9797 (N_9797,N_9741,N_9583);
nor U9798 (N_9798,N_9603,N_9656);
nand U9799 (N_9799,N_9737,N_9625);
xnor U9800 (N_9800,N_9678,N_9568);
nand U9801 (N_9801,N_9546,N_9721);
nand U9802 (N_9802,N_9606,N_9609);
xor U9803 (N_9803,N_9709,N_9538);
nor U9804 (N_9804,N_9577,N_9634);
nor U9805 (N_9805,N_9728,N_9619);
and U9806 (N_9806,N_9528,N_9608);
nor U9807 (N_9807,N_9509,N_9726);
and U9808 (N_9808,N_9573,N_9548);
and U9809 (N_9809,N_9611,N_9626);
nor U9810 (N_9810,N_9729,N_9527);
and U9811 (N_9811,N_9515,N_9664);
nor U9812 (N_9812,N_9556,N_9630);
nor U9813 (N_9813,N_9668,N_9628);
nand U9814 (N_9814,N_9715,N_9593);
nor U9815 (N_9815,N_9595,N_9542);
nand U9816 (N_9816,N_9604,N_9614);
nand U9817 (N_9817,N_9671,N_9748);
and U9818 (N_9818,N_9653,N_9720);
nor U9819 (N_9819,N_9650,N_9703);
nor U9820 (N_9820,N_9632,N_9537);
or U9821 (N_9821,N_9589,N_9502);
or U9822 (N_9822,N_9695,N_9702);
or U9823 (N_9823,N_9740,N_9733);
nand U9824 (N_9824,N_9615,N_9503);
nor U9825 (N_9825,N_9622,N_9559);
or U9826 (N_9826,N_9590,N_9676);
or U9827 (N_9827,N_9591,N_9526);
or U9828 (N_9828,N_9654,N_9581);
or U9829 (N_9829,N_9661,N_9518);
nor U9830 (N_9830,N_9522,N_9541);
nand U9831 (N_9831,N_9719,N_9744);
or U9832 (N_9832,N_9613,N_9631);
and U9833 (N_9833,N_9612,N_9710);
and U9834 (N_9834,N_9697,N_9620);
and U9835 (N_9835,N_9551,N_9529);
nor U9836 (N_9836,N_9602,N_9517);
xor U9837 (N_9837,N_9660,N_9707);
xor U9838 (N_9838,N_9536,N_9651);
and U9839 (N_9839,N_9574,N_9700);
or U9840 (N_9840,N_9743,N_9532);
and U9841 (N_9841,N_9747,N_9732);
xor U9842 (N_9842,N_9523,N_9716);
nor U9843 (N_9843,N_9500,N_9644);
or U9844 (N_9844,N_9641,N_9616);
and U9845 (N_9845,N_9507,N_9584);
or U9846 (N_9846,N_9585,N_9600);
xnor U9847 (N_9847,N_9657,N_9565);
nand U9848 (N_9848,N_9598,N_9683);
nand U9849 (N_9849,N_9566,N_9592);
or U9850 (N_9850,N_9567,N_9501);
or U9851 (N_9851,N_9663,N_9705);
and U9852 (N_9852,N_9677,N_9586);
nand U9853 (N_9853,N_9520,N_9543);
nand U9854 (N_9854,N_9724,N_9640);
xor U9855 (N_9855,N_9717,N_9699);
xor U9856 (N_9856,N_9696,N_9681);
or U9857 (N_9857,N_9629,N_9569);
xor U9858 (N_9858,N_9745,N_9648);
or U9859 (N_9859,N_9665,N_9535);
and U9860 (N_9860,N_9647,N_9739);
xnor U9861 (N_9861,N_9597,N_9708);
xnor U9862 (N_9862,N_9561,N_9698);
nor U9863 (N_9863,N_9662,N_9672);
nor U9864 (N_9864,N_9555,N_9531);
and U9865 (N_9865,N_9694,N_9539);
xnor U9866 (N_9866,N_9601,N_9658);
nor U9867 (N_9867,N_9727,N_9659);
nor U9868 (N_9868,N_9673,N_9713);
nor U9869 (N_9869,N_9704,N_9746);
and U9870 (N_9870,N_9570,N_9572);
or U9871 (N_9871,N_9512,N_9675);
xor U9872 (N_9872,N_9621,N_9734);
and U9873 (N_9873,N_9554,N_9510);
and U9874 (N_9874,N_9643,N_9687);
or U9875 (N_9875,N_9556,N_9705);
xnor U9876 (N_9876,N_9682,N_9732);
nor U9877 (N_9877,N_9536,N_9622);
nor U9878 (N_9878,N_9571,N_9503);
xor U9879 (N_9879,N_9596,N_9641);
xnor U9880 (N_9880,N_9561,N_9691);
or U9881 (N_9881,N_9699,N_9582);
nor U9882 (N_9882,N_9517,N_9699);
nand U9883 (N_9883,N_9620,N_9692);
nand U9884 (N_9884,N_9517,N_9656);
nor U9885 (N_9885,N_9607,N_9524);
or U9886 (N_9886,N_9626,N_9690);
or U9887 (N_9887,N_9612,N_9509);
nand U9888 (N_9888,N_9631,N_9649);
nor U9889 (N_9889,N_9614,N_9658);
and U9890 (N_9890,N_9633,N_9661);
or U9891 (N_9891,N_9658,N_9595);
nor U9892 (N_9892,N_9695,N_9599);
nor U9893 (N_9893,N_9623,N_9606);
and U9894 (N_9894,N_9707,N_9732);
nand U9895 (N_9895,N_9610,N_9578);
nor U9896 (N_9896,N_9521,N_9509);
and U9897 (N_9897,N_9624,N_9608);
nand U9898 (N_9898,N_9675,N_9502);
xnor U9899 (N_9899,N_9593,N_9576);
or U9900 (N_9900,N_9595,N_9581);
and U9901 (N_9901,N_9534,N_9543);
and U9902 (N_9902,N_9678,N_9712);
xor U9903 (N_9903,N_9513,N_9502);
nor U9904 (N_9904,N_9612,N_9630);
nand U9905 (N_9905,N_9513,N_9525);
nand U9906 (N_9906,N_9624,N_9611);
and U9907 (N_9907,N_9551,N_9723);
or U9908 (N_9908,N_9610,N_9524);
nor U9909 (N_9909,N_9627,N_9563);
xor U9910 (N_9910,N_9666,N_9658);
or U9911 (N_9911,N_9561,N_9643);
or U9912 (N_9912,N_9618,N_9518);
and U9913 (N_9913,N_9667,N_9528);
and U9914 (N_9914,N_9729,N_9735);
and U9915 (N_9915,N_9740,N_9543);
and U9916 (N_9916,N_9508,N_9626);
or U9917 (N_9917,N_9674,N_9655);
nand U9918 (N_9918,N_9586,N_9705);
or U9919 (N_9919,N_9716,N_9643);
and U9920 (N_9920,N_9638,N_9708);
and U9921 (N_9921,N_9566,N_9651);
nor U9922 (N_9922,N_9503,N_9576);
nand U9923 (N_9923,N_9654,N_9690);
and U9924 (N_9924,N_9599,N_9681);
xor U9925 (N_9925,N_9584,N_9561);
xnor U9926 (N_9926,N_9647,N_9615);
and U9927 (N_9927,N_9742,N_9601);
and U9928 (N_9928,N_9534,N_9523);
nor U9929 (N_9929,N_9515,N_9666);
xor U9930 (N_9930,N_9537,N_9739);
or U9931 (N_9931,N_9635,N_9738);
or U9932 (N_9932,N_9695,N_9650);
nor U9933 (N_9933,N_9550,N_9671);
nand U9934 (N_9934,N_9533,N_9646);
nand U9935 (N_9935,N_9738,N_9709);
or U9936 (N_9936,N_9540,N_9561);
xnor U9937 (N_9937,N_9675,N_9639);
xor U9938 (N_9938,N_9698,N_9730);
xnor U9939 (N_9939,N_9529,N_9723);
or U9940 (N_9940,N_9700,N_9646);
nor U9941 (N_9941,N_9548,N_9678);
nor U9942 (N_9942,N_9657,N_9624);
xor U9943 (N_9943,N_9606,N_9521);
nand U9944 (N_9944,N_9686,N_9656);
nor U9945 (N_9945,N_9711,N_9609);
or U9946 (N_9946,N_9590,N_9730);
or U9947 (N_9947,N_9531,N_9677);
or U9948 (N_9948,N_9621,N_9535);
nor U9949 (N_9949,N_9705,N_9537);
xor U9950 (N_9950,N_9719,N_9546);
nor U9951 (N_9951,N_9551,N_9675);
nand U9952 (N_9952,N_9534,N_9505);
nand U9953 (N_9953,N_9565,N_9525);
xor U9954 (N_9954,N_9570,N_9625);
or U9955 (N_9955,N_9518,N_9558);
xor U9956 (N_9956,N_9535,N_9722);
and U9957 (N_9957,N_9534,N_9710);
xor U9958 (N_9958,N_9557,N_9695);
or U9959 (N_9959,N_9639,N_9504);
xnor U9960 (N_9960,N_9639,N_9645);
or U9961 (N_9961,N_9603,N_9678);
xor U9962 (N_9962,N_9519,N_9627);
or U9963 (N_9963,N_9554,N_9711);
and U9964 (N_9964,N_9674,N_9673);
and U9965 (N_9965,N_9636,N_9549);
xnor U9966 (N_9966,N_9719,N_9688);
and U9967 (N_9967,N_9536,N_9738);
nand U9968 (N_9968,N_9575,N_9515);
nand U9969 (N_9969,N_9631,N_9591);
xnor U9970 (N_9970,N_9510,N_9670);
and U9971 (N_9971,N_9652,N_9573);
or U9972 (N_9972,N_9746,N_9707);
or U9973 (N_9973,N_9711,N_9589);
xor U9974 (N_9974,N_9717,N_9582);
or U9975 (N_9975,N_9533,N_9735);
nor U9976 (N_9976,N_9607,N_9582);
or U9977 (N_9977,N_9657,N_9632);
and U9978 (N_9978,N_9503,N_9556);
nand U9979 (N_9979,N_9615,N_9749);
and U9980 (N_9980,N_9739,N_9641);
xor U9981 (N_9981,N_9657,N_9630);
nand U9982 (N_9982,N_9524,N_9594);
nor U9983 (N_9983,N_9676,N_9546);
and U9984 (N_9984,N_9739,N_9688);
and U9985 (N_9985,N_9699,N_9516);
nor U9986 (N_9986,N_9597,N_9713);
nand U9987 (N_9987,N_9670,N_9553);
or U9988 (N_9988,N_9632,N_9647);
or U9989 (N_9989,N_9556,N_9598);
nor U9990 (N_9990,N_9658,N_9688);
or U9991 (N_9991,N_9727,N_9589);
nand U9992 (N_9992,N_9701,N_9665);
or U9993 (N_9993,N_9712,N_9619);
xor U9994 (N_9994,N_9595,N_9520);
xnor U9995 (N_9995,N_9577,N_9537);
nor U9996 (N_9996,N_9698,N_9555);
nand U9997 (N_9997,N_9594,N_9598);
nand U9998 (N_9998,N_9593,N_9511);
nand U9999 (N_9999,N_9594,N_9711);
xnor U10000 (N_10000,N_9848,N_9821);
or U10001 (N_10001,N_9789,N_9876);
and U10002 (N_10002,N_9830,N_9839);
nor U10003 (N_10003,N_9838,N_9938);
xnor U10004 (N_10004,N_9902,N_9953);
nand U10005 (N_10005,N_9842,N_9808);
nor U10006 (N_10006,N_9886,N_9810);
and U10007 (N_10007,N_9885,N_9792);
xor U10008 (N_10008,N_9807,N_9879);
nand U10009 (N_10009,N_9921,N_9864);
xnor U10010 (N_10010,N_9857,N_9954);
nor U10011 (N_10011,N_9892,N_9868);
nor U10012 (N_10012,N_9813,N_9793);
nor U10013 (N_10013,N_9777,N_9899);
xor U10014 (N_10014,N_9873,N_9918);
xnor U10015 (N_10015,N_9984,N_9795);
nand U10016 (N_10016,N_9968,N_9887);
or U10017 (N_10017,N_9890,N_9761);
nor U10018 (N_10018,N_9975,N_9904);
xor U10019 (N_10019,N_9782,N_9889);
nor U10020 (N_10020,N_9797,N_9962);
or U10021 (N_10021,N_9756,N_9880);
nor U10022 (N_10022,N_9751,N_9776);
or U10023 (N_10023,N_9866,N_9907);
or U10024 (N_10024,N_9897,N_9783);
nor U10025 (N_10025,N_9974,N_9773);
xnor U10026 (N_10026,N_9828,N_9949);
xnor U10027 (N_10027,N_9874,N_9977);
and U10028 (N_10028,N_9972,N_9896);
xor U10029 (N_10029,N_9869,N_9829);
nor U10030 (N_10030,N_9772,N_9779);
or U10031 (N_10031,N_9985,N_9774);
or U10032 (N_10032,N_9955,N_9911);
or U10033 (N_10033,N_9875,N_9894);
and U10034 (N_10034,N_9930,N_9946);
nor U10035 (N_10035,N_9958,N_9931);
nand U10036 (N_10036,N_9846,N_9941);
nand U10037 (N_10037,N_9816,N_9901);
and U10038 (N_10038,N_9820,N_9778);
nand U10039 (N_10039,N_9910,N_9883);
and U10040 (N_10040,N_9754,N_9979);
and U10041 (N_10041,N_9995,N_9815);
xor U10042 (N_10042,N_9814,N_9763);
or U10043 (N_10043,N_9944,N_9784);
or U10044 (N_10044,N_9960,N_9967);
xor U10045 (N_10045,N_9878,N_9964);
or U10046 (N_10046,N_9847,N_9852);
and U10047 (N_10047,N_9799,N_9798);
nor U10048 (N_10048,N_9835,N_9933);
nand U10049 (N_10049,N_9929,N_9981);
nor U10050 (N_10050,N_9822,N_9994);
nor U10051 (N_10051,N_9936,N_9914);
or U10052 (N_10052,N_9973,N_9831);
or U10053 (N_10053,N_9865,N_9861);
nor U10054 (N_10054,N_9856,N_9819);
and U10055 (N_10055,N_9983,N_9841);
or U10056 (N_10056,N_9766,N_9812);
xor U10057 (N_10057,N_9990,N_9917);
nor U10058 (N_10058,N_9752,N_9757);
xnor U10059 (N_10059,N_9895,N_9951);
xnor U10060 (N_10060,N_9826,N_9759);
xnor U10061 (N_10061,N_9755,N_9945);
and U10062 (N_10062,N_9859,N_9963);
nor U10063 (N_10063,N_9912,N_9855);
or U10064 (N_10064,N_9753,N_9800);
or U10065 (N_10065,N_9928,N_9872);
xnor U10066 (N_10066,N_9992,N_9934);
nand U10067 (N_10067,N_9854,N_9942);
nor U10068 (N_10068,N_9849,N_9827);
nor U10069 (N_10069,N_9957,N_9832);
xnor U10070 (N_10070,N_9833,N_9760);
and U10071 (N_10071,N_9862,N_9845);
nand U10072 (N_10072,N_9860,N_9959);
nand U10073 (N_10073,N_9966,N_9871);
xnor U10074 (N_10074,N_9775,N_9771);
xnor U10075 (N_10075,N_9870,N_9769);
xor U10076 (N_10076,N_9982,N_9785);
nand U10077 (N_10077,N_9758,N_9969);
or U10078 (N_10078,N_9988,N_9908);
and U10079 (N_10079,N_9956,N_9939);
xnor U10080 (N_10080,N_9888,N_9922);
xnor U10081 (N_10081,N_9987,N_9881);
nor U10082 (N_10082,N_9996,N_9867);
nor U10083 (N_10083,N_9844,N_9905);
nor U10084 (N_10084,N_9780,N_9937);
or U10085 (N_10085,N_9986,N_9843);
xor U10086 (N_10086,N_9786,N_9980);
nand U10087 (N_10087,N_9825,N_9919);
xnor U10088 (N_10088,N_9916,N_9767);
nand U10089 (N_10089,N_9851,N_9884);
nand U10090 (N_10090,N_9809,N_9850);
nor U10091 (N_10091,N_9787,N_9823);
and U10092 (N_10092,N_9909,N_9925);
or U10093 (N_10093,N_9882,N_9991);
nand U10094 (N_10094,N_9923,N_9840);
or U10095 (N_10095,N_9947,N_9811);
nand U10096 (N_10096,N_9858,N_9790);
xor U10097 (N_10097,N_9804,N_9961);
xnor U10098 (N_10098,N_9915,N_9998);
and U10099 (N_10099,N_9927,N_9971);
xnor U10100 (N_10100,N_9762,N_9970);
and U10101 (N_10101,N_9781,N_9853);
or U10102 (N_10102,N_9818,N_9900);
or U10103 (N_10103,N_9997,N_9836);
xnor U10104 (N_10104,N_9950,N_9794);
nor U10105 (N_10105,N_9805,N_9999);
and U10106 (N_10106,N_9898,N_9926);
nand U10107 (N_10107,N_9796,N_9943);
nor U10108 (N_10108,N_9834,N_9877);
and U10109 (N_10109,N_9791,N_9802);
and U10110 (N_10110,N_9770,N_9765);
xor U10111 (N_10111,N_9932,N_9906);
and U10112 (N_10112,N_9863,N_9837);
xor U10113 (N_10113,N_9989,N_9993);
nand U10114 (N_10114,N_9893,N_9788);
nor U10115 (N_10115,N_9978,N_9965);
nor U10116 (N_10116,N_9891,N_9920);
and U10117 (N_10117,N_9948,N_9924);
xnor U10118 (N_10118,N_9913,N_9764);
or U10119 (N_10119,N_9903,N_9801);
and U10120 (N_10120,N_9768,N_9976);
or U10121 (N_10121,N_9952,N_9940);
xnor U10122 (N_10122,N_9803,N_9750);
or U10123 (N_10123,N_9935,N_9824);
nor U10124 (N_10124,N_9806,N_9817);
and U10125 (N_10125,N_9760,N_9834);
xnor U10126 (N_10126,N_9999,N_9971);
nor U10127 (N_10127,N_9885,N_9752);
nand U10128 (N_10128,N_9982,N_9926);
nand U10129 (N_10129,N_9872,N_9873);
nand U10130 (N_10130,N_9774,N_9900);
nand U10131 (N_10131,N_9908,N_9998);
or U10132 (N_10132,N_9857,N_9831);
and U10133 (N_10133,N_9843,N_9996);
or U10134 (N_10134,N_9787,N_9791);
nand U10135 (N_10135,N_9977,N_9986);
xor U10136 (N_10136,N_9822,N_9999);
or U10137 (N_10137,N_9978,N_9891);
and U10138 (N_10138,N_9896,N_9792);
or U10139 (N_10139,N_9770,N_9777);
xnor U10140 (N_10140,N_9921,N_9915);
nor U10141 (N_10141,N_9866,N_9931);
nand U10142 (N_10142,N_9826,N_9812);
nand U10143 (N_10143,N_9850,N_9896);
nand U10144 (N_10144,N_9816,N_9953);
xnor U10145 (N_10145,N_9972,N_9992);
and U10146 (N_10146,N_9993,N_9988);
nand U10147 (N_10147,N_9843,N_9756);
and U10148 (N_10148,N_9809,N_9776);
xnor U10149 (N_10149,N_9765,N_9773);
nand U10150 (N_10150,N_9979,N_9936);
or U10151 (N_10151,N_9774,N_9990);
nor U10152 (N_10152,N_9794,N_9877);
xnor U10153 (N_10153,N_9753,N_9932);
nand U10154 (N_10154,N_9793,N_9834);
nor U10155 (N_10155,N_9869,N_9785);
nand U10156 (N_10156,N_9827,N_9807);
and U10157 (N_10157,N_9771,N_9861);
xor U10158 (N_10158,N_9906,N_9953);
nand U10159 (N_10159,N_9758,N_9871);
nand U10160 (N_10160,N_9827,N_9776);
and U10161 (N_10161,N_9813,N_9951);
nor U10162 (N_10162,N_9935,N_9806);
or U10163 (N_10163,N_9782,N_9771);
and U10164 (N_10164,N_9988,N_9832);
nor U10165 (N_10165,N_9799,N_9758);
nor U10166 (N_10166,N_9842,N_9943);
and U10167 (N_10167,N_9798,N_9807);
or U10168 (N_10168,N_9886,N_9894);
and U10169 (N_10169,N_9989,N_9753);
and U10170 (N_10170,N_9786,N_9837);
nand U10171 (N_10171,N_9996,N_9764);
nand U10172 (N_10172,N_9887,N_9839);
or U10173 (N_10173,N_9871,N_9769);
and U10174 (N_10174,N_9775,N_9806);
nor U10175 (N_10175,N_9989,N_9778);
and U10176 (N_10176,N_9790,N_9957);
xor U10177 (N_10177,N_9852,N_9750);
xor U10178 (N_10178,N_9978,N_9924);
xnor U10179 (N_10179,N_9985,N_9858);
nor U10180 (N_10180,N_9976,N_9808);
or U10181 (N_10181,N_9821,N_9774);
nor U10182 (N_10182,N_9779,N_9879);
or U10183 (N_10183,N_9814,N_9957);
or U10184 (N_10184,N_9790,N_9876);
and U10185 (N_10185,N_9859,N_9884);
xnor U10186 (N_10186,N_9987,N_9764);
xnor U10187 (N_10187,N_9972,N_9983);
xor U10188 (N_10188,N_9999,N_9769);
nand U10189 (N_10189,N_9750,N_9926);
nor U10190 (N_10190,N_9856,N_9807);
and U10191 (N_10191,N_9855,N_9950);
xor U10192 (N_10192,N_9781,N_9983);
nor U10193 (N_10193,N_9943,N_9878);
or U10194 (N_10194,N_9955,N_9917);
nand U10195 (N_10195,N_9874,N_9787);
nand U10196 (N_10196,N_9871,N_9787);
xor U10197 (N_10197,N_9754,N_9915);
or U10198 (N_10198,N_9793,N_9854);
and U10199 (N_10199,N_9761,N_9998);
nor U10200 (N_10200,N_9991,N_9863);
xnor U10201 (N_10201,N_9882,N_9927);
xnor U10202 (N_10202,N_9840,N_9812);
nor U10203 (N_10203,N_9959,N_9945);
or U10204 (N_10204,N_9873,N_9840);
or U10205 (N_10205,N_9806,N_9814);
nor U10206 (N_10206,N_9976,N_9940);
or U10207 (N_10207,N_9950,N_9978);
nand U10208 (N_10208,N_9918,N_9799);
nor U10209 (N_10209,N_9823,N_9758);
nand U10210 (N_10210,N_9869,N_9972);
or U10211 (N_10211,N_9833,N_9870);
or U10212 (N_10212,N_9849,N_9886);
nand U10213 (N_10213,N_9991,N_9999);
nor U10214 (N_10214,N_9961,N_9844);
or U10215 (N_10215,N_9896,N_9836);
nand U10216 (N_10216,N_9825,N_9868);
and U10217 (N_10217,N_9857,N_9882);
xnor U10218 (N_10218,N_9819,N_9976);
nor U10219 (N_10219,N_9962,N_9801);
and U10220 (N_10220,N_9897,N_9768);
xnor U10221 (N_10221,N_9938,N_9887);
and U10222 (N_10222,N_9955,N_9836);
and U10223 (N_10223,N_9951,N_9836);
nor U10224 (N_10224,N_9978,N_9776);
and U10225 (N_10225,N_9929,N_9913);
nor U10226 (N_10226,N_9883,N_9845);
xnor U10227 (N_10227,N_9876,N_9829);
and U10228 (N_10228,N_9885,N_9765);
nand U10229 (N_10229,N_9822,N_9966);
xor U10230 (N_10230,N_9990,N_9925);
nand U10231 (N_10231,N_9945,N_9876);
or U10232 (N_10232,N_9754,N_9882);
and U10233 (N_10233,N_9997,N_9757);
and U10234 (N_10234,N_9941,N_9781);
and U10235 (N_10235,N_9964,N_9761);
nor U10236 (N_10236,N_9850,N_9994);
nor U10237 (N_10237,N_9882,N_9764);
xnor U10238 (N_10238,N_9787,N_9872);
xor U10239 (N_10239,N_9784,N_9978);
and U10240 (N_10240,N_9809,N_9800);
nor U10241 (N_10241,N_9892,N_9780);
and U10242 (N_10242,N_9961,N_9771);
and U10243 (N_10243,N_9782,N_9891);
or U10244 (N_10244,N_9969,N_9982);
nand U10245 (N_10245,N_9854,N_9945);
nand U10246 (N_10246,N_9856,N_9964);
nand U10247 (N_10247,N_9817,N_9819);
nand U10248 (N_10248,N_9990,N_9936);
and U10249 (N_10249,N_9824,N_9782);
nor U10250 (N_10250,N_10012,N_10150);
or U10251 (N_10251,N_10225,N_10154);
xor U10252 (N_10252,N_10042,N_10103);
nor U10253 (N_10253,N_10246,N_10096);
or U10254 (N_10254,N_10056,N_10186);
xor U10255 (N_10255,N_10060,N_10112);
or U10256 (N_10256,N_10067,N_10038);
nand U10257 (N_10257,N_10242,N_10137);
nor U10258 (N_10258,N_10200,N_10066);
nor U10259 (N_10259,N_10172,N_10220);
nand U10260 (N_10260,N_10245,N_10239);
nand U10261 (N_10261,N_10053,N_10197);
and U10262 (N_10262,N_10212,N_10247);
xnor U10263 (N_10263,N_10173,N_10130);
xor U10264 (N_10264,N_10010,N_10182);
nand U10265 (N_10265,N_10037,N_10055);
xnor U10266 (N_10266,N_10223,N_10085);
nand U10267 (N_10267,N_10205,N_10122);
xnor U10268 (N_10268,N_10104,N_10021);
and U10269 (N_10269,N_10132,N_10213);
or U10270 (N_10270,N_10115,N_10093);
xor U10271 (N_10271,N_10126,N_10176);
or U10272 (N_10272,N_10167,N_10027);
or U10273 (N_10273,N_10035,N_10206);
xor U10274 (N_10274,N_10168,N_10183);
and U10275 (N_10275,N_10041,N_10028);
xor U10276 (N_10276,N_10057,N_10036);
xnor U10277 (N_10277,N_10171,N_10054);
or U10278 (N_10278,N_10236,N_10159);
or U10279 (N_10279,N_10240,N_10233);
and U10280 (N_10280,N_10047,N_10118);
nor U10281 (N_10281,N_10086,N_10189);
xnor U10282 (N_10282,N_10204,N_10123);
and U10283 (N_10283,N_10083,N_10025);
nand U10284 (N_10284,N_10065,N_10022);
nor U10285 (N_10285,N_10068,N_10217);
xor U10286 (N_10286,N_10165,N_10148);
or U10287 (N_10287,N_10109,N_10019);
xnor U10288 (N_10288,N_10194,N_10144);
xor U10289 (N_10289,N_10113,N_10032);
nand U10290 (N_10290,N_10237,N_10023);
xnor U10291 (N_10291,N_10040,N_10076);
xnor U10292 (N_10292,N_10029,N_10070);
xor U10293 (N_10293,N_10039,N_10151);
xor U10294 (N_10294,N_10181,N_10218);
nand U10295 (N_10295,N_10108,N_10134);
nor U10296 (N_10296,N_10013,N_10044);
nor U10297 (N_10297,N_10102,N_10015);
and U10298 (N_10298,N_10088,N_10228);
xnor U10299 (N_10299,N_10156,N_10138);
nor U10300 (N_10300,N_10203,N_10091);
xor U10301 (N_10301,N_10090,N_10110);
or U10302 (N_10302,N_10024,N_10146);
and U10303 (N_10303,N_10097,N_10064);
or U10304 (N_10304,N_10195,N_10111);
nand U10305 (N_10305,N_10034,N_10219);
xnor U10306 (N_10306,N_10187,N_10198);
or U10307 (N_10307,N_10177,N_10241);
or U10308 (N_10308,N_10133,N_10106);
and U10309 (N_10309,N_10081,N_10094);
nand U10310 (N_10310,N_10002,N_10179);
nor U10311 (N_10311,N_10058,N_10100);
nand U10312 (N_10312,N_10141,N_10117);
nor U10313 (N_10313,N_10149,N_10201);
and U10314 (N_10314,N_10059,N_10188);
xnor U10315 (N_10315,N_10005,N_10196);
or U10316 (N_10316,N_10008,N_10107);
and U10317 (N_10317,N_10001,N_10229);
nand U10318 (N_10318,N_10071,N_10114);
xor U10319 (N_10319,N_10006,N_10208);
xor U10320 (N_10320,N_10244,N_10062);
nor U10321 (N_10321,N_10216,N_10017);
and U10322 (N_10322,N_10243,N_10128);
nor U10323 (N_10323,N_10184,N_10248);
and U10324 (N_10324,N_10215,N_10072);
nand U10325 (N_10325,N_10222,N_10080);
xnor U10326 (N_10326,N_10221,N_10193);
xor U10327 (N_10327,N_10119,N_10190);
xor U10328 (N_10328,N_10069,N_10046);
nor U10329 (N_10329,N_10031,N_10143);
xor U10330 (N_10330,N_10147,N_10045);
nand U10331 (N_10331,N_10166,N_10026);
nor U10332 (N_10332,N_10178,N_10077);
or U10333 (N_10333,N_10227,N_10009);
nand U10334 (N_10334,N_10000,N_10089);
nor U10335 (N_10335,N_10140,N_10139);
nor U10336 (N_10336,N_10180,N_10136);
and U10337 (N_10337,N_10235,N_10135);
nor U10338 (N_10338,N_10210,N_10098);
nor U10339 (N_10339,N_10157,N_10105);
and U10340 (N_10340,N_10158,N_10142);
xor U10341 (N_10341,N_10016,N_10230);
nor U10342 (N_10342,N_10011,N_10169);
nor U10343 (N_10343,N_10020,N_10249);
and U10344 (N_10344,N_10101,N_10185);
xor U10345 (N_10345,N_10164,N_10078);
nor U10346 (N_10346,N_10153,N_10211);
nand U10347 (N_10347,N_10129,N_10174);
xnor U10348 (N_10348,N_10127,N_10199);
and U10349 (N_10349,N_10063,N_10074);
nor U10350 (N_10350,N_10124,N_10202);
or U10351 (N_10351,N_10207,N_10175);
or U10352 (N_10352,N_10214,N_10099);
nor U10353 (N_10353,N_10162,N_10030);
and U10354 (N_10354,N_10051,N_10234);
nor U10355 (N_10355,N_10018,N_10007);
or U10356 (N_10356,N_10163,N_10238);
and U10357 (N_10357,N_10121,N_10120);
nand U10358 (N_10358,N_10152,N_10073);
nand U10359 (N_10359,N_10050,N_10231);
and U10360 (N_10360,N_10079,N_10191);
nand U10361 (N_10361,N_10095,N_10004);
xnor U10362 (N_10362,N_10043,N_10049);
and U10363 (N_10363,N_10092,N_10160);
nor U10364 (N_10364,N_10087,N_10125);
and U10365 (N_10365,N_10192,N_10014);
nor U10366 (N_10366,N_10161,N_10003);
xnor U10367 (N_10367,N_10052,N_10033);
xnor U10368 (N_10368,N_10145,N_10075);
nor U10369 (N_10369,N_10170,N_10155);
and U10370 (N_10370,N_10131,N_10082);
nor U10371 (N_10371,N_10224,N_10061);
or U10372 (N_10372,N_10226,N_10232);
xor U10373 (N_10373,N_10048,N_10209);
nand U10374 (N_10374,N_10084,N_10116);
nand U10375 (N_10375,N_10245,N_10224);
and U10376 (N_10376,N_10128,N_10203);
and U10377 (N_10377,N_10229,N_10246);
nor U10378 (N_10378,N_10021,N_10144);
or U10379 (N_10379,N_10169,N_10119);
xor U10380 (N_10380,N_10225,N_10105);
or U10381 (N_10381,N_10238,N_10157);
nand U10382 (N_10382,N_10026,N_10211);
xnor U10383 (N_10383,N_10242,N_10192);
nor U10384 (N_10384,N_10079,N_10233);
xnor U10385 (N_10385,N_10154,N_10157);
xnor U10386 (N_10386,N_10033,N_10053);
nand U10387 (N_10387,N_10077,N_10055);
xor U10388 (N_10388,N_10049,N_10064);
nand U10389 (N_10389,N_10020,N_10076);
nand U10390 (N_10390,N_10149,N_10166);
nand U10391 (N_10391,N_10234,N_10244);
nand U10392 (N_10392,N_10153,N_10205);
or U10393 (N_10393,N_10029,N_10112);
nand U10394 (N_10394,N_10241,N_10060);
or U10395 (N_10395,N_10207,N_10191);
or U10396 (N_10396,N_10130,N_10216);
and U10397 (N_10397,N_10130,N_10058);
nand U10398 (N_10398,N_10217,N_10136);
and U10399 (N_10399,N_10145,N_10197);
nor U10400 (N_10400,N_10170,N_10246);
xnor U10401 (N_10401,N_10159,N_10244);
xnor U10402 (N_10402,N_10193,N_10231);
xnor U10403 (N_10403,N_10219,N_10109);
nor U10404 (N_10404,N_10221,N_10220);
or U10405 (N_10405,N_10156,N_10031);
nand U10406 (N_10406,N_10213,N_10161);
xor U10407 (N_10407,N_10210,N_10010);
xor U10408 (N_10408,N_10242,N_10143);
and U10409 (N_10409,N_10212,N_10115);
or U10410 (N_10410,N_10201,N_10221);
or U10411 (N_10411,N_10005,N_10106);
nor U10412 (N_10412,N_10019,N_10063);
or U10413 (N_10413,N_10037,N_10031);
and U10414 (N_10414,N_10071,N_10099);
and U10415 (N_10415,N_10068,N_10159);
xnor U10416 (N_10416,N_10120,N_10227);
and U10417 (N_10417,N_10180,N_10091);
nand U10418 (N_10418,N_10046,N_10075);
nand U10419 (N_10419,N_10090,N_10123);
xor U10420 (N_10420,N_10069,N_10095);
xnor U10421 (N_10421,N_10013,N_10203);
nor U10422 (N_10422,N_10070,N_10074);
nor U10423 (N_10423,N_10020,N_10108);
and U10424 (N_10424,N_10034,N_10000);
and U10425 (N_10425,N_10049,N_10038);
or U10426 (N_10426,N_10237,N_10135);
or U10427 (N_10427,N_10190,N_10062);
and U10428 (N_10428,N_10029,N_10172);
or U10429 (N_10429,N_10218,N_10114);
or U10430 (N_10430,N_10190,N_10132);
xnor U10431 (N_10431,N_10111,N_10168);
and U10432 (N_10432,N_10024,N_10071);
or U10433 (N_10433,N_10115,N_10081);
and U10434 (N_10434,N_10236,N_10104);
and U10435 (N_10435,N_10010,N_10109);
and U10436 (N_10436,N_10242,N_10122);
and U10437 (N_10437,N_10054,N_10066);
and U10438 (N_10438,N_10003,N_10042);
nand U10439 (N_10439,N_10004,N_10080);
xor U10440 (N_10440,N_10196,N_10193);
nor U10441 (N_10441,N_10214,N_10085);
xnor U10442 (N_10442,N_10153,N_10021);
and U10443 (N_10443,N_10092,N_10064);
nor U10444 (N_10444,N_10131,N_10053);
nor U10445 (N_10445,N_10130,N_10069);
nor U10446 (N_10446,N_10175,N_10050);
nand U10447 (N_10447,N_10193,N_10019);
and U10448 (N_10448,N_10211,N_10139);
and U10449 (N_10449,N_10226,N_10210);
or U10450 (N_10450,N_10242,N_10207);
nor U10451 (N_10451,N_10151,N_10186);
nor U10452 (N_10452,N_10037,N_10230);
or U10453 (N_10453,N_10057,N_10000);
or U10454 (N_10454,N_10233,N_10241);
xor U10455 (N_10455,N_10067,N_10232);
xor U10456 (N_10456,N_10082,N_10164);
nor U10457 (N_10457,N_10182,N_10174);
xnor U10458 (N_10458,N_10184,N_10243);
nor U10459 (N_10459,N_10079,N_10219);
xor U10460 (N_10460,N_10179,N_10248);
nor U10461 (N_10461,N_10246,N_10167);
or U10462 (N_10462,N_10051,N_10237);
or U10463 (N_10463,N_10201,N_10156);
nand U10464 (N_10464,N_10031,N_10104);
and U10465 (N_10465,N_10134,N_10034);
nand U10466 (N_10466,N_10054,N_10151);
xor U10467 (N_10467,N_10195,N_10050);
and U10468 (N_10468,N_10239,N_10043);
nor U10469 (N_10469,N_10067,N_10015);
xnor U10470 (N_10470,N_10245,N_10151);
and U10471 (N_10471,N_10102,N_10111);
and U10472 (N_10472,N_10008,N_10064);
and U10473 (N_10473,N_10098,N_10088);
or U10474 (N_10474,N_10228,N_10022);
or U10475 (N_10475,N_10012,N_10199);
nand U10476 (N_10476,N_10023,N_10170);
nand U10477 (N_10477,N_10094,N_10020);
xnor U10478 (N_10478,N_10236,N_10188);
nand U10479 (N_10479,N_10070,N_10208);
or U10480 (N_10480,N_10014,N_10027);
nor U10481 (N_10481,N_10202,N_10117);
xnor U10482 (N_10482,N_10028,N_10221);
and U10483 (N_10483,N_10193,N_10172);
or U10484 (N_10484,N_10178,N_10115);
nand U10485 (N_10485,N_10060,N_10098);
nor U10486 (N_10486,N_10183,N_10238);
nand U10487 (N_10487,N_10174,N_10134);
nor U10488 (N_10488,N_10091,N_10116);
nand U10489 (N_10489,N_10226,N_10042);
xnor U10490 (N_10490,N_10080,N_10063);
nand U10491 (N_10491,N_10013,N_10064);
nor U10492 (N_10492,N_10209,N_10218);
xnor U10493 (N_10493,N_10100,N_10050);
or U10494 (N_10494,N_10201,N_10169);
or U10495 (N_10495,N_10165,N_10069);
and U10496 (N_10496,N_10243,N_10029);
nand U10497 (N_10497,N_10037,N_10008);
nand U10498 (N_10498,N_10043,N_10015);
nand U10499 (N_10499,N_10160,N_10040);
nor U10500 (N_10500,N_10344,N_10431);
nand U10501 (N_10501,N_10472,N_10496);
and U10502 (N_10502,N_10339,N_10429);
nand U10503 (N_10503,N_10267,N_10368);
or U10504 (N_10504,N_10343,N_10308);
or U10505 (N_10505,N_10309,N_10325);
xor U10506 (N_10506,N_10361,N_10345);
nor U10507 (N_10507,N_10439,N_10485);
nand U10508 (N_10508,N_10314,N_10294);
nand U10509 (N_10509,N_10434,N_10328);
xor U10510 (N_10510,N_10357,N_10283);
nand U10511 (N_10511,N_10480,N_10385);
or U10512 (N_10512,N_10404,N_10486);
nor U10513 (N_10513,N_10287,N_10256);
xnor U10514 (N_10514,N_10278,N_10280);
nor U10515 (N_10515,N_10396,N_10377);
or U10516 (N_10516,N_10493,N_10448);
xnor U10517 (N_10517,N_10380,N_10461);
or U10518 (N_10518,N_10484,N_10464);
xor U10519 (N_10519,N_10335,N_10438);
xnor U10520 (N_10520,N_10497,N_10382);
nor U10521 (N_10521,N_10450,N_10250);
nand U10522 (N_10522,N_10299,N_10384);
and U10523 (N_10523,N_10435,N_10351);
or U10524 (N_10524,N_10410,N_10268);
and U10525 (N_10525,N_10284,N_10254);
nand U10526 (N_10526,N_10266,N_10264);
nand U10527 (N_10527,N_10282,N_10499);
or U10528 (N_10528,N_10370,N_10323);
and U10529 (N_10529,N_10457,N_10436);
and U10530 (N_10530,N_10408,N_10394);
and U10531 (N_10531,N_10476,N_10258);
nand U10532 (N_10532,N_10257,N_10298);
xnor U10533 (N_10533,N_10275,N_10333);
nor U10534 (N_10534,N_10399,N_10358);
and U10535 (N_10535,N_10467,N_10288);
nand U10536 (N_10536,N_10271,N_10261);
and U10537 (N_10537,N_10400,N_10419);
nor U10538 (N_10538,N_10468,N_10341);
or U10539 (N_10539,N_10348,N_10273);
and U10540 (N_10540,N_10255,N_10423);
nand U10541 (N_10541,N_10393,N_10455);
nor U10542 (N_10542,N_10313,N_10312);
and U10543 (N_10543,N_10379,N_10277);
xor U10544 (N_10544,N_10458,N_10296);
or U10545 (N_10545,N_10383,N_10405);
or U10546 (N_10546,N_10318,N_10303);
xor U10547 (N_10547,N_10445,N_10425);
xor U10548 (N_10548,N_10432,N_10437);
or U10549 (N_10549,N_10477,N_10494);
or U10550 (N_10550,N_10286,N_10409);
or U10551 (N_10551,N_10490,N_10498);
nand U10552 (N_10552,N_10363,N_10305);
and U10553 (N_10553,N_10320,N_10465);
xnor U10554 (N_10554,N_10362,N_10371);
nand U10555 (N_10555,N_10412,N_10297);
nand U10556 (N_10556,N_10413,N_10406);
or U10557 (N_10557,N_10420,N_10386);
and U10558 (N_10558,N_10260,N_10418);
xnor U10559 (N_10559,N_10359,N_10291);
nor U10560 (N_10560,N_10392,N_10442);
and U10561 (N_10561,N_10475,N_10454);
nand U10562 (N_10562,N_10466,N_10263);
and U10563 (N_10563,N_10331,N_10471);
and U10564 (N_10564,N_10346,N_10366);
nor U10565 (N_10565,N_10430,N_10272);
and U10566 (N_10566,N_10456,N_10274);
nor U10567 (N_10567,N_10381,N_10342);
and U10568 (N_10568,N_10462,N_10350);
xnor U10569 (N_10569,N_10451,N_10424);
xor U10570 (N_10570,N_10428,N_10495);
nor U10571 (N_10571,N_10302,N_10355);
xor U10572 (N_10572,N_10460,N_10444);
and U10573 (N_10573,N_10478,N_10353);
xnor U10574 (N_10574,N_10492,N_10337);
nor U10575 (N_10575,N_10321,N_10292);
nor U10576 (N_10576,N_10415,N_10372);
nand U10577 (N_10577,N_10293,N_10262);
xnor U10578 (N_10578,N_10452,N_10483);
and U10579 (N_10579,N_10446,N_10447);
and U10580 (N_10580,N_10290,N_10369);
nand U10581 (N_10581,N_10301,N_10365);
and U10582 (N_10582,N_10375,N_10440);
and U10583 (N_10583,N_10334,N_10367);
or U10584 (N_10584,N_10364,N_10330);
or U10585 (N_10585,N_10417,N_10388);
xor U10586 (N_10586,N_10402,N_10403);
and U10587 (N_10587,N_10398,N_10326);
nand U10588 (N_10588,N_10253,N_10397);
and U10589 (N_10589,N_10259,N_10387);
xor U10590 (N_10590,N_10269,N_10481);
nor U10591 (N_10591,N_10307,N_10354);
nand U10592 (N_10592,N_10443,N_10470);
nor U10593 (N_10593,N_10395,N_10374);
or U10594 (N_10594,N_10352,N_10251);
nand U10595 (N_10595,N_10304,N_10252);
or U10596 (N_10596,N_10449,N_10306);
and U10597 (N_10597,N_10391,N_10347);
nand U10598 (N_10598,N_10285,N_10279);
or U10599 (N_10599,N_10427,N_10336);
and U10600 (N_10600,N_10376,N_10289);
nor U10601 (N_10601,N_10340,N_10401);
or U10602 (N_10602,N_10389,N_10329);
or U10603 (N_10603,N_10373,N_10300);
nand U10604 (N_10604,N_10473,N_10421);
or U10605 (N_10605,N_10360,N_10265);
or U10606 (N_10606,N_10317,N_10414);
or U10607 (N_10607,N_10378,N_10407);
nand U10608 (N_10608,N_10482,N_10441);
nor U10609 (N_10609,N_10327,N_10433);
and U10610 (N_10610,N_10479,N_10319);
xnor U10611 (N_10611,N_10422,N_10488);
and U10612 (N_10612,N_10453,N_10281);
nor U10613 (N_10613,N_10487,N_10349);
and U10614 (N_10614,N_10459,N_10356);
or U10615 (N_10615,N_10474,N_10390);
and U10616 (N_10616,N_10310,N_10316);
nand U10617 (N_10617,N_10426,N_10270);
or U10618 (N_10618,N_10411,N_10469);
and U10619 (N_10619,N_10463,N_10295);
or U10620 (N_10620,N_10324,N_10276);
and U10621 (N_10621,N_10491,N_10311);
nand U10622 (N_10622,N_10338,N_10315);
nor U10623 (N_10623,N_10332,N_10416);
or U10624 (N_10624,N_10489,N_10322);
nand U10625 (N_10625,N_10300,N_10335);
xor U10626 (N_10626,N_10282,N_10399);
xor U10627 (N_10627,N_10287,N_10408);
or U10628 (N_10628,N_10465,N_10484);
or U10629 (N_10629,N_10325,N_10384);
and U10630 (N_10630,N_10359,N_10341);
xor U10631 (N_10631,N_10252,N_10272);
xnor U10632 (N_10632,N_10365,N_10316);
nand U10633 (N_10633,N_10315,N_10480);
or U10634 (N_10634,N_10476,N_10499);
xnor U10635 (N_10635,N_10264,N_10418);
xnor U10636 (N_10636,N_10366,N_10371);
xor U10637 (N_10637,N_10295,N_10438);
and U10638 (N_10638,N_10317,N_10339);
nand U10639 (N_10639,N_10445,N_10327);
nand U10640 (N_10640,N_10477,N_10355);
or U10641 (N_10641,N_10477,N_10318);
nor U10642 (N_10642,N_10394,N_10284);
xnor U10643 (N_10643,N_10431,N_10301);
nor U10644 (N_10644,N_10285,N_10275);
xnor U10645 (N_10645,N_10480,N_10327);
and U10646 (N_10646,N_10360,N_10316);
and U10647 (N_10647,N_10341,N_10371);
nand U10648 (N_10648,N_10465,N_10391);
xnor U10649 (N_10649,N_10363,N_10410);
nand U10650 (N_10650,N_10493,N_10276);
xor U10651 (N_10651,N_10253,N_10405);
or U10652 (N_10652,N_10316,N_10333);
nor U10653 (N_10653,N_10456,N_10463);
or U10654 (N_10654,N_10298,N_10393);
xor U10655 (N_10655,N_10255,N_10410);
or U10656 (N_10656,N_10467,N_10270);
and U10657 (N_10657,N_10288,N_10463);
or U10658 (N_10658,N_10439,N_10279);
nand U10659 (N_10659,N_10309,N_10411);
xor U10660 (N_10660,N_10300,N_10304);
and U10661 (N_10661,N_10467,N_10343);
or U10662 (N_10662,N_10343,N_10348);
and U10663 (N_10663,N_10382,N_10366);
nor U10664 (N_10664,N_10355,N_10335);
and U10665 (N_10665,N_10257,N_10275);
nor U10666 (N_10666,N_10300,N_10449);
nand U10667 (N_10667,N_10499,N_10369);
nand U10668 (N_10668,N_10286,N_10272);
or U10669 (N_10669,N_10304,N_10348);
or U10670 (N_10670,N_10415,N_10282);
or U10671 (N_10671,N_10402,N_10373);
xnor U10672 (N_10672,N_10302,N_10388);
xnor U10673 (N_10673,N_10495,N_10298);
nand U10674 (N_10674,N_10404,N_10490);
nor U10675 (N_10675,N_10471,N_10475);
and U10676 (N_10676,N_10346,N_10385);
and U10677 (N_10677,N_10403,N_10279);
nor U10678 (N_10678,N_10496,N_10498);
or U10679 (N_10679,N_10496,N_10387);
nor U10680 (N_10680,N_10322,N_10419);
or U10681 (N_10681,N_10428,N_10270);
and U10682 (N_10682,N_10468,N_10414);
xor U10683 (N_10683,N_10312,N_10463);
nor U10684 (N_10684,N_10485,N_10427);
nand U10685 (N_10685,N_10340,N_10344);
nand U10686 (N_10686,N_10262,N_10264);
and U10687 (N_10687,N_10327,N_10383);
and U10688 (N_10688,N_10312,N_10250);
nand U10689 (N_10689,N_10436,N_10283);
nand U10690 (N_10690,N_10496,N_10331);
and U10691 (N_10691,N_10258,N_10397);
nor U10692 (N_10692,N_10456,N_10305);
xor U10693 (N_10693,N_10399,N_10318);
nand U10694 (N_10694,N_10283,N_10267);
nand U10695 (N_10695,N_10479,N_10492);
xor U10696 (N_10696,N_10459,N_10312);
xor U10697 (N_10697,N_10463,N_10265);
and U10698 (N_10698,N_10486,N_10471);
nand U10699 (N_10699,N_10263,N_10273);
nand U10700 (N_10700,N_10447,N_10457);
xnor U10701 (N_10701,N_10413,N_10423);
nor U10702 (N_10702,N_10316,N_10267);
xor U10703 (N_10703,N_10482,N_10418);
or U10704 (N_10704,N_10431,N_10406);
and U10705 (N_10705,N_10387,N_10295);
or U10706 (N_10706,N_10483,N_10485);
and U10707 (N_10707,N_10422,N_10433);
xor U10708 (N_10708,N_10355,N_10304);
nor U10709 (N_10709,N_10344,N_10437);
and U10710 (N_10710,N_10447,N_10385);
nand U10711 (N_10711,N_10431,N_10469);
nand U10712 (N_10712,N_10439,N_10418);
nor U10713 (N_10713,N_10380,N_10383);
or U10714 (N_10714,N_10312,N_10335);
nand U10715 (N_10715,N_10272,N_10315);
xor U10716 (N_10716,N_10339,N_10466);
nand U10717 (N_10717,N_10264,N_10378);
nor U10718 (N_10718,N_10340,N_10338);
xnor U10719 (N_10719,N_10411,N_10385);
and U10720 (N_10720,N_10254,N_10426);
and U10721 (N_10721,N_10331,N_10451);
nand U10722 (N_10722,N_10443,N_10257);
nand U10723 (N_10723,N_10467,N_10329);
and U10724 (N_10724,N_10315,N_10287);
nand U10725 (N_10725,N_10456,N_10453);
and U10726 (N_10726,N_10419,N_10250);
or U10727 (N_10727,N_10335,N_10367);
nand U10728 (N_10728,N_10256,N_10285);
and U10729 (N_10729,N_10341,N_10283);
and U10730 (N_10730,N_10262,N_10276);
or U10731 (N_10731,N_10326,N_10377);
or U10732 (N_10732,N_10411,N_10281);
nand U10733 (N_10733,N_10252,N_10448);
or U10734 (N_10734,N_10323,N_10274);
nor U10735 (N_10735,N_10320,N_10396);
or U10736 (N_10736,N_10318,N_10269);
and U10737 (N_10737,N_10415,N_10303);
nand U10738 (N_10738,N_10405,N_10302);
nand U10739 (N_10739,N_10387,N_10461);
nor U10740 (N_10740,N_10433,N_10401);
nand U10741 (N_10741,N_10450,N_10316);
nand U10742 (N_10742,N_10265,N_10465);
nor U10743 (N_10743,N_10460,N_10326);
or U10744 (N_10744,N_10495,N_10304);
and U10745 (N_10745,N_10471,N_10443);
nand U10746 (N_10746,N_10257,N_10485);
nor U10747 (N_10747,N_10388,N_10407);
xor U10748 (N_10748,N_10290,N_10388);
nand U10749 (N_10749,N_10345,N_10463);
nand U10750 (N_10750,N_10667,N_10593);
nand U10751 (N_10751,N_10562,N_10500);
nor U10752 (N_10752,N_10529,N_10651);
xor U10753 (N_10753,N_10618,N_10739);
and U10754 (N_10754,N_10502,N_10583);
or U10755 (N_10755,N_10708,N_10705);
or U10756 (N_10756,N_10700,N_10533);
nand U10757 (N_10757,N_10539,N_10512);
xor U10758 (N_10758,N_10588,N_10697);
nor U10759 (N_10759,N_10702,N_10590);
xor U10760 (N_10760,N_10693,N_10725);
and U10761 (N_10761,N_10535,N_10622);
nor U10762 (N_10762,N_10706,N_10517);
nand U10763 (N_10763,N_10654,N_10532);
nor U10764 (N_10764,N_10666,N_10672);
and U10765 (N_10765,N_10582,N_10735);
or U10766 (N_10766,N_10515,N_10731);
nor U10767 (N_10767,N_10685,N_10552);
nor U10768 (N_10768,N_10748,N_10668);
nand U10769 (N_10769,N_10686,N_10629);
and U10770 (N_10770,N_10743,N_10508);
nand U10771 (N_10771,N_10570,N_10712);
xnor U10772 (N_10772,N_10589,N_10594);
nand U10773 (N_10773,N_10558,N_10546);
nor U10774 (N_10774,N_10548,N_10742);
or U10775 (N_10775,N_10726,N_10604);
xor U10776 (N_10776,N_10691,N_10701);
nor U10777 (N_10777,N_10577,N_10692);
or U10778 (N_10778,N_10641,N_10608);
nor U10779 (N_10779,N_10660,N_10631);
nand U10780 (N_10780,N_10528,N_10613);
xor U10781 (N_10781,N_10607,N_10520);
nand U10782 (N_10782,N_10741,N_10513);
or U10783 (N_10783,N_10661,N_10561);
nor U10784 (N_10784,N_10531,N_10547);
nor U10785 (N_10785,N_10650,N_10713);
and U10786 (N_10786,N_10602,N_10614);
or U10787 (N_10787,N_10678,N_10524);
and U10788 (N_10788,N_10656,N_10521);
nand U10789 (N_10789,N_10597,N_10573);
or U10790 (N_10790,N_10703,N_10628);
nand U10791 (N_10791,N_10567,N_10633);
xor U10792 (N_10792,N_10550,N_10537);
xor U10793 (N_10793,N_10530,N_10647);
xor U10794 (N_10794,N_10584,N_10673);
nor U10795 (N_10795,N_10665,N_10729);
nand U10796 (N_10796,N_10715,N_10684);
or U10797 (N_10797,N_10542,N_10511);
and U10798 (N_10798,N_10683,N_10732);
xnor U10799 (N_10799,N_10566,N_10527);
xnor U10800 (N_10800,N_10695,N_10698);
xor U10801 (N_10801,N_10676,N_10572);
or U10802 (N_10802,N_10749,N_10643);
and U10803 (N_10803,N_10663,N_10620);
and U10804 (N_10804,N_10579,N_10564);
nand U10805 (N_10805,N_10525,N_10574);
or U10806 (N_10806,N_10680,N_10687);
nor U10807 (N_10807,N_10596,N_10545);
xor U10808 (N_10808,N_10734,N_10501);
xnor U10809 (N_10809,N_10670,N_10689);
and U10810 (N_10810,N_10506,N_10675);
and U10811 (N_10811,N_10642,N_10523);
nor U10812 (N_10812,N_10503,N_10627);
nand U10813 (N_10813,N_10541,N_10709);
xnor U10814 (N_10814,N_10728,N_10612);
nand U10815 (N_10815,N_10640,N_10652);
xnor U10816 (N_10816,N_10679,N_10635);
and U10817 (N_10817,N_10720,N_10690);
nand U10818 (N_10818,N_10704,N_10624);
xor U10819 (N_10819,N_10518,N_10578);
nor U10820 (N_10820,N_10677,N_10625);
nand U10821 (N_10821,N_10718,N_10601);
xor U10822 (N_10822,N_10540,N_10587);
or U10823 (N_10823,N_10509,N_10544);
or U10824 (N_10824,N_10747,N_10580);
and U10825 (N_10825,N_10559,N_10738);
or U10826 (N_10826,N_10662,N_10626);
and U10827 (N_10827,N_10658,N_10504);
and U10828 (N_10828,N_10674,N_10609);
xor U10829 (N_10829,N_10681,N_10611);
and U10830 (N_10830,N_10534,N_10737);
or U10831 (N_10831,N_10745,N_10645);
xor U10832 (N_10832,N_10505,N_10727);
nor U10833 (N_10833,N_10543,N_10616);
and U10834 (N_10834,N_10716,N_10646);
and U10835 (N_10835,N_10733,N_10638);
or U10836 (N_10836,N_10740,N_10600);
nand U10837 (N_10837,N_10710,N_10581);
or U10838 (N_10838,N_10610,N_10514);
nor U10839 (N_10839,N_10746,N_10551);
or U10840 (N_10840,N_10636,N_10526);
nand U10841 (N_10841,N_10592,N_10507);
or U10842 (N_10842,N_10717,N_10571);
nor U10843 (N_10843,N_10595,N_10659);
nand U10844 (N_10844,N_10724,N_10553);
and U10845 (N_10845,N_10634,N_10591);
nand U10846 (N_10846,N_10696,N_10707);
or U10847 (N_10847,N_10619,N_10669);
xnor U10848 (N_10848,N_10598,N_10730);
and U10849 (N_10849,N_10555,N_10694);
and U10850 (N_10850,N_10621,N_10575);
xor U10851 (N_10851,N_10671,N_10556);
and U10852 (N_10852,N_10576,N_10519);
nand U10853 (N_10853,N_10639,N_10649);
xor U10854 (N_10854,N_10653,N_10719);
or U10855 (N_10855,N_10599,N_10565);
nor U10856 (N_10856,N_10699,N_10615);
and U10857 (N_10857,N_10569,N_10585);
and U10858 (N_10858,N_10632,N_10688);
nand U10859 (N_10859,N_10722,N_10736);
nand U10860 (N_10860,N_10648,N_10554);
xor U10861 (N_10861,N_10657,N_10644);
xnor U10862 (N_10862,N_10721,N_10617);
and U10863 (N_10863,N_10603,N_10723);
nand U10864 (N_10864,N_10557,N_10560);
xor U10865 (N_10865,N_10605,N_10606);
and U10866 (N_10866,N_10563,N_10664);
or U10867 (N_10867,N_10549,N_10637);
and U10868 (N_10868,N_10586,N_10630);
nor U10869 (N_10869,N_10516,N_10744);
nand U10870 (N_10870,N_10536,N_10538);
or U10871 (N_10871,N_10714,N_10623);
xor U10872 (N_10872,N_10711,N_10655);
and U10873 (N_10873,N_10568,N_10682);
nand U10874 (N_10874,N_10510,N_10522);
and U10875 (N_10875,N_10725,N_10731);
xnor U10876 (N_10876,N_10577,N_10735);
and U10877 (N_10877,N_10701,N_10714);
nand U10878 (N_10878,N_10666,N_10728);
or U10879 (N_10879,N_10547,N_10726);
xor U10880 (N_10880,N_10583,N_10506);
xor U10881 (N_10881,N_10556,N_10525);
nor U10882 (N_10882,N_10727,N_10541);
or U10883 (N_10883,N_10667,N_10599);
nand U10884 (N_10884,N_10619,N_10738);
nand U10885 (N_10885,N_10736,N_10711);
nor U10886 (N_10886,N_10625,N_10516);
xor U10887 (N_10887,N_10678,N_10525);
and U10888 (N_10888,N_10535,N_10506);
xnor U10889 (N_10889,N_10551,N_10560);
and U10890 (N_10890,N_10649,N_10728);
or U10891 (N_10891,N_10677,N_10534);
and U10892 (N_10892,N_10739,N_10733);
nand U10893 (N_10893,N_10510,N_10736);
nand U10894 (N_10894,N_10681,N_10679);
and U10895 (N_10895,N_10557,N_10574);
and U10896 (N_10896,N_10654,N_10548);
nor U10897 (N_10897,N_10595,N_10744);
nor U10898 (N_10898,N_10660,N_10550);
or U10899 (N_10899,N_10662,N_10584);
or U10900 (N_10900,N_10612,N_10596);
or U10901 (N_10901,N_10699,N_10584);
xor U10902 (N_10902,N_10593,N_10531);
xor U10903 (N_10903,N_10619,N_10555);
nand U10904 (N_10904,N_10625,N_10699);
nor U10905 (N_10905,N_10640,N_10585);
or U10906 (N_10906,N_10539,N_10604);
nor U10907 (N_10907,N_10508,N_10629);
nor U10908 (N_10908,N_10573,N_10577);
nor U10909 (N_10909,N_10601,N_10674);
xor U10910 (N_10910,N_10590,N_10701);
nor U10911 (N_10911,N_10624,N_10711);
or U10912 (N_10912,N_10734,N_10624);
xor U10913 (N_10913,N_10611,N_10618);
nor U10914 (N_10914,N_10560,N_10513);
xor U10915 (N_10915,N_10544,N_10700);
nor U10916 (N_10916,N_10503,N_10718);
nand U10917 (N_10917,N_10691,N_10596);
nand U10918 (N_10918,N_10578,N_10659);
nor U10919 (N_10919,N_10692,N_10646);
or U10920 (N_10920,N_10564,N_10655);
or U10921 (N_10921,N_10647,N_10625);
and U10922 (N_10922,N_10639,N_10578);
nand U10923 (N_10923,N_10687,N_10554);
nand U10924 (N_10924,N_10729,N_10599);
and U10925 (N_10925,N_10648,N_10626);
xor U10926 (N_10926,N_10553,N_10554);
and U10927 (N_10927,N_10542,N_10745);
and U10928 (N_10928,N_10520,N_10706);
and U10929 (N_10929,N_10541,N_10519);
or U10930 (N_10930,N_10729,N_10662);
nor U10931 (N_10931,N_10526,N_10606);
or U10932 (N_10932,N_10553,N_10715);
or U10933 (N_10933,N_10610,N_10727);
nand U10934 (N_10934,N_10561,N_10531);
and U10935 (N_10935,N_10723,N_10703);
nor U10936 (N_10936,N_10674,N_10519);
xnor U10937 (N_10937,N_10516,N_10671);
and U10938 (N_10938,N_10517,N_10625);
or U10939 (N_10939,N_10721,N_10664);
xor U10940 (N_10940,N_10535,N_10655);
and U10941 (N_10941,N_10543,N_10713);
nor U10942 (N_10942,N_10539,N_10629);
or U10943 (N_10943,N_10620,N_10662);
nand U10944 (N_10944,N_10605,N_10662);
nor U10945 (N_10945,N_10705,N_10510);
or U10946 (N_10946,N_10580,N_10581);
and U10947 (N_10947,N_10618,N_10733);
and U10948 (N_10948,N_10564,N_10502);
nand U10949 (N_10949,N_10582,N_10550);
nor U10950 (N_10950,N_10638,N_10630);
xnor U10951 (N_10951,N_10671,N_10692);
xnor U10952 (N_10952,N_10662,N_10744);
xnor U10953 (N_10953,N_10533,N_10505);
or U10954 (N_10954,N_10696,N_10670);
or U10955 (N_10955,N_10644,N_10689);
nor U10956 (N_10956,N_10518,N_10654);
nand U10957 (N_10957,N_10616,N_10696);
and U10958 (N_10958,N_10532,N_10710);
nor U10959 (N_10959,N_10598,N_10602);
xnor U10960 (N_10960,N_10527,N_10617);
nand U10961 (N_10961,N_10527,N_10563);
nor U10962 (N_10962,N_10516,N_10528);
and U10963 (N_10963,N_10533,N_10696);
and U10964 (N_10964,N_10579,N_10640);
nand U10965 (N_10965,N_10624,N_10589);
and U10966 (N_10966,N_10721,N_10719);
xor U10967 (N_10967,N_10512,N_10545);
nand U10968 (N_10968,N_10511,N_10571);
nand U10969 (N_10969,N_10663,N_10528);
or U10970 (N_10970,N_10505,N_10611);
or U10971 (N_10971,N_10663,N_10638);
xor U10972 (N_10972,N_10713,N_10517);
or U10973 (N_10973,N_10562,N_10566);
and U10974 (N_10974,N_10742,N_10545);
nor U10975 (N_10975,N_10624,N_10596);
xor U10976 (N_10976,N_10592,N_10699);
nor U10977 (N_10977,N_10622,N_10637);
xnor U10978 (N_10978,N_10583,N_10637);
nand U10979 (N_10979,N_10746,N_10527);
nor U10980 (N_10980,N_10665,N_10529);
or U10981 (N_10981,N_10630,N_10518);
or U10982 (N_10982,N_10695,N_10550);
or U10983 (N_10983,N_10575,N_10733);
nand U10984 (N_10984,N_10676,N_10517);
xor U10985 (N_10985,N_10711,N_10627);
and U10986 (N_10986,N_10736,N_10665);
nor U10987 (N_10987,N_10671,N_10666);
nand U10988 (N_10988,N_10732,N_10725);
nor U10989 (N_10989,N_10533,N_10655);
and U10990 (N_10990,N_10703,N_10575);
and U10991 (N_10991,N_10546,N_10743);
or U10992 (N_10992,N_10543,N_10715);
nor U10993 (N_10993,N_10570,N_10616);
xor U10994 (N_10994,N_10621,N_10707);
nor U10995 (N_10995,N_10614,N_10594);
xor U10996 (N_10996,N_10542,N_10667);
xnor U10997 (N_10997,N_10691,N_10539);
xor U10998 (N_10998,N_10661,N_10508);
or U10999 (N_10999,N_10555,N_10500);
nand U11000 (N_11000,N_10898,N_10809);
nor U11001 (N_11001,N_10967,N_10916);
and U11002 (N_11002,N_10975,N_10751);
xor U11003 (N_11003,N_10804,N_10991);
nor U11004 (N_11004,N_10905,N_10919);
and U11005 (N_11005,N_10912,N_10911);
xnor U11006 (N_11006,N_10946,N_10777);
nand U11007 (N_11007,N_10846,N_10948);
nand U11008 (N_11008,N_10845,N_10873);
and U11009 (N_11009,N_10821,N_10936);
xnor U11010 (N_11010,N_10836,N_10806);
nand U11011 (N_11011,N_10763,N_10790);
xor U11012 (N_11012,N_10849,N_10909);
nand U11013 (N_11013,N_10833,N_10877);
nor U11014 (N_11014,N_10997,N_10918);
nor U11015 (N_11015,N_10866,N_10860);
and U11016 (N_11016,N_10856,N_10828);
and U11017 (N_11017,N_10843,N_10965);
nor U11018 (N_11018,N_10811,N_10867);
nand U11019 (N_11019,N_10782,N_10779);
and U11020 (N_11020,N_10889,N_10924);
or U11021 (N_11021,N_10830,N_10848);
or U11022 (N_11022,N_10935,N_10954);
and U11023 (N_11023,N_10978,N_10944);
and U11024 (N_11024,N_10875,N_10953);
xor U11025 (N_11025,N_10966,N_10945);
or U11026 (N_11026,N_10955,N_10926);
and U11027 (N_11027,N_10835,N_10832);
nor U11028 (N_11028,N_10847,N_10915);
nor U11029 (N_11029,N_10893,N_10801);
or U11030 (N_11030,N_10822,N_10864);
nor U11031 (N_11031,N_10794,N_10810);
or U11032 (N_11032,N_10755,N_10929);
or U11033 (N_11033,N_10921,N_10939);
nor U11034 (N_11034,N_10983,N_10901);
and U11035 (N_11035,N_10895,N_10899);
nand U11036 (N_11036,N_10831,N_10827);
or U11037 (N_11037,N_10976,N_10994);
nand U11038 (N_11038,N_10868,N_10979);
xor U11039 (N_11039,N_10778,N_10813);
or U11040 (N_11040,N_10840,N_10906);
nand U11041 (N_11041,N_10816,N_10995);
nor U11042 (N_11042,N_10753,N_10826);
and U11043 (N_11043,N_10904,N_10869);
nand U11044 (N_11044,N_10781,N_10784);
or U11045 (N_11045,N_10783,N_10770);
and U11046 (N_11046,N_10817,N_10964);
and U11047 (N_11047,N_10787,N_10850);
xnor U11048 (N_11048,N_10851,N_10934);
xor U11049 (N_11049,N_10780,N_10768);
nor U11050 (N_11050,N_10969,N_10892);
and U11051 (N_11051,N_10758,N_10807);
xnor U11052 (N_11052,N_10880,N_10957);
or U11053 (N_11053,N_10890,N_10818);
and U11054 (N_11054,N_10928,N_10881);
nor U11055 (N_11055,N_10852,N_10886);
or U11056 (N_11056,N_10960,N_10767);
and U11057 (N_11057,N_10891,N_10762);
or U11058 (N_11058,N_10839,N_10878);
nand U11059 (N_11059,N_10764,N_10981);
nand U11060 (N_11060,N_10756,N_10863);
or U11061 (N_11061,N_10773,N_10925);
xor U11062 (N_11062,N_10883,N_10861);
nor U11063 (N_11063,N_10894,N_10799);
xor U11064 (N_11064,N_10797,N_10865);
xnor U11065 (N_11065,N_10927,N_10876);
xor U11066 (N_11066,N_10973,N_10859);
xor U11067 (N_11067,N_10952,N_10940);
or U11068 (N_11068,N_10949,N_10992);
or U11069 (N_11069,N_10998,N_10897);
or U11070 (N_11070,N_10943,N_10908);
xnor U11071 (N_11071,N_10947,N_10795);
and U11072 (N_11072,N_10750,N_10988);
and U11073 (N_11073,N_10792,N_10844);
or U11074 (N_11074,N_10942,N_10814);
nor U11075 (N_11075,N_10772,N_10841);
nand U11076 (N_11076,N_10999,N_10900);
nand U11077 (N_11077,N_10803,N_10775);
and U11078 (N_11078,N_10958,N_10815);
or U11079 (N_11079,N_10902,N_10785);
xor U11080 (N_11080,N_10879,N_10996);
xor U11081 (N_11081,N_10956,N_10903);
nand U11082 (N_11082,N_10941,N_10823);
or U11083 (N_11083,N_10808,N_10771);
or U11084 (N_11084,N_10788,N_10882);
nand U11085 (N_11085,N_10951,N_10933);
nand U11086 (N_11086,N_10987,N_10907);
nand U11087 (N_11087,N_10761,N_10950);
nand U11088 (N_11088,N_10990,N_10800);
xnor U11089 (N_11089,N_10855,N_10765);
nor U11090 (N_11090,N_10885,N_10805);
and U11091 (N_11091,N_10962,N_10989);
and U11092 (N_11092,N_10910,N_10970);
xnor U11093 (N_11093,N_10872,N_10963);
and U11094 (N_11094,N_10874,N_10824);
and U11095 (N_11095,N_10798,N_10774);
xor U11096 (N_11096,N_10793,N_10853);
xor U11097 (N_11097,N_10789,N_10884);
nor U11098 (N_11098,N_10791,N_10854);
nand U11099 (N_11099,N_10932,N_10959);
nor U11100 (N_11100,N_10862,N_10972);
nor U11101 (N_11101,N_10982,N_10838);
nand U11102 (N_11102,N_10837,N_10819);
xnor U11103 (N_11103,N_10796,N_10977);
nor U11104 (N_11104,N_10974,N_10993);
and U11105 (N_11105,N_10887,N_10812);
xnor U11106 (N_11106,N_10923,N_10985);
nand U11107 (N_11107,N_10786,N_10829);
or U11108 (N_11108,N_10769,N_10984);
xnor U11109 (N_11109,N_10931,N_10820);
and U11110 (N_11110,N_10757,N_10914);
xor U11111 (N_11111,N_10760,N_10986);
nand U11112 (N_11112,N_10870,N_10825);
nor U11113 (N_11113,N_10922,N_10896);
nor U11114 (N_11114,N_10759,N_10968);
xnor U11115 (N_11115,N_10913,N_10920);
nand U11116 (N_11116,N_10858,N_10971);
nor U11117 (N_11117,N_10917,N_10776);
or U11118 (N_11118,N_10871,N_10752);
xor U11119 (N_11119,N_10857,N_10961);
xor U11120 (N_11120,N_10980,N_10842);
or U11121 (N_11121,N_10766,N_10834);
nor U11122 (N_11122,N_10802,N_10754);
xor U11123 (N_11123,N_10930,N_10888);
or U11124 (N_11124,N_10937,N_10938);
and U11125 (N_11125,N_10784,N_10852);
and U11126 (N_11126,N_10912,N_10941);
and U11127 (N_11127,N_10879,N_10987);
or U11128 (N_11128,N_10750,N_10862);
and U11129 (N_11129,N_10845,N_10821);
nor U11130 (N_11130,N_10998,N_10754);
nor U11131 (N_11131,N_10961,N_10835);
nand U11132 (N_11132,N_10846,N_10873);
nor U11133 (N_11133,N_10793,N_10941);
or U11134 (N_11134,N_10849,N_10869);
nor U11135 (N_11135,N_10771,N_10827);
and U11136 (N_11136,N_10945,N_10900);
xnor U11137 (N_11137,N_10959,N_10803);
nand U11138 (N_11138,N_10844,N_10806);
nor U11139 (N_11139,N_10913,N_10955);
or U11140 (N_11140,N_10933,N_10998);
and U11141 (N_11141,N_10848,N_10872);
nor U11142 (N_11142,N_10767,N_10912);
nand U11143 (N_11143,N_10921,N_10908);
nand U11144 (N_11144,N_10825,N_10837);
xnor U11145 (N_11145,N_10998,N_10766);
and U11146 (N_11146,N_10781,N_10976);
nand U11147 (N_11147,N_10985,N_10760);
or U11148 (N_11148,N_10803,N_10878);
or U11149 (N_11149,N_10856,N_10937);
nand U11150 (N_11150,N_10829,N_10938);
and U11151 (N_11151,N_10757,N_10878);
and U11152 (N_11152,N_10950,N_10795);
or U11153 (N_11153,N_10816,N_10965);
nand U11154 (N_11154,N_10934,N_10976);
xnor U11155 (N_11155,N_10980,N_10912);
nor U11156 (N_11156,N_10893,N_10865);
nand U11157 (N_11157,N_10846,N_10830);
nand U11158 (N_11158,N_10811,N_10949);
or U11159 (N_11159,N_10866,N_10851);
and U11160 (N_11160,N_10908,N_10800);
and U11161 (N_11161,N_10957,N_10868);
xnor U11162 (N_11162,N_10887,N_10927);
or U11163 (N_11163,N_10881,N_10771);
or U11164 (N_11164,N_10932,N_10869);
or U11165 (N_11165,N_10831,N_10956);
nor U11166 (N_11166,N_10969,N_10962);
nand U11167 (N_11167,N_10950,N_10952);
nand U11168 (N_11168,N_10877,N_10983);
nor U11169 (N_11169,N_10854,N_10814);
and U11170 (N_11170,N_10973,N_10884);
and U11171 (N_11171,N_10757,N_10840);
nor U11172 (N_11172,N_10829,N_10899);
and U11173 (N_11173,N_10792,N_10892);
nand U11174 (N_11174,N_10825,N_10816);
nor U11175 (N_11175,N_10798,N_10870);
xnor U11176 (N_11176,N_10879,N_10939);
and U11177 (N_11177,N_10856,N_10763);
xnor U11178 (N_11178,N_10845,N_10947);
xnor U11179 (N_11179,N_10851,N_10964);
nor U11180 (N_11180,N_10954,N_10811);
xor U11181 (N_11181,N_10990,N_10892);
or U11182 (N_11182,N_10945,N_10932);
nor U11183 (N_11183,N_10961,N_10868);
or U11184 (N_11184,N_10788,N_10837);
nand U11185 (N_11185,N_10880,N_10750);
and U11186 (N_11186,N_10951,N_10926);
xor U11187 (N_11187,N_10773,N_10996);
nor U11188 (N_11188,N_10951,N_10752);
xnor U11189 (N_11189,N_10853,N_10935);
or U11190 (N_11190,N_10803,N_10958);
or U11191 (N_11191,N_10903,N_10887);
or U11192 (N_11192,N_10865,N_10841);
xnor U11193 (N_11193,N_10791,N_10886);
nand U11194 (N_11194,N_10874,N_10997);
nand U11195 (N_11195,N_10870,N_10845);
nand U11196 (N_11196,N_10989,N_10898);
nand U11197 (N_11197,N_10828,N_10887);
or U11198 (N_11198,N_10840,N_10927);
nand U11199 (N_11199,N_10951,N_10902);
xor U11200 (N_11200,N_10767,N_10873);
xnor U11201 (N_11201,N_10783,N_10985);
xor U11202 (N_11202,N_10817,N_10865);
and U11203 (N_11203,N_10811,N_10927);
and U11204 (N_11204,N_10990,N_10865);
xnor U11205 (N_11205,N_10831,N_10955);
and U11206 (N_11206,N_10832,N_10859);
nor U11207 (N_11207,N_10986,N_10964);
xor U11208 (N_11208,N_10797,N_10781);
nor U11209 (N_11209,N_10904,N_10830);
nor U11210 (N_11210,N_10884,N_10978);
and U11211 (N_11211,N_10915,N_10957);
and U11212 (N_11212,N_10988,N_10937);
xnor U11213 (N_11213,N_10991,N_10874);
nand U11214 (N_11214,N_10925,N_10998);
or U11215 (N_11215,N_10773,N_10985);
or U11216 (N_11216,N_10884,N_10938);
or U11217 (N_11217,N_10762,N_10830);
xnor U11218 (N_11218,N_10956,N_10933);
nor U11219 (N_11219,N_10849,N_10950);
nor U11220 (N_11220,N_10863,N_10768);
nor U11221 (N_11221,N_10841,N_10906);
xnor U11222 (N_11222,N_10758,N_10954);
nand U11223 (N_11223,N_10883,N_10994);
nand U11224 (N_11224,N_10909,N_10770);
or U11225 (N_11225,N_10825,N_10875);
xor U11226 (N_11226,N_10810,N_10873);
xnor U11227 (N_11227,N_10989,N_10968);
nand U11228 (N_11228,N_10814,N_10786);
nor U11229 (N_11229,N_10977,N_10836);
or U11230 (N_11230,N_10779,N_10806);
and U11231 (N_11231,N_10955,N_10813);
nor U11232 (N_11232,N_10852,N_10793);
nand U11233 (N_11233,N_10967,N_10804);
or U11234 (N_11234,N_10959,N_10789);
nor U11235 (N_11235,N_10941,N_10980);
nor U11236 (N_11236,N_10982,N_10925);
or U11237 (N_11237,N_10758,N_10940);
and U11238 (N_11238,N_10799,N_10939);
nand U11239 (N_11239,N_10964,N_10898);
or U11240 (N_11240,N_10754,N_10797);
nand U11241 (N_11241,N_10777,N_10897);
and U11242 (N_11242,N_10790,N_10935);
xnor U11243 (N_11243,N_10756,N_10835);
nand U11244 (N_11244,N_10816,N_10990);
and U11245 (N_11245,N_10768,N_10773);
nand U11246 (N_11246,N_10989,N_10897);
or U11247 (N_11247,N_10904,N_10907);
nand U11248 (N_11248,N_10987,N_10966);
nand U11249 (N_11249,N_10809,N_10751);
nor U11250 (N_11250,N_11211,N_11166);
or U11251 (N_11251,N_11153,N_11231);
xnor U11252 (N_11252,N_11239,N_11040);
and U11253 (N_11253,N_11070,N_11057);
nor U11254 (N_11254,N_11140,N_11125);
xor U11255 (N_11255,N_11074,N_11111);
and U11256 (N_11256,N_11178,N_11236);
and U11257 (N_11257,N_11158,N_11234);
nor U11258 (N_11258,N_11007,N_11180);
and U11259 (N_11259,N_11008,N_11096);
nand U11260 (N_11260,N_11184,N_11089);
xor U11261 (N_11261,N_11064,N_11109);
or U11262 (N_11262,N_11152,N_11077);
nand U11263 (N_11263,N_11208,N_11058);
xor U11264 (N_11264,N_11138,N_11018);
or U11265 (N_11265,N_11047,N_11122);
nor U11266 (N_11266,N_11176,N_11029);
xnor U11267 (N_11267,N_11151,N_11078);
xnor U11268 (N_11268,N_11145,N_11173);
or U11269 (N_11269,N_11130,N_11023);
xnor U11270 (N_11270,N_11225,N_11101);
nor U11271 (N_11271,N_11220,N_11126);
or U11272 (N_11272,N_11160,N_11249);
and U11273 (N_11273,N_11168,N_11226);
nand U11274 (N_11274,N_11033,N_11146);
xor U11275 (N_11275,N_11072,N_11024);
and U11276 (N_11276,N_11161,N_11013);
nand U11277 (N_11277,N_11043,N_11201);
or U11278 (N_11278,N_11035,N_11051);
or U11279 (N_11279,N_11190,N_11167);
nor U11280 (N_11280,N_11171,N_11163);
nand U11281 (N_11281,N_11149,N_11221);
or U11282 (N_11282,N_11091,N_11147);
and U11283 (N_11283,N_11244,N_11229);
nand U11284 (N_11284,N_11192,N_11009);
nor U11285 (N_11285,N_11218,N_11105);
nor U11286 (N_11286,N_11039,N_11195);
nand U11287 (N_11287,N_11162,N_11174);
xor U11288 (N_11288,N_11045,N_11020);
nand U11289 (N_11289,N_11059,N_11079);
nand U11290 (N_11290,N_11081,N_11127);
nor U11291 (N_11291,N_11238,N_11183);
xnor U11292 (N_11292,N_11002,N_11011);
or U11293 (N_11293,N_11215,N_11112);
nand U11294 (N_11294,N_11247,N_11200);
or U11295 (N_11295,N_11102,N_11015);
nand U11296 (N_11296,N_11243,N_11054);
and U11297 (N_11297,N_11068,N_11005);
and U11298 (N_11298,N_11000,N_11099);
xnor U11299 (N_11299,N_11141,N_11155);
and U11300 (N_11300,N_11212,N_11085);
xnor U11301 (N_11301,N_11094,N_11139);
xnor U11302 (N_11302,N_11165,N_11114);
nor U11303 (N_11303,N_11022,N_11026);
or U11304 (N_11304,N_11076,N_11044);
xor U11305 (N_11305,N_11093,N_11108);
or U11306 (N_11306,N_11073,N_11038);
nor U11307 (N_11307,N_11242,N_11027);
or U11308 (N_11308,N_11062,N_11144);
and U11309 (N_11309,N_11087,N_11071);
xnor U11310 (N_11310,N_11082,N_11206);
and U11311 (N_11311,N_11150,N_11143);
nand U11312 (N_11312,N_11197,N_11217);
nor U11313 (N_11313,N_11034,N_11124);
xor U11314 (N_11314,N_11003,N_11100);
and U11315 (N_11315,N_11010,N_11154);
or U11316 (N_11316,N_11121,N_11188);
and U11317 (N_11317,N_11028,N_11025);
xnor U11318 (N_11318,N_11065,N_11001);
nand U11319 (N_11319,N_11240,N_11129);
and U11320 (N_11320,N_11187,N_11063);
xnor U11321 (N_11321,N_11032,N_11169);
nor U11322 (N_11322,N_11230,N_11223);
or U11323 (N_11323,N_11050,N_11086);
and U11324 (N_11324,N_11172,N_11056);
nand U11325 (N_11325,N_11136,N_11104);
nor U11326 (N_11326,N_11128,N_11041);
and U11327 (N_11327,N_11170,N_11157);
and U11328 (N_11328,N_11060,N_11014);
nor U11329 (N_11329,N_11019,N_11103);
xor U11330 (N_11330,N_11012,N_11098);
nand U11331 (N_11331,N_11030,N_11132);
xor U11332 (N_11332,N_11037,N_11235);
nor U11333 (N_11333,N_11092,N_11049);
nor U11334 (N_11334,N_11042,N_11036);
and U11335 (N_11335,N_11069,N_11232);
and U11336 (N_11336,N_11194,N_11189);
or U11337 (N_11337,N_11216,N_11181);
nand U11338 (N_11338,N_11248,N_11135);
nand U11339 (N_11339,N_11237,N_11137);
nand U11340 (N_11340,N_11116,N_11210);
and U11341 (N_11341,N_11193,N_11052);
nor U11342 (N_11342,N_11066,N_11241);
or U11343 (N_11343,N_11118,N_11205);
xor U11344 (N_11344,N_11134,N_11090);
and U11345 (N_11345,N_11227,N_11246);
or U11346 (N_11346,N_11083,N_11016);
nand U11347 (N_11347,N_11075,N_11055);
nor U11348 (N_11348,N_11107,N_11115);
or U11349 (N_11349,N_11209,N_11061);
nand U11350 (N_11350,N_11133,N_11123);
and U11351 (N_11351,N_11175,N_11204);
or U11352 (N_11352,N_11021,N_11080);
xor U11353 (N_11353,N_11191,N_11095);
nor U11354 (N_11354,N_11048,N_11031);
or U11355 (N_11355,N_11214,N_11017);
xor U11356 (N_11356,N_11159,N_11233);
nand U11357 (N_11357,N_11179,N_11119);
and U11358 (N_11358,N_11113,N_11120);
and U11359 (N_11359,N_11142,N_11198);
and U11360 (N_11360,N_11156,N_11164);
nand U11361 (N_11361,N_11182,N_11110);
and U11362 (N_11362,N_11245,N_11228);
nand U11363 (N_11363,N_11117,N_11004);
nor U11364 (N_11364,N_11046,N_11053);
nor U11365 (N_11365,N_11203,N_11219);
nand U11366 (N_11366,N_11006,N_11088);
or U11367 (N_11367,N_11106,N_11148);
or U11368 (N_11368,N_11202,N_11084);
nor U11369 (N_11369,N_11222,N_11199);
xor U11370 (N_11370,N_11186,N_11196);
nand U11371 (N_11371,N_11177,N_11067);
or U11372 (N_11372,N_11097,N_11185);
nand U11373 (N_11373,N_11207,N_11213);
nor U11374 (N_11374,N_11131,N_11224);
or U11375 (N_11375,N_11093,N_11138);
nor U11376 (N_11376,N_11152,N_11244);
xnor U11377 (N_11377,N_11215,N_11037);
and U11378 (N_11378,N_11097,N_11243);
and U11379 (N_11379,N_11084,N_11222);
xor U11380 (N_11380,N_11080,N_11067);
nor U11381 (N_11381,N_11062,N_11180);
or U11382 (N_11382,N_11168,N_11138);
nand U11383 (N_11383,N_11006,N_11060);
and U11384 (N_11384,N_11066,N_11029);
and U11385 (N_11385,N_11073,N_11174);
or U11386 (N_11386,N_11090,N_11160);
nor U11387 (N_11387,N_11221,N_11006);
nand U11388 (N_11388,N_11175,N_11075);
or U11389 (N_11389,N_11211,N_11148);
nand U11390 (N_11390,N_11024,N_11111);
or U11391 (N_11391,N_11137,N_11045);
xnor U11392 (N_11392,N_11089,N_11050);
xor U11393 (N_11393,N_11163,N_11027);
xnor U11394 (N_11394,N_11062,N_11147);
xor U11395 (N_11395,N_11212,N_11131);
or U11396 (N_11396,N_11025,N_11034);
xnor U11397 (N_11397,N_11017,N_11019);
and U11398 (N_11398,N_11118,N_11171);
nor U11399 (N_11399,N_11133,N_11240);
or U11400 (N_11400,N_11005,N_11229);
or U11401 (N_11401,N_11185,N_11013);
or U11402 (N_11402,N_11152,N_11105);
or U11403 (N_11403,N_11160,N_11168);
nand U11404 (N_11404,N_11059,N_11053);
or U11405 (N_11405,N_11228,N_11188);
and U11406 (N_11406,N_11072,N_11092);
xor U11407 (N_11407,N_11188,N_11034);
nand U11408 (N_11408,N_11163,N_11214);
nand U11409 (N_11409,N_11204,N_11201);
nand U11410 (N_11410,N_11191,N_11073);
and U11411 (N_11411,N_11165,N_11147);
nor U11412 (N_11412,N_11232,N_11249);
xnor U11413 (N_11413,N_11166,N_11069);
nand U11414 (N_11414,N_11188,N_11203);
or U11415 (N_11415,N_11239,N_11179);
nand U11416 (N_11416,N_11132,N_11028);
or U11417 (N_11417,N_11041,N_11118);
or U11418 (N_11418,N_11061,N_11086);
nand U11419 (N_11419,N_11229,N_11249);
and U11420 (N_11420,N_11143,N_11236);
xor U11421 (N_11421,N_11038,N_11134);
nor U11422 (N_11422,N_11054,N_11114);
xnor U11423 (N_11423,N_11161,N_11117);
nor U11424 (N_11424,N_11046,N_11067);
nor U11425 (N_11425,N_11028,N_11192);
and U11426 (N_11426,N_11046,N_11043);
nor U11427 (N_11427,N_11095,N_11063);
and U11428 (N_11428,N_11090,N_11148);
or U11429 (N_11429,N_11006,N_11007);
or U11430 (N_11430,N_11146,N_11002);
nor U11431 (N_11431,N_11082,N_11146);
or U11432 (N_11432,N_11039,N_11140);
nand U11433 (N_11433,N_11099,N_11030);
and U11434 (N_11434,N_11241,N_11194);
and U11435 (N_11435,N_11243,N_11077);
and U11436 (N_11436,N_11224,N_11129);
and U11437 (N_11437,N_11185,N_11239);
xor U11438 (N_11438,N_11186,N_11165);
and U11439 (N_11439,N_11030,N_11234);
or U11440 (N_11440,N_11004,N_11186);
nor U11441 (N_11441,N_11171,N_11110);
nor U11442 (N_11442,N_11115,N_11056);
nor U11443 (N_11443,N_11010,N_11209);
nand U11444 (N_11444,N_11055,N_11192);
nand U11445 (N_11445,N_11231,N_11063);
or U11446 (N_11446,N_11147,N_11172);
and U11447 (N_11447,N_11248,N_11237);
xnor U11448 (N_11448,N_11225,N_11019);
xor U11449 (N_11449,N_11249,N_11134);
nor U11450 (N_11450,N_11245,N_11060);
xnor U11451 (N_11451,N_11050,N_11155);
nor U11452 (N_11452,N_11190,N_11078);
and U11453 (N_11453,N_11162,N_11202);
or U11454 (N_11454,N_11217,N_11059);
or U11455 (N_11455,N_11089,N_11107);
nor U11456 (N_11456,N_11138,N_11247);
xnor U11457 (N_11457,N_11194,N_11228);
nor U11458 (N_11458,N_11136,N_11192);
xnor U11459 (N_11459,N_11095,N_11116);
and U11460 (N_11460,N_11167,N_11076);
and U11461 (N_11461,N_11061,N_11089);
or U11462 (N_11462,N_11202,N_11128);
xnor U11463 (N_11463,N_11206,N_11067);
and U11464 (N_11464,N_11181,N_11021);
xor U11465 (N_11465,N_11032,N_11216);
or U11466 (N_11466,N_11122,N_11195);
and U11467 (N_11467,N_11093,N_11064);
nand U11468 (N_11468,N_11107,N_11094);
nand U11469 (N_11469,N_11188,N_11107);
and U11470 (N_11470,N_11065,N_11202);
nor U11471 (N_11471,N_11035,N_11012);
nor U11472 (N_11472,N_11208,N_11136);
xnor U11473 (N_11473,N_11003,N_11208);
xor U11474 (N_11474,N_11176,N_11143);
xor U11475 (N_11475,N_11183,N_11205);
xnor U11476 (N_11476,N_11061,N_11165);
nor U11477 (N_11477,N_11119,N_11154);
nand U11478 (N_11478,N_11026,N_11202);
and U11479 (N_11479,N_11073,N_11199);
and U11480 (N_11480,N_11080,N_11238);
nand U11481 (N_11481,N_11054,N_11092);
nand U11482 (N_11482,N_11143,N_11179);
nand U11483 (N_11483,N_11196,N_11036);
nor U11484 (N_11484,N_11131,N_11106);
nand U11485 (N_11485,N_11197,N_11225);
and U11486 (N_11486,N_11087,N_11214);
or U11487 (N_11487,N_11000,N_11184);
xor U11488 (N_11488,N_11166,N_11000);
and U11489 (N_11489,N_11199,N_11182);
xnor U11490 (N_11490,N_11237,N_11202);
xnor U11491 (N_11491,N_11236,N_11243);
xor U11492 (N_11492,N_11165,N_11193);
nor U11493 (N_11493,N_11016,N_11033);
xnor U11494 (N_11494,N_11034,N_11239);
and U11495 (N_11495,N_11218,N_11130);
nand U11496 (N_11496,N_11008,N_11071);
nor U11497 (N_11497,N_11129,N_11011);
nand U11498 (N_11498,N_11040,N_11029);
or U11499 (N_11499,N_11106,N_11058);
xor U11500 (N_11500,N_11317,N_11277);
nor U11501 (N_11501,N_11489,N_11424);
xnor U11502 (N_11502,N_11404,N_11493);
or U11503 (N_11503,N_11367,N_11454);
nor U11504 (N_11504,N_11430,N_11423);
nand U11505 (N_11505,N_11322,N_11390);
xnor U11506 (N_11506,N_11415,N_11378);
and U11507 (N_11507,N_11302,N_11336);
nor U11508 (N_11508,N_11333,N_11250);
nand U11509 (N_11509,N_11288,N_11449);
or U11510 (N_11510,N_11309,N_11492);
and U11511 (N_11511,N_11431,N_11366);
xor U11512 (N_11512,N_11330,N_11439);
and U11513 (N_11513,N_11436,N_11371);
and U11514 (N_11514,N_11414,N_11381);
xor U11515 (N_11515,N_11346,N_11455);
xnor U11516 (N_11516,N_11282,N_11268);
nand U11517 (N_11517,N_11375,N_11458);
and U11518 (N_11518,N_11457,N_11286);
and U11519 (N_11519,N_11410,N_11486);
and U11520 (N_11520,N_11283,N_11276);
nor U11521 (N_11521,N_11442,N_11447);
nor U11522 (N_11522,N_11324,N_11318);
nor U11523 (N_11523,N_11327,N_11320);
and U11524 (N_11524,N_11360,N_11344);
and U11525 (N_11525,N_11352,N_11355);
nor U11526 (N_11526,N_11398,N_11391);
nor U11527 (N_11527,N_11498,N_11316);
or U11528 (N_11528,N_11497,N_11402);
nand U11529 (N_11529,N_11293,N_11401);
xor U11530 (N_11530,N_11496,N_11358);
nor U11531 (N_11531,N_11345,N_11262);
nor U11532 (N_11532,N_11359,N_11406);
nand U11533 (N_11533,N_11263,N_11350);
nand U11534 (N_11534,N_11343,N_11321);
nand U11535 (N_11535,N_11475,N_11453);
xor U11536 (N_11536,N_11467,N_11269);
xnor U11537 (N_11537,N_11452,N_11429);
or U11538 (N_11538,N_11433,N_11335);
nand U11539 (N_11539,N_11259,N_11490);
xor U11540 (N_11540,N_11388,N_11304);
and U11541 (N_11541,N_11369,N_11361);
nor U11542 (N_11542,N_11334,N_11471);
nand U11543 (N_11543,N_11434,N_11351);
or U11544 (N_11544,N_11370,N_11264);
or U11545 (N_11545,N_11267,N_11257);
and U11546 (N_11546,N_11379,N_11484);
and U11547 (N_11547,N_11465,N_11303);
nand U11548 (N_11548,N_11308,N_11311);
nor U11549 (N_11549,N_11272,N_11461);
xnor U11550 (N_11550,N_11403,N_11495);
or U11551 (N_11551,N_11323,N_11418);
nor U11552 (N_11552,N_11413,N_11435);
or U11553 (N_11553,N_11255,N_11385);
or U11554 (N_11554,N_11332,N_11412);
xnor U11555 (N_11555,N_11298,N_11450);
and U11556 (N_11556,N_11290,N_11329);
nor U11557 (N_11557,N_11340,N_11494);
nor U11558 (N_11558,N_11397,N_11279);
xor U11559 (N_11559,N_11278,N_11491);
nand U11560 (N_11560,N_11432,N_11382);
or U11561 (N_11561,N_11353,N_11380);
nor U11562 (N_11562,N_11384,N_11438);
nor U11563 (N_11563,N_11488,N_11376);
and U11564 (N_11564,N_11300,N_11407);
nor U11565 (N_11565,N_11427,N_11297);
nor U11566 (N_11566,N_11325,N_11287);
xor U11567 (N_11567,N_11472,N_11291);
nand U11568 (N_11568,N_11393,N_11373);
xnor U11569 (N_11569,N_11312,N_11301);
nor U11570 (N_11570,N_11314,N_11299);
nor U11571 (N_11571,N_11348,N_11273);
xor U11572 (N_11572,N_11374,N_11356);
nand U11573 (N_11573,N_11252,N_11387);
nor U11574 (N_11574,N_11459,N_11428);
or U11575 (N_11575,N_11307,N_11499);
nor U11576 (N_11576,N_11271,N_11411);
nor U11577 (N_11577,N_11482,N_11463);
nand U11578 (N_11578,N_11478,N_11261);
nand U11579 (N_11579,N_11394,N_11313);
xor U11580 (N_11580,N_11481,N_11477);
and U11581 (N_11581,N_11294,N_11365);
nor U11582 (N_11582,N_11275,N_11425);
nor U11583 (N_11583,N_11341,N_11400);
xor U11584 (N_11584,N_11437,N_11285);
and U11585 (N_11585,N_11260,N_11354);
xnor U11586 (N_11586,N_11405,N_11456);
nor U11587 (N_11587,N_11392,N_11395);
xor U11588 (N_11588,N_11469,N_11445);
nor U11589 (N_11589,N_11483,N_11295);
nor U11590 (N_11590,N_11451,N_11256);
and U11591 (N_11591,N_11470,N_11416);
nor U11592 (N_11592,N_11466,N_11296);
or U11593 (N_11593,N_11349,N_11364);
and U11594 (N_11594,N_11362,N_11383);
and U11595 (N_11595,N_11446,N_11426);
nor U11596 (N_11596,N_11389,N_11274);
nand U11597 (N_11597,N_11399,N_11468);
nor U11598 (N_11598,N_11266,N_11377);
nand U11599 (N_11599,N_11479,N_11292);
xor U11600 (N_11600,N_11289,N_11281);
or U11601 (N_11601,N_11422,N_11280);
nand U11602 (N_11602,N_11441,N_11396);
nand U11603 (N_11603,N_11409,N_11339);
xor U11604 (N_11604,N_11270,N_11310);
nor U11605 (N_11605,N_11328,N_11347);
nor U11606 (N_11606,N_11420,N_11342);
or U11607 (N_11607,N_11326,N_11305);
nor U11608 (N_11608,N_11474,N_11357);
nand U11609 (N_11609,N_11440,N_11315);
nor U11610 (N_11610,N_11444,N_11480);
nand U11611 (N_11611,N_11448,N_11421);
or U11612 (N_11612,N_11464,N_11460);
and U11613 (N_11613,N_11319,N_11443);
and U11614 (N_11614,N_11251,N_11368);
and U11615 (N_11615,N_11265,N_11485);
and U11616 (N_11616,N_11337,N_11417);
or U11617 (N_11617,N_11363,N_11473);
xnor U11618 (N_11618,N_11284,N_11306);
nand U11619 (N_11619,N_11408,N_11253);
nand U11620 (N_11620,N_11462,N_11258);
nor U11621 (N_11621,N_11372,N_11338);
and U11622 (N_11622,N_11331,N_11476);
xnor U11623 (N_11623,N_11254,N_11487);
and U11624 (N_11624,N_11386,N_11419);
nand U11625 (N_11625,N_11476,N_11347);
nand U11626 (N_11626,N_11294,N_11337);
xnor U11627 (N_11627,N_11319,N_11379);
nand U11628 (N_11628,N_11262,N_11466);
or U11629 (N_11629,N_11446,N_11256);
xnor U11630 (N_11630,N_11436,N_11467);
or U11631 (N_11631,N_11274,N_11306);
nor U11632 (N_11632,N_11335,N_11283);
xnor U11633 (N_11633,N_11338,N_11339);
or U11634 (N_11634,N_11360,N_11357);
nand U11635 (N_11635,N_11466,N_11388);
xnor U11636 (N_11636,N_11275,N_11350);
nor U11637 (N_11637,N_11277,N_11398);
and U11638 (N_11638,N_11344,N_11287);
or U11639 (N_11639,N_11337,N_11486);
or U11640 (N_11640,N_11373,N_11408);
nand U11641 (N_11641,N_11269,N_11432);
or U11642 (N_11642,N_11392,N_11406);
nand U11643 (N_11643,N_11377,N_11285);
nand U11644 (N_11644,N_11493,N_11495);
and U11645 (N_11645,N_11405,N_11382);
or U11646 (N_11646,N_11499,N_11273);
and U11647 (N_11647,N_11457,N_11353);
nand U11648 (N_11648,N_11250,N_11453);
xor U11649 (N_11649,N_11273,N_11378);
nor U11650 (N_11650,N_11412,N_11481);
and U11651 (N_11651,N_11378,N_11363);
and U11652 (N_11652,N_11477,N_11487);
or U11653 (N_11653,N_11274,N_11446);
and U11654 (N_11654,N_11454,N_11480);
and U11655 (N_11655,N_11282,N_11465);
nor U11656 (N_11656,N_11362,N_11381);
or U11657 (N_11657,N_11350,N_11449);
nor U11658 (N_11658,N_11481,N_11445);
and U11659 (N_11659,N_11352,N_11380);
and U11660 (N_11660,N_11455,N_11439);
nor U11661 (N_11661,N_11257,N_11345);
and U11662 (N_11662,N_11414,N_11370);
and U11663 (N_11663,N_11292,N_11280);
and U11664 (N_11664,N_11459,N_11468);
nand U11665 (N_11665,N_11394,N_11314);
nor U11666 (N_11666,N_11315,N_11464);
or U11667 (N_11667,N_11373,N_11470);
or U11668 (N_11668,N_11312,N_11342);
and U11669 (N_11669,N_11444,N_11262);
and U11670 (N_11670,N_11293,N_11367);
nand U11671 (N_11671,N_11259,N_11394);
or U11672 (N_11672,N_11330,N_11488);
nand U11673 (N_11673,N_11478,N_11464);
nor U11674 (N_11674,N_11281,N_11459);
nand U11675 (N_11675,N_11316,N_11344);
or U11676 (N_11676,N_11430,N_11299);
nand U11677 (N_11677,N_11308,N_11389);
or U11678 (N_11678,N_11362,N_11348);
nand U11679 (N_11679,N_11348,N_11488);
nor U11680 (N_11680,N_11322,N_11276);
and U11681 (N_11681,N_11484,N_11470);
nor U11682 (N_11682,N_11355,N_11341);
nor U11683 (N_11683,N_11490,N_11355);
and U11684 (N_11684,N_11449,N_11313);
nor U11685 (N_11685,N_11498,N_11415);
and U11686 (N_11686,N_11379,N_11282);
nor U11687 (N_11687,N_11330,N_11498);
and U11688 (N_11688,N_11438,N_11428);
nor U11689 (N_11689,N_11450,N_11300);
nand U11690 (N_11690,N_11386,N_11395);
nor U11691 (N_11691,N_11383,N_11265);
and U11692 (N_11692,N_11289,N_11393);
or U11693 (N_11693,N_11365,N_11396);
or U11694 (N_11694,N_11374,N_11436);
and U11695 (N_11695,N_11462,N_11374);
nor U11696 (N_11696,N_11308,N_11282);
and U11697 (N_11697,N_11305,N_11323);
and U11698 (N_11698,N_11437,N_11250);
or U11699 (N_11699,N_11361,N_11413);
xnor U11700 (N_11700,N_11495,N_11289);
or U11701 (N_11701,N_11295,N_11482);
xor U11702 (N_11702,N_11281,N_11395);
nor U11703 (N_11703,N_11451,N_11434);
xnor U11704 (N_11704,N_11407,N_11361);
nor U11705 (N_11705,N_11274,N_11295);
nand U11706 (N_11706,N_11336,N_11413);
xor U11707 (N_11707,N_11454,N_11312);
nand U11708 (N_11708,N_11363,N_11325);
xnor U11709 (N_11709,N_11330,N_11419);
nand U11710 (N_11710,N_11437,N_11436);
and U11711 (N_11711,N_11259,N_11318);
or U11712 (N_11712,N_11441,N_11407);
nor U11713 (N_11713,N_11417,N_11254);
and U11714 (N_11714,N_11486,N_11424);
nand U11715 (N_11715,N_11461,N_11333);
and U11716 (N_11716,N_11310,N_11482);
nor U11717 (N_11717,N_11412,N_11298);
and U11718 (N_11718,N_11305,N_11409);
nand U11719 (N_11719,N_11307,N_11290);
or U11720 (N_11720,N_11468,N_11275);
nand U11721 (N_11721,N_11364,N_11438);
and U11722 (N_11722,N_11311,N_11390);
or U11723 (N_11723,N_11253,N_11330);
nor U11724 (N_11724,N_11438,N_11369);
nor U11725 (N_11725,N_11487,N_11253);
xnor U11726 (N_11726,N_11328,N_11394);
nand U11727 (N_11727,N_11440,N_11415);
nand U11728 (N_11728,N_11331,N_11466);
nor U11729 (N_11729,N_11253,N_11335);
and U11730 (N_11730,N_11341,N_11405);
and U11731 (N_11731,N_11380,N_11441);
nor U11732 (N_11732,N_11290,N_11435);
and U11733 (N_11733,N_11328,N_11381);
nand U11734 (N_11734,N_11362,N_11269);
xor U11735 (N_11735,N_11258,N_11319);
or U11736 (N_11736,N_11449,N_11338);
and U11737 (N_11737,N_11447,N_11420);
and U11738 (N_11738,N_11320,N_11477);
or U11739 (N_11739,N_11252,N_11274);
or U11740 (N_11740,N_11348,N_11271);
and U11741 (N_11741,N_11283,N_11447);
and U11742 (N_11742,N_11320,N_11287);
nand U11743 (N_11743,N_11482,N_11251);
nand U11744 (N_11744,N_11474,N_11312);
and U11745 (N_11745,N_11412,N_11250);
nor U11746 (N_11746,N_11329,N_11497);
nor U11747 (N_11747,N_11290,N_11432);
xor U11748 (N_11748,N_11421,N_11274);
xor U11749 (N_11749,N_11494,N_11428);
or U11750 (N_11750,N_11641,N_11695);
and U11751 (N_11751,N_11712,N_11525);
nand U11752 (N_11752,N_11543,N_11574);
or U11753 (N_11753,N_11542,N_11572);
xnor U11754 (N_11754,N_11521,N_11639);
xnor U11755 (N_11755,N_11737,N_11689);
and U11756 (N_11756,N_11513,N_11708);
or U11757 (N_11757,N_11656,N_11597);
nor U11758 (N_11758,N_11558,N_11511);
nand U11759 (N_11759,N_11744,N_11575);
nand U11760 (N_11760,N_11600,N_11675);
or U11761 (N_11761,N_11523,N_11514);
nand U11762 (N_11762,N_11520,N_11577);
xnor U11763 (N_11763,N_11537,N_11637);
nand U11764 (N_11764,N_11563,N_11701);
or U11765 (N_11765,N_11539,N_11646);
nand U11766 (N_11766,N_11591,N_11562);
xnor U11767 (N_11767,N_11655,N_11593);
nor U11768 (N_11768,N_11732,N_11601);
nor U11769 (N_11769,N_11584,N_11748);
nand U11770 (N_11770,N_11681,N_11614);
or U11771 (N_11771,N_11590,N_11711);
and U11772 (N_11772,N_11571,N_11682);
nor U11773 (N_11773,N_11657,N_11532);
or U11774 (N_11774,N_11727,N_11619);
nor U11775 (N_11775,N_11587,N_11557);
and U11776 (N_11776,N_11680,N_11569);
nor U11777 (N_11777,N_11726,N_11650);
or U11778 (N_11778,N_11545,N_11503);
xnor U11779 (N_11779,N_11615,N_11533);
xor U11780 (N_11780,N_11653,N_11559);
xor U11781 (N_11781,N_11556,N_11583);
and U11782 (N_11782,N_11705,N_11747);
xnor U11783 (N_11783,N_11723,N_11683);
and U11784 (N_11784,N_11638,N_11731);
xnor U11785 (N_11785,N_11596,N_11631);
xor U11786 (N_11786,N_11738,N_11546);
nand U11787 (N_11787,N_11606,N_11500);
xnor U11788 (N_11788,N_11635,N_11709);
xnor U11789 (N_11789,N_11612,N_11707);
nand U11790 (N_11790,N_11714,N_11516);
nor U11791 (N_11791,N_11671,N_11629);
nor U11792 (N_11792,N_11550,N_11628);
nand U11793 (N_11793,N_11673,N_11551);
and U11794 (N_11794,N_11538,N_11534);
or U11795 (N_11795,N_11724,N_11634);
nand U11796 (N_11796,N_11718,N_11664);
nand U11797 (N_11797,N_11685,N_11688);
xor U11798 (N_11798,N_11652,N_11715);
xnor U11799 (N_11799,N_11733,N_11648);
or U11800 (N_11800,N_11734,N_11725);
and U11801 (N_11801,N_11651,N_11686);
nand U11802 (N_11802,N_11610,N_11622);
nand U11803 (N_11803,N_11547,N_11519);
xor U11804 (N_11804,N_11560,N_11706);
and U11805 (N_11805,N_11504,N_11522);
and U11806 (N_11806,N_11554,N_11549);
xor U11807 (N_11807,N_11676,N_11697);
or U11808 (N_11808,N_11735,N_11586);
and U11809 (N_11809,N_11721,N_11626);
nor U11810 (N_11810,N_11643,N_11555);
nand U11811 (N_11811,N_11698,N_11527);
and U11812 (N_11812,N_11728,N_11674);
or U11813 (N_11813,N_11588,N_11576);
and U11814 (N_11814,N_11508,N_11509);
and U11815 (N_11815,N_11578,N_11529);
and U11816 (N_11816,N_11564,N_11579);
and U11817 (N_11817,N_11605,N_11722);
nor U11818 (N_11818,N_11589,N_11618);
xnor U11819 (N_11819,N_11699,N_11608);
nand U11820 (N_11820,N_11568,N_11599);
nor U11821 (N_11821,N_11613,N_11602);
xor U11822 (N_11822,N_11541,N_11566);
nor U11823 (N_11823,N_11710,N_11505);
and U11824 (N_11824,N_11561,N_11630);
nor U11825 (N_11825,N_11647,N_11611);
nand U11826 (N_11826,N_11524,N_11745);
xnor U11827 (N_11827,N_11544,N_11703);
nand U11828 (N_11828,N_11592,N_11620);
and U11829 (N_11829,N_11694,N_11739);
or U11830 (N_11830,N_11716,N_11654);
and U11831 (N_11831,N_11510,N_11669);
nor U11832 (N_11832,N_11582,N_11530);
and U11833 (N_11833,N_11581,N_11603);
or U11834 (N_11834,N_11515,N_11616);
and U11835 (N_11835,N_11668,N_11649);
and U11836 (N_11836,N_11729,N_11518);
nor U11837 (N_11837,N_11502,N_11570);
nor U11838 (N_11838,N_11609,N_11506);
or U11839 (N_11839,N_11741,N_11666);
and U11840 (N_11840,N_11730,N_11742);
xnor U11841 (N_11841,N_11512,N_11736);
nor U11842 (N_11842,N_11667,N_11565);
nor U11843 (N_11843,N_11693,N_11644);
or U11844 (N_11844,N_11580,N_11632);
xnor U11845 (N_11845,N_11702,N_11692);
xor U11846 (N_11846,N_11624,N_11659);
and U11847 (N_11847,N_11604,N_11696);
and U11848 (N_11848,N_11684,N_11535);
xor U11849 (N_11849,N_11640,N_11670);
xor U11850 (N_11850,N_11528,N_11713);
and U11851 (N_11851,N_11690,N_11553);
nand U11852 (N_11852,N_11623,N_11540);
nor U11853 (N_11853,N_11749,N_11720);
or U11854 (N_11854,N_11660,N_11665);
xor U11855 (N_11855,N_11662,N_11598);
or U11856 (N_11856,N_11717,N_11617);
and U11857 (N_11857,N_11573,N_11526);
nand U11858 (N_11858,N_11531,N_11548);
nand U11859 (N_11859,N_11567,N_11743);
or U11860 (N_11860,N_11642,N_11663);
nor U11861 (N_11861,N_11700,N_11607);
and U11862 (N_11862,N_11552,N_11633);
nor U11863 (N_11863,N_11595,N_11658);
or U11864 (N_11864,N_11645,N_11672);
nand U11865 (N_11865,N_11704,N_11621);
or U11866 (N_11866,N_11691,N_11679);
and U11867 (N_11867,N_11594,N_11740);
nand U11868 (N_11868,N_11719,N_11625);
nand U11869 (N_11869,N_11501,N_11536);
xor U11870 (N_11870,N_11687,N_11746);
nor U11871 (N_11871,N_11507,N_11585);
nand U11872 (N_11872,N_11661,N_11677);
xor U11873 (N_11873,N_11636,N_11517);
nand U11874 (N_11874,N_11678,N_11627);
nand U11875 (N_11875,N_11558,N_11538);
and U11876 (N_11876,N_11745,N_11591);
nor U11877 (N_11877,N_11654,N_11628);
nand U11878 (N_11878,N_11689,N_11652);
or U11879 (N_11879,N_11540,N_11611);
nand U11880 (N_11880,N_11659,N_11581);
xor U11881 (N_11881,N_11598,N_11731);
or U11882 (N_11882,N_11573,N_11502);
and U11883 (N_11883,N_11570,N_11659);
or U11884 (N_11884,N_11658,N_11572);
nand U11885 (N_11885,N_11674,N_11718);
nor U11886 (N_11886,N_11742,N_11711);
nand U11887 (N_11887,N_11730,N_11644);
and U11888 (N_11888,N_11669,N_11683);
nand U11889 (N_11889,N_11606,N_11555);
nand U11890 (N_11890,N_11581,N_11573);
and U11891 (N_11891,N_11646,N_11662);
xor U11892 (N_11892,N_11527,N_11695);
nand U11893 (N_11893,N_11524,N_11556);
nor U11894 (N_11894,N_11712,N_11521);
or U11895 (N_11895,N_11703,N_11684);
xor U11896 (N_11896,N_11632,N_11619);
nor U11897 (N_11897,N_11662,N_11657);
and U11898 (N_11898,N_11662,N_11658);
xnor U11899 (N_11899,N_11559,N_11601);
nand U11900 (N_11900,N_11505,N_11708);
nand U11901 (N_11901,N_11681,N_11643);
and U11902 (N_11902,N_11506,N_11670);
and U11903 (N_11903,N_11689,N_11518);
or U11904 (N_11904,N_11710,N_11741);
nand U11905 (N_11905,N_11529,N_11745);
and U11906 (N_11906,N_11719,N_11640);
nand U11907 (N_11907,N_11731,N_11671);
or U11908 (N_11908,N_11616,N_11670);
nor U11909 (N_11909,N_11628,N_11622);
xnor U11910 (N_11910,N_11557,N_11678);
or U11911 (N_11911,N_11574,N_11634);
nand U11912 (N_11912,N_11513,N_11545);
and U11913 (N_11913,N_11702,N_11516);
and U11914 (N_11914,N_11701,N_11564);
xnor U11915 (N_11915,N_11632,N_11726);
nand U11916 (N_11916,N_11580,N_11642);
or U11917 (N_11917,N_11504,N_11627);
nand U11918 (N_11918,N_11634,N_11587);
nand U11919 (N_11919,N_11577,N_11501);
or U11920 (N_11920,N_11611,N_11616);
nor U11921 (N_11921,N_11546,N_11717);
xnor U11922 (N_11922,N_11500,N_11515);
nand U11923 (N_11923,N_11547,N_11692);
nand U11924 (N_11924,N_11617,N_11689);
and U11925 (N_11925,N_11568,N_11666);
xor U11926 (N_11926,N_11691,N_11553);
nor U11927 (N_11927,N_11532,N_11634);
xor U11928 (N_11928,N_11575,N_11707);
xnor U11929 (N_11929,N_11724,N_11727);
xor U11930 (N_11930,N_11584,N_11630);
and U11931 (N_11931,N_11548,N_11512);
nor U11932 (N_11932,N_11638,N_11552);
nor U11933 (N_11933,N_11676,N_11598);
or U11934 (N_11934,N_11519,N_11523);
nor U11935 (N_11935,N_11583,N_11680);
or U11936 (N_11936,N_11584,N_11560);
or U11937 (N_11937,N_11607,N_11685);
nor U11938 (N_11938,N_11675,N_11583);
and U11939 (N_11939,N_11741,N_11517);
and U11940 (N_11940,N_11677,N_11719);
or U11941 (N_11941,N_11668,N_11524);
nand U11942 (N_11942,N_11608,N_11738);
and U11943 (N_11943,N_11580,N_11685);
and U11944 (N_11944,N_11603,N_11633);
nor U11945 (N_11945,N_11527,N_11505);
nand U11946 (N_11946,N_11581,N_11545);
or U11947 (N_11947,N_11509,N_11514);
or U11948 (N_11948,N_11648,N_11634);
nor U11949 (N_11949,N_11551,N_11525);
or U11950 (N_11950,N_11732,N_11633);
nand U11951 (N_11951,N_11696,N_11598);
xor U11952 (N_11952,N_11645,N_11523);
nor U11953 (N_11953,N_11523,N_11579);
or U11954 (N_11954,N_11634,N_11729);
or U11955 (N_11955,N_11559,N_11718);
nor U11956 (N_11956,N_11704,N_11557);
nand U11957 (N_11957,N_11741,N_11501);
xnor U11958 (N_11958,N_11689,N_11557);
or U11959 (N_11959,N_11693,N_11709);
nand U11960 (N_11960,N_11527,N_11572);
and U11961 (N_11961,N_11573,N_11536);
and U11962 (N_11962,N_11510,N_11638);
nand U11963 (N_11963,N_11700,N_11578);
nor U11964 (N_11964,N_11609,N_11525);
xor U11965 (N_11965,N_11746,N_11608);
nand U11966 (N_11966,N_11699,N_11596);
nor U11967 (N_11967,N_11694,N_11552);
or U11968 (N_11968,N_11610,N_11512);
or U11969 (N_11969,N_11731,N_11739);
or U11970 (N_11970,N_11668,N_11582);
xnor U11971 (N_11971,N_11542,N_11707);
xor U11972 (N_11972,N_11656,N_11659);
nand U11973 (N_11973,N_11631,N_11730);
nor U11974 (N_11974,N_11588,N_11525);
nor U11975 (N_11975,N_11749,N_11607);
and U11976 (N_11976,N_11640,N_11724);
or U11977 (N_11977,N_11674,N_11526);
nor U11978 (N_11978,N_11655,N_11721);
and U11979 (N_11979,N_11628,N_11514);
nor U11980 (N_11980,N_11570,N_11722);
or U11981 (N_11981,N_11717,N_11715);
and U11982 (N_11982,N_11519,N_11521);
xor U11983 (N_11983,N_11634,N_11557);
or U11984 (N_11984,N_11721,N_11570);
or U11985 (N_11985,N_11686,N_11598);
xnor U11986 (N_11986,N_11671,N_11708);
and U11987 (N_11987,N_11548,N_11572);
xnor U11988 (N_11988,N_11654,N_11743);
or U11989 (N_11989,N_11573,N_11696);
nand U11990 (N_11990,N_11564,N_11569);
nor U11991 (N_11991,N_11732,N_11505);
nand U11992 (N_11992,N_11678,N_11734);
nand U11993 (N_11993,N_11628,N_11637);
xnor U11994 (N_11994,N_11694,N_11541);
xor U11995 (N_11995,N_11512,N_11629);
xor U11996 (N_11996,N_11544,N_11629);
nor U11997 (N_11997,N_11700,N_11635);
nand U11998 (N_11998,N_11594,N_11558);
nor U11999 (N_11999,N_11652,N_11534);
or U12000 (N_12000,N_11888,N_11886);
or U12001 (N_12001,N_11813,N_11810);
xor U12002 (N_12002,N_11840,N_11850);
nand U12003 (N_12003,N_11923,N_11773);
or U12004 (N_12004,N_11869,N_11814);
or U12005 (N_12005,N_11936,N_11829);
and U12006 (N_12006,N_11753,N_11825);
xor U12007 (N_12007,N_11974,N_11986);
and U12008 (N_12008,N_11946,N_11839);
and U12009 (N_12009,N_11890,N_11849);
or U12010 (N_12010,N_11953,N_11812);
xor U12011 (N_12011,N_11938,N_11957);
nand U12012 (N_12012,N_11898,N_11821);
nand U12013 (N_12013,N_11949,N_11868);
or U12014 (N_12014,N_11940,N_11921);
nor U12015 (N_12015,N_11916,N_11950);
and U12016 (N_12016,N_11899,N_11955);
nand U12017 (N_12017,N_11934,N_11928);
nor U12018 (N_12018,N_11914,N_11807);
nor U12019 (N_12019,N_11878,N_11942);
xor U12020 (N_12020,N_11769,N_11901);
and U12021 (N_12021,N_11980,N_11788);
nor U12022 (N_12022,N_11766,N_11960);
or U12023 (N_12023,N_11817,N_11779);
xnor U12024 (N_12024,N_11751,N_11771);
xor U12025 (N_12025,N_11776,N_11881);
nor U12026 (N_12026,N_11845,N_11802);
xnor U12027 (N_12027,N_11952,N_11828);
nand U12028 (N_12028,N_11913,N_11896);
or U12029 (N_12029,N_11801,N_11857);
nor U12030 (N_12030,N_11922,N_11978);
and U12031 (N_12031,N_11907,N_11885);
nand U12032 (N_12032,N_11789,N_11854);
nand U12033 (N_12033,N_11893,N_11969);
nor U12034 (N_12034,N_11924,N_11847);
nor U12035 (N_12035,N_11932,N_11783);
nor U12036 (N_12036,N_11872,N_11965);
xnor U12037 (N_12037,N_11754,N_11834);
and U12038 (N_12038,N_11761,N_11757);
nor U12039 (N_12039,N_11822,N_11894);
xnor U12040 (N_12040,N_11875,N_11989);
nor U12041 (N_12041,N_11785,N_11837);
nand U12042 (N_12042,N_11851,N_11909);
or U12043 (N_12043,N_11871,N_11879);
nand U12044 (N_12044,N_11844,N_11985);
nand U12045 (N_12045,N_11992,N_11824);
nor U12046 (N_12046,N_11859,N_11959);
xor U12047 (N_12047,N_11937,N_11767);
or U12048 (N_12048,N_11910,N_11818);
xor U12049 (N_12049,N_11904,N_11999);
nand U12050 (N_12050,N_11760,N_11911);
nand U12051 (N_12051,N_11993,N_11948);
xor U12052 (N_12052,N_11846,N_11780);
xnor U12053 (N_12053,N_11756,N_11892);
or U12054 (N_12054,N_11981,N_11983);
nor U12055 (N_12055,N_11873,N_11838);
nor U12056 (N_12056,N_11973,N_11797);
or U12057 (N_12057,N_11791,N_11963);
xor U12058 (N_12058,N_11935,N_11793);
xor U12059 (N_12059,N_11795,N_11770);
xor U12060 (N_12060,N_11887,N_11996);
and U12061 (N_12061,N_11800,N_11815);
nand U12062 (N_12062,N_11843,N_11891);
or U12063 (N_12063,N_11926,N_11778);
and U12064 (N_12064,N_11866,N_11918);
nand U12065 (N_12065,N_11929,N_11763);
nor U12066 (N_12066,N_11995,N_11962);
and U12067 (N_12067,N_11968,N_11865);
xor U12068 (N_12068,N_11841,N_11880);
nand U12069 (N_12069,N_11772,N_11804);
xnor U12070 (N_12070,N_11764,N_11750);
xor U12071 (N_12071,N_11930,N_11768);
nor U12072 (N_12072,N_11874,N_11933);
xnor U12073 (N_12073,N_11765,N_11755);
xnor U12074 (N_12074,N_11964,N_11997);
nand U12075 (N_12075,N_11855,N_11944);
xnor U12076 (N_12076,N_11848,N_11906);
xor U12077 (N_12077,N_11777,N_11842);
and U12078 (N_12078,N_11990,N_11792);
and U12079 (N_12079,N_11951,N_11794);
nand U12080 (N_12080,N_11803,N_11931);
and U12081 (N_12081,N_11823,N_11941);
and U12082 (N_12082,N_11862,N_11939);
nor U12083 (N_12083,N_11858,N_11860);
nor U12084 (N_12084,N_11808,N_11920);
nand U12085 (N_12085,N_11861,N_11994);
and U12086 (N_12086,N_11833,N_11897);
and U12087 (N_12087,N_11863,N_11805);
and U12088 (N_12088,N_11816,N_11979);
or U12089 (N_12089,N_11966,N_11835);
or U12090 (N_12090,N_11806,N_11947);
nor U12091 (N_12091,N_11927,N_11925);
or U12092 (N_12092,N_11961,N_11902);
and U12093 (N_12093,N_11852,N_11972);
and U12094 (N_12094,N_11889,N_11775);
or U12095 (N_12095,N_11877,N_11998);
and U12096 (N_12096,N_11919,N_11809);
nand U12097 (N_12097,N_11956,N_11988);
nand U12098 (N_12098,N_11908,N_11984);
xor U12099 (N_12099,N_11870,N_11900);
nor U12100 (N_12100,N_11883,N_11832);
xnor U12101 (N_12101,N_11752,N_11971);
nor U12102 (N_12102,N_11970,N_11798);
nor U12103 (N_12103,N_11912,N_11987);
or U12104 (N_12104,N_11782,N_11915);
or U12105 (N_12105,N_11905,N_11836);
or U12106 (N_12106,N_11867,N_11856);
or U12107 (N_12107,N_11786,N_11774);
nor U12108 (N_12108,N_11762,N_11758);
xor U12109 (N_12109,N_11876,N_11976);
nand U12110 (N_12110,N_11958,N_11954);
nand U12111 (N_12111,N_11945,N_11903);
or U12112 (N_12112,N_11967,N_11831);
xor U12113 (N_12113,N_11830,N_11977);
nor U12114 (N_12114,N_11790,N_11864);
and U12115 (N_12115,N_11943,N_11884);
nor U12116 (N_12116,N_11759,N_11895);
xnor U12117 (N_12117,N_11991,N_11799);
nand U12118 (N_12118,N_11787,N_11781);
or U12119 (N_12119,N_11975,N_11982);
nand U12120 (N_12120,N_11811,N_11827);
or U12121 (N_12121,N_11917,N_11819);
nor U12122 (N_12122,N_11796,N_11820);
or U12123 (N_12123,N_11826,N_11882);
or U12124 (N_12124,N_11853,N_11784);
or U12125 (N_12125,N_11868,N_11933);
nand U12126 (N_12126,N_11783,N_11926);
or U12127 (N_12127,N_11951,N_11827);
xnor U12128 (N_12128,N_11850,N_11937);
and U12129 (N_12129,N_11949,N_11978);
nand U12130 (N_12130,N_11785,N_11989);
nand U12131 (N_12131,N_11775,N_11777);
nor U12132 (N_12132,N_11773,N_11894);
or U12133 (N_12133,N_11931,N_11920);
nand U12134 (N_12134,N_11826,N_11926);
and U12135 (N_12135,N_11901,N_11850);
xor U12136 (N_12136,N_11848,N_11905);
nand U12137 (N_12137,N_11890,N_11835);
xnor U12138 (N_12138,N_11919,N_11881);
xor U12139 (N_12139,N_11949,N_11857);
xnor U12140 (N_12140,N_11841,N_11891);
and U12141 (N_12141,N_11822,N_11969);
nor U12142 (N_12142,N_11839,N_11781);
nor U12143 (N_12143,N_11817,N_11780);
and U12144 (N_12144,N_11978,N_11896);
xor U12145 (N_12145,N_11948,N_11801);
and U12146 (N_12146,N_11967,N_11950);
nand U12147 (N_12147,N_11973,N_11786);
and U12148 (N_12148,N_11916,N_11974);
xor U12149 (N_12149,N_11966,N_11827);
and U12150 (N_12150,N_11944,N_11958);
xnor U12151 (N_12151,N_11895,N_11987);
and U12152 (N_12152,N_11966,N_11871);
nor U12153 (N_12153,N_11815,N_11751);
and U12154 (N_12154,N_11948,N_11925);
xnor U12155 (N_12155,N_11980,N_11965);
nand U12156 (N_12156,N_11984,N_11898);
and U12157 (N_12157,N_11958,N_11933);
xor U12158 (N_12158,N_11946,N_11960);
or U12159 (N_12159,N_11775,N_11751);
xnor U12160 (N_12160,N_11764,N_11996);
xor U12161 (N_12161,N_11989,N_11814);
nand U12162 (N_12162,N_11756,N_11904);
or U12163 (N_12163,N_11998,N_11941);
xnor U12164 (N_12164,N_11914,N_11923);
nor U12165 (N_12165,N_11858,N_11772);
nor U12166 (N_12166,N_11799,N_11794);
xor U12167 (N_12167,N_11832,N_11978);
nor U12168 (N_12168,N_11854,N_11899);
nand U12169 (N_12169,N_11864,N_11857);
and U12170 (N_12170,N_11943,N_11947);
or U12171 (N_12171,N_11752,N_11923);
xnor U12172 (N_12172,N_11808,N_11790);
and U12173 (N_12173,N_11970,N_11967);
and U12174 (N_12174,N_11921,N_11983);
xnor U12175 (N_12175,N_11893,N_11758);
or U12176 (N_12176,N_11755,N_11781);
nor U12177 (N_12177,N_11945,N_11996);
nand U12178 (N_12178,N_11844,N_11891);
xnor U12179 (N_12179,N_11879,N_11977);
nand U12180 (N_12180,N_11885,N_11924);
nor U12181 (N_12181,N_11981,N_11858);
xor U12182 (N_12182,N_11808,N_11919);
nor U12183 (N_12183,N_11796,N_11948);
nand U12184 (N_12184,N_11883,N_11903);
nand U12185 (N_12185,N_11899,N_11945);
and U12186 (N_12186,N_11824,N_11881);
nand U12187 (N_12187,N_11754,N_11865);
nor U12188 (N_12188,N_11761,N_11910);
or U12189 (N_12189,N_11758,N_11976);
or U12190 (N_12190,N_11782,N_11814);
xor U12191 (N_12191,N_11805,N_11770);
nor U12192 (N_12192,N_11972,N_11771);
nor U12193 (N_12193,N_11986,N_11914);
and U12194 (N_12194,N_11977,N_11850);
nor U12195 (N_12195,N_11990,N_11779);
nand U12196 (N_12196,N_11940,N_11846);
nor U12197 (N_12197,N_11990,N_11890);
and U12198 (N_12198,N_11891,N_11830);
nor U12199 (N_12199,N_11939,N_11846);
xor U12200 (N_12200,N_11987,N_11955);
xnor U12201 (N_12201,N_11789,N_11972);
nor U12202 (N_12202,N_11862,N_11881);
nor U12203 (N_12203,N_11938,N_11840);
xnor U12204 (N_12204,N_11965,N_11865);
xor U12205 (N_12205,N_11899,N_11803);
or U12206 (N_12206,N_11855,N_11880);
nand U12207 (N_12207,N_11967,N_11900);
nor U12208 (N_12208,N_11761,N_11896);
or U12209 (N_12209,N_11968,N_11857);
nor U12210 (N_12210,N_11879,N_11818);
nor U12211 (N_12211,N_11866,N_11811);
or U12212 (N_12212,N_11932,N_11850);
or U12213 (N_12213,N_11813,N_11790);
nor U12214 (N_12214,N_11783,N_11809);
nor U12215 (N_12215,N_11927,N_11903);
xor U12216 (N_12216,N_11801,N_11918);
nand U12217 (N_12217,N_11959,N_11997);
nor U12218 (N_12218,N_11964,N_11810);
xnor U12219 (N_12219,N_11894,N_11858);
nand U12220 (N_12220,N_11999,N_11772);
or U12221 (N_12221,N_11912,N_11911);
nor U12222 (N_12222,N_11820,N_11750);
xor U12223 (N_12223,N_11847,N_11952);
or U12224 (N_12224,N_11998,N_11868);
nor U12225 (N_12225,N_11828,N_11842);
or U12226 (N_12226,N_11785,N_11846);
nor U12227 (N_12227,N_11909,N_11865);
nand U12228 (N_12228,N_11896,N_11915);
and U12229 (N_12229,N_11945,N_11832);
xor U12230 (N_12230,N_11852,N_11969);
or U12231 (N_12231,N_11861,N_11787);
nand U12232 (N_12232,N_11822,N_11907);
nor U12233 (N_12233,N_11931,N_11834);
and U12234 (N_12234,N_11975,N_11897);
and U12235 (N_12235,N_11901,N_11807);
nor U12236 (N_12236,N_11912,N_11797);
nand U12237 (N_12237,N_11918,N_11755);
xnor U12238 (N_12238,N_11833,N_11938);
nor U12239 (N_12239,N_11879,N_11807);
or U12240 (N_12240,N_11910,N_11881);
and U12241 (N_12241,N_11923,N_11820);
nand U12242 (N_12242,N_11943,N_11786);
or U12243 (N_12243,N_11975,N_11910);
and U12244 (N_12244,N_11921,N_11782);
and U12245 (N_12245,N_11828,N_11982);
and U12246 (N_12246,N_11909,N_11945);
nand U12247 (N_12247,N_11916,N_11961);
nor U12248 (N_12248,N_11942,N_11781);
nand U12249 (N_12249,N_11801,N_11763);
or U12250 (N_12250,N_12056,N_12019);
and U12251 (N_12251,N_12119,N_12145);
and U12252 (N_12252,N_12241,N_12203);
xor U12253 (N_12253,N_12064,N_12130);
or U12254 (N_12254,N_12006,N_12157);
xnor U12255 (N_12255,N_12178,N_12181);
xor U12256 (N_12256,N_12030,N_12108);
xor U12257 (N_12257,N_12089,N_12135);
and U12258 (N_12258,N_12243,N_12068);
and U12259 (N_12259,N_12153,N_12021);
and U12260 (N_12260,N_12212,N_12054);
xor U12261 (N_12261,N_12100,N_12106);
xor U12262 (N_12262,N_12042,N_12000);
or U12263 (N_12263,N_12236,N_12142);
or U12264 (N_12264,N_12229,N_12245);
or U12265 (N_12265,N_12041,N_12063);
or U12266 (N_12266,N_12171,N_12080);
nor U12267 (N_12267,N_12095,N_12082);
nor U12268 (N_12268,N_12028,N_12225);
or U12269 (N_12269,N_12066,N_12183);
nand U12270 (N_12270,N_12158,N_12046);
nand U12271 (N_12271,N_12079,N_12073);
and U12272 (N_12272,N_12016,N_12248);
nor U12273 (N_12273,N_12085,N_12115);
or U12274 (N_12274,N_12086,N_12008);
xnor U12275 (N_12275,N_12051,N_12031);
xor U12276 (N_12276,N_12122,N_12092);
xnor U12277 (N_12277,N_12215,N_12062);
nand U12278 (N_12278,N_12099,N_12103);
xor U12279 (N_12279,N_12206,N_12118);
and U12280 (N_12280,N_12034,N_12218);
or U12281 (N_12281,N_12093,N_12104);
xor U12282 (N_12282,N_12039,N_12144);
and U12283 (N_12283,N_12094,N_12173);
nor U12284 (N_12284,N_12110,N_12175);
nor U12285 (N_12285,N_12214,N_12221);
nand U12286 (N_12286,N_12163,N_12043);
or U12287 (N_12287,N_12155,N_12090);
xor U12288 (N_12288,N_12139,N_12211);
nand U12289 (N_12289,N_12184,N_12015);
or U12290 (N_12290,N_12022,N_12105);
nand U12291 (N_12291,N_12190,N_12151);
and U12292 (N_12292,N_12117,N_12060);
nor U12293 (N_12293,N_12045,N_12192);
or U12294 (N_12294,N_12189,N_12058);
nor U12295 (N_12295,N_12065,N_12111);
nand U12296 (N_12296,N_12087,N_12159);
or U12297 (N_12297,N_12088,N_12007);
and U12298 (N_12298,N_12123,N_12071);
nand U12299 (N_12299,N_12249,N_12098);
and U12300 (N_12300,N_12097,N_12053);
and U12301 (N_12301,N_12120,N_12003);
xnor U12302 (N_12302,N_12240,N_12113);
or U12303 (N_12303,N_12017,N_12109);
or U12304 (N_12304,N_12128,N_12027);
xor U12305 (N_12305,N_12172,N_12025);
or U12306 (N_12306,N_12004,N_12197);
or U12307 (N_12307,N_12233,N_12029);
nand U12308 (N_12308,N_12055,N_12036);
nand U12309 (N_12309,N_12074,N_12199);
nand U12310 (N_12310,N_12057,N_12083);
xnor U12311 (N_12311,N_12180,N_12010);
nor U12312 (N_12312,N_12001,N_12005);
and U12313 (N_12313,N_12148,N_12235);
nor U12314 (N_12314,N_12138,N_12129);
nor U12315 (N_12315,N_12012,N_12147);
nand U12316 (N_12316,N_12107,N_12076);
nand U12317 (N_12317,N_12136,N_12132);
or U12318 (N_12318,N_12152,N_12037);
xor U12319 (N_12319,N_12165,N_12164);
and U12320 (N_12320,N_12047,N_12137);
and U12321 (N_12321,N_12223,N_12131);
or U12322 (N_12322,N_12141,N_12072);
and U12323 (N_12323,N_12170,N_12193);
xor U12324 (N_12324,N_12166,N_12191);
nor U12325 (N_12325,N_12140,N_12040);
xor U12326 (N_12326,N_12023,N_12247);
nor U12327 (N_12327,N_12244,N_12146);
xnor U12328 (N_12328,N_12200,N_12112);
nor U12329 (N_12329,N_12239,N_12125);
or U12330 (N_12330,N_12126,N_12230);
nand U12331 (N_12331,N_12081,N_12150);
and U12332 (N_12332,N_12024,N_12185);
nand U12333 (N_12333,N_12224,N_12156);
nor U12334 (N_12334,N_12011,N_12014);
xor U12335 (N_12335,N_12127,N_12116);
xor U12336 (N_12336,N_12143,N_12188);
xnor U12337 (N_12337,N_12222,N_12205);
and U12338 (N_12338,N_12038,N_12219);
xor U12339 (N_12339,N_12167,N_12169);
nand U12340 (N_12340,N_12202,N_12009);
nand U12341 (N_12341,N_12162,N_12070);
nand U12342 (N_12342,N_12195,N_12231);
or U12343 (N_12343,N_12114,N_12196);
and U12344 (N_12344,N_12084,N_12101);
or U12345 (N_12345,N_12177,N_12020);
or U12346 (N_12346,N_12091,N_12044);
xor U12347 (N_12347,N_12059,N_12035);
nand U12348 (N_12348,N_12075,N_12204);
nand U12349 (N_12349,N_12124,N_12186);
or U12350 (N_12350,N_12174,N_12061);
nand U12351 (N_12351,N_12102,N_12133);
nor U12352 (N_12352,N_12237,N_12242);
or U12353 (N_12353,N_12050,N_12002);
nand U12354 (N_12354,N_12033,N_12052);
and U12355 (N_12355,N_12238,N_12096);
nand U12356 (N_12356,N_12210,N_12154);
xnor U12357 (N_12357,N_12067,N_12209);
or U12358 (N_12358,N_12121,N_12208);
nand U12359 (N_12359,N_12026,N_12201);
nand U12360 (N_12360,N_12187,N_12049);
nand U12361 (N_12361,N_12160,N_12179);
nor U12362 (N_12362,N_12198,N_12228);
nand U12363 (N_12363,N_12226,N_12234);
nand U12364 (N_12364,N_12246,N_12013);
or U12365 (N_12365,N_12216,N_12227);
and U12366 (N_12366,N_12176,N_12232);
nor U12367 (N_12367,N_12018,N_12048);
or U12368 (N_12368,N_12220,N_12069);
nand U12369 (N_12369,N_12161,N_12168);
or U12370 (N_12370,N_12217,N_12078);
nand U12371 (N_12371,N_12182,N_12213);
nor U12372 (N_12372,N_12194,N_12149);
nor U12373 (N_12373,N_12134,N_12077);
nand U12374 (N_12374,N_12207,N_12032);
nor U12375 (N_12375,N_12202,N_12124);
or U12376 (N_12376,N_12014,N_12100);
nand U12377 (N_12377,N_12163,N_12023);
xor U12378 (N_12378,N_12117,N_12174);
and U12379 (N_12379,N_12152,N_12171);
or U12380 (N_12380,N_12074,N_12075);
xnor U12381 (N_12381,N_12094,N_12089);
or U12382 (N_12382,N_12163,N_12231);
or U12383 (N_12383,N_12087,N_12044);
nor U12384 (N_12384,N_12067,N_12048);
nor U12385 (N_12385,N_12203,N_12179);
and U12386 (N_12386,N_12027,N_12078);
or U12387 (N_12387,N_12045,N_12189);
xnor U12388 (N_12388,N_12079,N_12193);
nor U12389 (N_12389,N_12075,N_12028);
xnor U12390 (N_12390,N_12147,N_12002);
nor U12391 (N_12391,N_12198,N_12027);
and U12392 (N_12392,N_12049,N_12124);
nand U12393 (N_12393,N_12040,N_12131);
and U12394 (N_12394,N_12009,N_12059);
and U12395 (N_12395,N_12231,N_12199);
or U12396 (N_12396,N_12224,N_12159);
nor U12397 (N_12397,N_12127,N_12099);
xor U12398 (N_12398,N_12129,N_12002);
nand U12399 (N_12399,N_12093,N_12157);
and U12400 (N_12400,N_12021,N_12076);
nor U12401 (N_12401,N_12142,N_12012);
nor U12402 (N_12402,N_12187,N_12160);
nor U12403 (N_12403,N_12019,N_12007);
nor U12404 (N_12404,N_12005,N_12078);
nand U12405 (N_12405,N_12077,N_12022);
nand U12406 (N_12406,N_12065,N_12042);
and U12407 (N_12407,N_12144,N_12220);
nor U12408 (N_12408,N_12102,N_12249);
and U12409 (N_12409,N_12106,N_12239);
or U12410 (N_12410,N_12024,N_12039);
nor U12411 (N_12411,N_12186,N_12057);
nand U12412 (N_12412,N_12112,N_12116);
nand U12413 (N_12413,N_12009,N_12037);
and U12414 (N_12414,N_12087,N_12207);
nand U12415 (N_12415,N_12014,N_12139);
or U12416 (N_12416,N_12130,N_12207);
or U12417 (N_12417,N_12221,N_12249);
and U12418 (N_12418,N_12092,N_12195);
nor U12419 (N_12419,N_12089,N_12041);
and U12420 (N_12420,N_12093,N_12020);
xnor U12421 (N_12421,N_12047,N_12082);
nand U12422 (N_12422,N_12206,N_12147);
and U12423 (N_12423,N_12168,N_12146);
and U12424 (N_12424,N_12198,N_12096);
nand U12425 (N_12425,N_12082,N_12146);
and U12426 (N_12426,N_12124,N_12153);
xor U12427 (N_12427,N_12051,N_12193);
or U12428 (N_12428,N_12047,N_12168);
nand U12429 (N_12429,N_12212,N_12238);
nor U12430 (N_12430,N_12236,N_12053);
nor U12431 (N_12431,N_12180,N_12194);
nand U12432 (N_12432,N_12047,N_12208);
nor U12433 (N_12433,N_12186,N_12203);
nor U12434 (N_12434,N_12136,N_12087);
and U12435 (N_12435,N_12041,N_12222);
and U12436 (N_12436,N_12166,N_12146);
or U12437 (N_12437,N_12163,N_12221);
xnor U12438 (N_12438,N_12018,N_12165);
nand U12439 (N_12439,N_12146,N_12135);
xor U12440 (N_12440,N_12144,N_12239);
and U12441 (N_12441,N_12053,N_12089);
nand U12442 (N_12442,N_12070,N_12111);
xor U12443 (N_12443,N_12058,N_12191);
nand U12444 (N_12444,N_12031,N_12071);
nor U12445 (N_12445,N_12245,N_12195);
nand U12446 (N_12446,N_12057,N_12107);
or U12447 (N_12447,N_12093,N_12002);
and U12448 (N_12448,N_12185,N_12210);
xnor U12449 (N_12449,N_12224,N_12214);
and U12450 (N_12450,N_12117,N_12146);
and U12451 (N_12451,N_12219,N_12151);
and U12452 (N_12452,N_12163,N_12166);
xnor U12453 (N_12453,N_12143,N_12150);
or U12454 (N_12454,N_12131,N_12202);
nor U12455 (N_12455,N_12239,N_12149);
nand U12456 (N_12456,N_12174,N_12203);
nand U12457 (N_12457,N_12232,N_12110);
nor U12458 (N_12458,N_12131,N_12068);
xor U12459 (N_12459,N_12124,N_12142);
xor U12460 (N_12460,N_12125,N_12074);
or U12461 (N_12461,N_12101,N_12096);
and U12462 (N_12462,N_12173,N_12021);
nand U12463 (N_12463,N_12169,N_12249);
or U12464 (N_12464,N_12120,N_12148);
nand U12465 (N_12465,N_12240,N_12102);
nor U12466 (N_12466,N_12249,N_12033);
nand U12467 (N_12467,N_12022,N_12024);
nand U12468 (N_12468,N_12075,N_12044);
xor U12469 (N_12469,N_12199,N_12125);
xor U12470 (N_12470,N_12237,N_12213);
or U12471 (N_12471,N_12049,N_12103);
and U12472 (N_12472,N_12016,N_12059);
nand U12473 (N_12473,N_12154,N_12170);
nand U12474 (N_12474,N_12139,N_12114);
or U12475 (N_12475,N_12191,N_12209);
nand U12476 (N_12476,N_12160,N_12104);
or U12477 (N_12477,N_12044,N_12104);
and U12478 (N_12478,N_12246,N_12177);
or U12479 (N_12479,N_12182,N_12180);
nand U12480 (N_12480,N_12109,N_12232);
nand U12481 (N_12481,N_12184,N_12199);
nand U12482 (N_12482,N_12200,N_12164);
xnor U12483 (N_12483,N_12057,N_12209);
xor U12484 (N_12484,N_12054,N_12066);
nor U12485 (N_12485,N_12075,N_12079);
or U12486 (N_12486,N_12022,N_12164);
nor U12487 (N_12487,N_12190,N_12096);
or U12488 (N_12488,N_12179,N_12018);
or U12489 (N_12489,N_12218,N_12181);
xor U12490 (N_12490,N_12168,N_12113);
and U12491 (N_12491,N_12079,N_12041);
xnor U12492 (N_12492,N_12036,N_12091);
xor U12493 (N_12493,N_12230,N_12072);
and U12494 (N_12494,N_12145,N_12125);
nand U12495 (N_12495,N_12198,N_12220);
or U12496 (N_12496,N_12203,N_12248);
xnor U12497 (N_12497,N_12088,N_12173);
and U12498 (N_12498,N_12212,N_12003);
nor U12499 (N_12499,N_12224,N_12136);
nor U12500 (N_12500,N_12302,N_12339);
or U12501 (N_12501,N_12385,N_12379);
xnor U12502 (N_12502,N_12348,N_12380);
xnor U12503 (N_12503,N_12257,N_12285);
and U12504 (N_12504,N_12481,N_12449);
and U12505 (N_12505,N_12414,N_12251);
or U12506 (N_12506,N_12398,N_12286);
and U12507 (N_12507,N_12358,N_12471);
and U12508 (N_12508,N_12483,N_12420);
or U12509 (N_12509,N_12296,N_12405);
nor U12510 (N_12510,N_12455,N_12493);
and U12511 (N_12511,N_12354,N_12349);
nor U12512 (N_12512,N_12320,N_12368);
xnor U12513 (N_12513,N_12280,N_12419);
nor U12514 (N_12514,N_12315,N_12317);
or U12515 (N_12515,N_12276,N_12431);
nor U12516 (N_12516,N_12273,N_12259);
xor U12517 (N_12517,N_12332,N_12258);
nor U12518 (N_12518,N_12347,N_12353);
xnor U12519 (N_12519,N_12433,N_12355);
nand U12520 (N_12520,N_12328,N_12340);
xor U12521 (N_12521,N_12497,N_12308);
xor U12522 (N_12522,N_12312,N_12452);
nand U12523 (N_12523,N_12334,N_12350);
or U12524 (N_12524,N_12445,N_12463);
and U12525 (N_12525,N_12459,N_12443);
xnor U12526 (N_12526,N_12313,N_12441);
or U12527 (N_12527,N_12279,N_12485);
or U12528 (N_12528,N_12451,N_12408);
and U12529 (N_12529,N_12428,N_12399);
and U12530 (N_12530,N_12266,N_12395);
or U12531 (N_12531,N_12322,N_12382);
nor U12532 (N_12532,N_12432,N_12298);
nor U12533 (N_12533,N_12396,N_12316);
or U12534 (N_12534,N_12498,N_12400);
xnor U12535 (N_12535,N_12287,N_12410);
nand U12536 (N_12536,N_12264,N_12477);
nand U12537 (N_12537,N_12299,N_12486);
nor U12538 (N_12538,N_12482,N_12422);
and U12539 (N_12539,N_12364,N_12326);
xnor U12540 (N_12540,N_12458,N_12331);
or U12541 (N_12541,N_12475,N_12479);
nand U12542 (N_12542,N_12288,N_12499);
or U12543 (N_12543,N_12278,N_12440);
or U12544 (N_12544,N_12284,N_12427);
or U12545 (N_12545,N_12492,N_12268);
or U12546 (N_12546,N_12387,N_12424);
and U12547 (N_12547,N_12423,N_12310);
nor U12548 (N_12548,N_12270,N_12436);
and U12549 (N_12549,N_12469,N_12415);
or U12550 (N_12550,N_12404,N_12437);
and U12551 (N_12551,N_12304,N_12359);
nand U12552 (N_12552,N_12417,N_12373);
nor U12553 (N_12553,N_12450,N_12457);
xor U12554 (N_12554,N_12335,N_12426);
or U12555 (N_12555,N_12438,N_12321);
and U12556 (N_12556,N_12374,N_12394);
and U12557 (N_12557,N_12429,N_12372);
nand U12558 (N_12558,N_12327,N_12383);
xnor U12559 (N_12559,N_12388,N_12378);
or U12560 (N_12560,N_12392,N_12289);
and U12561 (N_12561,N_12314,N_12352);
or U12562 (N_12562,N_12351,N_12384);
xnor U12563 (N_12563,N_12301,N_12411);
nor U12564 (N_12564,N_12323,N_12324);
nand U12565 (N_12565,N_12361,N_12442);
nor U12566 (N_12566,N_12435,N_12478);
nor U12567 (N_12567,N_12356,N_12283);
xnor U12568 (N_12568,N_12490,N_12267);
nor U12569 (N_12569,N_12467,N_12495);
or U12570 (N_12570,N_12447,N_12260);
xor U12571 (N_12571,N_12472,N_12446);
and U12572 (N_12572,N_12430,N_12305);
and U12573 (N_12573,N_12338,N_12494);
nor U12574 (N_12574,N_12377,N_12297);
or U12575 (N_12575,N_12330,N_12376);
xor U12576 (N_12576,N_12465,N_12360);
and U12577 (N_12577,N_12474,N_12253);
nor U12578 (N_12578,N_12397,N_12367);
and U12579 (N_12579,N_12274,N_12391);
or U12580 (N_12580,N_12318,N_12484);
xor U12581 (N_12581,N_12291,N_12263);
nand U12582 (N_12582,N_12293,N_12456);
or U12583 (N_12583,N_12434,N_12343);
and U12584 (N_12584,N_12386,N_12269);
nor U12585 (N_12585,N_12346,N_12487);
nor U12586 (N_12586,N_12290,N_12462);
and U12587 (N_12587,N_12295,N_12370);
or U12588 (N_12588,N_12333,N_12381);
xor U12589 (N_12589,N_12375,N_12262);
xor U12590 (N_12590,N_12275,N_12345);
and U12591 (N_12591,N_12403,N_12491);
nor U12592 (N_12592,N_12337,N_12336);
nor U12593 (N_12593,N_12294,N_12281);
xnor U12594 (N_12594,N_12282,N_12461);
nand U12595 (N_12595,N_12480,N_12476);
xor U12596 (N_12596,N_12329,N_12473);
xnor U12597 (N_12597,N_12371,N_12416);
and U12598 (N_12598,N_12453,N_12271);
and U12599 (N_12599,N_12300,N_12448);
or U12600 (N_12600,N_12489,N_12307);
or U12601 (N_12601,N_12466,N_12418);
nand U12602 (N_12602,N_12250,N_12393);
or U12603 (N_12603,N_12401,N_12464);
xor U12604 (N_12604,N_12256,N_12292);
or U12605 (N_12605,N_12309,N_12342);
nand U12606 (N_12606,N_12303,N_12254);
and U12607 (N_12607,N_12341,N_12454);
xnor U12608 (N_12608,N_12470,N_12306);
and U12609 (N_12609,N_12272,N_12468);
and U12610 (N_12610,N_12425,N_12407);
xnor U12611 (N_12611,N_12252,N_12311);
or U12612 (N_12612,N_12365,N_12344);
and U12613 (N_12613,N_12421,N_12261);
nand U12614 (N_12614,N_12488,N_12496);
xor U12615 (N_12615,N_12389,N_12412);
nor U12616 (N_12616,N_12362,N_12255);
xnor U12617 (N_12617,N_12439,N_12413);
or U12618 (N_12618,N_12265,N_12409);
nor U12619 (N_12619,N_12460,N_12277);
xor U12620 (N_12620,N_12319,N_12366);
xor U12621 (N_12621,N_12325,N_12363);
xnor U12622 (N_12622,N_12444,N_12369);
xnor U12623 (N_12623,N_12390,N_12357);
or U12624 (N_12624,N_12406,N_12402);
xor U12625 (N_12625,N_12404,N_12328);
or U12626 (N_12626,N_12335,N_12373);
nand U12627 (N_12627,N_12493,N_12414);
and U12628 (N_12628,N_12277,N_12274);
and U12629 (N_12629,N_12330,N_12464);
xnor U12630 (N_12630,N_12310,N_12318);
xnor U12631 (N_12631,N_12442,N_12335);
or U12632 (N_12632,N_12399,N_12469);
nor U12633 (N_12633,N_12258,N_12381);
nor U12634 (N_12634,N_12277,N_12309);
nor U12635 (N_12635,N_12278,N_12407);
nor U12636 (N_12636,N_12333,N_12456);
xnor U12637 (N_12637,N_12404,N_12308);
nand U12638 (N_12638,N_12376,N_12368);
nand U12639 (N_12639,N_12293,N_12271);
or U12640 (N_12640,N_12472,N_12304);
or U12641 (N_12641,N_12257,N_12302);
or U12642 (N_12642,N_12306,N_12389);
nor U12643 (N_12643,N_12338,N_12490);
xnor U12644 (N_12644,N_12395,N_12453);
xor U12645 (N_12645,N_12499,N_12400);
and U12646 (N_12646,N_12253,N_12469);
and U12647 (N_12647,N_12315,N_12345);
and U12648 (N_12648,N_12313,N_12292);
and U12649 (N_12649,N_12273,N_12287);
and U12650 (N_12650,N_12411,N_12404);
nor U12651 (N_12651,N_12402,N_12391);
nor U12652 (N_12652,N_12348,N_12342);
or U12653 (N_12653,N_12403,N_12484);
nand U12654 (N_12654,N_12319,N_12344);
and U12655 (N_12655,N_12426,N_12423);
xnor U12656 (N_12656,N_12367,N_12492);
or U12657 (N_12657,N_12429,N_12431);
xnor U12658 (N_12658,N_12408,N_12436);
and U12659 (N_12659,N_12323,N_12284);
or U12660 (N_12660,N_12315,N_12309);
nand U12661 (N_12661,N_12268,N_12457);
xnor U12662 (N_12662,N_12424,N_12279);
or U12663 (N_12663,N_12377,N_12369);
xnor U12664 (N_12664,N_12301,N_12252);
nand U12665 (N_12665,N_12267,N_12376);
nand U12666 (N_12666,N_12313,N_12465);
and U12667 (N_12667,N_12311,N_12283);
nor U12668 (N_12668,N_12265,N_12405);
or U12669 (N_12669,N_12409,N_12463);
and U12670 (N_12670,N_12417,N_12289);
or U12671 (N_12671,N_12480,N_12423);
nor U12672 (N_12672,N_12481,N_12332);
xor U12673 (N_12673,N_12257,N_12314);
nor U12674 (N_12674,N_12336,N_12457);
xnor U12675 (N_12675,N_12407,N_12329);
xor U12676 (N_12676,N_12486,N_12354);
xnor U12677 (N_12677,N_12473,N_12317);
and U12678 (N_12678,N_12481,N_12267);
nand U12679 (N_12679,N_12450,N_12267);
nor U12680 (N_12680,N_12276,N_12285);
xnor U12681 (N_12681,N_12287,N_12271);
or U12682 (N_12682,N_12394,N_12313);
or U12683 (N_12683,N_12267,N_12353);
xnor U12684 (N_12684,N_12439,N_12330);
or U12685 (N_12685,N_12416,N_12398);
xor U12686 (N_12686,N_12398,N_12423);
nand U12687 (N_12687,N_12476,N_12322);
and U12688 (N_12688,N_12360,N_12445);
or U12689 (N_12689,N_12479,N_12464);
nand U12690 (N_12690,N_12371,N_12413);
xnor U12691 (N_12691,N_12279,N_12261);
or U12692 (N_12692,N_12416,N_12280);
nand U12693 (N_12693,N_12414,N_12353);
nand U12694 (N_12694,N_12321,N_12320);
nor U12695 (N_12695,N_12402,N_12333);
xor U12696 (N_12696,N_12481,N_12329);
or U12697 (N_12697,N_12417,N_12410);
nand U12698 (N_12698,N_12259,N_12465);
nor U12699 (N_12699,N_12266,N_12347);
nand U12700 (N_12700,N_12275,N_12388);
nand U12701 (N_12701,N_12286,N_12320);
nor U12702 (N_12702,N_12431,N_12414);
nor U12703 (N_12703,N_12459,N_12409);
or U12704 (N_12704,N_12321,N_12476);
nand U12705 (N_12705,N_12272,N_12347);
nor U12706 (N_12706,N_12320,N_12494);
nor U12707 (N_12707,N_12481,N_12496);
xnor U12708 (N_12708,N_12263,N_12280);
nor U12709 (N_12709,N_12342,N_12268);
and U12710 (N_12710,N_12378,N_12264);
nand U12711 (N_12711,N_12412,N_12349);
or U12712 (N_12712,N_12277,N_12444);
xor U12713 (N_12713,N_12492,N_12373);
or U12714 (N_12714,N_12497,N_12338);
nand U12715 (N_12715,N_12269,N_12476);
xor U12716 (N_12716,N_12280,N_12405);
nor U12717 (N_12717,N_12476,N_12288);
or U12718 (N_12718,N_12270,N_12378);
and U12719 (N_12719,N_12470,N_12414);
xor U12720 (N_12720,N_12494,N_12478);
or U12721 (N_12721,N_12449,N_12337);
or U12722 (N_12722,N_12292,N_12261);
xor U12723 (N_12723,N_12366,N_12312);
and U12724 (N_12724,N_12253,N_12313);
nand U12725 (N_12725,N_12491,N_12298);
nand U12726 (N_12726,N_12274,N_12359);
xor U12727 (N_12727,N_12308,N_12492);
nand U12728 (N_12728,N_12363,N_12498);
nor U12729 (N_12729,N_12365,N_12332);
xor U12730 (N_12730,N_12317,N_12451);
nor U12731 (N_12731,N_12492,N_12385);
nand U12732 (N_12732,N_12306,N_12384);
or U12733 (N_12733,N_12257,N_12359);
or U12734 (N_12734,N_12343,N_12254);
or U12735 (N_12735,N_12370,N_12433);
nor U12736 (N_12736,N_12440,N_12432);
nor U12737 (N_12737,N_12350,N_12283);
nor U12738 (N_12738,N_12431,N_12298);
and U12739 (N_12739,N_12360,N_12437);
xor U12740 (N_12740,N_12374,N_12450);
and U12741 (N_12741,N_12429,N_12438);
nor U12742 (N_12742,N_12431,N_12422);
nand U12743 (N_12743,N_12260,N_12359);
nand U12744 (N_12744,N_12308,N_12344);
nand U12745 (N_12745,N_12264,N_12254);
or U12746 (N_12746,N_12481,N_12289);
xor U12747 (N_12747,N_12472,N_12349);
xnor U12748 (N_12748,N_12437,N_12367);
and U12749 (N_12749,N_12463,N_12461);
or U12750 (N_12750,N_12692,N_12562);
nand U12751 (N_12751,N_12690,N_12716);
xor U12752 (N_12752,N_12681,N_12542);
xor U12753 (N_12753,N_12703,N_12616);
xnor U12754 (N_12754,N_12666,N_12515);
or U12755 (N_12755,N_12531,N_12675);
xor U12756 (N_12756,N_12748,N_12576);
xnor U12757 (N_12757,N_12551,N_12604);
and U12758 (N_12758,N_12505,N_12737);
and U12759 (N_12759,N_12525,N_12660);
or U12760 (N_12760,N_12655,N_12521);
and U12761 (N_12761,N_12652,N_12570);
and U12762 (N_12762,N_12644,N_12746);
nor U12763 (N_12763,N_12718,N_12583);
or U12764 (N_12764,N_12595,N_12640);
nor U12765 (N_12765,N_12739,N_12621);
or U12766 (N_12766,N_12671,N_12512);
nand U12767 (N_12767,N_12687,N_12665);
or U12768 (N_12768,N_12609,N_12518);
nand U12769 (N_12769,N_12627,N_12566);
nor U12770 (N_12770,N_12734,N_12573);
or U12771 (N_12771,N_12552,N_12610);
or U12772 (N_12772,N_12569,N_12749);
xor U12773 (N_12773,N_12568,N_12704);
nor U12774 (N_12774,N_12538,N_12741);
and U12775 (N_12775,N_12637,N_12585);
and U12776 (N_12776,N_12500,N_12557);
nor U12777 (N_12777,N_12633,N_12678);
or U12778 (N_12778,N_12672,N_12722);
and U12779 (N_12779,N_12727,N_12636);
or U12780 (N_12780,N_12527,N_12624);
or U12781 (N_12781,N_12558,N_12594);
xnor U12782 (N_12782,N_12601,N_12508);
and U12783 (N_12783,N_12723,N_12528);
nand U12784 (N_12784,N_12625,N_12642);
nand U12785 (N_12785,N_12641,N_12700);
or U12786 (N_12786,N_12548,N_12685);
nand U12787 (N_12787,N_12539,N_12617);
xnor U12788 (N_12788,N_12667,N_12683);
and U12789 (N_12789,N_12541,N_12688);
nor U12790 (N_12790,N_12743,N_12731);
xor U12791 (N_12791,N_12684,N_12717);
nand U12792 (N_12792,N_12674,N_12584);
nand U12793 (N_12793,N_12579,N_12649);
xor U12794 (N_12794,N_12648,N_12673);
and U12795 (N_12795,N_12608,N_12619);
and U12796 (N_12796,N_12588,N_12645);
nor U12797 (N_12797,N_12698,N_12517);
nand U12798 (N_12798,N_12546,N_12598);
or U12799 (N_12799,N_12707,N_12524);
nand U12800 (N_12800,N_12606,N_12695);
and U12801 (N_12801,N_12599,N_12689);
xnor U12802 (N_12802,N_12693,N_12547);
nor U12803 (N_12803,N_12618,N_12607);
nor U12804 (N_12804,N_12520,N_12581);
nand U12805 (N_12805,N_12677,N_12503);
nor U12806 (N_12806,N_12733,N_12522);
nor U12807 (N_12807,N_12535,N_12744);
and U12808 (N_12808,N_12589,N_12549);
nand U12809 (N_12809,N_12669,N_12555);
and U12810 (N_12810,N_12519,N_12600);
and U12811 (N_12811,N_12691,N_12738);
and U12812 (N_12812,N_12715,N_12597);
or U12813 (N_12813,N_12514,N_12736);
and U12814 (N_12814,N_12676,N_12565);
nor U12815 (N_12815,N_12501,N_12602);
nor U12816 (N_12816,N_12511,N_12507);
nor U12817 (N_12817,N_12593,N_12613);
nor U12818 (N_12818,N_12638,N_12592);
or U12819 (N_12819,N_12596,N_12590);
xor U12820 (N_12820,N_12543,N_12575);
nor U12821 (N_12821,N_12702,N_12571);
nor U12822 (N_12822,N_12726,N_12635);
or U12823 (N_12823,N_12556,N_12620);
or U12824 (N_12824,N_12587,N_12670);
nand U12825 (N_12825,N_12559,N_12577);
nor U12826 (N_12826,N_12537,N_12574);
and U12827 (N_12827,N_12605,N_12651);
nand U12828 (N_12828,N_12664,N_12696);
and U12829 (N_12829,N_12647,N_12626);
xnor U12830 (N_12830,N_12632,N_12639);
xor U12831 (N_12831,N_12612,N_12536);
xnor U12832 (N_12832,N_12740,N_12561);
xnor U12833 (N_12833,N_12530,N_12586);
or U12834 (N_12834,N_12709,N_12630);
nor U12835 (N_12835,N_12694,N_12614);
nor U12836 (N_12836,N_12653,N_12725);
or U12837 (N_12837,N_12567,N_12719);
nor U12838 (N_12838,N_12701,N_12591);
and U12839 (N_12839,N_12680,N_12705);
xor U12840 (N_12840,N_12628,N_12682);
nor U12841 (N_12841,N_12611,N_12720);
and U12842 (N_12842,N_12578,N_12603);
and U12843 (N_12843,N_12550,N_12710);
nand U12844 (N_12844,N_12659,N_12513);
or U12845 (N_12845,N_12582,N_12545);
and U12846 (N_12846,N_12686,N_12742);
and U12847 (N_12847,N_12526,N_12563);
or U12848 (N_12848,N_12544,N_12747);
nor U12849 (N_12849,N_12504,N_12745);
and U12850 (N_12850,N_12650,N_12510);
nor U12851 (N_12851,N_12631,N_12706);
xor U12852 (N_12852,N_12564,N_12656);
and U12853 (N_12853,N_12623,N_12712);
and U12854 (N_12854,N_12735,N_12711);
or U12855 (N_12855,N_12533,N_12529);
or U12856 (N_12856,N_12572,N_12657);
or U12857 (N_12857,N_12532,N_12729);
xnor U12858 (N_12858,N_12540,N_12732);
nor U12859 (N_12859,N_12654,N_12509);
or U12860 (N_12860,N_12534,N_12730);
nand U12861 (N_12861,N_12714,N_12629);
xnor U12862 (N_12862,N_12615,N_12697);
xnor U12863 (N_12863,N_12516,N_12663);
nor U12864 (N_12864,N_12502,N_12708);
or U12865 (N_12865,N_12721,N_12580);
or U12866 (N_12866,N_12661,N_12713);
and U12867 (N_12867,N_12728,N_12523);
and U12868 (N_12868,N_12699,N_12662);
xnor U12869 (N_12869,N_12646,N_12668);
xor U12870 (N_12870,N_12643,N_12622);
nor U12871 (N_12871,N_12553,N_12679);
nor U12872 (N_12872,N_12724,N_12634);
xor U12873 (N_12873,N_12554,N_12506);
xor U12874 (N_12874,N_12658,N_12560);
or U12875 (N_12875,N_12696,N_12585);
or U12876 (N_12876,N_12622,N_12630);
and U12877 (N_12877,N_12675,N_12710);
nand U12878 (N_12878,N_12665,N_12703);
or U12879 (N_12879,N_12539,N_12658);
and U12880 (N_12880,N_12653,N_12625);
or U12881 (N_12881,N_12710,N_12544);
nand U12882 (N_12882,N_12719,N_12727);
nand U12883 (N_12883,N_12627,N_12510);
nor U12884 (N_12884,N_12509,N_12634);
xor U12885 (N_12885,N_12555,N_12550);
and U12886 (N_12886,N_12516,N_12575);
nand U12887 (N_12887,N_12644,N_12721);
nor U12888 (N_12888,N_12645,N_12683);
or U12889 (N_12889,N_12602,N_12507);
and U12890 (N_12890,N_12515,N_12662);
or U12891 (N_12891,N_12522,N_12598);
or U12892 (N_12892,N_12631,N_12548);
nand U12893 (N_12893,N_12649,N_12520);
nor U12894 (N_12894,N_12622,N_12614);
or U12895 (N_12895,N_12698,N_12682);
xnor U12896 (N_12896,N_12696,N_12528);
and U12897 (N_12897,N_12572,N_12721);
and U12898 (N_12898,N_12693,N_12521);
nor U12899 (N_12899,N_12509,N_12628);
nor U12900 (N_12900,N_12654,N_12534);
xnor U12901 (N_12901,N_12616,N_12558);
xor U12902 (N_12902,N_12579,N_12694);
xor U12903 (N_12903,N_12743,N_12668);
nor U12904 (N_12904,N_12707,N_12552);
nand U12905 (N_12905,N_12722,N_12594);
nand U12906 (N_12906,N_12582,N_12504);
and U12907 (N_12907,N_12690,N_12661);
nand U12908 (N_12908,N_12558,N_12593);
or U12909 (N_12909,N_12627,N_12539);
xnor U12910 (N_12910,N_12554,N_12590);
xnor U12911 (N_12911,N_12690,N_12624);
xor U12912 (N_12912,N_12553,N_12742);
or U12913 (N_12913,N_12543,N_12733);
nor U12914 (N_12914,N_12638,N_12539);
and U12915 (N_12915,N_12655,N_12548);
xnor U12916 (N_12916,N_12557,N_12624);
xor U12917 (N_12917,N_12546,N_12610);
nor U12918 (N_12918,N_12630,N_12518);
nor U12919 (N_12919,N_12719,N_12626);
or U12920 (N_12920,N_12504,N_12680);
or U12921 (N_12921,N_12624,N_12741);
and U12922 (N_12922,N_12599,N_12605);
xor U12923 (N_12923,N_12528,N_12535);
nor U12924 (N_12924,N_12554,N_12743);
nand U12925 (N_12925,N_12659,N_12506);
or U12926 (N_12926,N_12600,N_12636);
or U12927 (N_12927,N_12598,N_12569);
nand U12928 (N_12928,N_12746,N_12672);
or U12929 (N_12929,N_12721,N_12570);
nor U12930 (N_12930,N_12501,N_12634);
and U12931 (N_12931,N_12639,N_12538);
xnor U12932 (N_12932,N_12520,N_12604);
nor U12933 (N_12933,N_12671,N_12647);
nand U12934 (N_12934,N_12627,N_12669);
nand U12935 (N_12935,N_12586,N_12552);
and U12936 (N_12936,N_12658,N_12592);
xnor U12937 (N_12937,N_12664,N_12644);
and U12938 (N_12938,N_12502,N_12696);
nand U12939 (N_12939,N_12640,N_12662);
nand U12940 (N_12940,N_12628,N_12716);
or U12941 (N_12941,N_12716,N_12501);
and U12942 (N_12942,N_12583,N_12697);
or U12943 (N_12943,N_12547,N_12698);
xor U12944 (N_12944,N_12563,N_12737);
and U12945 (N_12945,N_12555,N_12530);
or U12946 (N_12946,N_12537,N_12524);
and U12947 (N_12947,N_12553,N_12663);
and U12948 (N_12948,N_12514,N_12662);
nor U12949 (N_12949,N_12611,N_12672);
and U12950 (N_12950,N_12681,N_12590);
nand U12951 (N_12951,N_12545,N_12670);
xnor U12952 (N_12952,N_12721,N_12522);
and U12953 (N_12953,N_12686,N_12584);
or U12954 (N_12954,N_12578,N_12637);
and U12955 (N_12955,N_12711,N_12597);
nor U12956 (N_12956,N_12655,N_12526);
or U12957 (N_12957,N_12545,N_12673);
xnor U12958 (N_12958,N_12623,N_12692);
nor U12959 (N_12959,N_12556,N_12573);
or U12960 (N_12960,N_12734,N_12510);
nor U12961 (N_12961,N_12559,N_12638);
xnor U12962 (N_12962,N_12627,N_12561);
and U12963 (N_12963,N_12617,N_12743);
or U12964 (N_12964,N_12515,N_12697);
xor U12965 (N_12965,N_12573,N_12676);
nand U12966 (N_12966,N_12552,N_12574);
nor U12967 (N_12967,N_12677,N_12716);
and U12968 (N_12968,N_12660,N_12670);
and U12969 (N_12969,N_12531,N_12545);
xor U12970 (N_12970,N_12596,N_12568);
nand U12971 (N_12971,N_12736,N_12641);
nand U12972 (N_12972,N_12514,N_12576);
nor U12973 (N_12973,N_12645,N_12613);
and U12974 (N_12974,N_12539,N_12669);
and U12975 (N_12975,N_12550,N_12577);
and U12976 (N_12976,N_12606,N_12623);
or U12977 (N_12977,N_12685,N_12739);
and U12978 (N_12978,N_12505,N_12544);
nand U12979 (N_12979,N_12563,N_12674);
xor U12980 (N_12980,N_12548,N_12593);
nand U12981 (N_12981,N_12665,N_12642);
and U12982 (N_12982,N_12607,N_12714);
or U12983 (N_12983,N_12537,N_12618);
xor U12984 (N_12984,N_12534,N_12713);
or U12985 (N_12985,N_12616,N_12528);
nand U12986 (N_12986,N_12602,N_12541);
or U12987 (N_12987,N_12672,N_12623);
xor U12988 (N_12988,N_12747,N_12727);
nor U12989 (N_12989,N_12521,N_12697);
or U12990 (N_12990,N_12546,N_12558);
nand U12991 (N_12991,N_12598,N_12722);
and U12992 (N_12992,N_12531,N_12601);
nor U12993 (N_12993,N_12683,N_12573);
nor U12994 (N_12994,N_12532,N_12636);
or U12995 (N_12995,N_12654,N_12555);
and U12996 (N_12996,N_12526,N_12524);
and U12997 (N_12997,N_12719,N_12588);
nor U12998 (N_12998,N_12721,N_12515);
or U12999 (N_12999,N_12522,N_12535);
xor U13000 (N_13000,N_12808,N_12832);
nand U13001 (N_13001,N_12884,N_12870);
nor U13002 (N_13002,N_12776,N_12789);
nand U13003 (N_13003,N_12887,N_12754);
xor U13004 (N_13004,N_12911,N_12795);
and U13005 (N_13005,N_12907,N_12914);
nor U13006 (N_13006,N_12793,N_12852);
nor U13007 (N_13007,N_12949,N_12984);
xor U13008 (N_13008,N_12751,N_12962);
nand U13009 (N_13009,N_12883,N_12916);
or U13010 (N_13010,N_12845,N_12903);
or U13011 (N_13011,N_12902,N_12941);
or U13012 (N_13012,N_12975,N_12805);
or U13013 (N_13013,N_12928,N_12792);
or U13014 (N_13014,N_12950,N_12995);
or U13015 (N_13015,N_12920,N_12945);
or U13016 (N_13016,N_12953,N_12858);
nand U13017 (N_13017,N_12806,N_12872);
and U13018 (N_13018,N_12861,N_12804);
and U13019 (N_13019,N_12900,N_12819);
or U13020 (N_13020,N_12823,N_12769);
and U13021 (N_13021,N_12809,N_12818);
and U13022 (N_13022,N_12882,N_12763);
and U13023 (N_13023,N_12951,N_12948);
nor U13024 (N_13024,N_12915,N_12932);
nand U13025 (N_13025,N_12865,N_12770);
nand U13026 (N_13026,N_12943,N_12844);
xor U13027 (N_13027,N_12968,N_12997);
xor U13028 (N_13028,N_12912,N_12874);
or U13029 (N_13029,N_12802,N_12825);
and U13030 (N_13030,N_12843,N_12952);
nand U13031 (N_13031,N_12781,N_12775);
xnor U13032 (N_13032,N_12862,N_12933);
nand U13033 (N_13033,N_12764,N_12773);
xnor U13034 (N_13034,N_12859,N_12752);
xor U13035 (N_13035,N_12803,N_12979);
or U13036 (N_13036,N_12813,N_12886);
or U13037 (N_13037,N_12836,N_12982);
or U13038 (N_13038,N_12904,N_12753);
xnor U13039 (N_13039,N_12972,N_12991);
nand U13040 (N_13040,N_12855,N_12937);
nand U13041 (N_13041,N_12787,N_12992);
nand U13042 (N_13042,N_12924,N_12959);
nor U13043 (N_13043,N_12847,N_12799);
or U13044 (N_13044,N_12934,N_12956);
nor U13045 (N_13045,N_12822,N_12983);
and U13046 (N_13046,N_12910,N_12864);
and U13047 (N_13047,N_12891,N_12827);
and U13048 (N_13048,N_12878,N_12810);
and U13049 (N_13049,N_12797,N_12899);
xnor U13050 (N_13050,N_12867,N_12919);
xor U13051 (N_13051,N_12758,N_12767);
and U13052 (N_13052,N_12977,N_12963);
nor U13053 (N_13053,N_12927,N_12851);
and U13054 (N_13054,N_12888,N_12971);
nand U13055 (N_13055,N_12930,N_12926);
or U13056 (N_13056,N_12811,N_12925);
xnor U13057 (N_13057,N_12976,N_12957);
and U13058 (N_13058,N_12909,N_12942);
or U13059 (N_13059,N_12893,N_12794);
xor U13060 (N_13060,N_12829,N_12966);
and U13061 (N_13061,N_12774,N_12828);
nor U13062 (N_13062,N_12881,N_12820);
nor U13063 (N_13063,N_12771,N_12834);
xnor U13064 (N_13064,N_12961,N_12783);
and U13065 (N_13065,N_12964,N_12885);
xor U13066 (N_13066,N_12777,N_12922);
and U13067 (N_13067,N_12929,N_12816);
nor U13068 (N_13068,N_12880,N_12955);
nand U13069 (N_13069,N_12866,N_12760);
and U13070 (N_13070,N_12894,N_12850);
nor U13071 (N_13071,N_12821,N_12798);
or U13072 (N_13072,N_12938,N_12940);
xor U13073 (N_13073,N_12838,N_12897);
nand U13074 (N_13074,N_12766,N_12840);
nor U13075 (N_13075,N_12833,N_12762);
nor U13076 (N_13076,N_12796,N_12863);
nand U13077 (N_13077,N_12994,N_12784);
nand U13078 (N_13078,N_12875,N_12842);
nor U13079 (N_13079,N_12755,N_12987);
or U13080 (N_13080,N_12785,N_12998);
and U13081 (N_13081,N_12935,N_12898);
nor U13082 (N_13082,N_12826,N_12757);
xor U13083 (N_13083,N_12978,N_12879);
nand U13084 (N_13084,N_12849,N_12780);
nor U13085 (N_13085,N_12947,N_12814);
and U13086 (N_13086,N_12989,N_12750);
nand U13087 (N_13087,N_12901,N_12846);
and U13088 (N_13088,N_12986,N_12981);
or U13089 (N_13089,N_12958,N_12812);
nand U13090 (N_13090,N_12969,N_12890);
nor U13091 (N_13091,N_12918,N_12939);
nand U13092 (N_13092,N_12860,N_12815);
nand U13093 (N_13093,N_12954,N_12848);
nor U13094 (N_13094,N_12768,N_12807);
and U13095 (N_13095,N_12782,N_12923);
nor U13096 (N_13096,N_12996,N_12801);
and U13097 (N_13097,N_12817,N_12868);
xor U13098 (N_13098,N_12869,N_12973);
or U13099 (N_13099,N_12856,N_12970);
xnor U13100 (N_13100,N_12936,N_12965);
and U13101 (N_13101,N_12837,N_12908);
xor U13102 (N_13102,N_12974,N_12854);
nand U13103 (N_13103,N_12857,N_12960);
or U13104 (N_13104,N_12985,N_12830);
or U13105 (N_13105,N_12788,N_12779);
nand U13106 (N_13106,N_12993,N_12917);
xnor U13107 (N_13107,N_12877,N_12946);
or U13108 (N_13108,N_12931,N_12791);
nand U13109 (N_13109,N_12873,N_12765);
and U13110 (N_13110,N_12921,N_12999);
xor U13111 (N_13111,N_12831,N_12853);
xnor U13112 (N_13112,N_12876,N_12790);
nand U13113 (N_13113,N_12841,N_12896);
nor U13114 (N_13114,N_12905,N_12944);
nand U13115 (N_13115,N_12800,N_12824);
or U13116 (N_13116,N_12990,N_12759);
and U13117 (N_13117,N_12889,N_12967);
and U13118 (N_13118,N_12980,N_12761);
nor U13119 (N_13119,N_12772,N_12906);
and U13120 (N_13120,N_12988,N_12786);
nand U13121 (N_13121,N_12778,N_12835);
and U13122 (N_13122,N_12871,N_12892);
xnor U13123 (N_13123,N_12913,N_12895);
nor U13124 (N_13124,N_12839,N_12756);
nor U13125 (N_13125,N_12752,N_12763);
xnor U13126 (N_13126,N_12865,N_12930);
xor U13127 (N_13127,N_12888,N_12766);
or U13128 (N_13128,N_12849,N_12948);
or U13129 (N_13129,N_12894,N_12815);
and U13130 (N_13130,N_12890,N_12878);
nand U13131 (N_13131,N_12932,N_12908);
nand U13132 (N_13132,N_12762,N_12943);
nor U13133 (N_13133,N_12806,N_12906);
nor U13134 (N_13134,N_12952,N_12944);
xnor U13135 (N_13135,N_12909,N_12870);
or U13136 (N_13136,N_12941,N_12753);
nor U13137 (N_13137,N_12834,N_12901);
xnor U13138 (N_13138,N_12889,N_12992);
and U13139 (N_13139,N_12888,N_12755);
and U13140 (N_13140,N_12792,N_12885);
nand U13141 (N_13141,N_12947,N_12966);
xnor U13142 (N_13142,N_12811,N_12993);
nor U13143 (N_13143,N_12835,N_12908);
or U13144 (N_13144,N_12905,N_12958);
and U13145 (N_13145,N_12764,N_12974);
and U13146 (N_13146,N_12955,N_12933);
nand U13147 (N_13147,N_12884,N_12913);
xor U13148 (N_13148,N_12751,N_12936);
xnor U13149 (N_13149,N_12891,N_12997);
or U13150 (N_13150,N_12813,N_12955);
or U13151 (N_13151,N_12909,N_12865);
nand U13152 (N_13152,N_12911,N_12979);
xor U13153 (N_13153,N_12990,N_12960);
nor U13154 (N_13154,N_12889,N_12931);
nand U13155 (N_13155,N_12817,N_12934);
xor U13156 (N_13156,N_12971,N_12798);
and U13157 (N_13157,N_12809,N_12787);
and U13158 (N_13158,N_12760,N_12997);
nor U13159 (N_13159,N_12787,N_12849);
xor U13160 (N_13160,N_12904,N_12807);
or U13161 (N_13161,N_12848,N_12793);
nand U13162 (N_13162,N_12870,N_12751);
nor U13163 (N_13163,N_12988,N_12936);
and U13164 (N_13164,N_12814,N_12911);
or U13165 (N_13165,N_12909,N_12913);
or U13166 (N_13166,N_12909,N_12762);
or U13167 (N_13167,N_12949,N_12994);
and U13168 (N_13168,N_12991,N_12914);
nor U13169 (N_13169,N_12750,N_12802);
or U13170 (N_13170,N_12900,N_12874);
nand U13171 (N_13171,N_12842,N_12823);
nand U13172 (N_13172,N_12863,N_12787);
nor U13173 (N_13173,N_12926,N_12980);
nor U13174 (N_13174,N_12901,N_12862);
xnor U13175 (N_13175,N_12897,N_12765);
nor U13176 (N_13176,N_12998,N_12750);
nor U13177 (N_13177,N_12830,N_12976);
and U13178 (N_13178,N_12878,N_12947);
or U13179 (N_13179,N_12798,N_12947);
and U13180 (N_13180,N_12795,N_12923);
or U13181 (N_13181,N_12994,N_12921);
or U13182 (N_13182,N_12919,N_12801);
nand U13183 (N_13183,N_12754,N_12936);
nor U13184 (N_13184,N_12888,N_12901);
nor U13185 (N_13185,N_12994,N_12801);
or U13186 (N_13186,N_12781,N_12966);
nor U13187 (N_13187,N_12933,N_12847);
and U13188 (N_13188,N_12898,N_12971);
nand U13189 (N_13189,N_12773,N_12900);
and U13190 (N_13190,N_12970,N_12796);
nand U13191 (N_13191,N_12943,N_12938);
xor U13192 (N_13192,N_12997,N_12819);
nand U13193 (N_13193,N_12799,N_12773);
nor U13194 (N_13194,N_12926,N_12833);
nor U13195 (N_13195,N_12879,N_12860);
nor U13196 (N_13196,N_12950,N_12965);
nand U13197 (N_13197,N_12750,N_12764);
xor U13198 (N_13198,N_12863,N_12858);
nor U13199 (N_13199,N_12938,N_12945);
or U13200 (N_13200,N_12878,N_12828);
and U13201 (N_13201,N_12925,N_12819);
and U13202 (N_13202,N_12974,N_12922);
nor U13203 (N_13203,N_12926,N_12869);
xnor U13204 (N_13204,N_12864,N_12789);
nand U13205 (N_13205,N_12759,N_12755);
and U13206 (N_13206,N_12809,N_12997);
xor U13207 (N_13207,N_12928,N_12893);
nor U13208 (N_13208,N_12764,N_12909);
xor U13209 (N_13209,N_12890,N_12756);
xnor U13210 (N_13210,N_12903,N_12959);
nor U13211 (N_13211,N_12899,N_12874);
xor U13212 (N_13212,N_12975,N_12823);
or U13213 (N_13213,N_12962,N_12961);
or U13214 (N_13214,N_12791,N_12985);
xnor U13215 (N_13215,N_12924,N_12792);
or U13216 (N_13216,N_12845,N_12849);
nor U13217 (N_13217,N_12908,N_12986);
xnor U13218 (N_13218,N_12963,N_12914);
or U13219 (N_13219,N_12830,N_12775);
and U13220 (N_13220,N_12831,N_12827);
or U13221 (N_13221,N_12905,N_12868);
xor U13222 (N_13222,N_12784,N_12938);
xor U13223 (N_13223,N_12800,N_12880);
and U13224 (N_13224,N_12831,N_12820);
or U13225 (N_13225,N_12937,N_12780);
and U13226 (N_13226,N_12785,N_12875);
or U13227 (N_13227,N_12973,N_12802);
and U13228 (N_13228,N_12855,N_12851);
nor U13229 (N_13229,N_12810,N_12968);
xor U13230 (N_13230,N_12771,N_12882);
and U13231 (N_13231,N_12902,N_12812);
nand U13232 (N_13232,N_12990,N_12926);
and U13233 (N_13233,N_12870,N_12831);
nor U13234 (N_13234,N_12851,N_12760);
nand U13235 (N_13235,N_12865,N_12960);
nand U13236 (N_13236,N_12826,N_12943);
or U13237 (N_13237,N_12869,N_12813);
nor U13238 (N_13238,N_12860,N_12841);
nor U13239 (N_13239,N_12783,N_12884);
and U13240 (N_13240,N_12773,N_12762);
xnor U13241 (N_13241,N_12926,N_12978);
xnor U13242 (N_13242,N_12926,N_12880);
xnor U13243 (N_13243,N_12903,N_12789);
nand U13244 (N_13244,N_12879,N_12867);
and U13245 (N_13245,N_12879,N_12903);
nand U13246 (N_13246,N_12870,N_12756);
or U13247 (N_13247,N_12793,N_12824);
and U13248 (N_13248,N_12986,N_12833);
or U13249 (N_13249,N_12852,N_12954);
nand U13250 (N_13250,N_13004,N_13058);
nand U13251 (N_13251,N_13142,N_13036);
or U13252 (N_13252,N_13071,N_13165);
nand U13253 (N_13253,N_13126,N_13236);
xor U13254 (N_13254,N_13180,N_13013);
nand U13255 (N_13255,N_13108,N_13211);
nor U13256 (N_13256,N_13124,N_13100);
nor U13257 (N_13257,N_13215,N_13105);
xnor U13258 (N_13258,N_13009,N_13096);
nor U13259 (N_13259,N_13040,N_13000);
or U13260 (N_13260,N_13187,N_13116);
nand U13261 (N_13261,N_13195,N_13148);
or U13262 (N_13262,N_13169,N_13183);
and U13263 (N_13263,N_13133,N_13177);
xor U13264 (N_13264,N_13098,N_13055);
and U13265 (N_13265,N_13225,N_13045);
and U13266 (N_13266,N_13086,N_13031);
nor U13267 (N_13267,N_13011,N_13172);
or U13268 (N_13268,N_13216,N_13151);
xor U13269 (N_13269,N_13099,N_13175);
and U13270 (N_13270,N_13022,N_13028);
and U13271 (N_13271,N_13076,N_13164);
and U13272 (N_13272,N_13041,N_13034);
and U13273 (N_13273,N_13242,N_13107);
xnor U13274 (N_13274,N_13176,N_13209);
xnor U13275 (N_13275,N_13042,N_13219);
or U13276 (N_13276,N_13154,N_13057);
nand U13277 (N_13277,N_13199,N_13248);
nand U13278 (N_13278,N_13155,N_13162);
nor U13279 (N_13279,N_13080,N_13049);
nor U13280 (N_13280,N_13005,N_13050);
nand U13281 (N_13281,N_13025,N_13149);
nor U13282 (N_13282,N_13051,N_13249);
nand U13283 (N_13283,N_13019,N_13048);
or U13284 (N_13284,N_13246,N_13145);
and U13285 (N_13285,N_13137,N_13161);
xor U13286 (N_13286,N_13212,N_13044);
nor U13287 (N_13287,N_13113,N_13073);
xnor U13288 (N_13288,N_13127,N_13224);
or U13289 (N_13289,N_13132,N_13115);
nand U13290 (N_13290,N_13181,N_13208);
nand U13291 (N_13291,N_13245,N_13141);
xnor U13292 (N_13292,N_13217,N_13231);
or U13293 (N_13293,N_13012,N_13170);
nor U13294 (N_13294,N_13066,N_13078);
nor U13295 (N_13295,N_13119,N_13146);
nand U13296 (N_13296,N_13026,N_13092);
and U13297 (N_13297,N_13232,N_13226);
xor U13298 (N_13298,N_13082,N_13110);
nand U13299 (N_13299,N_13213,N_13056);
xor U13300 (N_13300,N_13241,N_13106);
nand U13301 (N_13301,N_13240,N_13160);
xnor U13302 (N_13302,N_13139,N_13191);
and U13303 (N_13303,N_13001,N_13182);
nor U13304 (N_13304,N_13196,N_13239);
xor U13305 (N_13305,N_13143,N_13220);
and U13306 (N_13306,N_13010,N_13035);
nand U13307 (N_13307,N_13024,N_13184);
nor U13308 (N_13308,N_13186,N_13152);
or U13309 (N_13309,N_13174,N_13074);
nor U13310 (N_13310,N_13083,N_13136);
and U13311 (N_13311,N_13059,N_13179);
xnor U13312 (N_13312,N_13079,N_13192);
or U13313 (N_13313,N_13085,N_13144);
nand U13314 (N_13314,N_13157,N_13065);
nor U13315 (N_13315,N_13054,N_13037);
and U13316 (N_13316,N_13068,N_13244);
or U13317 (N_13317,N_13029,N_13150);
nand U13318 (N_13318,N_13128,N_13084);
nor U13319 (N_13319,N_13189,N_13077);
nand U13320 (N_13320,N_13193,N_13023);
or U13321 (N_13321,N_13178,N_13061);
and U13322 (N_13322,N_13147,N_13006);
nand U13323 (N_13323,N_13102,N_13003);
nor U13324 (N_13324,N_13104,N_13043);
nand U13325 (N_13325,N_13087,N_13093);
nor U13326 (N_13326,N_13218,N_13221);
nor U13327 (N_13327,N_13016,N_13168);
and U13328 (N_13328,N_13038,N_13138);
xor U13329 (N_13329,N_13122,N_13117);
nor U13330 (N_13330,N_13018,N_13135);
and U13331 (N_13331,N_13053,N_13046);
and U13332 (N_13332,N_13089,N_13047);
xnor U13333 (N_13333,N_13101,N_13069);
xnor U13334 (N_13334,N_13072,N_13230);
nor U13335 (N_13335,N_13112,N_13198);
nand U13336 (N_13336,N_13238,N_13062);
and U13337 (N_13337,N_13091,N_13064);
nand U13338 (N_13338,N_13134,N_13033);
or U13339 (N_13339,N_13233,N_13167);
nand U13340 (N_13340,N_13114,N_13123);
or U13341 (N_13341,N_13008,N_13039);
xor U13342 (N_13342,N_13166,N_13094);
nand U13343 (N_13343,N_13159,N_13190);
nor U13344 (N_13344,N_13197,N_13021);
xnor U13345 (N_13345,N_13125,N_13204);
nor U13346 (N_13346,N_13120,N_13163);
nand U13347 (N_13347,N_13081,N_13130);
and U13348 (N_13348,N_13227,N_13030);
nor U13349 (N_13349,N_13171,N_13229);
nor U13350 (N_13350,N_13235,N_13103);
and U13351 (N_13351,N_13158,N_13185);
xor U13352 (N_13352,N_13140,N_13243);
xor U13353 (N_13353,N_13194,N_13247);
nand U13354 (N_13354,N_13060,N_13111);
xor U13355 (N_13355,N_13207,N_13007);
nand U13356 (N_13356,N_13090,N_13205);
xnor U13357 (N_13357,N_13052,N_13156);
or U13358 (N_13358,N_13131,N_13017);
and U13359 (N_13359,N_13067,N_13201);
xor U13360 (N_13360,N_13203,N_13210);
nor U13361 (N_13361,N_13129,N_13222);
xnor U13362 (N_13362,N_13118,N_13020);
or U13363 (N_13363,N_13075,N_13032);
and U13364 (N_13364,N_13121,N_13237);
or U13365 (N_13365,N_13095,N_13109);
or U13366 (N_13366,N_13214,N_13200);
and U13367 (N_13367,N_13027,N_13202);
xnor U13368 (N_13368,N_13070,N_13088);
nand U13369 (N_13369,N_13173,N_13206);
or U13370 (N_13370,N_13063,N_13002);
nor U13371 (N_13371,N_13097,N_13223);
or U13372 (N_13372,N_13188,N_13014);
or U13373 (N_13373,N_13228,N_13015);
nand U13374 (N_13374,N_13153,N_13234);
and U13375 (N_13375,N_13016,N_13061);
and U13376 (N_13376,N_13072,N_13024);
xnor U13377 (N_13377,N_13075,N_13198);
and U13378 (N_13378,N_13231,N_13235);
or U13379 (N_13379,N_13199,N_13042);
nor U13380 (N_13380,N_13155,N_13103);
xor U13381 (N_13381,N_13085,N_13231);
and U13382 (N_13382,N_13195,N_13136);
xor U13383 (N_13383,N_13208,N_13206);
xnor U13384 (N_13384,N_13070,N_13008);
nor U13385 (N_13385,N_13146,N_13007);
nor U13386 (N_13386,N_13001,N_13106);
nor U13387 (N_13387,N_13101,N_13003);
and U13388 (N_13388,N_13090,N_13142);
xor U13389 (N_13389,N_13131,N_13146);
and U13390 (N_13390,N_13041,N_13229);
or U13391 (N_13391,N_13013,N_13052);
xor U13392 (N_13392,N_13186,N_13166);
or U13393 (N_13393,N_13000,N_13017);
xnor U13394 (N_13394,N_13074,N_13203);
or U13395 (N_13395,N_13191,N_13199);
nor U13396 (N_13396,N_13228,N_13035);
nor U13397 (N_13397,N_13016,N_13067);
nand U13398 (N_13398,N_13093,N_13225);
and U13399 (N_13399,N_13034,N_13125);
nor U13400 (N_13400,N_13056,N_13034);
nand U13401 (N_13401,N_13064,N_13111);
and U13402 (N_13402,N_13092,N_13038);
nand U13403 (N_13403,N_13028,N_13168);
xor U13404 (N_13404,N_13107,N_13177);
or U13405 (N_13405,N_13176,N_13220);
nor U13406 (N_13406,N_13179,N_13211);
or U13407 (N_13407,N_13168,N_13228);
or U13408 (N_13408,N_13237,N_13077);
or U13409 (N_13409,N_13035,N_13023);
and U13410 (N_13410,N_13059,N_13145);
or U13411 (N_13411,N_13096,N_13189);
nand U13412 (N_13412,N_13074,N_13103);
xor U13413 (N_13413,N_13248,N_13131);
xor U13414 (N_13414,N_13163,N_13207);
or U13415 (N_13415,N_13207,N_13048);
nor U13416 (N_13416,N_13083,N_13167);
or U13417 (N_13417,N_13244,N_13144);
nor U13418 (N_13418,N_13139,N_13126);
nand U13419 (N_13419,N_13107,N_13058);
nor U13420 (N_13420,N_13033,N_13177);
or U13421 (N_13421,N_13187,N_13068);
xor U13422 (N_13422,N_13220,N_13190);
and U13423 (N_13423,N_13076,N_13204);
nor U13424 (N_13424,N_13063,N_13226);
or U13425 (N_13425,N_13116,N_13017);
and U13426 (N_13426,N_13025,N_13078);
nand U13427 (N_13427,N_13074,N_13028);
and U13428 (N_13428,N_13004,N_13095);
nand U13429 (N_13429,N_13170,N_13081);
nand U13430 (N_13430,N_13150,N_13096);
and U13431 (N_13431,N_13066,N_13163);
or U13432 (N_13432,N_13003,N_13067);
xor U13433 (N_13433,N_13172,N_13106);
nor U13434 (N_13434,N_13199,N_13116);
nor U13435 (N_13435,N_13133,N_13233);
or U13436 (N_13436,N_13055,N_13179);
nor U13437 (N_13437,N_13100,N_13047);
nor U13438 (N_13438,N_13231,N_13224);
and U13439 (N_13439,N_13023,N_13194);
and U13440 (N_13440,N_13061,N_13241);
nor U13441 (N_13441,N_13076,N_13087);
xnor U13442 (N_13442,N_13037,N_13137);
or U13443 (N_13443,N_13220,N_13237);
xor U13444 (N_13444,N_13136,N_13056);
and U13445 (N_13445,N_13230,N_13115);
and U13446 (N_13446,N_13108,N_13188);
nand U13447 (N_13447,N_13112,N_13173);
xnor U13448 (N_13448,N_13005,N_13231);
nand U13449 (N_13449,N_13100,N_13125);
xor U13450 (N_13450,N_13109,N_13216);
nor U13451 (N_13451,N_13007,N_13198);
nand U13452 (N_13452,N_13032,N_13222);
and U13453 (N_13453,N_13000,N_13120);
nor U13454 (N_13454,N_13196,N_13134);
nand U13455 (N_13455,N_13034,N_13192);
and U13456 (N_13456,N_13128,N_13132);
xnor U13457 (N_13457,N_13215,N_13244);
xor U13458 (N_13458,N_13048,N_13121);
nor U13459 (N_13459,N_13204,N_13005);
or U13460 (N_13460,N_13136,N_13166);
and U13461 (N_13461,N_13019,N_13102);
and U13462 (N_13462,N_13192,N_13133);
and U13463 (N_13463,N_13158,N_13055);
nor U13464 (N_13464,N_13151,N_13192);
nand U13465 (N_13465,N_13036,N_13169);
or U13466 (N_13466,N_13237,N_13214);
and U13467 (N_13467,N_13223,N_13230);
and U13468 (N_13468,N_13041,N_13145);
and U13469 (N_13469,N_13006,N_13171);
nor U13470 (N_13470,N_13136,N_13139);
nor U13471 (N_13471,N_13179,N_13196);
and U13472 (N_13472,N_13014,N_13167);
or U13473 (N_13473,N_13137,N_13059);
xor U13474 (N_13474,N_13198,N_13216);
xor U13475 (N_13475,N_13028,N_13186);
xor U13476 (N_13476,N_13127,N_13161);
nand U13477 (N_13477,N_13233,N_13159);
or U13478 (N_13478,N_13205,N_13082);
nand U13479 (N_13479,N_13006,N_13150);
or U13480 (N_13480,N_13162,N_13172);
nand U13481 (N_13481,N_13230,N_13244);
nor U13482 (N_13482,N_13210,N_13110);
xnor U13483 (N_13483,N_13178,N_13186);
nand U13484 (N_13484,N_13124,N_13038);
nor U13485 (N_13485,N_13093,N_13195);
nor U13486 (N_13486,N_13045,N_13015);
nand U13487 (N_13487,N_13163,N_13147);
nand U13488 (N_13488,N_13195,N_13240);
or U13489 (N_13489,N_13008,N_13196);
xor U13490 (N_13490,N_13225,N_13008);
xor U13491 (N_13491,N_13100,N_13128);
nand U13492 (N_13492,N_13019,N_13010);
nand U13493 (N_13493,N_13021,N_13128);
or U13494 (N_13494,N_13068,N_13039);
nand U13495 (N_13495,N_13111,N_13027);
xor U13496 (N_13496,N_13107,N_13002);
and U13497 (N_13497,N_13062,N_13064);
nand U13498 (N_13498,N_13078,N_13067);
nor U13499 (N_13499,N_13096,N_13032);
xor U13500 (N_13500,N_13252,N_13420);
and U13501 (N_13501,N_13403,N_13250);
and U13502 (N_13502,N_13475,N_13337);
xnor U13503 (N_13503,N_13363,N_13412);
or U13504 (N_13504,N_13479,N_13357);
xor U13505 (N_13505,N_13466,N_13306);
xnor U13506 (N_13506,N_13325,N_13279);
and U13507 (N_13507,N_13369,N_13387);
and U13508 (N_13508,N_13326,N_13285);
xnor U13509 (N_13509,N_13333,N_13267);
or U13510 (N_13510,N_13347,N_13254);
or U13511 (N_13511,N_13471,N_13410);
nor U13512 (N_13512,N_13472,N_13436);
nor U13513 (N_13513,N_13257,N_13274);
and U13514 (N_13514,N_13276,N_13344);
xnor U13515 (N_13515,N_13486,N_13413);
nor U13516 (N_13516,N_13314,N_13409);
xnor U13517 (N_13517,N_13497,N_13275);
and U13518 (N_13518,N_13284,N_13353);
and U13519 (N_13519,N_13414,N_13376);
or U13520 (N_13520,N_13312,N_13434);
xnor U13521 (N_13521,N_13457,N_13321);
and U13522 (N_13522,N_13291,N_13322);
nor U13523 (N_13523,N_13378,N_13340);
nor U13524 (N_13524,N_13401,N_13308);
nand U13525 (N_13525,N_13271,N_13473);
nor U13526 (N_13526,N_13263,N_13330);
xor U13527 (N_13527,N_13418,N_13426);
nand U13528 (N_13528,N_13290,N_13411);
or U13529 (N_13529,N_13354,N_13341);
or U13530 (N_13530,N_13358,N_13361);
or U13531 (N_13531,N_13327,N_13262);
nor U13532 (N_13532,N_13251,N_13311);
xor U13533 (N_13533,N_13281,N_13295);
or U13534 (N_13534,N_13255,N_13421);
xor U13535 (N_13535,N_13296,N_13382);
and U13536 (N_13536,N_13294,N_13396);
nand U13537 (N_13537,N_13392,N_13364);
nor U13538 (N_13538,N_13261,N_13459);
nor U13539 (N_13539,N_13343,N_13456);
nand U13540 (N_13540,N_13366,N_13370);
xor U13541 (N_13541,N_13367,N_13423);
nand U13542 (N_13542,N_13407,N_13338);
nand U13543 (N_13543,N_13277,N_13336);
nand U13544 (N_13544,N_13481,N_13352);
nor U13545 (N_13545,N_13297,N_13480);
nand U13546 (N_13546,N_13298,N_13304);
xor U13547 (N_13547,N_13455,N_13339);
nand U13548 (N_13548,N_13345,N_13394);
nand U13549 (N_13549,N_13381,N_13334);
nor U13550 (N_13550,N_13299,N_13342);
nor U13551 (N_13551,N_13493,N_13417);
nand U13552 (N_13552,N_13498,N_13273);
nand U13553 (N_13553,N_13406,N_13402);
xnor U13554 (N_13554,N_13292,N_13470);
xnor U13555 (N_13555,N_13391,N_13408);
and U13556 (N_13556,N_13443,N_13303);
or U13557 (N_13557,N_13465,N_13260);
nand U13558 (N_13558,N_13454,N_13464);
nand U13559 (N_13559,N_13383,N_13256);
and U13560 (N_13560,N_13368,N_13259);
xnor U13561 (N_13561,N_13258,N_13458);
nor U13562 (N_13562,N_13395,N_13490);
and U13563 (N_13563,N_13390,N_13425);
or U13564 (N_13564,N_13483,N_13374);
or U13565 (N_13565,N_13415,N_13346);
and U13566 (N_13566,N_13315,N_13451);
or U13567 (N_13567,N_13307,N_13269);
or U13568 (N_13568,N_13253,N_13373);
and U13569 (N_13569,N_13301,N_13404);
nor U13570 (N_13570,N_13355,N_13427);
nand U13571 (N_13571,N_13265,N_13323);
xor U13572 (N_13572,N_13380,N_13362);
xor U13573 (N_13573,N_13416,N_13468);
nand U13574 (N_13574,N_13313,N_13293);
or U13575 (N_13575,N_13283,N_13328);
or U13576 (N_13576,N_13499,N_13492);
or U13577 (N_13577,N_13371,N_13300);
xor U13578 (N_13578,N_13460,N_13309);
xor U13579 (N_13579,N_13316,N_13289);
or U13580 (N_13580,N_13446,N_13440);
nor U13581 (N_13581,N_13282,N_13442);
nand U13582 (N_13582,N_13445,N_13450);
nand U13583 (N_13583,N_13431,N_13422);
nand U13584 (N_13584,N_13437,N_13424);
xor U13585 (N_13585,N_13288,N_13305);
xnor U13586 (N_13586,N_13287,N_13485);
nor U13587 (N_13587,N_13432,N_13452);
or U13588 (N_13588,N_13439,N_13435);
xor U13589 (N_13589,N_13482,N_13329);
or U13590 (N_13590,N_13385,N_13487);
and U13591 (N_13591,N_13428,N_13474);
xor U13592 (N_13592,N_13320,N_13441);
nor U13593 (N_13593,N_13270,N_13398);
and U13594 (N_13594,N_13429,N_13356);
or U13595 (N_13595,N_13377,N_13318);
nor U13596 (N_13596,N_13433,N_13419);
nor U13597 (N_13597,N_13266,N_13463);
and U13598 (N_13598,N_13389,N_13365);
nand U13599 (N_13599,N_13268,N_13324);
nor U13600 (N_13600,N_13310,N_13286);
nand U13601 (N_13601,N_13384,N_13484);
nor U13602 (N_13602,N_13400,N_13453);
nor U13603 (N_13603,N_13438,N_13278);
nand U13604 (N_13604,N_13388,N_13280);
or U13605 (N_13605,N_13386,N_13462);
and U13606 (N_13606,N_13469,N_13495);
nor U13607 (N_13607,N_13397,N_13379);
and U13608 (N_13608,N_13444,N_13359);
or U13609 (N_13609,N_13489,N_13476);
nor U13610 (N_13610,N_13448,N_13494);
or U13611 (N_13611,N_13477,N_13488);
nand U13612 (N_13612,N_13360,N_13496);
xor U13613 (N_13613,N_13375,N_13351);
or U13614 (N_13614,N_13399,N_13335);
nand U13615 (N_13615,N_13491,N_13430);
or U13616 (N_13616,N_13461,N_13393);
nor U13617 (N_13617,N_13319,N_13332);
or U13618 (N_13618,N_13302,N_13272);
or U13619 (N_13619,N_13264,N_13372);
or U13620 (N_13620,N_13467,N_13405);
nor U13621 (N_13621,N_13350,N_13349);
or U13622 (N_13622,N_13478,N_13447);
xor U13623 (N_13623,N_13348,N_13331);
or U13624 (N_13624,N_13449,N_13317);
xnor U13625 (N_13625,N_13422,N_13377);
nor U13626 (N_13626,N_13371,N_13339);
or U13627 (N_13627,N_13415,N_13350);
nand U13628 (N_13628,N_13336,N_13321);
xnor U13629 (N_13629,N_13325,N_13439);
nor U13630 (N_13630,N_13372,N_13448);
xor U13631 (N_13631,N_13267,N_13417);
or U13632 (N_13632,N_13461,N_13368);
xnor U13633 (N_13633,N_13382,N_13352);
and U13634 (N_13634,N_13303,N_13419);
nand U13635 (N_13635,N_13453,N_13313);
nor U13636 (N_13636,N_13482,N_13411);
and U13637 (N_13637,N_13395,N_13349);
nand U13638 (N_13638,N_13301,N_13250);
nand U13639 (N_13639,N_13265,N_13470);
and U13640 (N_13640,N_13402,N_13432);
xnor U13641 (N_13641,N_13461,N_13444);
xnor U13642 (N_13642,N_13322,N_13376);
nand U13643 (N_13643,N_13299,N_13391);
and U13644 (N_13644,N_13250,N_13305);
nor U13645 (N_13645,N_13283,N_13364);
xor U13646 (N_13646,N_13445,N_13256);
and U13647 (N_13647,N_13396,N_13486);
or U13648 (N_13648,N_13421,N_13347);
nand U13649 (N_13649,N_13321,N_13374);
or U13650 (N_13650,N_13390,N_13427);
or U13651 (N_13651,N_13343,N_13374);
xor U13652 (N_13652,N_13460,N_13302);
and U13653 (N_13653,N_13301,N_13255);
nor U13654 (N_13654,N_13477,N_13482);
nand U13655 (N_13655,N_13294,N_13464);
or U13656 (N_13656,N_13470,N_13476);
nand U13657 (N_13657,N_13285,N_13397);
and U13658 (N_13658,N_13342,N_13280);
nor U13659 (N_13659,N_13374,N_13477);
or U13660 (N_13660,N_13467,N_13327);
xor U13661 (N_13661,N_13497,N_13287);
xor U13662 (N_13662,N_13416,N_13470);
nor U13663 (N_13663,N_13412,N_13480);
nor U13664 (N_13664,N_13487,N_13366);
xor U13665 (N_13665,N_13335,N_13296);
xor U13666 (N_13666,N_13323,N_13334);
and U13667 (N_13667,N_13325,N_13269);
nand U13668 (N_13668,N_13478,N_13319);
xnor U13669 (N_13669,N_13404,N_13251);
or U13670 (N_13670,N_13367,N_13352);
nand U13671 (N_13671,N_13328,N_13395);
and U13672 (N_13672,N_13415,N_13492);
nand U13673 (N_13673,N_13445,N_13392);
nand U13674 (N_13674,N_13264,N_13379);
xnor U13675 (N_13675,N_13486,N_13375);
or U13676 (N_13676,N_13374,N_13452);
nor U13677 (N_13677,N_13264,N_13351);
or U13678 (N_13678,N_13254,N_13448);
or U13679 (N_13679,N_13338,N_13455);
xnor U13680 (N_13680,N_13318,N_13435);
xnor U13681 (N_13681,N_13488,N_13321);
xor U13682 (N_13682,N_13377,N_13343);
or U13683 (N_13683,N_13389,N_13427);
xnor U13684 (N_13684,N_13287,N_13289);
nand U13685 (N_13685,N_13484,N_13326);
xor U13686 (N_13686,N_13469,N_13446);
and U13687 (N_13687,N_13482,N_13393);
nor U13688 (N_13688,N_13499,N_13307);
nand U13689 (N_13689,N_13323,N_13446);
xor U13690 (N_13690,N_13407,N_13493);
xor U13691 (N_13691,N_13495,N_13337);
or U13692 (N_13692,N_13391,N_13399);
xor U13693 (N_13693,N_13282,N_13285);
nor U13694 (N_13694,N_13495,N_13318);
nand U13695 (N_13695,N_13287,N_13311);
or U13696 (N_13696,N_13261,N_13429);
nand U13697 (N_13697,N_13311,N_13303);
xnor U13698 (N_13698,N_13449,N_13397);
nand U13699 (N_13699,N_13251,N_13264);
and U13700 (N_13700,N_13454,N_13366);
nor U13701 (N_13701,N_13434,N_13422);
nand U13702 (N_13702,N_13325,N_13336);
and U13703 (N_13703,N_13274,N_13464);
or U13704 (N_13704,N_13444,N_13451);
nand U13705 (N_13705,N_13362,N_13488);
or U13706 (N_13706,N_13437,N_13464);
or U13707 (N_13707,N_13383,N_13307);
or U13708 (N_13708,N_13480,N_13286);
nand U13709 (N_13709,N_13258,N_13473);
or U13710 (N_13710,N_13252,N_13293);
or U13711 (N_13711,N_13442,N_13451);
xnor U13712 (N_13712,N_13402,N_13449);
and U13713 (N_13713,N_13323,N_13281);
nand U13714 (N_13714,N_13412,N_13350);
nand U13715 (N_13715,N_13382,N_13321);
nor U13716 (N_13716,N_13375,N_13267);
xnor U13717 (N_13717,N_13390,N_13393);
or U13718 (N_13718,N_13372,N_13387);
and U13719 (N_13719,N_13435,N_13342);
nor U13720 (N_13720,N_13497,N_13385);
xor U13721 (N_13721,N_13435,N_13316);
xnor U13722 (N_13722,N_13388,N_13269);
nor U13723 (N_13723,N_13299,N_13315);
and U13724 (N_13724,N_13265,N_13480);
nand U13725 (N_13725,N_13426,N_13450);
xnor U13726 (N_13726,N_13276,N_13335);
nor U13727 (N_13727,N_13497,N_13282);
nand U13728 (N_13728,N_13355,N_13408);
or U13729 (N_13729,N_13332,N_13435);
or U13730 (N_13730,N_13483,N_13389);
or U13731 (N_13731,N_13317,N_13469);
nor U13732 (N_13732,N_13330,N_13276);
nand U13733 (N_13733,N_13311,N_13425);
and U13734 (N_13734,N_13284,N_13332);
nand U13735 (N_13735,N_13363,N_13419);
nor U13736 (N_13736,N_13318,N_13373);
or U13737 (N_13737,N_13475,N_13272);
and U13738 (N_13738,N_13457,N_13361);
or U13739 (N_13739,N_13462,N_13343);
and U13740 (N_13740,N_13411,N_13399);
xnor U13741 (N_13741,N_13467,N_13316);
and U13742 (N_13742,N_13334,N_13324);
nor U13743 (N_13743,N_13443,N_13329);
and U13744 (N_13744,N_13339,N_13338);
xnor U13745 (N_13745,N_13256,N_13381);
nand U13746 (N_13746,N_13325,N_13323);
nand U13747 (N_13747,N_13402,N_13472);
nor U13748 (N_13748,N_13419,N_13279);
or U13749 (N_13749,N_13386,N_13342);
and U13750 (N_13750,N_13559,N_13513);
nand U13751 (N_13751,N_13586,N_13566);
xor U13752 (N_13752,N_13505,N_13656);
nand U13753 (N_13753,N_13530,N_13585);
or U13754 (N_13754,N_13556,N_13717);
or U13755 (N_13755,N_13652,N_13744);
and U13756 (N_13756,N_13736,N_13662);
nand U13757 (N_13757,N_13592,N_13682);
nand U13758 (N_13758,N_13548,N_13683);
or U13759 (N_13759,N_13723,N_13713);
nor U13760 (N_13760,N_13712,N_13634);
xor U13761 (N_13761,N_13646,N_13573);
nand U13762 (N_13762,N_13577,N_13593);
or U13763 (N_13763,N_13678,N_13549);
nand U13764 (N_13764,N_13668,N_13676);
nand U13765 (N_13765,N_13605,N_13720);
xnor U13766 (N_13766,N_13677,N_13655);
nand U13767 (N_13767,N_13700,N_13747);
and U13768 (N_13768,N_13533,N_13689);
nand U13769 (N_13769,N_13738,N_13580);
or U13770 (N_13770,N_13614,N_13638);
xor U13771 (N_13771,N_13635,N_13616);
nand U13772 (N_13772,N_13623,N_13708);
and U13773 (N_13773,N_13613,N_13532);
or U13774 (N_13774,N_13698,N_13692);
and U13775 (N_13775,N_13597,N_13546);
or U13776 (N_13776,N_13749,N_13693);
nand U13777 (N_13777,N_13551,N_13604);
xor U13778 (N_13778,N_13620,N_13695);
xnor U13779 (N_13779,N_13732,N_13507);
and U13780 (N_13780,N_13598,N_13557);
or U13781 (N_13781,N_13517,N_13528);
and U13782 (N_13782,N_13748,N_13608);
nand U13783 (N_13783,N_13703,N_13624);
nand U13784 (N_13784,N_13603,N_13569);
xor U13785 (N_13785,N_13511,N_13726);
xnor U13786 (N_13786,N_13576,N_13628);
or U13787 (N_13787,N_13591,N_13588);
and U13788 (N_13788,N_13639,N_13550);
and U13789 (N_13789,N_13632,N_13705);
nand U13790 (N_13790,N_13711,N_13663);
xor U13791 (N_13791,N_13706,N_13694);
or U13792 (N_13792,N_13515,N_13534);
nand U13793 (N_13793,N_13718,N_13615);
nand U13794 (N_13794,N_13699,N_13640);
nand U13795 (N_13795,N_13607,N_13503);
or U13796 (N_13796,N_13696,N_13554);
or U13797 (N_13797,N_13527,N_13673);
nand U13798 (N_13798,N_13715,N_13645);
xor U13799 (N_13799,N_13649,N_13724);
or U13800 (N_13800,N_13589,N_13571);
nor U13801 (N_13801,N_13508,N_13667);
nand U13802 (N_13802,N_13562,N_13567);
or U13803 (N_13803,N_13594,N_13704);
nand U13804 (N_13804,N_13502,N_13596);
xor U13805 (N_13805,N_13519,N_13583);
nor U13806 (N_13806,N_13581,N_13669);
nand U13807 (N_13807,N_13545,N_13619);
nor U13808 (N_13808,N_13627,N_13524);
or U13809 (N_13809,N_13670,N_13741);
nor U13810 (N_13810,N_13686,N_13504);
and U13811 (N_13811,N_13540,N_13609);
and U13812 (N_13812,N_13709,N_13500);
nor U13813 (N_13813,N_13531,N_13730);
and U13814 (N_13814,N_13561,N_13737);
nor U13815 (N_13815,N_13553,N_13740);
xor U13816 (N_13816,N_13538,N_13707);
and U13817 (N_13817,N_13743,N_13629);
xor U13818 (N_13818,N_13701,N_13688);
nor U13819 (N_13819,N_13525,N_13637);
nor U13820 (N_13820,N_13539,N_13582);
nand U13821 (N_13821,N_13560,N_13716);
xor U13822 (N_13822,N_13735,N_13660);
nand U13823 (N_13823,N_13684,N_13512);
and U13824 (N_13824,N_13636,N_13685);
nor U13825 (N_13825,N_13612,N_13610);
and U13826 (N_13826,N_13690,N_13579);
nor U13827 (N_13827,N_13568,N_13552);
and U13828 (N_13828,N_13746,N_13602);
or U13829 (N_13829,N_13520,N_13675);
or U13830 (N_13830,N_13570,N_13651);
and U13831 (N_13831,N_13563,N_13555);
nor U13832 (N_13832,N_13537,N_13714);
nand U13833 (N_13833,N_13543,N_13681);
or U13834 (N_13834,N_13697,N_13745);
and U13835 (N_13835,N_13742,N_13691);
xor U13836 (N_13836,N_13565,N_13587);
and U13837 (N_13837,N_13666,N_13642);
or U13838 (N_13838,N_13510,N_13572);
nand U13839 (N_13839,N_13626,N_13659);
nand U13840 (N_13840,N_13687,N_13725);
nor U13841 (N_13841,N_13647,N_13535);
nand U13842 (N_13842,N_13518,N_13575);
nor U13843 (N_13843,N_13542,N_13661);
nor U13844 (N_13844,N_13618,N_13536);
or U13845 (N_13845,N_13643,N_13633);
nor U13846 (N_13846,N_13621,N_13727);
and U13847 (N_13847,N_13558,N_13617);
xnor U13848 (N_13848,N_13710,N_13599);
or U13849 (N_13849,N_13529,N_13731);
nand U13850 (N_13850,N_13657,N_13679);
and U13851 (N_13851,N_13648,N_13547);
and U13852 (N_13852,N_13721,N_13590);
and U13853 (N_13853,N_13650,N_13672);
xnor U13854 (N_13854,N_13664,N_13541);
and U13855 (N_13855,N_13641,N_13653);
nor U13856 (N_13856,N_13578,N_13584);
xor U13857 (N_13857,N_13521,N_13671);
nand U13858 (N_13858,N_13523,N_13526);
nand U13859 (N_13859,N_13631,N_13654);
nor U13860 (N_13860,N_13644,N_13622);
or U13861 (N_13861,N_13564,N_13522);
xor U13862 (N_13862,N_13606,N_13702);
and U13863 (N_13863,N_13509,N_13601);
and U13864 (N_13864,N_13516,N_13595);
xor U13865 (N_13865,N_13600,N_13734);
and U13866 (N_13866,N_13501,N_13514);
nor U13867 (N_13867,N_13630,N_13611);
and U13868 (N_13868,N_13739,N_13574);
nand U13869 (N_13869,N_13733,N_13658);
or U13870 (N_13870,N_13665,N_13674);
or U13871 (N_13871,N_13719,N_13729);
and U13872 (N_13872,N_13625,N_13506);
and U13873 (N_13873,N_13722,N_13544);
nor U13874 (N_13874,N_13680,N_13728);
and U13875 (N_13875,N_13565,N_13549);
nand U13876 (N_13876,N_13649,N_13696);
nor U13877 (N_13877,N_13557,N_13665);
nor U13878 (N_13878,N_13609,N_13710);
nand U13879 (N_13879,N_13625,N_13503);
xor U13880 (N_13880,N_13625,N_13631);
xnor U13881 (N_13881,N_13714,N_13584);
and U13882 (N_13882,N_13661,N_13573);
or U13883 (N_13883,N_13509,N_13597);
nand U13884 (N_13884,N_13650,N_13735);
nor U13885 (N_13885,N_13718,N_13523);
xnor U13886 (N_13886,N_13691,N_13528);
xor U13887 (N_13887,N_13710,N_13566);
xnor U13888 (N_13888,N_13579,N_13536);
or U13889 (N_13889,N_13526,N_13655);
nand U13890 (N_13890,N_13737,N_13688);
nand U13891 (N_13891,N_13503,N_13639);
and U13892 (N_13892,N_13615,N_13618);
xnor U13893 (N_13893,N_13674,N_13675);
or U13894 (N_13894,N_13713,N_13699);
or U13895 (N_13895,N_13615,N_13745);
nand U13896 (N_13896,N_13733,N_13588);
nand U13897 (N_13897,N_13541,N_13625);
nand U13898 (N_13898,N_13522,N_13602);
or U13899 (N_13899,N_13681,N_13604);
xnor U13900 (N_13900,N_13662,N_13598);
or U13901 (N_13901,N_13529,N_13616);
or U13902 (N_13902,N_13665,N_13660);
nand U13903 (N_13903,N_13682,N_13686);
xnor U13904 (N_13904,N_13585,N_13608);
nor U13905 (N_13905,N_13681,N_13695);
nand U13906 (N_13906,N_13549,N_13532);
and U13907 (N_13907,N_13623,N_13654);
xnor U13908 (N_13908,N_13667,N_13512);
and U13909 (N_13909,N_13588,N_13721);
and U13910 (N_13910,N_13662,N_13569);
or U13911 (N_13911,N_13624,N_13597);
or U13912 (N_13912,N_13673,N_13666);
and U13913 (N_13913,N_13522,N_13519);
nor U13914 (N_13914,N_13531,N_13608);
and U13915 (N_13915,N_13536,N_13508);
xor U13916 (N_13916,N_13547,N_13572);
xor U13917 (N_13917,N_13692,N_13594);
nor U13918 (N_13918,N_13693,N_13544);
or U13919 (N_13919,N_13737,N_13552);
nor U13920 (N_13920,N_13594,N_13556);
nor U13921 (N_13921,N_13733,N_13628);
nand U13922 (N_13922,N_13641,N_13650);
nand U13923 (N_13923,N_13603,N_13709);
or U13924 (N_13924,N_13503,N_13668);
xnor U13925 (N_13925,N_13644,N_13606);
nand U13926 (N_13926,N_13548,N_13518);
nand U13927 (N_13927,N_13605,N_13598);
nor U13928 (N_13928,N_13588,N_13533);
xor U13929 (N_13929,N_13551,N_13687);
and U13930 (N_13930,N_13733,N_13655);
and U13931 (N_13931,N_13629,N_13748);
xor U13932 (N_13932,N_13664,N_13565);
xnor U13933 (N_13933,N_13745,N_13568);
xor U13934 (N_13934,N_13652,N_13710);
or U13935 (N_13935,N_13615,N_13735);
nor U13936 (N_13936,N_13630,N_13657);
nor U13937 (N_13937,N_13621,N_13513);
nor U13938 (N_13938,N_13717,N_13719);
or U13939 (N_13939,N_13748,N_13631);
and U13940 (N_13940,N_13523,N_13577);
xnor U13941 (N_13941,N_13681,N_13667);
or U13942 (N_13942,N_13689,N_13618);
and U13943 (N_13943,N_13645,N_13565);
nor U13944 (N_13944,N_13653,N_13730);
xnor U13945 (N_13945,N_13732,N_13682);
xor U13946 (N_13946,N_13612,N_13723);
nor U13947 (N_13947,N_13744,N_13639);
and U13948 (N_13948,N_13706,N_13595);
xnor U13949 (N_13949,N_13573,N_13743);
or U13950 (N_13950,N_13720,N_13633);
nor U13951 (N_13951,N_13716,N_13678);
nand U13952 (N_13952,N_13510,N_13553);
or U13953 (N_13953,N_13733,N_13626);
xnor U13954 (N_13954,N_13549,N_13566);
nand U13955 (N_13955,N_13516,N_13593);
nor U13956 (N_13956,N_13552,N_13607);
nor U13957 (N_13957,N_13616,N_13739);
or U13958 (N_13958,N_13686,N_13589);
xnor U13959 (N_13959,N_13710,N_13679);
nor U13960 (N_13960,N_13729,N_13693);
and U13961 (N_13961,N_13606,N_13558);
nand U13962 (N_13962,N_13731,N_13630);
nand U13963 (N_13963,N_13649,N_13705);
and U13964 (N_13964,N_13590,N_13586);
or U13965 (N_13965,N_13519,N_13559);
or U13966 (N_13966,N_13554,N_13710);
and U13967 (N_13967,N_13674,N_13528);
xnor U13968 (N_13968,N_13659,N_13621);
xnor U13969 (N_13969,N_13575,N_13719);
and U13970 (N_13970,N_13690,N_13655);
xor U13971 (N_13971,N_13693,N_13638);
or U13972 (N_13972,N_13649,N_13539);
or U13973 (N_13973,N_13715,N_13553);
nor U13974 (N_13974,N_13535,N_13704);
and U13975 (N_13975,N_13545,N_13568);
nand U13976 (N_13976,N_13539,N_13747);
nand U13977 (N_13977,N_13638,N_13548);
nor U13978 (N_13978,N_13689,N_13560);
or U13979 (N_13979,N_13630,N_13555);
and U13980 (N_13980,N_13607,N_13528);
xnor U13981 (N_13981,N_13614,N_13653);
or U13982 (N_13982,N_13521,N_13511);
nand U13983 (N_13983,N_13748,N_13684);
nor U13984 (N_13984,N_13727,N_13743);
xnor U13985 (N_13985,N_13637,N_13683);
xor U13986 (N_13986,N_13601,N_13646);
nor U13987 (N_13987,N_13572,N_13556);
or U13988 (N_13988,N_13679,N_13687);
xor U13989 (N_13989,N_13585,N_13565);
nand U13990 (N_13990,N_13728,N_13515);
and U13991 (N_13991,N_13508,N_13697);
nor U13992 (N_13992,N_13508,N_13599);
or U13993 (N_13993,N_13736,N_13680);
or U13994 (N_13994,N_13749,N_13725);
nor U13995 (N_13995,N_13611,N_13595);
and U13996 (N_13996,N_13510,N_13645);
and U13997 (N_13997,N_13556,N_13526);
and U13998 (N_13998,N_13523,N_13726);
and U13999 (N_13999,N_13672,N_13513);
or U14000 (N_14000,N_13891,N_13890);
nor U14001 (N_14001,N_13866,N_13928);
nor U14002 (N_14002,N_13926,N_13804);
or U14003 (N_14003,N_13852,N_13843);
or U14004 (N_14004,N_13964,N_13805);
nand U14005 (N_14005,N_13946,N_13836);
nor U14006 (N_14006,N_13865,N_13908);
nor U14007 (N_14007,N_13953,N_13932);
nor U14008 (N_14008,N_13832,N_13871);
xnor U14009 (N_14009,N_13905,N_13767);
and U14010 (N_14010,N_13861,N_13800);
or U14011 (N_14011,N_13878,N_13984);
and U14012 (N_14012,N_13787,N_13780);
or U14013 (N_14013,N_13753,N_13825);
xor U14014 (N_14014,N_13976,N_13837);
or U14015 (N_14015,N_13783,N_13988);
and U14016 (N_14016,N_13770,N_13876);
or U14017 (N_14017,N_13824,N_13779);
or U14018 (N_14018,N_13846,N_13809);
nand U14019 (N_14019,N_13808,N_13751);
or U14020 (N_14020,N_13909,N_13991);
nor U14021 (N_14021,N_13790,N_13941);
or U14022 (N_14022,N_13803,N_13955);
or U14023 (N_14023,N_13880,N_13833);
or U14024 (N_14024,N_13918,N_13786);
and U14025 (N_14025,N_13962,N_13872);
xnor U14026 (N_14026,N_13999,N_13792);
or U14027 (N_14027,N_13813,N_13951);
and U14028 (N_14028,N_13914,N_13952);
xor U14029 (N_14029,N_13784,N_13823);
nand U14030 (N_14030,N_13930,N_13933);
or U14031 (N_14031,N_13752,N_13882);
and U14032 (N_14032,N_13993,N_13820);
xnor U14033 (N_14033,N_13750,N_13987);
nor U14034 (N_14034,N_13915,N_13958);
nor U14035 (N_14035,N_13947,N_13996);
nand U14036 (N_14036,N_13769,N_13757);
or U14037 (N_14037,N_13845,N_13887);
or U14038 (N_14038,N_13835,N_13869);
or U14039 (N_14039,N_13791,N_13916);
xor U14040 (N_14040,N_13806,N_13983);
and U14041 (N_14041,N_13898,N_13768);
and U14042 (N_14042,N_13816,N_13998);
xnor U14043 (N_14043,N_13818,N_13885);
nor U14044 (N_14044,N_13756,N_13788);
nand U14045 (N_14045,N_13839,N_13960);
nor U14046 (N_14046,N_13799,N_13797);
and U14047 (N_14047,N_13766,N_13798);
and U14048 (N_14048,N_13877,N_13771);
nor U14049 (N_14049,N_13944,N_13957);
nor U14050 (N_14050,N_13873,N_13919);
or U14051 (N_14051,N_13985,N_13969);
and U14052 (N_14052,N_13764,N_13966);
or U14053 (N_14053,N_13870,N_13795);
nand U14054 (N_14054,N_13826,N_13936);
nand U14055 (N_14055,N_13992,N_13862);
nand U14056 (N_14056,N_13970,N_13886);
nand U14057 (N_14057,N_13989,N_13939);
and U14058 (N_14058,N_13902,N_13945);
and U14059 (N_14059,N_13844,N_13903);
and U14060 (N_14060,N_13828,N_13774);
nand U14061 (N_14061,N_13830,N_13840);
nand U14062 (N_14062,N_13978,N_13785);
nand U14063 (N_14063,N_13973,N_13773);
and U14064 (N_14064,N_13812,N_13807);
xor U14065 (N_14065,N_13810,N_13974);
nor U14066 (N_14066,N_13889,N_13949);
and U14067 (N_14067,N_13943,N_13777);
nand U14068 (N_14068,N_13981,N_13923);
nand U14069 (N_14069,N_13948,N_13847);
nor U14070 (N_14070,N_13831,N_13789);
and U14071 (N_14071,N_13841,N_13879);
nor U14072 (N_14072,N_13971,N_13986);
or U14073 (N_14073,N_13863,N_13796);
or U14074 (N_14074,N_13917,N_13935);
or U14075 (N_14075,N_13778,N_13896);
or U14076 (N_14076,N_13929,N_13821);
nand U14077 (N_14077,N_13811,N_13895);
and U14078 (N_14078,N_13758,N_13963);
xor U14079 (N_14079,N_13848,N_13892);
xor U14080 (N_14080,N_13920,N_13940);
and U14081 (N_14081,N_13829,N_13906);
nor U14082 (N_14082,N_13762,N_13913);
nor U14083 (N_14083,N_13793,N_13858);
nand U14084 (N_14084,N_13893,N_13860);
or U14085 (N_14085,N_13838,N_13781);
xor U14086 (N_14086,N_13997,N_13794);
nand U14087 (N_14087,N_13875,N_13934);
xnor U14088 (N_14088,N_13931,N_13901);
and U14089 (N_14089,N_13888,N_13856);
and U14090 (N_14090,N_13782,N_13965);
nand U14091 (N_14091,N_13763,N_13765);
nor U14092 (N_14092,N_13990,N_13851);
nand U14093 (N_14093,N_13925,N_13859);
nand U14094 (N_14094,N_13822,N_13854);
and U14095 (N_14095,N_13897,N_13883);
and U14096 (N_14096,N_13942,N_13834);
nor U14097 (N_14097,N_13759,N_13853);
nand U14098 (N_14098,N_13775,N_13995);
or U14099 (N_14099,N_13849,N_13954);
or U14100 (N_14100,N_13857,N_13907);
and U14101 (N_14101,N_13904,N_13842);
nor U14102 (N_14102,N_13922,N_13956);
and U14103 (N_14103,N_13761,N_13772);
or U14104 (N_14104,N_13968,N_13801);
nor U14105 (N_14105,N_13924,N_13760);
or U14106 (N_14106,N_13994,N_13921);
nand U14107 (N_14107,N_13864,N_13911);
xor U14108 (N_14108,N_13894,N_13910);
and U14109 (N_14109,N_13900,N_13884);
nand U14110 (N_14110,N_13938,N_13819);
nand U14111 (N_14111,N_13827,N_13817);
nor U14112 (N_14112,N_13980,N_13868);
nor U14113 (N_14113,N_13881,N_13874);
and U14114 (N_14114,N_13815,N_13776);
and U14115 (N_14115,N_13967,N_13982);
nand U14116 (N_14116,N_13979,N_13975);
or U14117 (N_14117,N_13937,N_13754);
and U14118 (N_14118,N_13814,N_13977);
nor U14119 (N_14119,N_13899,N_13959);
and U14120 (N_14120,N_13755,N_13972);
xor U14121 (N_14121,N_13855,N_13850);
or U14122 (N_14122,N_13950,N_13802);
xor U14123 (N_14123,N_13912,N_13867);
nand U14124 (N_14124,N_13927,N_13961);
nand U14125 (N_14125,N_13789,N_13857);
xnor U14126 (N_14126,N_13960,N_13835);
and U14127 (N_14127,N_13824,N_13806);
nand U14128 (N_14128,N_13999,N_13756);
or U14129 (N_14129,N_13774,N_13980);
nand U14130 (N_14130,N_13931,N_13762);
xor U14131 (N_14131,N_13999,N_13774);
and U14132 (N_14132,N_13777,N_13754);
or U14133 (N_14133,N_13806,N_13848);
and U14134 (N_14134,N_13819,N_13923);
nor U14135 (N_14135,N_13966,N_13806);
xnor U14136 (N_14136,N_13911,N_13950);
xnor U14137 (N_14137,N_13838,N_13989);
nand U14138 (N_14138,N_13921,N_13810);
xor U14139 (N_14139,N_13959,N_13977);
nand U14140 (N_14140,N_13887,N_13997);
and U14141 (N_14141,N_13872,N_13929);
nand U14142 (N_14142,N_13835,N_13973);
and U14143 (N_14143,N_13853,N_13911);
and U14144 (N_14144,N_13999,N_13968);
and U14145 (N_14145,N_13803,N_13927);
and U14146 (N_14146,N_13968,N_13888);
xor U14147 (N_14147,N_13922,N_13938);
xor U14148 (N_14148,N_13930,N_13875);
xor U14149 (N_14149,N_13843,N_13763);
xnor U14150 (N_14150,N_13806,N_13852);
or U14151 (N_14151,N_13939,N_13856);
nor U14152 (N_14152,N_13964,N_13811);
or U14153 (N_14153,N_13844,N_13794);
xor U14154 (N_14154,N_13979,N_13818);
or U14155 (N_14155,N_13880,N_13786);
and U14156 (N_14156,N_13885,N_13978);
or U14157 (N_14157,N_13887,N_13865);
nor U14158 (N_14158,N_13929,N_13915);
and U14159 (N_14159,N_13976,N_13884);
nor U14160 (N_14160,N_13914,N_13779);
and U14161 (N_14161,N_13967,N_13780);
or U14162 (N_14162,N_13909,N_13961);
xor U14163 (N_14163,N_13761,N_13964);
nand U14164 (N_14164,N_13808,N_13842);
or U14165 (N_14165,N_13868,N_13869);
xor U14166 (N_14166,N_13960,N_13842);
or U14167 (N_14167,N_13942,N_13789);
or U14168 (N_14168,N_13981,N_13937);
nor U14169 (N_14169,N_13888,N_13862);
xnor U14170 (N_14170,N_13763,N_13906);
and U14171 (N_14171,N_13863,N_13853);
xor U14172 (N_14172,N_13768,N_13926);
and U14173 (N_14173,N_13817,N_13988);
and U14174 (N_14174,N_13992,N_13988);
nand U14175 (N_14175,N_13963,N_13778);
or U14176 (N_14176,N_13872,N_13986);
nor U14177 (N_14177,N_13772,N_13903);
and U14178 (N_14178,N_13956,N_13808);
nand U14179 (N_14179,N_13907,N_13788);
nor U14180 (N_14180,N_13976,N_13821);
and U14181 (N_14181,N_13859,N_13874);
or U14182 (N_14182,N_13979,N_13843);
nor U14183 (N_14183,N_13954,N_13818);
xnor U14184 (N_14184,N_13787,N_13918);
nand U14185 (N_14185,N_13805,N_13861);
and U14186 (N_14186,N_13858,N_13829);
and U14187 (N_14187,N_13923,N_13879);
or U14188 (N_14188,N_13939,N_13992);
or U14189 (N_14189,N_13914,N_13844);
nor U14190 (N_14190,N_13981,N_13803);
nand U14191 (N_14191,N_13864,N_13947);
nand U14192 (N_14192,N_13885,N_13912);
or U14193 (N_14193,N_13982,N_13980);
or U14194 (N_14194,N_13917,N_13919);
and U14195 (N_14195,N_13948,N_13870);
nor U14196 (N_14196,N_13875,N_13757);
nor U14197 (N_14197,N_13827,N_13754);
or U14198 (N_14198,N_13824,N_13786);
nand U14199 (N_14199,N_13781,N_13917);
and U14200 (N_14200,N_13811,N_13922);
or U14201 (N_14201,N_13824,N_13767);
and U14202 (N_14202,N_13936,N_13995);
and U14203 (N_14203,N_13906,N_13800);
xor U14204 (N_14204,N_13817,N_13803);
xor U14205 (N_14205,N_13765,N_13937);
nor U14206 (N_14206,N_13824,N_13762);
nor U14207 (N_14207,N_13897,N_13919);
nor U14208 (N_14208,N_13979,N_13938);
xor U14209 (N_14209,N_13906,N_13891);
and U14210 (N_14210,N_13886,N_13762);
nand U14211 (N_14211,N_13799,N_13783);
or U14212 (N_14212,N_13937,N_13873);
or U14213 (N_14213,N_13765,N_13973);
or U14214 (N_14214,N_13991,N_13855);
or U14215 (N_14215,N_13900,N_13851);
and U14216 (N_14216,N_13823,N_13853);
and U14217 (N_14217,N_13900,N_13868);
nor U14218 (N_14218,N_13850,N_13851);
nand U14219 (N_14219,N_13999,N_13802);
xor U14220 (N_14220,N_13955,N_13911);
or U14221 (N_14221,N_13770,N_13918);
or U14222 (N_14222,N_13973,N_13934);
or U14223 (N_14223,N_13898,N_13991);
or U14224 (N_14224,N_13943,N_13976);
or U14225 (N_14225,N_13799,N_13913);
and U14226 (N_14226,N_13753,N_13823);
or U14227 (N_14227,N_13895,N_13864);
or U14228 (N_14228,N_13972,N_13928);
or U14229 (N_14229,N_13930,N_13937);
nand U14230 (N_14230,N_13934,N_13763);
nand U14231 (N_14231,N_13977,N_13782);
nand U14232 (N_14232,N_13921,N_13968);
nand U14233 (N_14233,N_13880,N_13914);
nand U14234 (N_14234,N_13860,N_13854);
xor U14235 (N_14235,N_13797,N_13764);
xor U14236 (N_14236,N_13888,N_13812);
nor U14237 (N_14237,N_13986,N_13945);
or U14238 (N_14238,N_13893,N_13844);
and U14239 (N_14239,N_13983,N_13965);
xor U14240 (N_14240,N_13912,N_13813);
nor U14241 (N_14241,N_13879,N_13944);
nor U14242 (N_14242,N_13987,N_13817);
nor U14243 (N_14243,N_13872,N_13870);
xnor U14244 (N_14244,N_13801,N_13847);
xor U14245 (N_14245,N_13758,N_13766);
or U14246 (N_14246,N_13902,N_13873);
nor U14247 (N_14247,N_13909,N_13835);
or U14248 (N_14248,N_13945,N_13910);
xnor U14249 (N_14249,N_13923,N_13757);
and U14250 (N_14250,N_14172,N_14146);
or U14251 (N_14251,N_14113,N_14173);
and U14252 (N_14252,N_14137,N_14095);
or U14253 (N_14253,N_14110,N_14241);
nor U14254 (N_14254,N_14231,N_14052);
and U14255 (N_14255,N_14078,N_14029);
nand U14256 (N_14256,N_14125,N_14012);
nand U14257 (N_14257,N_14072,N_14120);
nand U14258 (N_14258,N_14077,N_14067);
xor U14259 (N_14259,N_14188,N_14183);
nor U14260 (N_14260,N_14056,N_14061);
nand U14261 (N_14261,N_14036,N_14060);
xnor U14262 (N_14262,N_14090,N_14022);
nor U14263 (N_14263,N_14082,N_14195);
or U14264 (N_14264,N_14074,N_14218);
nor U14265 (N_14265,N_14084,N_14194);
nor U14266 (N_14266,N_14073,N_14122);
and U14267 (N_14267,N_14013,N_14203);
or U14268 (N_14268,N_14180,N_14225);
nor U14269 (N_14269,N_14049,N_14042);
and U14270 (N_14270,N_14004,N_14031);
xor U14271 (N_14271,N_14071,N_14069);
nor U14272 (N_14272,N_14002,N_14210);
nand U14273 (N_14273,N_14048,N_14102);
nor U14274 (N_14274,N_14000,N_14026);
xnor U14275 (N_14275,N_14123,N_14010);
or U14276 (N_14276,N_14190,N_14141);
xnor U14277 (N_14277,N_14205,N_14015);
nor U14278 (N_14278,N_14237,N_14175);
nor U14279 (N_14279,N_14089,N_14181);
nor U14280 (N_14280,N_14219,N_14033);
or U14281 (N_14281,N_14213,N_14105);
and U14282 (N_14282,N_14150,N_14126);
or U14283 (N_14283,N_14005,N_14234);
xor U14284 (N_14284,N_14116,N_14041);
xor U14285 (N_14285,N_14206,N_14235);
and U14286 (N_14286,N_14130,N_14151);
and U14287 (N_14287,N_14001,N_14006);
and U14288 (N_14288,N_14230,N_14014);
nand U14289 (N_14289,N_14220,N_14139);
nand U14290 (N_14290,N_14112,N_14140);
xor U14291 (N_14291,N_14035,N_14045);
xnor U14292 (N_14292,N_14059,N_14162);
nor U14293 (N_14293,N_14008,N_14103);
xor U14294 (N_14294,N_14009,N_14228);
and U14295 (N_14295,N_14243,N_14065);
and U14296 (N_14296,N_14003,N_14165);
nand U14297 (N_14297,N_14104,N_14158);
and U14298 (N_14298,N_14196,N_14199);
nor U14299 (N_14299,N_14136,N_14086);
and U14300 (N_14300,N_14092,N_14053);
or U14301 (N_14301,N_14211,N_14197);
nand U14302 (N_14302,N_14046,N_14083);
xor U14303 (N_14303,N_14020,N_14106);
xor U14304 (N_14304,N_14244,N_14186);
or U14305 (N_14305,N_14249,N_14018);
and U14306 (N_14306,N_14027,N_14118);
nand U14307 (N_14307,N_14044,N_14128);
and U14308 (N_14308,N_14093,N_14233);
and U14309 (N_14309,N_14221,N_14057);
xor U14310 (N_14310,N_14238,N_14142);
nand U14311 (N_14311,N_14214,N_14064);
and U14312 (N_14312,N_14117,N_14163);
and U14313 (N_14313,N_14179,N_14068);
nor U14314 (N_14314,N_14070,N_14215);
and U14315 (N_14315,N_14127,N_14058);
and U14316 (N_14316,N_14170,N_14157);
nor U14317 (N_14317,N_14075,N_14138);
nand U14318 (N_14318,N_14025,N_14066);
xor U14319 (N_14319,N_14019,N_14246);
nand U14320 (N_14320,N_14047,N_14200);
and U14321 (N_14321,N_14152,N_14182);
or U14322 (N_14322,N_14201,N_14017);
xnor U14323 (N_14323,N_14129,N_14164);
nor U14324 (N_14324,N_14007,N_14087);
nor U14325 (N_14325,N_14242,N_14147);
and U14326 (N_14326,N_14155,N_14111);
or U14327 (N_14327,N_14134,N_14209);
and U14328 (N_14328,N_14156,N_14034);
and U14329 (N_14329,N_14132,N_14154);
nand U14330 (N_14330,N_14216,N_14198);
or U14331 (N_14331,N_14232,N_14101);
or U14332 (N_14332,N_14133,N_14114);
xnor U14333 (N_14333,N_14098,N_14051);
or U14334 (N_14334,N_14021,N_14148);
or U14335 (N_14335,N_14245,N_14174);
nor U14336 (N_14336,N_14191,N_14167);
nand U14337 (N_14337,N_14217,N_14176);
or U14338 (N_14338,N_14161,N_14109);
and U14339 (N_14339,N_14159,N_14085);
or U14340 (N_14340,N_14032,N_14171);
and U14341 (N_14341,N_14193,N_14229);
xnor U14342 (N_14342,N_14227,N_14119);
or U14343 (N_14343,N_14011,N_14121);
xnor U14344 (N_14344,N_14094,N_14208);
or U14345 (N_14345,N_14043,N_14160);
nand U14346 (N_14346,N_14039,N_14131);
and U14347 (N_14347,N_14076,N_14149);
nand U14348 (N_14348,N_14189,N_14038);
and U14349 (N_14349,N_14055,N_14023);
xor U14350 (N_14350,N_14050,N_14178);
xor U14351 (N_14351,N_14124,N_14212);
nor U14352 (N_14352,N_14016,N_14081);
nor U14353 (N_14353,N_14040,N_14239);
or U14354 (N_14354,N_14115,N_14240);
or U14355 (N_14355,N_14028,N_14145);
or U14356 (N_14356,N_14107,N_14192);
or U14357 (N_14357,N_14024,N_14100);
xnor U14358 (N_14358,N_14226,N_14247);
xor U14359 (N_14359,N_14202,N_14187);
or U14360 (N_14360,N_14222,N_14063);
and U14361 (N_14361,N_14166,N_14099);
and U14362 (N_14362,N_14062,N_14079);
xnor U14363 (N_14363,N_14054,N_14088);
nor U14364 (N_14364,N_14108,N_14144);
and U14365 (N_14365,N_14236,N_14096);
nor U14366 (N_14366,N_14097,N_14135);
and U14367 (N_14367,N_14080,N_14223);
nor U14368 (N_14368,N_14177,N_14184);
nand U14369 (N_14369,N_14168,N_14143);
and U14370 (N_14370,N_14207,N_14224);
xor U14371 (N_14371,N_14169,N_14204);
and U14372 (N_14372,N_14030,N_14091);
and U14373 (N_14373,N_14037,N_14153);
nor U14374 (N_14374,N_14248,N_14185);
nand U14375 (N_14375,N_14156,N_14246);
xnor U14376 (N_14376,N_14018,N_14236);
and U14377 (N_14377,N_14082,N_14090);
or U14378 (N_14378,N_14247,N_14097);
and U14379 (N_14379,N_14168,N_14163);
and U14380 (N_14380,N_14198,N_14044);
and U14381 (N_14381,N_14224,N_14123);
or U14382 (N_14382,N_14203,N_14170);
and U14383 (N_14383,N_14055,N_14240);
nand U14384 (N_14384,N_14151,N_14080);
nand U14385 (N_14385,N_14117,N_14194);
xnor U14386 (N_14386,N_14121,N_14088);
nor U14387 (N_14387,N_14173,N_14145);
or U14388 (N_14388,N_14157,N_14080);
and U14389 (N_14389,N_14245,N_14223);
and U14390 (N_14390,N_14071,N_14010);
and U14391 (N_14391,N_14230,N_14054);
xor U14392 (N_14392,N_14056,N_14149);
nor U14393 (N_14393,N_14097,N_14090);
nor U14394 (N_14394,N_14083,N_14066);
xnor U14395 (N_14395,N_14005,N_14204);
and U14396 (N_14396,N_14216,N_14137);
and U14397 (N_14397,N_14078,N_14022);
and U14398 (N_14398,N_14102,N_14165);
xnor U14399 (N_14399,N_14204,N_14110);
xnor U14400 (N_14400,N_14156,N_14152);
nor U14401 (N_14401,N_14060,N_14186);
or U14402 (N_14402,N_14084,N_14141);
nand U14403 (N_14403,N_14035,N_14230);
and U14404 (N_14404,N_14168,N_14026);
and U14405 (N_14405,N_14180,N_14077);
and U14406 (N_14406,N_14238,N_14205);
nand U14407 (N_14407,N_14102,N_14099);
nor U14408 (N_14408,N_14207,N_14129);
and U14409 (N_14409,N_14139,N_14108);
xor U14410 (N_14410,N_14136,N_14175);
xor U14411 (N_14411,N_14046,N_14094);
and U14412 (N_14412,N_14118,N_14192);
xnor U14413 (N_14413,N_14184,N_14013);
or U14414 (N_14414,N_14223,N_14133);
or U14415 (N_14415,N_14049,N_14090);
nand U14416 (N_14416,N_14109,N_14088);
and U14417 (N_14417,N_14153,N_14239);
or U14418 (N_14418,N_14050,N_14170);
nand U14419 (N_14419,N_14026,N_14212);
nand U14420 (N_14420,N_14238,N_14154);
nand U14421 (N_14421,N_14229,N_14083);
or U14422 (N_14422,N_14063,N_14093);
nand U14423 (N_14423,N_14099,N_14119);
nand U14424 (N_14424,N_14058,N_14193);
xnor U14425 (N_14425,N_14158,N_14091);
nor U14426 (N_14426,N_14216,N_14236);
nor U14427 (N_14427,N_14061,N_14069);
and U14428 (N_14428,N_14041,N_14227);
nand U14429 (N_14429,N_14098,N_14017);
nand U14430 (N_14430,N_14208,N_14198);
nand U14431 (N_14431,N_14184,N_14236);
xor U14432 (N_14432,N_14084,N_14105);
and U14433 (N_14433,N_14123,N_14132);
xnor U14434 (N_14434,N_14153,N_14005);
or U14435 (N_14435,N_14158,N_14176);
nor U14436 (N_14436,N_14235,N_14116);
or U14437 (N_14437,N_14120,N_14067);
nand U14438 (N_14438,N_14160,N_14207);
and U14439 (N_14439,N_14203,N_14112);
nand U14440 (N_14440,N_14156,N_14056);
xnor U14441 (N_14441,N_14138,N_14201);
nand U14442 (N_14442,N_14188,N_14174);
xnor U14443 (N_14443,N_14143,N_14041);
or U14444 (N_14444,N_14067,N_14116);
or U14445 (N_14445,N_14049,N_14074);
nor U14446 (N_14446,N_14011,N_14239);
or U14447 (N_14447,N_14107,N_14023);
nor U14448 (N_14448,N_14113,N_14084);
and U14449 (N_14449,N_14183,N_14012);
nor U14450 (N_14450,N_14086,N_14057);
nor U14451 (N_14451,N_14012,N_14080);
or U14452 (N_14452,N_14118,N_14130);
xnor U14453 (N_14453,N_14185,N_14088);
nand U14454 (N_14454,N_14217,N_14137);
and U14455 (N_14455,N_14135,N_14027);
or U14456 (N_14456,N_14235,N_14031);
nand U14457 (N_14457,N_14173,N_14011);
or U14458 (N_14458,N_14129,N_14136);
nor U14459 (N_14459,N_14027,N_14162);
nand U14460 (N_14460,N_14242,N_14155);
nand U14461 (N_14461,N_14027,N_14193);
nand U14462 (N_14462,N_14239,N_14211);
nand U14463 (N_14463,N_14118,N_14098);
and U14464 (N_14464,N_14202,N_14167);
xnor U14465 (N_14465,N_14192,N_14076);
or U14466 (N_14466,N_14216,N_14174);
xnor U14467 (N_14467,N_14008,N_14107);
xnor U14468 (N_14468,N_14214,N_14023);
xnor U14469 (N_14469,N_14029,N_14214);
and U14470 (N_14470,N_14055,N_14109);
and U14471 (N_14471,N_14179,N_14111);
or U14472 (N_14472,N_14180,N_14212);
nand U14473 (N_14473,N_14189,N_14044);
or U14474 (N_14474,N_14096,N_14114);
and U14475 (N_14475,N_14216,N_14066);
nor U14476 (N_14476,N_14200,N_14165);
nand U14477 (N_14477,N_14125,N_14165);
and U14478 (N_14478,N_14044,N_14203);
or U14479 (N_14479,N_14174,N_14004);
and U14480 (N_14480,N_14200,N_14020);
and U14481 (N_14481,N_14041,N_14104);
nor U14482 (N_14482,N_14188,N_14197);
or U14483 (N_14483,N_14113,N_14169);
and U14484 (N_14484,N_14024,N_14063);
and U14485 (N_14485,N_14182,N_14042);
nand U14486 (N_14486,N_14068,N_14149);
xor U14487 (N_14487,N_14084,N_14211);
nor U14488 (N_14488,N_14058,N_14136);
xor U14489 (N_14489,N_14212,N_14017);
nor U14490 (N_14490,N_14082,N_14154);
xnor U14491 (N_14491,N_14137,N_14229);
nand U14492 (N_14492,N_14242,N_14065);
nor U14493 (N_14493,N_14071,N_14074);
nor U14494 (N_14494,N_14156,N_14123);
nor U14495 (N_14495,N_14229,N_14152);
or U14496 (N_14496,N_14079,N_14213);
nor U14497 (N_14497,N_14016,N_14064);
and U14498 (N_14498,N_14148,N_14166);
xor U14499 (N_14499,N_14038,N_14072);
nor U14500 (N_14500,N_14454,N_14475);
and U14501 (N_14501,N_14344,N_14402);
or U14502 (N_14502,N_14488,N_14290);
and U14503 (N_14503,N_14367,N_14285);
and U14504 (N_14504,N_14343,N_14419);
and U14505 (N_14505,N_14494,N_14336);
nor U14506 (N_14506,N_14469,N_14349);
nand U14507 (N_14507,N_14445,N_14281);
and U14508 (N_14508,N_14371,N_14376);
nand U14509 (N_14509,N_14356,N_14299);
and U14510 (N_14510,N_14252,N_14312);
xor U14511 (N_14511,N_14263,N_14490);
nand U14512 (N_14512,N_14325,N_14401);
nand U14513 (N_14513,N_14258,N_14482);
nand U14514 (N_14514,N_14364,N_14440);
nor U14515 (N_14515,N_14394,N_14462);
and U14516 (N_14516,N_14363,N_14493);
xnor U14517 (N_14517,N_14470,N_14451);
and U14518 (N_14518,N_14426,N_14448);
xnor U14519 (N_14519,N_14381,N_14305);
or U14520 (N_14520,N_14329,N_14268);
or U14521 (N_14521,N_14358,N_14428);
and U14522 (N_14522,N_14279,N_14480);
nand U14523 (N_14523,N_14301,N_14271);
nand U14524 (N_14524,N_14395,N_14377);
nor U14525 (N_14525,N_14266,N_14277);
and U14526 (N_14526,N_14257,N_14467);
nand U14527 (N_14527,N_14284,N_14437);
nor U14528 (N_14528,N_14471,N_14452);
xnor U14529 (N_14529,N_14276,N_14302);
and U14530 (N_14530,N_14303,N_14286);
xor U14531 (N_14531,N_14464,N_14479);
and U14532 (N_14532,N_14379,N_14444);
xor U14533 (N_14533,N_14337,N_14365);
or U14534 (N_14534,N_14251,N_14407);
nor U14535 (N_14535,N_14422,N_14412);
and U14536 (N_14536,N_14273,N_14439);
nand U14537 (N_14537,N_14399,N_14347);
and U14538 (N_14538,N_14413,N_14432);
nand U14539 (N_14539,N_14418,N_14322);
nand U14540 (N_14540,N_14430,N_14373);
and U14541 (N_14541,N_14361,N_14328);
xnor U14542 (N_14542,N_14455,N_14438);
and U14543 (N_14543,N_14380,N_14435);
xor U14544 (N_14544,N_14282,N_14450);
and U14545 (N_14545,N_14264,N_14311);
and U14546 (N_14546,N_14324,N_14459);
xor U14547 (N_14547,N_14352,N_14476);
xor U14548 (N_14548,N_14259,N_14278);
xor U14549 (N_14549,N_14421,N_14327);
nand U14550 (N_14550,N_14353,N_14404);
and U14551 (N_14551,N_14387,N_14355);
or U14552 (N_14552,N_14345,N_14292);
nand U14553 (N_14553,N_14431,N_14420);
or U14554 (N_14554,N_14314,N_14427);
xnor U14555 (N_14555,N_14487,N_14293);
nor U14556 (N_14556,N_14375,N_14335);
nand U14557 (N_14557,N_14400,N_14256);
or U14558 (N_14558,N_14331,N_14318);
xnor U14559 (N_14559,N_14499,N_14265);
and U14560 (N_14560,N_14489,N_14348);
and U14561 (N_14561,N_14386,N_14274);
xnor U14562 (N_14562,N_14463,N_14416);
nor U14563 (N_14563,N_14410,N_14270);
nand U14564 (N_14564,N_14283,N_14309);
xnor U14565 (N_14565,N_14370,N_14457);
xnor U14566 (N_14566,N_14374,N_14313);
nand U14567 (N_14567,N_14368,N_14483);
xor U14568 (N_14568,N_14306,N_14403);
and U14569 (N_14569,N_14486,N_14316);
xor U14570 (N_14570,N_14498,N_14398);
nor U14571 (N_14571,N_14288,N_14425);
and U14572 (N_14572,N_14287,N_14497);
or U14573 (N_14573,N_14472,N_14423);
xnor U14574 (N_14574,N_14289,N_14466);
or U14575 (N_14575,N_14384,N_14275);
or U14576 (N_14576,N_14492,N_14383);
xnor U14577 (N_14577,N_14291,N_14414);
xnor U14578 (N_14578,N_14388,N_14272);
and U14579 (N_14579,N_14392,N_14350);
and U14580 (N_14580,N_14474,N_14409);
nand U14581 (N_14581,N_14389,N_14447);
or U14582 (N_14582,N_14405,N_14393);
nor U14583 (N_14583,N_14468,N_14304);
nor U14584 (N_14584,N_14296,N_14397);
xnor U14585 (N_14585,N_14346,N_14340);
xnor U14586 (N_14586,N_14357,N_14481);
xor U14587 (N_14587,N_14330,N_14320);
xor U14588 (N_14588,N_14477,N_14441);
and U14589 (N_14589,N_14267,N_14326);
nor U14590 (N_14590,N_14323,N_14443);
and U14591 (N_14591,N_14382,N_14369);
nand U14592 (N_14592,N_14446,N_14429);
nand U14593 (N_14593,N_14449,N_14351);
nand U14594 (N_14594,N_14461,N_14261);
xnor U14595 (N_14595,N_14411,N_14342);
nand U14596 (N_14596,N_14396,N_14436);
xor U14597 (N_14597,N_14255,N_14473);
xor U14598 (N_14598,N_14300,N_14298);
nor U14599 (N_14599,N_14310,N_14360);
nand U14600 (N_14600,N_14317,N_14491);
or U14601 (N_14601,N_14495,N_14253);
or U14602 (N_14602,N_14294,N_14391);
or U14603 (N_14603,N_14442,N_14372);
nor U14604 (N_14604,N_14339,N_14297);
nand U14605 (N_14605,N_14434,N_14460);
nor U14606 (N_14606,N_14250,N_14308);
nand U14607 (N_14607,N_14260,N_14307);
nor U14608 (N_14608,N_14378,N_14332);
or U14609 (N_14609,N_14319,N_14354);
nor U14610 (N_14610,N_14496,N_14366);
xnor U14611 (N_14611,N_14390,N_14295);
xnor U14612 (N_14612,N_14456,N_14362);
nand U14613 (N_14613,N_14359,N_14485);
or U14614 (N_14614,N_14458,N_14269);
nor U14615 (N_14615,N_14338,N_14417);
or U14616 (N_14616,N_14321,N_14262);
or U14617 (N_14617,N_14280,N_14406);
nand U14618 (N_14618,N_14408,N_14478);
or U14619 (N_14619,N_14433,N_14315);
xor U14620 (N_14620,N_14333,N_14453);
nor U14621 (N_14621,N_14424,N_14385);
xor U14622 (N_14622,N_14415,N_14341);
xor U14623 (N_14623,N_14465,N_14484);
xor U14624 (N_14624,N_14254,N_14334);
or U14625 (N_14625,N_14298,N_14332);
nand U14626 (N_14626,N_14444,N_14456);
nor U14627 (N_14627,N_14253,N_14297);
xnor U14628 (N_14628,N_14446,N_14408);
or U14629 (N_14629,N_14277,N_14430);
xor U14630 (N_14630,N_14303,N_14351);
or U14631 (N_14631,N_14354,N_14379);
nor U14632 (N_14632,N_14292,N_14497);
or U14633 (N_14633,N_14298,N_14486);
xnor U14634 (N_14634,N_14384,N_14264);
and U14635 (N_14635,N_14440,N_14482);
and U14636 (N_14636,N_14253,N_14386);
nand U14637 (N_14637,N_14453,N_14268);
and U14638 (N_14638,N_14418,N_14292);
nand U14639 (N_14639,N_14335,N_14497);
and U14640 (N_14640,N_14463,N_14292);
xnor U14641 (N_14641,N_14283,N_14364);
xor U14642 (N_14642,N_14456,N_14295);
and U14643 (N_14643,N_14484,N_14371);
xnor U14644 (N_14644,N_14340,N_14254);
nor U14645 (N_14645,N_14411,N_14266);
and U14646 (N_14646,N_14252,N_14417);
or U14647 (N_14647,N_14271,N_14264);
xor U14648 (N_14648,N_14449,N_14258);
and U14649 (N_14649,N_14286,N_14298);
xnor U14650 (N_14650,N_14391,N_14434);
or U14651 (N_14651,N_14375,N_14490);
xor U14652 (N_14652,N_14402,N_14323);
or U14653 (N_14653,N_14445,N_14432);
nor U14654 (N_14654,N_14316,N_14496);
and U14655 (N_14655,N_14398,N_14393);
xnor U14656 (N_14656,N_14453,N_14370);
and U14657 (N_14657,N_14334,N_14373);
or U14658 (N_14658,N_14352,N_14443);
xnor U14659 (N_14659,N_14440,N_14316);
nand U14660 (N_14660,N_14316,N_14428);
and U14661 (N_14661,N_14317,N_14313);
and U14662 (N_14662,N_14458,N_14261);
xnor U14663 (N_14663,N_14359,N_14477);
nand U14664 (N_14664,N_14404,N_14482);
and U14665 (N_14665,N_14329,N_14292);
xnor U14666 (N_14666,N_14404,N_14441);
xor U14667 (N_14667,N_14316,N_14434);
or U14668 (N_14668,N_14442,N_14331);
xor U14669 (N_14669,N_14484,N_14451);
nand U14670 (N_14670,N_14496,N_14256);
nand U14671 (N_14671,N_14279,N_14387);
and U14672 (N_14672,N_14493,N_14421);
or U14673 (N_14673,N_14417,N_14379);
nand U14674 (N_14674,N_14371,N_14444);
nor U14675 (N_14675,N_14277,N_14414);
and U14676 (N_14676,N_14428,N_14435);
nor U14677 (N_14677,N_14405,N_14387);
and U14678 (N_14678,N_14284,N_14391);
and U14679 (N_14679,N_14282,N_14298);
xnor U14680 (N_14680,N_14444,N_14398);
nand U14681 (N_14681,N_14319,N_14470);
xnor U14682 (N_14682,N_14351,N_14364);
or U14683 (N_14683,N_14438,N_14341);
nor U14684 (N_14684,N_14468,N_14315);
and U14685 (N_14685,N_14298,N_14420);
or U14686 (N_14686,N_14299,N_14448);
and U14687 (N_14687,N_14395,N_14487);
nand U14688 (N_14688,N_14398,N_14310);
nor U14689 (N_14689,N_14363,N_14326);
and U14690 (N_14690,N_14261,N_14298);
and U14691 (N_14691,N_14416,N_14408);
nor U14692 (N_14692,N_14350,N_14405);
and U14693 (N_14693,N_14306,N_14494);
and U14694 (N_14694,N_14487,N_14319);
nor U14695 (N_14695,N_14251,N_14426);
and U14696 (N_14696,N_14396,N_14418);
xnor U14697 (N_14697,N_14472,N_14377);
and U14698 (N_14698,N_14317,N_14459);
xor U14699 (N_14699,N_14398,N_14442);
and U14700 (N_14700,N_14461,N_14370);
and U14701 (N_14701,N_14352,N_14454);
and U14702 (N_14702,N_14257,N_14267);
xor U14703 (N_14703,N_14402,N_14358);
nor U14704 (N_14704,N_14366,N_14266);
xor U14705 (N_14705,N_14366,N_14359);
nand U14706 (N_14706,N_14293,N_14327);
nand U14707 (N_14707,N_14496,N_14328);
nor U14708 (N_14708,N_14417,N_14497);
or U14709 (N_14709,N_14380,N_14287);
and U14710 (N_14710,N_14444,N_14307);
xnor U14711 (N_14711,N_14372,N_14409);
and U14712 (N_14712,N_14497,N_14493);
and U14713 (N_14713,N_14446,N_14454);
or U14714 (N_14714,N_14262,N_14492);
and U14715 (N_14715,N_14392,N_14366);
and U14716 (N_14716,N_14387,N_14291);
xnor U14717 (N_14717,N_14489,N_14270);
or U14718 (N_14718,N_14322,N_14265);
or U14719 (N_14719,N_14415,N_14423);
xnor U14720 (N_14720,N_14451,N_14276);
nor U14721 (N_14721,N_14263,N_14363);
nor U14722 (N_14722,N_14452,N_14365);
and U14723 (N_14723,N_14309,N_14440);
or U14724 (N_14724,N_14399,N_14356);
and U14725 (N_14725,N_14312,N_14319);
and U14726 (N_14726,N_14482,N_14323);
nor U14727 (N_14727,N_14270,N_14265);
or U14728 (N_14728,N_14273,N_14331);
xnor U14729 (N_14729,N_14304,N_14394);
or U14730 (N_14730,N_14279,N_14255);
and U14731 (N_14731,N_14338,N_14499);
or U14732 (N_14732,N_14444,N_14323);
nand U14733 (N_14733,N_14277,N_14390);
nor U14734 (N_14734,N_14403,N_14441);
xnor U14735 (N_14735,N_14458,N_14253);
or U14736 (N_14736,N_14424,N_14475);
and U14737 (N_14737,N_14279,N_14482);
nand U14738 (N_14738,N_14253,N_14258);
nand U14739 (N_14739,N_14412,N_14473);
nand U14740 (N_14740,N_14330,N_14380);
nand U14741 (N_14741,N_14494,N_14344);
or U14742 (N_14742,N_14372,N_14472);
or U14743 (N_14743,N_14324,N_14290);
nand U14744 (N_14744,N_14326,N_14295);
nand U14745 (N_14745,N_14408,N_14345);
or U14746 (N_14746,N_14391,N_14361);
and U14747 (N_14747,N_14311,N_14251);
and U14748 (N_14748,N_14413,N_14388);
and U14749 (N_14749,N_14394,N_14251);
and U14750 (N_14750,N_14735,N_14503);
nor U14751 (N_14751,N_14719,N_14553);
nor U14752 (N_14752,N_14738,N_14641);
and U14753 (N_14753,N_14561,N_14565);
xnor U14754 (N_14754,N_14713,N_14642);
nor U14755 (N_14755,N_14726,N_14661);
or U14756 (N_14756,N_14607,N_14551);
nor U14757 (N_14757,N_14519,N_14574);
or U14758 (N_14758,N_14695,N_14690);
or U14759 (N_14759,N_14680,N_14567);
nor U14760 (N_14760,N_14688,N_14527);
nand U14761 (N_14761,N_14742,N_14546);
or U14762 (N_14762,N_14717,N_14655);
or U14763 (N_14763,N_14564,N_14727);
and U14764 (N_14764,N_14517,N_14600);
nor U14765 (N_14765,N_14530,N_14671);
nor U14766 (N_14766,N_14591,N_14711);
or U14767 (N_14767,N_14692,N_14634);
and U14768 (N_14768,N_14595,N_14603);
nand U14769 (N_14769,N_14552,N_14525);
xor U14770 (N_14770,N_14572,N_14612);
or U14771 (N_14771,N_14656,N_14507);
or U14772 (N_14772,N_14628,N_14644);
or U14773 (N_14773,N_14532,N_14544);
xnor U14774 (N_14774,N_14737,N_14508);
or U14775 (N_14775,N_14531,N_14706);
nor U14776 (N_14776,N_14685,N_14588);
and U14777 (N_14777,N_14635,N_14645);
nor U14778 (N_14778,N_14667,N_14707);
nor U14779 (N_14779,N_14675,N_14580);
nand U14780 (N_14780,N_14709,N_14678);
xnor U14781 (N_14781,N_14749,N_14657);
nand U14782 (N_14782,N_14577,N_14631);
or U14783 (N_14783,N_14558,N_14683);
nand U14784 (N_14784,N_14734,N_14694);
and U14785 (N_14785,N_14523,N_14528);
xor U14786 (N_14786,N_14677,N_14629);
xnor U14787 (N_14787,N_14548,N_14723);
or U14788 (N_14788,N_14718,N_14616);
and U14789 (N_14789,N_14543,N_14573);
xor U14790 (N_14790,N_14696,N_14686);
nand U14791 (N_14791,N_14668,N_14609);
nor U14792 (N_14792,N_14584,N_14672);
and U14793 (N_14793,N_14556,N_14563);
xnor U14794 (N_14794,N_14619,N_14625);
nor U14795 (N_14795,N_14559,N_14663);
xor U14796 (N_14796,N_14520,N_14693);
xnor U14797 (N_14797,N_14557,N_14512);
or U14798 (N_14798,N_14585,N_14647);
and U14799 (N_14799,N_14592,N_14502);
nor U14800 (N_14800,N_14504,N_14540);
nand U14801 (N_14801,N_14599,N_14582);
xor U14802 (N_14802,N_14575,N_14526);
and U14803 (N_14803,N_14571,N_14511);
nand U14804 (N_14804,N_14566,N_14699);
and U14805 (N_14805,N_14681,N_14715);
nand U14806 (N_14806,N_14518,N_14513);
nor U14807 (N_14807,N_14596,N_14716);
or U14808 (N_14808,N_14550,N_14691);
xor U14809 (N_14809,N_14714,N_14722);
or U14810 (N_14810,N_14594,N_14622);
nor U14811 (N_14811,N_14748,N_14606);
and U14812 (N_14812,N_14746,N_14537);
or U14813 (N_14813,N_14669,N_14665);
nand U14814 (N_14814,N_14682,N_14515);
or U14815 (N_14815,N_14636,N_14620);
nor U14816 (N_14816,N_14666,N_14651);
nand U14817 (N_14817,N_14615,N_14679);
xnor U14818 (N_14818,N_14522,N_14664);
or U14819 (N_14819,N_14587,N_14674);
nand U14820 (N_14820,N_14649,N_14630);
nor U14821 (N_14821,N_14633,N_14611);
and U14822 (N_14822,N_14662,N_14617);
nand U14823 (N_14823,N_14562,N_14560);
nand U14824 (N_14824,N_14654,N_14684);
nand U14825 (N_14825,N_14741,N_14621);
and U14826 (N_14826,N_14624,N_14689);
nand U14827 (N_14827,N_14730,N_14704);
nor U14828 (N_14828,N_14618,N_14632);
and U14829 (N_14829,N_14712,N_14589);
nor U14830 (N_14830,N_14524,N_14676);
or U14831 (N_14831,N_14658,N_14578);
or U14832 (N_14832,N_14613,N_14729);
xor U14833 (N_14833,N_14660,N_14721);
nand U14834 (N_14834,N_14602,N_14739);
and U14835 (N_14835,N_14733,N_14501);
and U14836 (N_14836,N_14538,N_14701);
and U14837 (N_14837,N_14627,N_14601);
and U14838 (N_14838,N_14509,N_14743);
nand U14839 (N_14839,N_14576,N_14541);
xnor U14840 (N_14840,N_14597,N_14650);
xor U14841 (N_14841,N_14614,N_14605);
nor U14842 (N_14842,N_14581,N_14623);
and U14843 (N_14843,N_14736,N_14542);
xor U14844 (N_14844,N_14539,N_14731);
and U14845 (N_14845,N_14700,N_14516);
nor U14846 (N_14846,N_14579,N_14593);
nor U14847 (N_14847,N_14568,N_14640);
nor U14848 (N_14848,N_14514,N_14708);
nor U14849 (N_14849,N_14653,N_14652);
nor U14850 (N_14850,N_14670,N_14724);
and U14851 (N_14851,N_14554,N_14745);
xor U14852 (N_14852,N_14626,N_14646);
or U14853 (N_14853,N_14702,N_14710);
xor U14854 (N_14854,N_14535,N_14648);
or U14855 (N_14855,N_14705,N_14569);
or U14856 (N_14856,N_14697,N_14604);
and U14857 (N_14857,N_14590,N_14728);
and U14858 (N_14858,N_14639,N_14570);
nor U14859 (N_14859,N_14643,N_14506);
and U14860 (N_14860,N_14740,N_14545);
nand U14861 (N_14861,N_14610,N_14698);
xnor U14862 (N_14862,N_14549,N_14687);
xnor U14863 (N_14863,N_14521,N_14547);
nor U14864 (N_14864,N_14533,N_14586);
and U14865 (N_14865,N_14505,N_14725);
and U14866 (N_14866,N_14598,N_14637);
nor U14867 (N_14867,N_14529,N_14555);
and U14868 (N_14868,N_14583,N_14744);
or U14869 (N_14869,N_14732,N_14747);
nand U14870 (N_14870,N_14720,N_14673);
xnor U14871 (N_14871,N_14500,N_14703);
xnor U14872 (N_14872,N_14659,N_14638);
and U14873 (N_14873,N_14608,N_14536);
and U14874 (N_14874,N_14534,N_14510);
nor U14875 (N_14875,N_14628,N_14745);
xor U14876 (N_14876,N_14604,N_14600);
nor U14877 (N_14877,N_14557,N_14509);
and U14878 (N_14878,N_14607,N_14615);
xor U14879 (N_14879,N_14583,N_14685);
and U14880 (N_14880,N_14717,N_14730);
or U14881 (N_14881,N_14653,N_14501);
nand U14882 (N_14882,N_14656,N_14708);
and U14883 (N_14883,N_14500,N_14639);
xnor U14884 (N_14884,N_14520,N_14551);
or U14885 (N_14885,N_14526,N_14711);
or U14886 (N_14886,N_14699,N_14507);
or U14887 (N_14887,N_14517,N_14644);
or U14888 (N_14888,N_14593,N_14515);
nand U14889 (N_14889,N_14692,N_14680);
or U14890 (N_14890,N_14598,N_14666);
xor U14891 (N_14891,N_14632,N_14583);
or U14892 (N_14892,N_14522,N_14623);
and U14893 (N_14893,N_14634,N_14622);
and U14894 (N_14894,N_14645,N_14736);
nor U14895 (N_14895,N_14674,N_14513);
or U14896 (N_14896,N_14553,N_14680);
nand U14897 (N_14897,N_14518,N_14600);
nand U14898 (N_14898,N_14553,N_14696);
xnor U14899 (N_14899,N_14566,N_14561);
nor U14900 (N_14900,N_14595,N_14617);
nor U14901 (N_14901,N_14684,N_14511);
nand U14902 (N_14902,N_14565,N_14682);
or U14903 (N_14903,N_14612,N_14607);
and U14904 (N_14904,N_14578,N_14613);
nor U14905 (N_14905,N_14635,N_14695);
nand U14906 (N_14906,N_14685,N_14557);
xnor U14907 (N_14907,N_14609,N_14582);
xor U14908 (N_14908,N_14588,N_14501);
or U14909 (N_14909,N_14536,N_14724);
or U14910 (N_14910,N_14511,N_14533);
nor U14911 (N_14911,N_14674,N_14740);
nor U14912 (N_14912,N_14747,N_14557);
nor U14913 (N_14913,N_14566,N_14546);
nand U14914 (N_14914,N_14665,N_14673);
and U14915 (N_14915,N_14599,N_14625);
and U14916 (N_14916,N_14535,N_14517);
or U14917 (N_14917,N_14599,N_14742);
nor U14918 (N_14918,N_14650,N_14525);
or U14919 (N_14919,N_14690,N_14738);
nand U14920 (N_14920,N_14605,N_14699);
nor U14921 (N_14921,N_14544,N_14746);
or U14922 (N_14922,N_14624,N_14648);
or U14923 (N_14923,N_14581,N_14546);
nor U14924 (N_14924,N_14662,N_14677);
and U14925 (N_14925,N_14567,N_14719);
or U14926 (N_14926,N_14706,N_14676);
or U14927 (N_14927,N_14684,N_14623);
nand U14928 (N_14928,N_14612,N_14513);
nand U14929 (N_14929,N_14710,N_14576);
and U14930 (N_14930,N_14731,N_14516);
xor U14931 (N_14931,N_14524,N_14503);
nor U14932 (N_14932,N_14714,N_14638);
nand U14933 (N_14933,N_14582,N_14517);
nand U14934 (N_14934,N_14721,N_14592);
nor U14935 (N_14935,N_14723,N_14732);
nor U14936 (N_14936,N_14513,N_14656);
or U14937 (N_14937,N_14709,N_14578);
nand U14938 (N_14938,N_14634,N_14588);
nor U14939 (N_14939,N_14545,N_14710);
nand U14940 (N_14940,N_14711,N_14646);
xnor U14941 (N_14941,N_14553,N_14548);
and U14942 (N_14942,N_14738,N_14656);
or U14943 (N_14943,N_14631,N_14685);
xor U14944 (N_14944,N_14664,N_14608);
and U14945 (N_14945,N_14527,N_14588);
nand U14946 (N_14946,N_14653,N_14680);
or U14947 (N_14947,N_14708,N_14515);
and U14948 (N_14948,N_14532,N_14615);
or U14949 (N_14949,N_14707,N_14538);
xnor U14950 (N_14950,N_14603,N_14531);
or U14951 (N_14951,N_14715,N_14684);
nand U14952 (N_14952,N_14692,N_14568);
and U14953 (N_14953,N_14687,N_14555);
nor U14954 (N_14954,N_14619,N_14593);
and U14955 (N_14955,N_14638,N_14621);
xor U14956 (N_14956,N_14669,N_14590);
xor U14957 (N_14957,N_14586,N_14687);
nand U14958 (N_14958,N_14500,N_14663);
nand U14959 (N_14959,N_14518,N_14687);
or U14960 (N_14960,N_14661,N_14591);
nand U14961 (N_14961,N_14528,N_14611);
nand U14962 (N_14962,N_14604,N_14630);
nor U14963 (N_14963,N_14556,N_14716);
nand U14964 (N_14964,N_14516,N_14693);
nand U14965 (N_14965,N_14623,N_14567);
and U14966 (N_14966,N_14595,N_14648);
xor U14967 (N_14967,N_14536,N_14504);
nand U14968 (N_14968,N_14664,N_14571);
or U14969 (N_14969,N_14562,N_14535);
xor U14970 (N_14970,N_14667,N_14544);
nor U14971 (N_14971,N_14749,N_14744);
nor U14972 (N_14972,N_14521,N_14568);
nor U14973 (N_14973,N_14593,N_14734);
nand U14974 (N_14974,N_14682,N_14505);
or U14975 (N_14975,N_14568,N_14523);
nor U14976 (N_14976,N_14580,N_14701);
nor U14977 (N_14977,N_14650,N_14530);
nor U14978 (N_14978,N_14662,N_14516);
and U14979 (N_14979,N_14693,N_14716);
and U14980 (N_14980,N_14530,N_14712);
and U14981 (N_14981,N_14619,N_14717);
xnor U14982 (N_14982,N_14521,N_14609);
and U14983 (N_14983,N_14718,N_14591);
nand U14984 (N_14984,N_14609,N_14688);
nand U14985 (N_14985,N_14597,N_14536);
and U14986 (N_14986,N_14707,N_14509);
nor U14987 (N_14987,N_14635,N_14687);
xor U14988 (N_14988,N_14611,N_14662);
xnor U14989 (N_14989,N_14645,N_14737);
xor U14990 (N_14990,N_14558,N_14706);
xnor U14991 (N_14991,N_14644,N_14720);
xor U14992 (N_14992,N_14500,N_14646);
xnor U14993 (N_14993,N_14714,N_14619);
xnor U14994 (N_14994,N_14528,N_14671);
xnor U14995 (N_14995,N_14532,N_14742);
and U14996 (N_14996,N_14692,N_14578);
nor U14997 (N_14997,N_14662,N_14514);
and U14998 (N_14998,N_14558,N_14588);
and U14999 (N_14999,N_14711,N_14726);
or UO_0 (O_0,N_14841,N_14790);
nand UO_1 (O_1,N_14928,N_14794);
nor UO_2 (O_2,N_14810,N_14856);
nand UO_3 (O_3,N_14912,N_14819);
nand UO_4 (O_4,N_14814,N_14767);
nand UO_5 (O_5,N_14880,N_14958);
nand UO_6 (O_6,N_14801,N_14861);
nor UO_7 (O_7,N_14782,N_14753);
nor UO_8 (O_8,N_14800,N_14891);
or UO_9 (O_9,N_14983,N_14972);
or UO_10 (O_10,N_14953,N_14837);
nor UO_11 (O_11,N_14942,N_14895);
nand UO_12 (O_12,N_14973,N_14916);
nor UO_13 (O_13,N_14905,N_14866);
or UO_14 (O_14,N_14902,N_14967);
nand UO_15 (O_15,N_14757,N_14795);
and UO_16 (O_16,N_14862,N_14915);
xor UO_17 (O_17,N_14934,N_14892);
xnor UO_18 (O_18,N_14952,N_14830);
nor UO_19 (O_19,N_14899,N_14930);
xnor UO_20 (O_20,N_14997,N_14765);
and UO_21 (O_21,N_14998,N_14760);
xnor UO_22 (O_22,N_14931,N_14940);
and UO_23 (O_23,N_14806,N_14846);
nand UO_24 (O_24,N_14761,N_14828);
xor UO_25 (O_25,N_14885,N_14957);
nand UO_26 (O_26,N_14909,N_14988);
and UO_27 (O_27,N_14871,N_14923);
or UO_28 (O_28,N_14787,N_14950);
xnor UO_29 (O_29,N_14775,N_14858);
xor UO_30 (O_30,N_14961,N_14829);
xnor UO_31 (O_31,N_14919,N_14850);
nand UO_32 (O_32,N_14750,N_14815);
or UO_33 (O_33,N_14857,N_14867);
xnor UO_34 (O_34,N_14981,N_14991);
nor UO_35 (O_35,N_14783,N_14881);
xor UO_36 (O_36,N_14977,N_14774);
and UO_37 (O_37,N_14766,N_14922);
xnor UO_38 (O_38,N_14852,N_14848);
or UO_39 (O_39,N_14808,N_14901);
or UO_40 (O_40,N_14821,N_14924);
and UO_41 (O_41,N_14859,N_14823);
nand UO_42 (O_42,N_14944,N_14799);
or UO_43 (O_43,N_14995,N_14763);
or UO_44 (O_44,N_14968,N_14978);
and UO_45 (O_45,N_14875,N_14836);
nor UO_46 (O_46,N_14752,N_14835);
nand UO_47 (O_47,N_14876,N_14863);
or UO_48 (O_48,N_14751,N_14869);
and UO_49 (O_49,N_14911,N_14807);
and UO_50 (O_50,N_14969,N_14793);
nor UO_51 (O_51,N_14938,N_14804);
nand UO_52 (O_52,N_14762,N_14965);
nor UO_53 (O_53,N_14847,N_14927);
or UO_54 (O_54,N_14888,N_14925);
and UO_55 (O_55,N_14985,N_14797);
and UO_56 (O_56,N_14879,N_14939);
nand UO_57 (O_57,N_14851,N_14975);
nor UO_58 (O_58,N_14853,N_14779);
nand UO_59 (O_59,N_14758,N_14755);
nor UO_60 (O_60,N_14894,N_14802);
xnor UO_61 (O_61,N_14865,N_14769);
and UO_62 (O_62,N_14898,N_14893);
and UO_63 (O_63,N_14951,N_14900);
and UO_64 (O_64,N_14897,N_14936);
nor UO_65 (O_65,N_14826,N_14780);
xnor UO_66 (O_66,N_14896,N_14812);
nand UO_67 (O_67,N_14976,N_14824);
xnor UO_68 (O_68,N_14887,N_14788);
nor UO_69 (O_69,N_14992,N_14822);
nand UO_70 (O_70,N_14868,N_14960);
nor UO_71 (O_71,N_14820,N_14993);
nor UO_72 (O_72,N_14831,N_14874);
or UO_73 (O_73,N_14979,N_14903);
nor UO_74 (O_74,N_14994,N_14918);
xnor UO_75 (O_75,N_14803,N_14791);
xnor UO_76 (O_76,N_14789,N_14945);
nand UO_77 (O_77,N_14770,N_14811);
or UO_78 (O_78,N_14864,N_14982);
or UO_79 (O_79,N_14827,N_14778);
or UO_80 (O_80,N_14785,N_14832);
nand UO_81 (O_81,N_14984,N_14920);
nand UO_82 (O_82,N_14825,N_14890);
and UO_83 (O_83,N_14781,N_14932);
xnor UO_84 (O_84,N_14870,N_14873);
nor UO_85 (O_85,N_14929,N_14882);
or UO_86 (O_86,N_14980,N_14809);
and UO_87 (O_87,N_14877,N_14817);
and UO_88 (O_88,N_14843,N_14948);
nand UO_89 (O_89,N_14844,N_14963);
and UO_90 (O_90,N_14756,N_14962);
or UO_91 (O_91,N_14816,N_14910);
nand UO_92 (O_92,N_14949,N_14933);
nand UO_93 (O_93,N_14926,N_14917);
nor UO_94 (O_94,N_14906,N_14845);
xnor UO_95 (O_95,N_14907,N_14908);
or UO_96 (O_96,N_14966,N_14798);
or UO_97 (O_97,N_14937,N_14889);
or UO_98 (O_98,N_14974,N_14834);
nand UO_99 (O_99,N_14784,N_14956);
nor UO_100 (O_100,N_14838,N_14792);
xnor UO_101 (O_101,N_14833,N_14860);
and UO_102 (O_102,N_14886,N_14754);
and UO_103 (O_103,N_14818,N_14935);
or UO_104 (O_104,N_14947,N_14839);
xnor UO_105 (O_105,N_14921,N_14954);
or UO_106 (O_106,N_14971,N_14996);
and UO_107 (O_107,N_14946,N_14773);
and UO_108 (O_108,N_14764,N_14796);
and UO_109 (O_109,N_14987,N_14854);
or UO_110 (O_110,N_14884,N_14990);
or UO_111 (O_111,N_14914,N_14786);
nor UO_112 (O_112,N_14759,N_14964);
nand UO_113 (O_113,N_14849,N_14878);
xor UO_114 (O_114,N_14904,N_14776);
or UO_115 (O_115,N_14986,N_14999);
xor UO_116 (O_116,N_14959,N_14772);
nand UO_117 (O_117,N_14840,N_14768);
xor UO_118 (O_118,N_14913,N_14941);
nor UO_119 (O_119,N_14842,N_14989);
and UO_120 (O_120,N_14813,N_14955);
nand UO_121 (O_121,N_14777,N_14771);
and UO_122 (O_122,N_14943,N_14805);
nand UO_123 (O_123,N_14970,N_14855);
nand UO_124 (O_124,N_14883,N_14872);
nand UO_125 (O_125,N_14822,N_14863);
and UO_126 (O_126,N_14983,N_14953);
xor UO_127 (O_127,N_14800,N_14755);
nand UO_128 (O_128,N_14872,N_14898);
nor UO_129 (O_129,N_14925,N_14895);
or UO_130 (O_130,N_14907,N_14999);
nor UO_131 (O_131,N_14876,N_14862);
nand UO_132 (O_132,N_14926,N_14815);
or UO_133 (O_133,N_14823,N_14973);
xor UO_134 (O_134,N_14878,N_14966);
or UO_135 (O_135,N_14816,N_14762);
or UO_136 (O_136,N_14934,N_14811);
and UO_137 (O_137,N_14786,N_14939);
nor UO_138 (O_138,N_14753,N_14883);
nor UO_139 (O_139,N_14796,N_14775);
and UO_140 (O_140,N_14805,N_14920);
xor UO_141 (O_141,N_14882,N_14797);
nor UO_142 (O_142,N_14885,N_14846);
nor UO_143 (O_143,N_14757,N_14900);
nand UO_144 (O_144,N_14756,N_14929);
nand UO_145 (O_145,N_14768,N_14898);
nor UO_146 (O_146,N_14822,N_14844);
xor UO_147 (O_147,N_14887,N_14829);
or UO_148 (O_148,N_14896,N_14999);
nor UO_149 (O_149,N_14877,N_14838);
and UO_150 (O_150,N_14922,N_14755);
and UO_151 (O_151,N_14858,N_14799);
and UO_152 (O_152,N_14834,N_14844);
and UO_153 (O_153,N_14994,N_14883);
and UO_154 (O_154,N_14775,N_14933);
xnor UO_155 (O_155,N_14980,N_14871);
or UO_156 (O_156,N_14970,N_14987);
nand UO_157 (O_157,N_14804,N_14970);
or UO_158 (O_158,N_14782,N_14910);
xor UO_159 (O_159,N_14888,N_14927);
nand UO_160 (O_160,N_14999,N_14884);
nand UO_161 (O_161,N_14791,N_14814);
nor UO_162 (O_162,N_14923,N_14942);
and UO_163 (O_163,N_14991,N_14939);
xor UO_164 (O_164,N_14830,N_14758);
nand UO_165 (O_165,N_14918,N_14874);
xor UO_166 (O_166,N_14819,N_14777);
and UO_167 (O_167,N_14876,N_14925);
or UO_168 (O_168,N_14902,N_14859);
or UO_169 (O_169,N_14987,N_14979);
or UO_170 (O_170,N_14987,N_14927);
or UO_171 (O_171,N_14899,N_14835);
or UO_172 (O_172,N_14907,N_14861);
or UO_173 (O_173,N_14762,N_14972);
and UO_174 (O_174,N_14856,N_14874);
or UO_175 (O_175,N_14823,N_14809);
and UO_176 (O_176,N_14896,N_14783);
or UO_177 (O_177,N_14916,N_14818);
nor UO_178 (O_178,N_14861,N_14982);
nand UO_179 (O_179,N_14831,N_14825);
nand UO_180 (O_180,N_14991,N_14767);
or UO_181 (O_181,N_14916,N_14784);
nor UO_182 (O_182,N_14877,N_14799);
and UO_183 (O_183,N_14795,N_14982);
nand UO_184 (O_184,N_14952,N_14779);
nor UO_185 (O_185,N_14755,N_14857);
xor UO_186 (O_186,N_14940,N_14832);
nor UO_187 (O_187,N_14758,N_14979);
nand UO_188 (O_188,N_14762,N_14899);
nor UO_189 (O_189,N_14959,N_14813);
or UO_190 (O_190,N_14885,N_14941);
nand UO_191 (O_191,N_14831,N_14757);
xnor UO_192 (O_192,N_14774,N_14779);
nor UO_193 (O_193,N_14977,N_14906);
nand UO_194 (O_194,N_14885,N_14908);
or UO_195 (O_195,N_14773,N_14903);
nor UO_196 (O_196,N_14753,N_14919);
xor UO_197 (O_197,N_14981,N_14947);
nor UO_198 (O_198,N_14877,N_14860);
xnor UO_199 (O_199,N_14787,N_14864);
nor UO_200 (O_200,N_14925,N_14860);
nor UO_201 (O_201,N_14803,N_14837);
nor UO_202 (O_202,N_14952,N_14984);
xnor UO_203 (O_203,N_14841,N_14817);
xor UO_204 (O_204,N_14866,N_14999);
nand UO_205 (O_205,N_14970,N_14833);
nand UO_206 (O_206,N_14791,N_14978);
nand UO_207 (O_207,N_14841,N_14968);
nor UO_208 (O_208,N_14966,N_14779);
and UO_209 (O_209,N_14967,N_14895);
or UO_210 (O_210,N_14961,N_14973);
and UO_211 (O_211,N_14758,N_14856);
or UO_212 (O_212,N_14944,N_14975);
nor UO_213 (O_213,N_14983,N_14999);
xnor UO_214 (O_214,N_14800,N_14887);
nand UO_215 (O_215,N_14898,N_14954);
and UO_216 (O_216,N_14795,N_14954);
and UO_217 (O_217,N_14861,N_14976);
or UO_218 (O_218,N_14908,N_14838);
nor UO_219 (O_219,N_14809,N_14931);
or UO_220 (O_220,N_14852,N_14799);
or UO_221 (O_221,N_14834,N_14972);
nor UO_222 (O_222,N_14828,N_14917);
nand UO_223 (O_223,N_14802,N_14804);
xnor UO_224 (O_224,N_14864,N_14921);
or UO_225 (O_225,N_14955,N_14832);
or UO_226 (O_226,N_14974,N_14907);
xnor UO_227 (O_227,N_14861,N_14753);
nor UO_228 (O_228,N_14895,N_14936);
nor UO_229 (O_229,N_14779,N_14874);
or UO_230 (O_230,N_14808,N_14875);
nand UO_231 (O_231,N_14764,N_14911);
xnor UO_232 (O_232,N_14893,N_14909);
and UO_233 (O_233,N_14831,N_14990);
or UO_234 (O_234,N_14783,N_14975);
or UO_235 (O_235,N_14925,N_14962);
nand UO_236 (O_236,N_14825,N_14906);
nor UO_237 (O_237,N_14854,N_14982);
nor UO_238 (O_238,N_14929,N_14927);
and UO_239 (O_239,N_14753,N_14979);
nand UO_240 (O_240,N_14769,N_14993);
xnor UO_241 (O_241,N_14847,N_14836);
and UO_242 (O_242,N_14911,N_14885);
xnor UO_243 (O_243,N_14923,N_14939);
or UO_244 (O_244,N_14768,N_14807);
nor UO_245 (O_245,N_14754,N_14796);
xnor UO_246 (O_246,N_14994,N_14897);
or UO_247 (O_247,N_14888,N_14796);
nand UO_248 (O_248,N_14781,N_14941);
or UO_249 (O_249,N_14981,N_14852);
nor UO_250 (O_250,N_14999,N_14818);
or UO_251 (O_251,N_14793,N_14792);
nor UO_252 (O_252,N_14992,N_14929);
and UO_253 (O_253,N_14871,N_14793);
nand UO_254 (O_254,N_14986,N_14757);
xnor UO_255 (O_255,N_14789,N_14797);
nand UO_256 (O_256,N_14762,N_14867);
or UO_257 (O_257,N_14804,N_14796);
and UO_258 (O_258,N_14823,N_14828);
or UO_259 (O_259,N_14851,N_14758);
nand UO_260 (O_260,N_14986,N_14851);
xor UO_261 (O_261,N_14834,N_14900);
or UO_262 (O_262,N_14865,N_14901);
and UO_263 (O_263,N_14847,N_14960);
and UO_264 (O_264,N_14912,N_14843);
nand UO_265 (O_265,N_14797,N_14957);
or UO_266 (O_266,N_14934,N_14841);
xnor UO_267 (O_267,N_14766,N_14883);
and UO_268 (O_268,N_14967,N_14751);
nor UO_269 (O_269,N_14944,N_14982);
nand UO_270 (O_270,N_14778,N_14842);
or UO_271 (O_271,N_14951,N_14819);
or UO_272 (O_272,N_14834,N_14994);
nor UO_273 (O_273,N_14767,N_14994);
and UO_274 (O_274,N_14764,N_14912);
nand UO_275 (O_275,N_14822,N_14930);
nor UO_276 (O_276,N_14851,N_14923);
xnor UO_277 (O_277,N_14874,N_14894);
nor UO_278 (O_278,N_14942,N_14786);
nor UO_279 (O_279,N_14916,N_14862);
nand UO_280 (O_280,N_14794,N_14898);
nor UO_281 (O_281,N_14935,N_14843);
nand UO_282 (O_282,N_14884,N_14880);
nand UO_283 (O_283,N_14754,N_14889);
xor UO_284 (O_284,N_14785,N_14882);
nand UO_285 (O_285,N_14907,N_14992);
xor UO_286 (O_286,N_14854,N_14955);
or UO_287 (O_287,N_14935,N_14856);
nand UO_288 (O_288,N_14843,N_14763);
nor UO_289 (O_289,N_14892,N_14873);
nor UO_290 (O_290,N_14911,N_14786);
and UO_291 (O_291,N_14845,N_14888);
or UO_292 (O_292,N_14893,N_14945);
nor UO_293 (O_293,N_14870,N_14766);
or UO_294 (O_294,N_14870,N_14832);
and UO_295 (O_295,N_14807,N_14797);
xnor UO_296 (O_296,N_14831,N_14907);
nor UO_297 (O_297,N_14859,N_14915);
and UO_298 (O_298,N_14995,N_14786);
xor UO_299 (O_299,N_14780,N_14806);
nand UO_300 (O_300,N_14806,N_14801);
xnor UO_301 (O_301,N_14840,N_14856);
nand UO_302 (O_302,N_14964,N_14913);
nand UO_303 (O_303,N_14828,N_14824);
nand UO_304 (O_304,N_14770,N_14983);
nand UO_305 (O_305,N_14919,N_14959);
xor UO_306 (O_306,N_14893,N_14774);
and UO_307 (O_307,N_14988,N_14955);
xnor UO_308 (O_308,N_14938,N_14819);
xor UO_309 (O_309,N_14850,N_14978);
nand UO_310 (O_310,N_14857,N_14946);
and UO_311 (O_311,N_14824,N_14893);
or UO_312 (O_312,N_14945,N_14925);
and UO_313 (O_313,N_14774,N_14813);
or UO_314 (O_314,N_14838,N_14968);
or UO_315 (O_315,N_14906,N_14946);
xor UO_316 (O_316,N_14991,N_14756);
xnor UO_317 (O_317,N_14802,N_14959);
xnor UO_318 (O_318,N_14790,N_14931);
xnor UO_319 (O_319,N_14757,N_14853);
nor UO_320 (O_320,N_14990,N_14762);
nand UO_321 (O_321,N_14810,N_14776);
nor UO_322 (O_322,N_14960,N_14888);
or UO_323 (O_323,N_14983,N_14887);
xor UO_324 (O_324,N_14751,N_14915);
nand UO_325 (O_325,N_14994,N_14763);
xnor UO_326 (O_326,N_14949,N_14945);
nand UO_327 (O_327,N_14804,N_14893);
or UO_328 (O_328,N_14935,N_14893);
nand UO_329 (O_329,N_14771,N_14969);
xnor UO_330 (O_330,N_14829,N_14891);
xnor UO_331 (O_331,N_14901,N_14985);
and UO_332 (O_332,N_14857,N_14814);
xor UO_333 (O_333,N_14980,N_14799);
and UO_334 (O_334,N_14828,N_14849);
or UO_335 (O_335,N_14933,N_14978);
and UO_336 (O_336,N_14807,N_14754);
nor UO_337 (O_337,N_14809,N_14793);
nor UO_338 (O_338,N_14781,N_14760);
nand UO_339 (O_339,N_14840,N_14830);
xor UO_340 (O_340,N_14850,N_14953);
xor UO_341 (O_341,N_14934,N_14961);
and UO_342 (O_342,N_14839,N_14787);
and UO_343 (O_343,N_14800,N_14935);
nor UO_344 (O_344,N_14900,N_14914);
and UO_345 (O_345,N_14760,N_14831);
xnor UO_346 (O_346,N_14876,N_14891);
xnor UO_347 (O_347,N_14911,N_14948);
nand UO_348 (O_348,N_14762,N_14797);
xor UO_349 (O_349,N_14846,N_14935);
and UO_350 (O_350,N_14781,N_14894);
or UO_351 (O_351,N_14823,N_14792);
or UO_352 (O_352,N_14888,N_14963);
nor UO_353 (O_353,N_14790,N_14779);
xor UO_354 (O_354,N_14947,N_14905);
and UO_355 (O_355,N_14821,N_14982);
or UO_356 (O_356,N_14973,N_14832);
nand UO_357 (O_357,N_14845,N_14838);
or UO_358 (O_358,N_14913,N_14938);
nor UO_359 (O_359,N_14860,N_14944);
nand UO_360 (O_360,N_14765,N_14863);
xor UO_361 (O_361,N_14910,N_14948);
xnor UO_362 (O_362,N_14817,N_14830);
or UO_363 (O_363,N_14794,N_14951);
xnor UO_364 (O_364,N_14905,N_14812);
and UO_365 (O_365,N_14913,N_14970);
nor UO_366 (O_366,N_14895,N_14974);
xor UO_367 (O_367,N_14963,N_14919);
or UO_368 (O_368,N_14877,N_14857);
and UO_369 (O_369,N_14794,N_14995);
or UO_370 (O_370,N_14757,N_14910);
xor UO_371 (O_371,N_14853,N_14807);
xor UO_372 (O_372,N_14856,N_14800);
xnor UO_373 (O_373,N_14804,N_14964);
xnor UO_374 (O_374,N_14803,N_14842);
nand UO_375 (O_375,N_14841,N_14831);
nor UO_376 (O_376,N_14932,N_14800);
nand UO_377 (O_377,N_14834,N_14775);
or UO_378 (O_378,N_14926,N_14887);
xor UO_379 (O_379,N_14819,N_14828);
nand UO_380 (O_380,N_14947,N_14893);
and UO_381 (O_381,N_14904,N_14841);
and UO_382 (O_382,N_14891,N_14849);
or UO_383 (O_383,N_14892,N_14803);
nand UO_384 (O_384,N_14792,N_14921);
nor UO_385 (O_385,N_14884,N_14946);
xor UO_386 (O_386,N_14970,N_14784);
nor UO_387 (O_387,N_14825,N_14915);
nor UO_388 (O_388,N_14848,N_14922);
xor UO_389 (O_389,N_14865,N_14884);
or UO_390 (O_390,N_14827,N_14909);
xnor UO_391 (O_391,N_14804,N_14894);
and UO_392 (O_392,N_14858,N_14878);
and UO_393 (O_393,N_14820,N_14834);
or UO_394 (O_394,N_14966,N_14847);
and UO_395 (O_395,N_14943,N_14950);
nand UO_396 (O_396,N_14961,N_14774);
nor UO_397 (O_397,N_14772,N_14837);
nor UO_398 (O_398,N_14895,N_14978);
or UO_399 (O_399,N_14992,N_14794);
or UO_400 (O_400,N_14929,N_14846);
nand UO_401 (O_401,N_14899,N_14801);
or UO_402 (O_402,N_14837,N_14987);
or UO_403 (O_403,N_14984,N_14854);
nand UO_404 (O_404,N_14887,N_14923);
or UO_405 (O_405,N_14897,N_14792);
or UO_406 (O_406,N_14880,N_14825);
or UO_407 (O_407,N_14969,N_14962);
xor UO_408 (O_408,N_14806,N_14805);
and UO_409 (O_409,N_14948,N_14811);
or UO_410 (O_410,N_14982,N_14827);
nand UO_411 (O_411,N_14798,N_14953);
and UO_412 (O_412,N_14806,N_14974);
nor UO_413 (O_413,N_14958,N_14901);
xor UO_414 (O_414,N_14852,N_14752);
and UO_415 (O_415,N_14882,N_14900);
nand UO_416 (O_416,N_14824,N_14807);
nand UO_417 (O_417,N_14855,N_14952);
xor UO_418 (O_418,N_14830,N_14969);
xor UO_419 (O_419,N_14882,N_14820);
or UO_420 (O_420,N_14996,N_14883);
nand UO_421 (O_421,N_14904,N_14871);
or UO_422 (O_422,N_14939,N_14894);
and UO_423 (O_423,N_14815,N_14975);
xor UO_424 (O_424,N_14845,N_14912);
nor UO_425 (O_425,N_14943,N_14833);
xor UO_426 (O_426,N_14882,N_14997);
nor UO_427 (O_427,N_14816,N_14962);
xor UO_428 (O_428,N_14796,N_14944);
xnor UO_429 (O_429,N_14997,N_14975);
and UO_430 (O_430,N_14889,N_14820);
nor UO_431 (O_431,N_14815,N_14962);
nand UO_432 (O_432,N_14837,N_14847);
nor UO_433 (O_433,N_14795,N_14817);
and UO_434 (O_434,N_14967,N_14817);
or UO_435 (O_435,N_14973,N_14908);
nor UO_436 (O_436,N_14873,N_14906);
xor UO_437 (O_437,N_14933,N_14787);
nor UO_438 (O_438,N_14899,N_14952);
or UO_439 (O_439,N_14794,N_14805);
nor UO_440 (O_440,N_14975,N_14856);
or UO_441 (O_441,N_14979,N_14782);
or UO_442 (O_442,N_14873,N_14902);
xnor UO_443 (O_443,N_14857,N_14873);
and UO_444 (O_444,N_14950,N_14854);
nand UO_445 (O_445,N_14876,N_14875);
and UO_446 (O_446,N_14786,N_14797);
or UO_447 (O_447,N_14892,N_14751);
and UO_448 (O_448,N_14884,N_14930);
nor UO_449 (O_449,N_14977,N_14807);
or UO_450 (O_450,N_14957,N_14854);
nor UO_451 (O_451,N_14845,N_14797);
nor UO_452 (O_452,N_14841,N_14889);
or UO_453 (O_453,N_14986,N_14905);
and UO_454 (O_454,N_14951,N_14929);
or UO_455 (O_455,N_14841,N_14852);
or UO_456 (O_456,N_14792,N_14886);
or UO_457 (O_457,N_14910,N_14867);
and UO_458 (O_458,N_14872,N_14773);
nor UO_459 (O_459,N_14879,N_14821);
xor UO_460 (O_460,N_14901,N_14774);
or UO_461 (O_461,N_14985,N_14995);
nand UO_462 (O_462,N_14778,N_14976);
or UO_463 (O_463,N_14972,N_14823);
nor UO_464 (O_464,N_14979,N_14834);
nor UO_465 (O_465,N_14768,N_14893);
nor UO_466 (O_466,N_14798,N_14758);
and UO_467 (O_467,N_14814,N_14858);
and UO_468 (O_468,N_14918,N_14930);
nand UO_469 (O_469,N_14946,N_14824);
and UO_470 (O_470,N_14915,N_14966);
or UO_471 (O_471,N_14837,N_14899);
and UO_472 (O_472,N_14901,N_14870);
nand UO_473 (O_473,N_14985,N_14827);
nor UO_474 (O_474,N_14959,N_14843);
and UO_475 (O_475,N_14999,N_14759);
nor UO_476 (O_476,N_14911,N_14773);
xor UO_477 (O_477,N_14991,N_14935);
or UO_478 (O_478,N_14775,N_14849);
nor UO_479 (O_479,N_14829,N_14856);
nand UO_480 (O_480,N_14862,N_14973);
and UO_481 (O_481,N_14833,N_14840);
or UO_482 (O_482,N_14787,N_14960);
nand UO_483 (O_483,N_14802,N_14781);
or UO_484 (O_484,N_14808,N_14877);
or UO_485 (O_485,N_14923,N_14777);
nand UO_486 (O_486,N_14971,N_14848);
nor UO_487 (O_487,N_14822,N_14888);
xnor UO_488 (O_488,N_14981,N_14758);
or UO_489 (O_489,N_14948,N_14929);
nand UO_490 (O_490,N_14845,N_14785);
xnor UO_491 (O_491,N_14977,N_14806);
and UO_492 (O_492,N_14821,N_14945);
or UO_493 (O_493,N_14758,N_14834);
and UO_494 (O_494,N_14809,N_14912);
or UO_495 (O_495,N_14987,N_14842);
xnor UO_496 (O_496,N_14840,N_14892);
xor UO_497 (O_497,N_14817,N_14943);
or UO_498 (O_498,N_14790,N_14830);
and UO_499 (O_499,N_14977,N_14770);
or UO_500 (O_500,N_14808,N_14852);
and UO_501 (O_501,N_14888,N_14945);
xor UO_502 (O_502,N_14929,N_14861);
nand UO_503 (O_503,N_14892,N_14777);
xnor UO_504 (O_504,N_14876,N_14877);
nor UO_505 (O_505,N_14768,N_14828);
nor UO_506 (O_506,N_14857,N_14888);
or UO_507 (O_507,N_14970,N_14916);
or UO_508 (O_508,N_14759,N_14790);
nor UO_509 (O_509,N_14761,N_14953);
or UO_510 (O_510,N_14898,N_14846);
xnor UO_511 (O_511,N_14937,N_14760);
and UO_512 (O_512,N_14832,N_14815);
nand UO_513 (O_513,N_14846,N_14942);
nor UO_514 (O_514,N_14843,N_14930);
or UO_515 (O_515,N_14993,N_14923);
nor UO_516 (O_516,N_14885,N_14929);
xor UO_517 (O_517,N_14811,N_14976);
nor UO_518 (O_518,N_14861,N_14780);
nand UO_519 (O_519,N_14839,N_14975);
and UO_520 (O_520,N_14852,N_14750);
xor UO_521 (O_521,N_14877,N_14790);
xnor UO_522 (O_522,N_14758,N_14914);
nand UO_523 (O_523,N_14865,N_14809);
or UO_524 (O_524,N_14753,N_14996);
nand UO_525 (O_525,N_14977,N_14933);
nor UO_526 (O_526,N_14986,N_14777);
xor UO_527 (O_527,N_14866,N_14851);
or UO_528 (O_528,N_14930,N_14960);
nor UO_529 (O_529,N_14899,N_14935);
nand UO_530 (O_530,N_14764,N_14915);
nand UO_531 (O_531,N_14975,N_14847);
or UO_532 (O_532,N_14937,N_14902);
and UO_533 (O_533,N_14912,N_14977);
nor UO_534 (O_534,N_14790,N_14777);
nor UO_535 (O_535,N_14885,N_14883);
nor UO_536 (O_536,N_14875,N_14993);
or UO_537 (O_537,N_14995,N_14925);
and UO_538 (O_538,N_14983,N_14955);
nor UO_539 (O_539,N_14846,N_14868);
xor UO_540 (O_540,N_14991,N_14819);
xor UO_541 (O_541,N_14766,N_14899);
nor UO_542 (O_542,N_14954,N_14775);
or UO_543 (O_543,N_14830,N_14943);
xnor UO_544 (O_544,N_14856,N_14947);
nand UO_545 (O_545,N_14947,N_14943);
nand UO_546 (O_546,N_14922,N_14754);
or UO_547 (O_547,N_14773,N_14953);
xnor UO_548 (O_548,N_14844,N_14976);
or UO_549 (O_549,N_14883,N_14799);
xor UO_550 (O_550,N_14862,N_14878);
xor UO_551 (O_551,N_14793,N_14902);
xor UO_552 (O_552,N_14967,N_14978);
xnor UO_553 (O_553,N_14954,N_14992);
nor UO_554 (O_554,N_14781,N_14993);
xor UO_555 (O_555,N_14956,N_14974);
and UO_556 (O_556,N_14808,N_14773);
or UO_557 (O_557,N_14928,N_14789);
nand UO_558 (O_558,N_14865,N_14797);
xor UO_559 (O_559,N_14943,N_14820);
or UO_560 (O_560,N_14753,N_14858);
nand UO_561 (O_561,N_14921,N_14951);
nand UO_562 (O_562,N_14826,N_14900);
xor UO_563 (O_563,N_14846,N_14945);
or UO_564 (O_564,N_14881,N_14753);
xnor UO_565 (O_565,N_14901,N_14978);
xnor UO_566 (O_566,N_14887,N_14864);
nor UO_567 (O_567,N_14972,N_14763);
and UO_568 (O_568,N_14823,N_14926);
or UO_569 (O_569,N_14940,N_14864);
nor UO_570 (O_570,N_14758,N_14768);
nand UO_571 (O_571,N_14761,N_14820);
nand UO_572 (O_572,N_14895,N_14880);
xor UO_573 (O_573,N_14895,N_14947);
and UO_574 (O_574,N_14865,N_14952);
nand UO_575 (O_575,N_14929,N_14998);
or UO_576 (O_576,N_14761,N_14843);
nand UO_577 (O_577,N_14818,N_14827);
or UO_578 (O_578,N_14924,N_14959);
xor UO_579 (O_579,N_14766,N_14901);
nor UO_580 (O_580,N_14807,N_14784);
xnor UO_581 (O_581,N_14902,N_14918);
or UO_582 (O_582,N_14905,N_14833);
and UO_583 (O_583,N_14842,N_14776);
or UO_584 (O_584,N_14914,N_14751);
nand UO_585 (O_585,N_14976,N_14859);
and UO_586 (O_586,N_14852,N_14851);
nand UO_587 (O_587,N_14903,N_14857);
nor UO_588 (O_588,N_14837,N_14836);
nor UO_589 (O_589,N_14774,N_14985);
nor UO_590 (O_590,N_14832,N_14920);
or UO_591 (O_591,N_14940,N_14754);
xor UO_592 (O_592,N_14834,N_14801);
or UO_593 (O_593,N_14848,N_14839);
and UO_594 (O_594,N_14862,N_14855);
nand UO_595 (O_595,N_14900,N_14853);
or UO_596 (O_596,N_14854,N_14978);
or UO_597 (O_597,N_14754,N_14794);
and UO_598 (O_598,N_14889,N_14860);
nand UO_599 (O_599,N_14927,N_14802);
and UO_600 (O_600,N_14808,N_14868);
nor UO_601 (O_601,N_14849,N_14769);
and UO_602 (O_602,N_14972,N_14985);
nand UO_603 (O_603,N_14766,N_14967);
nand UO_604 (O_604,N_14763,N_14866);
xor UO_605 (O_605,N_14904,N_14801);
nor UO_606 (O_606,N_14930,N_14956);
nor UO_607 (O_607,N_14760,N_14789);
or UO_608 (O_608,N_14996,N_14778);
and UO_609 (O_609,N_14915,N_14829);
and UO_610 (O_610,N_14979,N_14776);
nor UO_611 (O_611,N_14826,N_14888);
and UO_612 (O_612,N_14890,N_14946);
nor UO_613 (O_613,N_14926,N_14750);
xnor UO_614 (O_614,N_14895,N_14867);
and UO_615 (O_615,N_14782,N_14917);
nand UO_616 (O_616,N_14869,N_14786);
and UO_617 (O_617,N_14909,N_14854);
or UO_618 (O_618,N_14955,N_14984);
nand UO_619 (O_619,N_14837,N_14776);
nor UO_620 (O_620,N_14768,N_14904);
nor UO_621 (O_621,N_14876,N_14884);
or UO_622 (O_622,N_14908,N_14871);
xor UO_623 (O_623,N_14812,N_14900);
nor UO_624 (O_624,N_14937,N_14778);
or UO_625 (O_625,N_14756,N_14763);
nor UO_626 (O_626,N_14777,N_14803);
nor UO_627 (O_627,N_14923,N_14816);
and UO_628 (O_628,N_14798,N_14979);
xor UO_629 (O_629,N_14783,N_14957);
xnor UO_630 (O_630,N_14938,N_14791);
xnor UO_631 (O_631,N_14911,N_14772);
or UO_632 (O_632,N_14861,N_14996);
nor UO_633 (O_633,N_14876,N_14902);
and UO_634 (O_634,N_14983,N_14784);
xnor UO_635 (O_635,N_14819,N_14779);
or UO_636 (O_636,N_14862,N_14980);
or UO_637 (O_637,N_14791,N_14839);
and UO_638 (O_638,N_14879,N_14900);
xor UO_639 (O_639,N_14775,N_14824);
and UO_640 (O_640,N_14987,N_14988);
and UO_641 (O_641,N_14760,N_14959);
or UO_642 (O_642,N_14782,N_14958);
xnor UO_643 (O_643,N_14877,N_14958);
xnor UO_644 (O_644,N_14909,N_14766);
or UO_645 (O_645,N_14783,N_14879);
or UO_646 (O_646,N_14981,N_14799);
or UO_647 (O_647,N_14769,N_14991);
or UO_648 (O_648,N_14922,N_14820);
nor UO_649 (O_649,N_14915,N_14806);
or UO_650 (O_650,N_14958,N_14837);
nor UO_651 (O_651,N_14796,N_14793);
nand UO_652 (O_652,N_14918,N_14911);
or UO_653 (O_653,N_14788,N_14993);
or UO_654 (O_654,N_14967,N_14898);
nand UO_655 (O_655,N_14986,N_14874);
nor UO_656 (O_656,N_14872,N_14821);
or UO_657 (O_657,N_14857,N_14977);
and UO_658 (O_658,N_14914,N_14917);
and UO_659 (O_659,N_14940,N_14818);
and UO_660 (O_660,N_14968,N_14919);
xnor UO_661 (O_661,N_14826,N_14889);
nand UO_662 (O_662,N_14826,N_14921);
xnor UO_663 (O_663,N_14771,N_14772);
nand UO_664 (O_664,N_14969,N_14810);
nor UO_665 (O_665,N_14997,N_14793);
nand UO_666 (O_666,N_14884,N_14949);
and UO_667 (O_667,N_14977,N_14928);
nand UO_668 (O_668,N_14788,N_14865);
and UO_669 (O_669,N_14787,N_14944);
and UO_670 (O_670,N_14995,N_14856);
nor UO_671 (O_671,N_14889,N_14771);
nand UO_672 (O_672,N_14961,N_14965);
nor UO_673 (O_673,N_14839,N_14884);
xnor UO_674 (O_674,N_14782,N_14841);
xnor UO_675 (O_675,N_14802,N_14809);
xnor UO_676 (O_676,N_14780,N_14804);
and UO_677 (O_677,N_14953,N_14896);
nand UO_678 (O_678,N_14888,N_14984);
xnor UO_679 (O_679,N_14940,N_14889);
xnor UO_680 (O_680,N_14804,N_14900);
and UO_681 (O_681,N_14854,N_14792);
nor UO_682 (O_682,N_14819,N_14781);
and UO_683 (O_683,N_14893,N_14770);
and UO_684 (O_684,N_14970,N_14794);
and UO_685 (O_685,N_14785,N_14860);
and UO_686 (O_686,N_14860,N_14888);
nand UO_687 (O_687,N_14922,N_14750);
or UO_688 (O_688,N_14827,N_14782);
nand UO_689 (O_689,N_14845,N_14827);
nand UO_690 (O_690,N_14967,N_14816);
or UO_691 (O_691,N_14792,N_14966);
xnor UO_692 (O_692,N_14862,N_14893);
and UO_693 (O_693,N_14931,N_14984);
xnor UO_694 (O_694,N_14958,N_14873);
or UO_695 (O_695,N_14805,N_14957);
and UO_696 (O_696,N_14851,N_14972);
and UO_697 (O_697,N_14994,N_14911);
or UO_698 (O_698,N_14808,N_14959);
or UO_699 (O_699,N_14773,N_14793);
nor UO_700 (O_700,N_14963,N_14891);
and UO_701 (O_701,N_14900,N_14777);
nor UO_702 (O_702,N_14991,N_14924);
nand UO_703 (O_703,N_14959,N_14983);
and UO_704 (O_704,N_14954,N_14753);
nand UO_705 (O_705,N_14792,N_14799);
xor UO_706 (O_706,N_14872,N_14886);
and UO_707 (O_707,N_14782,N_14932);
and UO_708 (O_708,N_14860,N_14940);
nand UO_709 (O_709,N_14916,N_14808);
nand UO_710 (O_710,N_14808,N_14766);
or UO_711 (O_711,N_14915,N_14819);
nand UO_712 (O_712,N_14798,N_14807);
xor UO_713 (O_713,N_14939,N_14983);
xnor UO_714 (O_714,N_14915,N_14888);
nand UO_715 (O_715,N_14824,N_14903);
nor UO_716 (O_716,N_14805,N_14796);
xor UO_717 (O_717,N_14779,N_14943);
and UO_718 (O_718,N_14865,N_14883);
and UO_719 (O_719,N_14984,N_14769);
nand UO_720 (O_720,N_14827,N_14777);
nand UO_721 (O_721,N_14887,N_14786);
and UO_722 (O_722,N_14960,N_14962);
or UO_723 (O_723,N_14973,N_14903);
and UO_724 (O_724,N_14766,N_14794);
nor UO_725 (O_725,N_14992,N_14820);
nand UO_726 (O_726,N_14851,N_14774);
nor UO_727 (O_727,N_14881,N_14947);
xnor UO_728 (O_728,N_14836,N_14764);
and UO_729 (O_729,N_14882,N_14871);
nor UO_730 (O_730,N_14971,N_14896);
and UO_731 (O_731,N_14806,N_14858);
xor UO_732 (O_732,N_14806,N_14989);
nor UO_733 (O_733,N_14787,N_14762);
nor UO_734 (O_734,N_14901,N_14934);
and UO_735 (O_735,N_14954,N_14902);
nor UO_736 (O_736,N_14900,N_14779);
and UO_737 (O_737,N_14883,N_14849);
nand UO_738 (O_738,N_14832,N_14925);
and UO_739 (O_739,N_14971,N_14863);
or UO_740 (O_740,N_14993,N_14888);
xor UO_741 (O_741,N_14968,N_14918);
or UO_742 (O_742,N_14841,N_14981);
or UO_743 (O_743,N_14787,N_14911);
nor UO_744 (O_744,N_14861,N_14773);
nor UO_745 (O_745,N_14817,N_14931);
nand UO_746 (O_746,N_14982,N_14990);
or UO_747 (O_747,N_14860,N_14895);
xor UO_748 (O_748,N_14924,N_14893);
and UO_749 (O_749,N_14908,N_14761);
nor UO_750 (O_750,N_14806,N_14793);
xor UO_751 (O_751,N_14901,N_14917);
or UO_752 (O_752,N_14855,N_14752);
xnor UO_753 (O_753,N_14756,N_14764);
nor UO_754 (O_754,N_14969,N_14769);
nor UO_755 (O_755,N_14958,N_14803);
nor UO_756 (O_756,N_14845,N_14801);
nand UO_757 (O_757,N_14971,N_14794);
nand UO_758 (O_758,N_14887,N_14928);
nand UO_759 (O_759,N_14871,N_14932);
nand UO_760 (O_760,N_14790,N_14943);
nor UO_761 (O_761,N_14999,N_14872);
or UO_762 (O_762,N_14872,N_14944);
or UO_763 (O_763,N_14903,N_14789);
and UO_764 (O_764,N_14765,N_14977);
xor UO_765 (O_765,N_14808,N_14892);
and UO_766 (O_766,N_14889,N_14894);
nand UO_767 (O_767,N_14895,N_14788);
and UO_768 (O_768,N_14785,N_14976);
or UO_769 (O_769,N_14797,N_14852);
nand UO_770 (O_770,N_14791,N_14751);
nand UO_771 (O_771,N_14971,N_14985);
nand UO_772 (O_772,N_14852,N_14753);
xor UO_773 (O_773,N_14835,N_14834);
and UO_774 (O_774,N_14964,N_14805);
xor UO_775 (O_775,N_14911,N_14855);
and UO_776 (O_776,N_14764,N_14949);
nand UO_777 (O_777,N_14770,N_14853);
nor UO_778 (O_778,N_14860,N_14926);
and UO_779 (O_779,N_14960,N_14757);
or UO_780 (O_780,N_14961,N_14904);
and UO_781 (O_781,N_14987,N_14922);
and UO_782 (O_782,N_14935,N_14865);
or UO_783 (O_783,N_14811,N_14988);
xor UO_784 (O_784,N_14836,N_14808);
xnor UO_785 (O_785,N_14826,N_14918);
or UO_786 (O_786,N_14987,N_14770);
nor UO_787 (O_787,N_14954,N_14896);
xnor UO_788 (O_788,N_14823,N_14940);
nor UO_789 (O_789,N_14894,N_14774);
xnor UO_790 (O_790,N_14982,N_14969);
nand UO_791 (O_791,N_14832,N_14771);
nor UO_792 (O_792,N_14884,N_14829);
or UO_793 (O_793,N_14779,N_14958);
or UO_794 (O_794,N_14868,N_14908);
and UO_795 (O_795,N_14942,N_14838);
and UO_796 (O_796,N_14792,N_14888);
or UO_797 (O_797,N_14764,N_14898);
and UO_798 (O_798,N_14963,N_14977);
and UO_799 (O_799,N_14772,N_14784);
and UO_800 (O_800,N_14807,N_14781);
or UO_801 (O_801,N_14829,N_14978);
xor UO_802 (O_802,N_14781,N_14901);
nand UO_803 (O_803,N_14839,N_14883);
xor UO_804 (O_804,N_14973,N_14853);
and UO_805 (O_805,N_14880,N_14908);
and UO_806 (O_806,N_14824,N_14764);
nand UO_807 (O_807,N_14925,N_14773);
nand UO_808 (O_808,N_14963,N_14985);
xor UO_809 (O_809,N_14976,N_14912);
nand UO_810 (O_810,N_14846,N_14946);
nor UO_811 (O_811,N_14847,N_14888);
or UO_812 (O_812,N_14802,N_14770);
or UO_813 (O_813,N_14916,N_14768);
nand UO_814 (O_814,N_14843,N_14945);
or UO_815 (O_815,N_14884,N_14753);
or UO_816 (O_816,N_14774,N_14866);
and UO_817 (O_817,N_14949,N_14834);
and UO_818 (O_818,N_14921,N_14866);
nand UO_819 (O_819,N_14768,N_14761);
or UO_820 (O_820,N_14892,N_14770);
or UO_821 (O_821,N_14859,N_14964);
nand UO_822 (O_822,N_14846,N_14802);
or UO_823 (O_823,N_14857,N_14978);
nor UO_824 (O_824,N_14929,N_14833);
xnor UO_825 (O_825,N_14978,N_14794);
and UO_826 (O_826,N_14955,N_14802);
xnor UO_827 (O_827,N_14757,N_14911);
nand UO_828 (O_828,N_14934,N_14830);
or UO_829 (O_829,N_14920,N_14958);
or UO_830 (O_830,N_14750,N_14921);
nor UO_831 (O_831,N_14857,N_14798);
nand UO_832 (O_832,N_14943,N_14967);
nand UO_833 (O_833,N_14936,N_14998);
nor UO_834 (O_834,N_14850,N_14955);
nand UO_835 (O_835,N_14972,N_14901);
xor UO_836 (O_836,N_14863,N_14827);
and UO_837 (O_837,N_14871,N_14892);
xnor UO_838 (O_838,N_14931,N_14908);
nor UO_839 (O_839,N_14948,N_14920);
nand UO_840 (O_840,N_14873,N_14949);
nor UO_841 (O_841,N_14857,N_14883);
and UO_842 (O_842,N_14974,N_14760);
nand UO_843 (O_843,N_14850,N_14756);
nor UO_844 (O_844,N_14876,N_14906);
nor UO_845 (O_845,N_14842,N_14867);
xor UO_846 (O_846,N_14778,N_14934);
nand UO_847 (O_847,N_14802,N_14881);
nand UO_848 (O_848,N_14878,N_14954);
and UO_849 (O_849,N_14765,N_14994);
xnor UO_850 (O_850,N_14846,N_14840);
and UO_851 (O_851,N_14962,N_14934);
or UO_852 (O_852,N_14823,N_14751);
or UO_853 (O_853,N_14817,N_14996);
xor UO_854 (O_854,N_14924,N_14999);
nand UO_855 (O_855,N_14817,N_14834);
and UO_856 (O_856,N_14765,N_14797);
and UO_857 (O_857,N_14983,N_14755);
nand UO_858 (O_858,N_14885,N_14967);
or UO_859 (O_859,N_14984,N_14820);
nand UO_860 (O_860,N_14834,N_14990);
and UO_861 (O_861,N_14895,N_14981);
nand UO_862 (O_862,N_14849,N_14766);
and UO_863 (O_863,N_14799,N_14918);
xor UO_864 (O_864,N_14867,N_14773);
xnor UO_865 (O_865,N_14907,N_14967);
nor UO_866 (O_866,N_14848,N_14913);
nor UO_867 (O_867,N_14988,N_14759);
nand UO_868 (O_868,N_14905,N_14896);
nor UO_869 (O_869,N_14964,N_14809);
nand UO_870 (O_870,N_14934,N_14922);
nand UO_871 (O_871,N_14924,N_14768);
nor UO_872 (O_872,N_14890,N_14853);
xnor UO_873 (O_873,N_14886,N_14756);
nand UO_874 (O_874,N_14957,N_14852);
nand UO_875 (O_875,N_14834,N_14836);
nand UO_876 (O_876,N_14922,N_14761);
nor UO_877 (O_877,N_14966,N_14852);
nand UO_878 (O_878,N_14978,N_14760);
nand UO_879 (O_879,N_14817,N_14757);
nor UO_880 (O_880,N_14960,N_14904);
nor UO_881 (O_881,N_14959,N_14951);
and UO_882 (O_882,N_14965,N_14773);
and UO_883 (O_883,N_14873,N_14938);
and UO_884 (O_884,N_14820,N_14999);
xnor UO_885 (O_885,N_14821,N_14923);
or UO_886 (O_886,N_14962,N_14966);
nand UO_887 (O_887,N_14973,N_14970);
and UO_888 (O_888,N_14756,N_14798);
nor UO_889 (O_889,N_14898,N_14787);
and UO_890 (O_890,N_14981,N_14976);
xor UO_891 (O_891,N_14756,N_14922);
and UO_892 (O_892,N_14958,N_14810);
nor UO_893 (O_893,N_14818,N_14912);
xor UO_894 (O_894,N_14911,N_14998);
nor UO_895 (O_895,N_14830,N_14842);
and UO_896 (O_896,N_14851,N_14819);
nand UO_897 (O_897,N_14881,N_14997);
or UO_898 (O_898,N_14908,N_14828);
nand UO_899 (O_899,N_14998,N_14854);
xnor UO_900 (O_900,N_14894,N_14863);
nand UO_901 (O_901,N_14822,N_14780);
and UO_902 (O_902,N_14984,N_14997);
or UO_903 (O_903,N_14782,N_14978);
or UO_904 (O_904,N_14918,N_14952);
or UO_905 (O_905,N_14938,N_14866);
xor UO_906 (O_906,N_14947,N_14758);
nand UO_907 (O_907,N_14976,N_14894);
or UO_908 (O_908,N_14868,N_14995);
nor UO_909 (O_909,N_14798,N_14892);
xor UO_910 (O_910,N_14950,N_14772);
nor UO_911 (O_911,N_14804,N_14908);
or UO_912 (O_912,N_14811,N_14835);
nor UO_913 (O_913,N_14856,N_14811);
nor UO_914 (O_914,N_14817,N_14924);
nand UO_915 (O_915,N_14876,N_14846);
xor UO_916 (O_916,N_14764,N_14965);
and UO_917 (O_917,N_14875,N_14868);
nand UO_918 (O_918,N_14947,N_14870);
and UO_919 (O_919,N_14908,N_14977);
and UO_920 (O_920,N_14819,N_14783);
and UO_921 (O_921,N_14876,N_14801);
and UO_922 (O_922,N_14999,N_14811);
or UO_923 (O_923,N_14954,N_14918);
nor UO_924 (O_924,N_14852,N_14809);
and UO_925 (O_925,N_14814,N_14944);
nor UO_926 (O_926,N_14816,N_14999);
xnor UO_927 (O_927,N_14866,N_14810);
nand UO_928 (O_928,N_14952,N_14962);
nor UO_929 (O_929,N_14948,N_14914);
xnor UO_930 (O_930,N_14911,N_14775);
or UO_931 (O_931,N_14935,N_14902);
or UO_932 (O_932,N_14816,N_14847);
nand UO_933 (O_933,N_14885,N_14942);
and UO_934 (O_934,N_14941,N_14783);
and UO_935 (O_935,N_14765,N_14909);
nand UO_936 (O_936,N_14858,N_14801);
or UO_937 (O_937,N_14808,N_14879);
xor UO_938 (O_938,N_14898,N_14890);
nor UO_939 (O_939,N_14958,N_14867);
nor UO_940 (O_940,N_14922,N_14825);
nand UO_941 (O_941,N_14961,N_14803);
nand UO_942 (O_942,N_14764,N_14997);
and UO_943 (O_943,N_14823,N_14900);
xnor UO_944 (O_944,N_14885,N_14958);
and UO_945 (O_945,N_14933,N_14843);
nand UO_946 (O_946,N_14934,N_14798);
nor UO_947 (O_947,N_14925,N_14934);
and UO_948 (O_948,N_14809,N_14862);
or UO_949 (O_949,N_14973,N_14805);
and UO_950 (O_950,N_14922,N_14771);
xnor UO_951 (O_951,N_14963,N_14845);
or UO_952 (O_952,N_14849,N_14926);
nor UO_953 (O_953,N_14932,N_14797);
nand UO_954 (O_954,N_14840,N_14953);
nor UO_955 (O_955,N_14870,N_14910);
or UO_956 (O_956,N_14828,N_14756);
and UO_957 (O_957,N_14762,N_14861);
nand UO_958 (O_958,N_14752,N_14818);
or UO_959 (O_959,N_14833,N_14802);
nor UO_960 (O_960,N_14767,N_14878);
xor UO_961 (O_961,N_14992,N_14919);
nor UO_962 (O_962,N_14970,N_14908);
and UO_963 (O_963,N_14757,N_14828);
and UO_964 (O_964,N_14894,N_14983);
and UO_965 (O_965,N_14948,N_14988);
and UO_966 (O_966,N_14974,N_14802);
or UO_967 (O_967,N_14946,N_14783);
nand UO_968 (O_968,N_14946,N_14949);
or UO_969 (O_969,N_14904,N_14881);
and UO_970 (O_970,N_14813,N_14786);
and UO_971 (O_971,N_14924,N_14964);
or UO_972 (O_972,N_14906,N_14881);
xnor UO_973 (O_973,N_14966,N_14775);
and UO_974 (O_974,N_14911,N_14900);
nor UO_975 (O_975,N_14796,N_14778);
or UO_976 (O_976,N_14783,N_14840);
or UO_977 (O_977,N_14911,N_14954);
or UO_978 (O_978,N_14948,N_14791);
and UO_979 (O_979,N_14833,N_14966);
nor UO_980 (O_980,N_14874,N_14812);
xor UO_981 (O_981,N_14802,N_14855);
nand UO_982 (O_982,N_14921,N_14798);
nand UO_983 (O_983,N_14888,N_14969);
or UO_984 (O_984,N_14854,N_14988);
nor UO_985 (O_985,N_14923,N_14917);
and UO_986 (O_986,N_14978,N_14790);
or UO_987 (O_987,N_14930,N_14871);
nand UO_988 (O_988,N_14828,N_14887);
nor UO_989 (O_989,N_14788,N_14862);
or UO_990 (O_990,N_14813,N_14823);
nand UO_991 (O_991,N_14941,N_14924);
or UO_992 (O_992,N_14839,N_14959);
or UO_993 (O_993,N_14898,N_14762);
and UO_994 (O_994,N_14834,N_14872);
xnor UO_995 (O_995,N_14991,N_14917);
and UO_996 (O_996,N_14984,N_14948);
nor UO_997 (O_997,N_14804,N_14994);
nor UO_998 (O_998,N_14989,N_14793);
and UO_999 (O_999,N_14809,N_14864);
nor UO_1000 (O_1000,N_14943,N_14819);
or UO_1001 (O_1001,N_14868,N_14831);
nor UO_1002 (O_1002,N_14892,N_14946);
and UO_1003 (O_1003,N_14830,N_14887);
and UO_1004 (O_1004,N_14888,N_14982);
nand UO_1005 (O_1005,N_14929,N_14857);
xor UO_1006 (O_1006,N_14921,N_14823);
xor UO_1007 (O_1007,N_14867,N_14814);
and UO_1008 (O_1008,N_14851,N_14796);
xor UO_1009 (O_1009,N_14935,N_14787);
and UO_1010 (O_1010,N_14816,N_14891);
nand UO_1011 (O_1011,N_14771,N_14851);
xor UO_1012 (O_1012,N_14891,N_14856);
nand UO_1013 (O_1013,N_14815,N_14968);
xnor UO_1014 (O_1014,N_14846,N_14877);
nor UO_1015 (O_1015,N_14802,N_14926);
and UO_1016 (O_1016,N_14759,N_14871);
nand UO_1017 (O_1017,N_14932,N_14934);
nor UO_1018 (O_1018,N_14788,N_14845);
and UO_1019 (O_1019,N_14842,N_14977);
nand UO_1020 (O_1020,N_14790,N_14799);
nor UO_1021 (O_1021,N_14969,N_14970);
nand UO_1022 (O_1022,N_14887,N_14880);
and UO_1023 (O_1023,N_14838,N_14771);
nor UO_1024 (O_1024,N_14800,N_14906);
and UO_1025 (O_1025,N_14940,N_14979);
nand UO_1026 (O_1026,N_14889,N_14765);
and UO_1027 (O_1027,N_14952,N_14891);
or UO_1028 (O_1028,N_14892,N_14940);
or UO_1029 (O_1029,N_14938,N_14784);
xnor UO_1030 (O_1030,N_14804,N_14825);
and UO_1031 (O_1031,N_14974,N_14967);
and UO_1032 (O_1032,N_14757,N_14761);
nor UO_1033 (O_1033,N_14757,N_14751);
nor UO_1034 (O_1034,N_14862,N_14918);
nor UO_1035 (O_1035,N_14792,N_14833);
or UO_1036 (O_1036,N_14797,N_14758);
and UO_1037 (O_1037,N_14938,N_14885);
and UO_1038 (O_1038,N_14963,N_14864);
nand UO_1039 (O_1039,N_14838,N_14851);
nor UO_1040 (O_1040,N_14828,N_14930);
and UO_1041 (O_1041,N_14965,N_14966);
nor UO_1042 (O_1042,N_14929,N_14923);
or UO_1043 (O_1043,N_14990,N_14877);
nand UO_1044 (O_1044,N_14816,N_14907);
and UO_1045 (O_1045,N_14988,N_14797);
or UO_1046 (O_1046,N_14992,N_14897);
xor UO_1047 (O_1047,N_14808,N_14947);
xor UO_1048 (O_1048,N_14930,N_14807);
or UO_1049 (O_1049,N_14862,N_14958);
xnor UO_1050 (O_1050,N_14931,N_14805);
nand UO_1051 (O_1051,N_14844,N_14846);
and UO_1052 (O_1052,N_14780,N_14881);
nor UO_1053 (O_1053,N_14957,N_14992);
nor UO_1054 (O_1054,N_14919,N_14791);
and UO_1055 (O_1055,N_14811,N_14771);
nor UO_1056 (O_1056,N_14949,N_14899);
nand UO_1057 (O_1057,N_14830,N_14976);
or UO_1058 (O_1058,N_14821,N_14792);
xnor UO_1059 (O_1059,N_14993,N_14817);
nor UO_1060 (O_1060,N_14795,N_14943);
xnor UO_1061 (O_1061,N_14800,N_14909);
or UO_1062 (O_1062,N_14991,N_14763);
and UO_1063 (O_1063,N_14997,N_14828);
nand UO_1064 (O_1064,N_14892,N_14832);
and UO_1065 (O_1065,N_14968,N_14924);
or UO_1066 (O_1066,N_14867,N_14919);
nor UO_1067 (O_1067,N_14823,N_14853);
xnor UO_1068 (O_1068,N_14903,N_14760);
nor UO_1069 (O_1069,N_14821,N_14772);
or UO_1070 (O_1070,N_14945,N_14764);
or UO_1071 (O_1071,N_14973,N_14890);
nor UO_1072 (O_1072,N_14871,N_14969);
or UO_1073 (O_1073,N_14762,N_14955);
or UO_1074 (O_1074,N_14755,N_14789);
or UO_1075 (O_1075,N_14936,N_14799);
and UO_1076 (O_1076,N_14865,N_14994);
nor UO_1077 (O_1077,N_14780,N_14952);
or UO_1078 (O_1078,N_14793,N_14751);
nand UO_1079 (O_1079,N_14964,N_14799);
and UO_1080 (O_1080,N_14758,N_14863);
nand UO_1081 (O_1081,N_14819,N_14974);
xnor UO_1082 (O_1082,N_14905,N_14824);
or UO_1083 (O_1083,N_14811,N_14782);
and UO_1084 (O_1084,N_14875,N_14844);
nor UO_1085 (O_1085,N_14786,N_14958);
xnor UO_1086 (O_1086,N_14970,N_14978);
and UO_1087 (O_1087,N_14985,N_14982);
and UO_1088 (O_1088,N_14883,N_14969);
and UO_1089 (O_1089,N_14864,N_14911);
or UO_1090 (O_1090,N_14950,N_14778);
xnor UO_1091 (O_1091,N_14851,N_14834);
or UO_1092 (O_1092,N_14865,N_14768);
nor UO_1093 (O_1093,N_14834,N_14897);
nand UO_1094 (O_1094,N_14802,N_14983);
and UO_1095 (O_1095,N_14936,N_14941);
and UO_1096 (O_1096,N_14818,N_14868);
or UO_1097 (O_1097,N_14768,N_14813);
xor UO_1098 (O_1098,N_14831,N_14903);
nor UO_1099 (O_1099,N_14993,N_14860);
and UO_1100 (O_1100,N_14940,N_14973);
xor UO_1101 (O_1101,N_14964,N_14780);
xnor UO_1102 (O_1102,N_14805,N_14954);
and UO_1103 (O_1103,N_14762,N_14789);
nor UO_1104 (O_1104,N_14883,N_14960);
nand UO_1105 (O_1105,N_14919,N_14796);
or UO_1106 (O_1106,N_14864,N_14783);
nor UO_1107 (O_1107,N_14844,N_14818);
and UO_1108 (O_1108,N_14869,N_14785);
xnor UO_1109 (O_1109,N_14758,N_14829);
nand UO_1110 (O_1110,N_14905,N_14903);
nand UO_1111 (O_1111,N_14933,N_14837);
nand UO_1112 (O_1112,N_14911,N_14981);
and UO_1113 (O_1113,N_14852,N_14866);
and UO_1114 (O_1114,N_14932,N_14830);
nand UO_1115 (O_1115,N_14972,N_14910);
nor UO_1116 (O_1116,N_14764,N_14933);
xnor UO_1117 (O_1117,N_14906,N_14904);
nand UO_1118 (O_1118,N_14784,N_14849);
nand UO_1119 (O_1119,N_14971,N_14938);
and UO_1120 (O_1120,N_14982,N_14831);
nand UO_1121 (O_1121,N_14809,N_14944);
xnor UO_1122 (O_1122,N_14835,N_14926);
and UO_1123 (O_1123,N_14896,N_14921);
nor UO_1124 (O_1124,N_14864,N_14898);
and UO_1125 (O_1125,N_14796,N_14830);
nand UO_1126 (O_1126,N_14908,N_14816);
xor UO_1127 (O_1127,N_14774,N_14905);
xor UO_1128 (O_1128,N_14936,N_14837);
nor UO_1129 (O_1129,N_14945,N_14799);
nor UO_1130 (O_1130,N_14883,N_14936);
nand UO_1131 (O_1131,N_14758,N_14857);
nor UO_1132 (O_1132,N_14892,N_14882);
nand UO_1133 (O_1133,N_14926,N_14879);
or UO_1134 (O_1134,N_14949,N_14806);
xnor UO_1135 (O_1135,N_14790,N_14886);
nand UO_1136 (O_1136,N_14989,N_14871);
nand UO_1137 (O_1137,N_14832,N_14836);
and UO_1138 (O_1138,N_14971,N_14950);
nand UO_1139 (O_1139,N_14831,N_14971);
and UO_1140 (O_1140,N_14793,N_14916);
or UO_1141 (O_1141,N_14832,N_14800);
and UO_1142 (O_1142,N_14854,N_14817);
and UO_1143 (O_1143,N_14931,N_14937);
or UO_1144 (O_1144,N_14850,N_14912);
nand UO_1145 (O_1145,N_14899,N_14978);
or UO_1146 (O_1146,N_14904,N_14870);
and UO_1147 (O_1147,N_14987,N_14971);
and UO_1148 (O_1148,N_14948,N_14969);
nand UO_1149 (O_1149,N_14792,N_14834);
or UO_1150 (O_1150,N_14889,N_14971);
and UO_1151 (O_1151,N_14855,N_14918);
or UO_1152 (O_1152,N_14971,N_14841);
nand UO_1153 (O_1153,N_14796,N_14861);
and UO_1154 (O_1154,N_14764,N_14846);
nand UO_1155 (O_1155,N_14995,N_14981);
and UO_1156 (O_1156,N_14830,N_14845);
and UO_1157 (O_1157,N_14943,N_14912);
nor UO_1158 (O_1158,N_14855,N_14776);
xnor UO_1159 (O_1159,N_14963,N_14918);
and UO_1160 (O_1160,N_14773,N_14996);
nor UO_1161 (O_1161,N_14812,N_14907);
and UO_1162 (O_1162,N_14987,N_14943);
nor UO_1163 (O_1163,N_14803,N_14982);
xnor UO_1164 (O_1164,N_14793,N_14753);
nand UO_1165 (O_1165,N_14981,N_14959);
or UO_1166 (O_1166,N_14873,N_14954);
nor UO_1167 (O_1167,N_14757,N_14988);
and UO_1168 (O_1168,N_14862,N_14899);
xor UO_1169 (O_1169,N_14907,N_14842);
nor UO_1170 (O_1170,N_14899,N_14923);
or UO_1171 (O_1171,N_14896,N_14917);
nor UO_1172 (O_1172,N_14945,N_14849);
xor UO_1173 (O_1173,N_14898,N_14896);
nand UO_1174 (O_1174,N_14886,N_14773);
nand UO_1175 (O_1175,N_14905,N_14957);
and UO_1176 (O_1176,N_14901,N_14855);
nand UO_1177 (O_1177,N_14976,N_14776);
nor UO_1178 (O_1178,N_14825,N_14910);
xor UO_1179 (O_1179,N_14958,N_14988);
nand UO_1180 (O_1180,N_14993,N_14838);
or UO_1181 (O_1181,N_14795,N_14850);
nor UO_1182 (O_1182,N_14789,N_14940);
xnor UO_1183 (O_1183,N_14916,N_14831);
nand UO_1184 (O_1184,N_14861,N_14924);
nor UO_1185 (O_1185,N_14761,N_14877);
and UO_1186 (O_1186,N_14885,N_14758);
nor UO_1187 (O_1187,N_14773,N_14824);
nand UO_1188 (O_1188,N_14921,N_14882);
and UO_1189 (O_1189,N_14878,N_14785);
and UO_1190 (O_1190,N_14928,N_14945);
nand UO_1191 (O_1191,N_14830,N_14853);
or UO_1192 (O_1192,N_14951,N_14789);
nand UO_1193 (O_1193,N_14811,N_14967);
nor UO_1194 (O_1194,N_14881,N_14915);
nand UO_1195 (O_1195,N_14750,N_14765);
xor UO_1196 (O_1196,N_14811,N_14820);
nand UO_1197 (O_1197,N_14832,N_14899);
xor UO_1198 (O_1198,N_14823,N_14943);
and UO_1199 (O_1199,N_14787,N_14951);
nor UO_1200 (O_1200,N_14989,N_14877);
and UO_1201 (O_1201,N_14890,N_14914);
or UO_1202 (O_1202,N_14779,N_14862);
or UO_1203 (O_1203,N_14805,N_14886);
nor UO_1204 (O_1204,N_14865,N_14841);
and UO_1205 (O_1205,N_14764,N_14811);
nand UO_1206 (O_1206,N_14870,N_14807);
nand UO_1207 (O_1207,N_14964,N_14936);
nand UO_1208 (O_1208,N_14773,N_14897);
and UO_1209 (O_1209,N_14758,N_14802);
xnor UO_1210 (O_1210,N_14918,N_14831);
xor UO_1211 (O_1211,N_14979,N_14803);
or UO_1212 (O_1212,N_14775,N_14887);
nor UO_1213 (O_1213,N_14793,N_14872);
xor UO_1214 (O_1214,N_14946,N_14863);
nor UO_1215 (O_1215,N_14978,N_14931);
and UO_1216 (O_1216,N_14793,N_14910);
or UO_1217 (O_1217,N_14829,N_14941);
nand UO_1218 (O_1218,N_14903,N_14854);
xor UO_1219 (O_1219,N_14786,N_14891);
nand UO_1220 (O_1220,N_14842,N_14756);
nor UO_1221 (O_1221,N_14964,N_14842);
xnor UO_1222 (O_1222,N_14812,N_14878);
nor UO_1223 (O_1223,N_14891,N_14819);
xor UO_1224 (O_1224,N_14814,N_14849);
and UO_1225 (O_1225,N_14956,N_14865);
or UO_1226 (O_1226,N_14816,N_14827);
nor UO_1227 (O_1227,N_14827,N_14843);
or UO_1228 (O_1228,N_14923,N_14989);
or UO_1229 (O_1229,N_14850,N_14911);
xor UO_1230 (O_1230,N_14762,N_14904);
and UO_1231 (O_1231,N_14996,N_14905);
or UO_1232 (O_1232,N_14789,N_14804);
nand UO_1233 (O_1233,N_14988,N_14851);
xnor UO_1234 (O_1234,N_14926,N_14800);
xnor UO_1235 (O_1235,N_14961,N_14787);
nand UO_1236 (O_1236,N_14936,N_14867);
nand UO_1237 (O_1237,N_14756,N_14932);
and UO_1238 (O_1238,N_14899,N_14946);
nor UO_1239 (O_1239,N_14789,N_14846);
nand UO_1240 (O_1240,N_14806,N_14911);
xnor UO_1241 (O_1241,N_14960,N_14859);
nor UO_1242 (O_1242,N_14861,N_14928);
xor UO_1243 (O_1243,N_14897,N_14914);
and UO_1244 (O_1244,N_14823,N_14989);
or UO_1245 (O_1245,N_14804,N_14907);
nor UO_1246 (O_1246,N_14925,N_14903);
or UO_1247 (O_1247,N_14880,N_14934);
nor UO_1248 (O_1248,N_14979,N_14982);
and UO_1249 (O_1249,N_14960,N_14967);
nor UO_1250 (O_1250,N_14975,N_14934);
nand UO_1251 (O_1251,N_14819,N_14972);
nor UO_1252 (O_1252,N_14791,N_14914);
and UO_1253 (O_1253,N_14750,N_14889);
xor UO_1254 (O_1254,N_14820,N_14832);
xnor UO_1255 (O_1255,N_14823,N_14806);
or UO_1256 (O_1256,N_14879,N_14845);
and UO_1257 (O_1257,N_14782,N_14845);
xnor UO_1258 (O_1258,N_14872,N_14820);
and UO_1259 (O_1259,N_14767,N_14900);
nand UO_1260 (O_1260,N_14990,N_14892);
xnor UO_1261 (O_1261,N_14899,N_14920);
nand UO_1262 (O_1262,N_14974,N_14796);
nand UO_1263 (O_1263,N_14830,N_14958);
and UO_1264 (O_1264,N_14807,N_14922);
nand UO_1265 (O_1265,N_14927,N_14791);
nor UO_1266 (O_1266,N_14836,N_14841);
and UO_1267 (O_1267,N_14757,N_14946);
nand UO_1268 (O_1268,N_14800,N_14898);
nor UO_1269 (O_1269,N_14845,N_14971);
nor UO_1270 (O_1270,N_14845,N_14844);
xnor UO_1271 (O_1271,N_14887,N_14797);
xor UO_1272 (O_1272,N_14989,N_14825);
xnor UO_1273 (O_1273,N_14969,N_14899);
nand UO_1274 (O_1274,N_14979,N_14919);
nand UO_1275 (O_1275,N_14912,N_14798);
xor UO_1276 (O_1276,N_14828,N_14820);
nand UO_1277 (O_1277,N_14937,N_14899);
xor UO_1278 (O_1278,N_14811,N_14859);
nor UO_1279 (O_1279,N_14936,N_14917);
or UO_1280 (O_1280,N_14787,N_14927);
nor UO_1281 (O_1281,N_14767,N_14884);
or UO_1282 (O_1282,N_14915,N_14985);
nor UO_1283 (O_1283,N_14926,N_14875);
and UO_1284 (O_1284,N_14988,N_14976);
xnor UO_1285 (O_1285,N_14954,N_14975);
xnor UO_1286 (O_1286,N_14946,N_14996);
or UO_1287 (O_1287,N_14880,N_14816);
and UO_1288 (O_1288,N_14916,N_14866);
xnor UO_1289 (O_1289,N_14779,N_14824);
and UO_1290 (O_1290,N_14897,N_14982);
nor UO_1291 (O_1291,N_14950,N_14873);
nor UO_1292 (O_1292,N_14764,N_14787);
or UO_1293 (O_1293,N_14863,N_14771);
and UO_1294 (O_1294,N_14923,N_14778);
xor UO_1295 (O_1295,N_14815,N_14786);
nand UO_1296 (O_1296,N_14873,N_14781);
xor UO_1297 (O_1297,N_14801,N_14816);
nand UO_1298 (O_1298,N_14807,N_14893);
nor UO_1299 (O_1299,N_14834,N_14881);
or UO_1300 (O_1300,N_14894,N_14946);
xnor UO_1301 (O_1301,N_14971,N_14763);
and UO_1302 (O_1302,N_14865,N_14826);
or UO_1303 (O_1303,N_14904,N_14863);
and UO_1304 (O_1304,N_14752,N_14767);
or UO_1305 (O_1305,N_14865,N_14984);
xor UO_1306 (O_1306,N_14875,N_14802);
or UO_1307 (O_1307,N_14750,N_14864);
or UO_1308 (O_1308,N_14924,N_14862);
and UO_1309 (O_1309,N_14965,N_14905);
and UO_1310 (O_1310,N_14907,N_14928);
or UO_1311 (O_1311,N_14991,N_14965);
and UO_1312 (O_1312,N_14989,N_14904);
and UO_1313 (O_1313,N_14824,N_14961);
nor UO_1314 (O_1314,N_14770,N_14756);
xnor UO_1315 (O_1315,N_14871,N_14791);
nor UO_1316 (O_1316,N_14878,N_14803);
nand UO_1317 (O_1317,N_14934,N_14936);
xor UO_1318 (O_1318,N_14842,N_14889);
xnor UO_1319 (O_1319,N_14916,N_14960);
xor UO_1320 (O_1320,N_14828,N_14766);
and UO_1321 (O_1321,N_14785,N_14790);
nand UO_1322 (O_1322,N_14802,N_14832);
and UO_1323 (O_1323,N_14773,N_14874);
nand UO_1324 (O_1324,N_14999,N_14917);
or UO_1325 (O_1325,N_14807,N_14883);
xor UO_1326 (O_1326,N_14772,N_14811);
nor UO_1327 (O_1327,N_14808,N_14768);
and UO_1328 (O_1328,N_14852,N_14895);
and UO_1329 (O_1329,N_14963,N_14957);
nor UO_1330 (O_1330,N_14961,N_14812);
or UO_1331 (O_1331,N_14764,N_14932);
or UO_1332 (O_1332,N_14868,N_14909);
and UO_1333 (O_1333,N_14890,N_14817);
or UO_1334 (O_1334,N_14781,N_14996);
or UO_1335 (O_1335,N_14939,N_14906);
nor UO_1336 (O_1336,N_14849,N_14796);
and UO_1337 (O_1337,N_14944,N_14862);
nand UO_1338 (O_1338,N_14890,N_14798);
and UO_1339 (O_1339,N_14814,N_14975);
nor UO_1340 (O_1340,N_14892,N_14793);
and UO_1341 (O_1341,N_14899,N_14973);
xnor UO_1342 (O_1342,N_14842,N_14981);
or UO_1343 (O_1343,N_14757,N_14947);
or UO_1344 (O_1344,N_14862,N_14885);
nand UO_1345 (O_1345,N_14761,N_14797);
and UO_1346 (O_1346,N_14927,N_14958);
or UO_1347 (O_1347,N_14906,N_14866);
nand UO_1348 (O_1348,N_14941,N_14914);
xnor UO_1349 (O_1349,N_14798,N_14917);
nand UO_1350 (O_1350,N_14846,N_14852);
or UO_1351 (O_1351,N_14874,N_14819);
nand UO_1352 (O_1352,N_14869,N_14890);
xnor UO_1353 (O_1353,N_14842,N_14869);
or UO_1354 (O_1354,N_14954,N_14947);
nand UO_1355 (O_1355,N_14874,N_14891);
and UO_1356 (O_1356,N_14839,N_14898);
or UO_1357 (O_1357,N_14912,N_14851);
and UO_1358 (O_1358,N_14980,N_14830);
and UO_1359 (O_1359,N_14778,N_14781);
nor UO_1360 (O_1360,N_14871,N_14857);
nor UO_1361 (O_1361,N_14770,N_14773);
xnor UO_1362 (O_1362,N_14893,N_14866);
xor UO_1363 (O_1363,N_14780,N_14782);
xnor UO_1364 (O_1364,N_14759,N_14824);
and UO_1365 (O_1365,N_14927,N_14902);
and UO_1366 (O_1366,N_14841,N_14753);
xor UO_1367 (O_1367,N_14878,N_14962);
nor UO_1368 (O_1368,N_14886,N_14827);
and UO_1369 (O_1369,N_14857,N_14922);
xor UO_1370 (O_1370,N_14778,N_14958);
and UO_1371 (O_1371,N_14943,N_14941);
xnor UO_1372 (O_1372,N_14858,N_14977);
or UO_1373 (O_1373,N_14957,N_14975);
xor UO_1374 (O_1374,N_14794,N_14769);
or UO_1375 (O_1375,N_14985,N_14798);
and UO_1376 (O_1376,N_14833,N_14827);
or UO_1377 (O_1377,N_14803,N_14836);
nor UO_1378 (O_1378,N_14785,N_14991);
and UO_1379 (O_1379,N_14860,N_14779);
xnor UO_1380 (O_1380,N_14863,N_14953);
xnor UO_1381 (O_1381,N_14887,N_14932);
or UO_1382 (O_1382,N_14837,N_14827);
nor UO_1383 (O_1383,N_14963,N_14860);
and UO_1384 (O_1384,N_14859,N_14756);
xor UO_1385 (O_1385,N_14854,N_14862);
xnor UO_1386 (O_1386,N_14778,N_14859);
xnor UO_1387 (O_1387,N_14839,N_14976);
or UO_1388 (O_1388,N_14822,N_14870);
xnor UO_1389 (O_1389,N_14930,N_14824);
xnor UO_1390 (O_1390,N_14877,N_14869);
or UO_1391 (O_1391,N_14785,N_14918);
and UO_1392 (O_1392,N_14968,N_14867);
and UO_1393 (O_1393,N_14974,N_14950);
nand UO_1394 (O_1394,N_14975,N_14845);
nand UO_1395 (O_1395,N_14798,N_14945);
or UO_1396 (O_1396,N_14846,N_14861);
xor UO_1397 (O_1397,N_14911,N_14826);
nor UO_1398 (O_1398,N_14980,N_14982);
nand UO_1399 (O_1399,N_14856,N_14871);
and UO_1400 (O_1400,N_14790,N_14857);
xor UO_1401 (O_1401,N_14947,N_14843);
nand UO_1402 (O_1402,N_14868,N_14999);
nand UO_1403 (O_1403,N_14755,N_14855);
and UO_1404 (O_1404,N_14764,N_14954);
or UO_1405 (O_1405,N_14910,N_14892);
nand UO_1406 (O_1406,N_14789,N_14831);
nand UO_1407 (O_1407,N_14901,N_14758);
and UO_1408 (O_1408,N_14763,N_14906);
nor UO_1409 (O_1409,N_14819,N_14946);
and UO_1410 (O_1410,N_14897,N_14877);
xnor UO_1411 (O_1411,N_14814,N_14883);
nor UO_1412 (O_1412,N_14835,N_14911);
nor UO_1413 (O_1413,N_14819,N_14928);
and UO_1414 (O_1414,N_14844,N_14921);
and UO_1415 (O_1415,N_14989,N_14773);
nor UO_1416 (O_1416,N_14874,N_14848);
nor UO_1417 (O_1417,N_14898,N_14873);
or UO_1418 (O_1418,N_14988,N_14984);
xnor UO_1419 (O_1419,N_14803,N_14797);
nand UO_1420 (O_1420,N_14910,N_14754);
or UO_1421 (O_1421,N_14847,N_14922);
nand UO_1422 (O_1422,N_14827,N_14879);
nor UO_1423 (O_1423,N_14885,N_14879);
xor UO_1424 (O_1424,N_14972,N_14886);
xnor UO_1425 (O_1425,N_14987,N_14940);
and UO_1426 (O_1426,N_14767,N_14990);
and UO_1427 (O_1427,N_14956,N_14911);
or UO_1428 (O_1428,N_14780,N_14987);
or UO_1429 (O_1429,N_14985,N_14955);
nand UO_1430 (O_1430,N_14822,N_14818);
xor UO_1431 (O_1431,N_14793,N_14754);
xor UO_1432 (O_1432,N_14885,N_14910);
nand UO_1433 (O_1433,N_14992,N_14960);
or UO_1434 (O_1434,N_14991,N_14812);
xnor UO_1435 (O_1435,N_14827,N_14905);
xor UO_1436 (O_1436,N_14955,N_14779);
or UO_1437 (O_1437,N_14770,N_14938);
xor UO_1438 (O_1438,N_14813,N_14948);
or UO_1439 (O_1439,N_14830,N_14944);
nand UO_1440 (O_1440,N_14925,N_14787);
nor UO_1441 (O_1441,N_14945,N_14805);
nor UO_1442 (O_1442,N_14773,N_14950);
or UO_1443 (O_1443,N_14980,N_14986);
or UO_1444 (O_1444,N_14984,N_14899);
xor UO_1445 (O_1445,N_14905,N_14900);
nor UO_1446 (O_1446,N_14880,N_14882);
nand UO_1447 (O_1447,N_14904,N_14944);
nor UO_1448 (O_1448,N_14877,N_14813);
nand UO_1449 (O_1449,N_14781,N_14785);
nor UO_1450 (O_1450,N_14880,N_14964);
and UO_1451 (O_1451,N_14869,N_14935);
xor UO_1452 (O_1452,N_14952,N_14765);
or UO_1453 (O_1453,N_14755,N_14757);
xnor UO_1454 (O_1454,N_14877,N_14948);
nor UO_1455 (O_1455,N_14847,N_14807);
xor UO_1456 (O_1456,N_14949,N_14880);
or UO_1457 (O_1457,N_14996,N_14993);
nor UO_1458 (O_1458,N_14924,N_14972);
or UO_1459 (O_1459,N_14868,N_14894);
nand UO_1460 (O_1460,N_14828,N_14795);
nand UO_1461 (O_1461,N_14769,N_14812);
nor UO_1462 (O_1462,N_14975,N_14998);
or UO_1463 (O_1463,N_14838,N_14854);
xor UO_1464 (O_1464,N_14948,N_14993);
xnor UO_1465 (O_1465,N_14780,N_14811);
nand UO_1466 (O_1466,N_14920,N_14867);
nand UO_1467 (O_1467,N_14997,N_14808);
nand UO_1468 (O_1468,N_14827,N_14850);
nand UO_1469 (O_1469,N_14864,N_14759);
xor UO_1470 (O_1470,N_14794,N_14931);
nor UO_1471 (O_1471,N_14758,N_14984);
xor UO_1472 (O_1472,N_14915,N_14830);
xnor UO_1473 (O_1473,N_14919,N_14784);
xnor UO_1474 (O_1474,N_14959,N_14947);
nand UO_1475 (O_1475,N_14967,N_14849);
or UO_1476 (O_1476,N_14803,N_14951);
xor UO_1477 (O_1477,N_14856,N_14775);
and UO_1478 (O_1478,N_14850,N_14809);
xor UO_1479 (O_1479,N_14847,N_14949);
nor UO_1480 (O_1480,N_14910,N_14958);
and UO_1481 (O_1481,N_14917,N_14916);
nor UO_1482 (O_1482,N_14934,N_14978);
or UO_1483 (O_1483,N_14872,N_14880);
nand UO_1484 (O_1484,N_14834,N_14992);
or UO_1485 (O_1485,N_14938,N_14893);
or UO_1486 (O_1486,N_14890,N_14821);
nor UO_1487 (O_1487,N_14759,N_14926);
and UO_1488 (O_1488,N_14943,N_14873);
nand UO_1489 (O_1489,N_14838,N_14891);
and UO_1490 (O_1490,N_14816,N_14846);
or UO_1491 (O_1491,N_14923,N_14895);
nor UO_1492 (O_1492,N_14940,N_14790);
xor UO_1493 (O_1493,N_14802,N_14821);
or UO_1494 (O_1494,N_14827,N_14856);
nor UO_1495 (O_1495,N_14909,N_14955);
nor UO_1496 (O_1496,N_14920,N_14844);
or UO_1497 (O_1497,N_14969,N_14777);
nand UO_1498 (O_1498,N_14980,N_14863);
or UO_1499 (O_1499,N_14906,N_14764);
nand UO_1500 (O_1500,N_14879,N_14849);
or UO_1501 (O_1501,N_14833,N_14813);
or UO_1502 (O_1502,N_14914,N_14774);
or UO_1503 (O_1503,N_14811,N_14985);
nor UO_1504 (O_1504,N_14847,N_14978);
nor UO_1505 (O_1505,N_14894,N_14813);
nand UO_1506 (O_1506,N_14892,N_14801);
nand UO_1507 (O_1507,N_14878,N_14994);
or UO_1508 (O_1508,N_14870,N_14964);
xor UO_1509 (O_1509,N_14788,N_14986);
or UO_1510 (O_1510,N_14823,N_14899);
nor UO_1511 (O_1511,N_14773,N_14855);
and UO_1512 (O_1512,N_14834,N_14944);
nand UO_1513 (O_1513,N_14752,N_14895);
or UO_1514 (O_1514,N_14851,N_14873);
xor UO_1515 (O_1515,N_14839,N_14891);
or UO_1516 (O_1516,N_14772,N_14840);
nor UO_1517 (O_1517,N_14968,N_14975);
and UO_1518 (O_1518,N_14789,N_14926);
and UO_1519 (O_1519,N_14817,N_14882);
and UO_1520 (O_1520,N_14759,N_14861);
nor UO_1521 (O_1521,N_14757,N_14917);
nor UO_1522 (O_1522,N_14851,N_14891);
or UO_1523 (O_1523,N_14913,N_14968);
or UO_1524 (O_1524,N_14937,N_14892);
or UO_1525 (O_1525,N_14795,N_14883);
nand UO_1526 (O_1526,N_14851,N_14949);
nand UO_1527 (O_1527,N_14841,N_14977);
and UO_1528 (O_1528,N_14905,N_14906);
and UO_1529 (O_1529,N_14899,N_14775);
and UO_1530 (O_1530,N_14761,N_14840);
nor UO_1531 (O_1531,N_14884,N_14905);
or UO_1532 (O_1532,N_14803,N_14784);
nand UO_1533 (O_1533,N_14763,N_14750);
nand UO_1534 (O_1534,N_14837,N_14811);
or UO_1535 (O_1535,N_14919,N_14800);
and UO_1536 (O_1536,N_14862,N_14967);
and UO_1537 (O_1537,N_14997,N_14983);
or UO_1538 (O_1538,N_14772,N_14767);
nor UO_1539 (O_1539,N_14995,N_14908);
nor UO_1540 (O_1540,N_14929,N_14952);
nand UO_1541 (O_1541,N_14805,N_14951);
nor UO_1542 (O_1542,N_14852,N_14937);
xor UO_1543 (O_1543,N_14803,N_14906);
xor UO_1544 (O_1544,N_14881,N_14765);
xnor UO_1545 (O_1545,N_14834,N_14925);
and UO_1546 (O_1546,N_14811,N_14890);
or UO_1547 (O_1547,N_14999,N_14934);
nor UO_1548 (O_1548,N_14751,N_14818);
and UO_1549 (O_1549,N_14938,N_14848);
or UO_1550 (O_1550,N_14854,N_14837);
and UO_1551 (O_1551,N_14929,N_14830);
xnor UO_1552 (O_1552,N_14991,N_14908);
and UO_1553 (O_1553,N_14757,N_14839);
xnor UO_1554 (O_1554,N_14897,N_14802);
nor UO_1555 (O_1555,N_14891,N_14896);
nor UO_1556 (O_1556,N_14877,N_14873);
nor UO_1557 (O_1557,N_14964,N_14955);
or UO_1558 (O_1558,N_14908,N_14839);
nor UO_1559 (O_1559,N_14898,N_14886);
xor UO_1560 (O_1560,N_14794,N_14878);
xor UO_1561 (O_1561,N_14978,N_14841);
nand UO_1562 (O_1562,N_14960,N_14924);
xor UO_1563 (O_1563,N_14918,N_14834);
and UO_1564 (O_1564,N_14973,N_14958);
and UO_1565 (O_1565,N_14963,N_14879);
xor UO_1566 (O_1566,N_14771,N_14834);
or UO_1567 (O_1567,N_14978,N_14883);
or UO_1568 (O_1568,N_14815,N_14913);
and UO_1569 (O_1569,N_14759,N_14780);
nor UO_1570 (O_1570,N_14856,N_14883);
or UO_1571 (O_1571,N_14980,N_14949);
or UO_1572 (O_1572,N_14916,N_14948);
and UO_1573 (O_1573,N_14857,N_14779);
xor UO_1574 (O_1574,N_14842,N_14835);
nor UO_1575 (O_1575,N_14897,N_14873);
or UO_1576 (O_1576,N_14835,N_14943);
or UO_1577 (O_1577,N_14844,N_14991);
xnor UO_1578 (O_1578,N_14911,N_14795);
and UO_1579 (O_1579,N_14784,N_14752);
xnor UO_1580 (O_1580,N_14943,N_14866);
or UO_1581 (O_1581,N_14965,N_14834);
nor UO_1582 (O_1582,N_14840,N_14975);
nand UO_1583 (O_1583,N_14892,N_14797);
nand UO_1584 (O_1584,N_14790,N_14976);
or UO_1585 (O_1585,N_14894,N_14959);
nand UO_1586 (O_1586,N_14789,N_14919);
and UO_1587 (O_1587,N_14859,N_14868);
or UO_1588 (O_1588,N_14820,N_14989);
nor UO_1589 (O_1589,N_14988,N_14906);
nor UO_1590 (O_1590,N_14946,N_14958);
nor UO_1591 (O_1591,N_14759,N_14876);
nor UO_1592 (O_1592,N_14995,N_14944);
and UO_1593 (O_1593,N_14881,N_14846);
nor UO_1594 (O_1594,N_14888,N_14919);
or UO_1595 (O_1595,N_14804,N_14840);
nand UO_1596 (O_1596,N_14870,N_14767);
nor UO_1597 (O_1597,N_14916,N_14991);
and UO_1598 (O_1598,N_14934,N_14817);
or UO_1599 (O_1599,N_14857,N_14997);
xnor UO_1600 (O_1600,N_14827,N_14991);
or UO_1601 (O_1601,N_14880,N_14982);
or UO_1602 (O_1602,N_14974,N_14964);
nand UO_1603 (O_1603,N_14892,N_14856);
nor UO_1604 (O_1604,N_14868,N_14907);
xnor UO_1605 (O_1605,N_14764,N_14837);
nand UO_1606 (O_1606,N_14900,N_14875);
and UO_1607 (O_1607,N_14902,N_14952);
or UO_1608 (O_1608,N_14790,N_14818);
and UO_1609 (O_1609,N_14780,N_14808);
nand UO_1610 (O_1610,N_14911,N_14923);
or UO_1611 (O_1611,N_14833,N_14764);
nor UO_1612 (O_1612,N_14882,N_14923);
or UO_1613 (O_1613,N_14806,N_14961);
and UO_1614 (O_1614,N_14980,N_14828);
and UO_1615 (O_1615,N_14884,N_14860);
xnor UO_1616 (O_1616,N_14867,N_14951);
and UO_1617 (O_1617,N_14791,N_14936);
and UO_1618 (O_1618,N_14978,N_14860);
and UO_1619 (O_1619,N_14888,N_14985);
and UO_1620 (O_1620,N_14969,N_14998);
xor UO_1621 (O_1621,N_14772,N_14886);
nand UO_1622 (O_1622,N_14848,N_14771);
and UO_1623 (O_1623,N_14902,N_14787);
nor UO_1624 (O_1624,N_14961,N_14799);
nand UO_1625 (O_1625,N_14971,N_14776);
or UO_1626 (O_1626,N_14808,N_14940);
or UO_1627 (O_1627,N_14877,N_14849);
xnor UO_1628 (O_1628,N_14770,N_14794);
nor UO_1629 (O_1629,N_14982,N_14940);
and UO_1630 (O_1630,N_14859,N_14924);
xor UO_1631 (O_1631,N_14829,N_14973);
nand UO_1632 (O_1632,N_14898,N_14889);
or UO_1633 (O_1633,N_14803,N_14908);
nor UO_1634 (O_1634,N_14913,N_14777);
nand UO_1635 (O_1635,N_14832,N_14935);
nand UO_1636 (O_1636,N_14803,N_14964);
and UO_1637 (O_1637,N_14834,N_14754);
nand UO_1638 (O_1638,N_14924,N_14784);
nor UO_1639 (O_1639,N_14999,N_14977);
nor UO_1640 (O_1640,N_14842,N_14910);
or UO_1641 (O_1641,N_14758,N_14878);
nand UO_1642 (O_1642,N_14785,N_14964);
nor UO_1643 (O_1643,N_14945,N_14754);
nor UO_1644 (O_1644,N_14862,N_14853);
nor UO_1645 (O_1645,N_14991,N_14836);
nor UO_1646 (O_1646,N_14852,N_14872);
xnor UO_1647 (O_1647,N_14893,N_14759);
nand UO_1648 (O_1648,N_14959,N_14949);
nor UO_1649 (O_1649,N_14908,N_14889);
and UO_1650 (O_1650,N_14755,N_14866);
nor UO_1651 (O_1651,N_14899,N_14761);
nand UO_1652 (O_1652,N_14948,N_14781);
nand UO_1653 (O_1653,N_14884,N_14944);
and UO_1654 (O_1654,N_14849,N_14910);
xor UO_1655 (O_1655,N_14837,N_14800);
and UO_1656 (O_1656,N_14857,N_14813);
or UO_1657 (O_1657,N_14806,N_14898);
nor UO_1658 (O_1658,N_14796,N_14997);
or UO_1659 (O_1659,N_14900,N_14954);
nor UO_1660 (O_1660,N_14788,N_14958);
and UO_1661 (O_1661,N_14939,N_14805);
nand UO_1662 (O_1662,N_14772,N_14987);
or UO_1663 (O_1663,N_14932,N_14824);
xnor UO_1664 (O_1664,N_14953,N_14789);
and UO_1665 (O_1665,N_14927,N_14878);
nand UO_1666 (O_1666,N_14973,N_14814);
nor UO_1667 (O_1667,N_14780,N_14819);
or UO_1668 (O_1668,N_14849,N_14765);
xnor UO_1669 (O_1669,N_14975,N_14959);
xor UO_1670 (O_1670,N_14899,N_14924);
and UO_1671 (O_1671,N_14900,N_14912);
or UO_1672 (O_1672,N_14900,N_14924);
or UO_1673 (O_1673,N_14757,N_14906);
nor UO_1674 (O_1674,N_14759,N_14925);
nor UO_1675 (O_1675,N_14805,N_14871);
or UO_1676 (O_1676,N_14993,N_14988);
or UO_1677 (O_1677,N_14835,N_14912);
and UO_1678 (O_1678,N_14923,N_14885);
and UO_1679 (O_1679,N_14762,N_14984);
and UO_1680 (O_1680,N_14905,N_14788);
xor UO_1681 (O_1681,N_14818,N_14909);
nor UO_1682 (O_1682,N_14796,N_14820);
nor UO_1683 (O_1683,N_14992,N_14774);
nand UO_1684 (O_1684,N_14909,N_14761);
nor UO_1685 (O_1685,N_14819,N_14970);
and UO_1686 (O_1686,N_14862,N_14776);
or UO_1687 (O_1687,N_14896,N_14803);
xor UO_1688 (O_1688,N_14779,N_14848);
or UO_1689 (O_1689,N_14834,N_14947);
or UO_1690 (O_1690,N_14995,N_14988);
xnor UO_1691 (O_1691,N_14929,N_14837);
or UO_1692 (O_1692,N_14878,N_14889);
xor UO_1693 (O_1693,N_14909,N_14946);
or UO_1694 (O_1694,N_14869,N_14880);
and UO_1695 (O_1695,N_14895,N_14836);
nor UO_1696 (O_1696,N_14856,N_14931);
nand UO_1697 (O_1697,N_14964,N_14943);
nor UO_1698 (O_1698,N_14879,N_14814);
nand UO_1699 (O_1699,N_14847,N_14757);
nand UO_1700 (O_1700,N_14925,N_14839);
and UO_1701 (O_1701,N_14763,N_14878);
xnor UO_1702 (O_1702,N_14858,N_14958);
and UO_1703 (O_1703,N_14987,N_14880);
or UO_1704 (O_1704,N_14875,N_14811);
or UO_1705 (O_1705,N_14897,N_14812);
and UO_1706 (O_1706,N_14911,N_14852);
or UO_1707 (O_1707,N_14898,N_14932);
nand UO_1708 (O_1708,N_14914,N_14760);
or UO_1709 (O_1709,N_14920,N_14828);
nand UO_1710 (O_1710,N_14958,N_14895);
xnor UO_1711 (O_1711,N_14957,N_14943);
xor UO_1712 (O_1712,N_14988,N_14957);
and UO_1713 (O_1713,N_14861,N_14949);
and UO_1714 (O_1714,N_14924,N_14926);
nand UO_1715 (O_1715,N_14978,N_14825);
or UO_1716 (O_1716,N_14755,N_14764);
nand UO_1717 (O_1717,N_14853,N_14917);
nor UO_1718 (O_1718,N_14802,N_14794);
or UO_1719 (O_1719,N_14793,N_14795);
or UO_1720 (O_1720,N_14984,N_14967);
or UO_1721 (O_1721,N_14768,N_14842);
and UO_1722 (O_1722,N_14780,N_14977);
and UO_1723 (O_1723,N_14950,N_14777);
xnor UO_1724 (O_1724,N_14876,N_14784);
nor UO_1725 (O_1725,N_14856,N_14921);
xor UO_1726 (O_1726,N_14954,N_14867);
nor UO_1727 (O_1727,N_14834,N_14968);
and UO_1728 (O_1728,N_14833,N_14930);
and UO_1729 (O_1729,N_14767,N_14804);
or UO_1730 (O_1730,N_14769,N_14971);
xnor UO_1731 (O_1731,N_14958,N_14994);
and UO_1732 (O_1732,N_14915,N_14978);
and UO_1733 (O_1733,N_14829,N_14794);
and UO_1734 (O_1734,N_14922,N_14966);
xor UO_1735 (O_1735,N_14887,N_14920);
or UO_1736 (O_1736,N_14821,N_14773);
xor UO_1737 (O_1737,N_14760,N_14972);
nand UO_1738 (O_1738,N_14788,N_14870);
and UO_1739 (O_1739,N_14866,N_14948);
xnor UO_1740 (O_1740,N_14910,N_14893);
nand UO_1741 (O_1741,N_14970,N_14882);
xnor UO_1742 (O_1742,N_14883,N_14800);
or UO_1743 (O_1743,N_14882,N_14931);
nor UO_1744 (O_1744,N_14790,N_14774);
xor UO_1745 (O_1745,N_14810,N_14919);
nand UO_1746 (O_1746,N_14849,N_14993);
or UO_1747 (O_1747,N_14947,N_14766);
and UO_1748 (O_1748,N_14759,N_14986);
and UO_1749 (O_1749,N_14939,N_14757);
nor UO_1750 (O_1750,N_14791,N_14860);
and UO_1751 (O_1751,N_14947,N_14793);
or UO_1752 (O_1752,N_14938,N_14805);
and UO_1753 (O_1753,N_14941,N_14987);
or UO_1754 (O_1754,N_14829,N_14868);
xor UO_1755 (O_1755,N_14871,N_14870);
and UO_1756 (O_1756,N_14767,N_14880);
xnor UO_1757 (O_1757,N_14752,N_14937);
and UO_1758 (O_1758,N_14792,N_14976);
or UO_1759 (O_1759,N_14940,N_14774);
nand UO_1760 (O_1760,N_14780,N_14995);
nor UO_1761 (O_1761,N_14794,N_14800);
or UO_1762 (O_1762,N_14868,N_14958);
or UO_1763 (O_1763,N_14786,N_14846);
and UO_1764 (O_1764,N_14914,N_14750);
nand UO_1765 (O_1765,N_14943,N_14768);
nor UO_1766 (O_1766,N_14773,N_14891);
or UO_1767 (O_1767,N_14824,N_14835);
and UO_1768 (O_1768,N_14892,N_14780);
nor UO_1769 (O_1769,N_14997,N_14777);
or UO_1770 (O_1770,N_14921,N_14805);
nand UO_1771 (O_1771,N_14906,N_14942);
nand UO_1772 (O_1772,N_14846,N_14790);
nor UO_1773 (O_1773,N_14921,N_14911);
nor UO_1774 (O_1774,N_14928,N_14773);
nand UO_1775 (O_1775,N_14791,N_14979);
or UO_1776 (O_1776,N_14987,N_14936);
and UO_1777 (O_1777,N_14803,N_14959);
and UO_1778 (O_1778,N_14968,N_14781);
xor UO_1779 (O_1779,N_14927,N_14879);
nor UO_1780 (O_1780,N_14987,N_14844);
or UO_1781 (O_1781,N_14912,N_14905);
xnor UO_1782 (O_1782,N_14879,N_14950);
and UO_1783 (O_1783,N_14755,N_14781);
and UO_1784 (O_1784,N_14956,N_14757);
and UO_1785 (O_1785,N_14969,N_14804);
xnor UO_1786 (O_1786,N_14896,N_14771);
nor UO_1787 (O_1787,N_14838,N_14962);
nor UO_1788 (O_1788,N_14757,N_14843);
and UO_1789 (O_1789,N_14878,N_14764);
nor UO_1790 (O_1790,N_14895,N_14953);
and UO_1791 (O_1791,N_14851,N_14854);
nor UO_1792 (O_1792,N_14811,N_14769);
nand UO_1793 (O_1793,N_14752,N_14914);
nand UO_1794 (O_1794,N_14998,N_14910);
xor UO_1795 (O_1795,N_14777,N_14861);
and UO_1796 (O_1796,N_14991,N_14820);
nor UO_1797 (O_1797,N_14816,N_14976);
and UO_1798 (O_1798,N_14881,N_14898);
xor UO_1799 (O_1799,N_14819,N_14808);
and UO_1800 (O_1800,N_14941,N_14843);
and UO_1801 (O_1801,N_14922,N_14885);
xor UO_1802 (O_1802,N_14969,N_14782);
or UO_1803 (O_1803,N_14885,N_14974);
nand UO_1804 (O_1804,N_14771,N_14788);
xor UO_1805 (O_1805,N_14815,N_14964);
xor UO_1806 (O_1806,N_14854,N_14812);
nor UO_1807 (O_1807,N_14981,N_14978);
xnor UO_1808 (O_1808,N_14867,N_14953);
nand UO_1809 (O_1809,N_14995,N_14927);
xor UO_1810 (O_1810,N_14949,N_14997);
nor UO_1811 (O_1811,N_14863,N_14773);
or UO_1812 (O_1812,N_14973,N_14977);
nand UO_1813 (O_1813,N_14753,N_14984);
nand UO_1814 (O_1814,N_14976,N_14756);
xnor UO_1815 (O_1815,N_14990,N_14773);
or UO_1816 (O_1816,N_14867,N_14901);
xnor UO_1817 (O_1817,N_14936,N_14863);
or UO_1818 (O_1818,N_14956,N_14860);
or UO_1819 (O_1819,N_14897,N_14755);
nor UO_1820 (O_1820,N_14910,N_14963);
or UO_1821 (O_1821,N_14984,N_14850);
xor UO_1822 (O_1822,N_14832,N_14817);
xor UO_1823 (O_1823,N_14849,N_14984);
and UO_1824 (O_1824,N_14991,N_14786);
xnor UO_1825 (O_1825,N_14813,N_14929);
xnor UO_1826 (O_1826,N_14833,N_14845);
nand UO_1827 (O_1827,N_14947,N_14971);
nand UO_1828 (O_1828,N_14886,N_14954);
or UO_1829 (O_1829,N_14821,N_14949);
nor UO_1830 (O_1830,N_14977,N_14777);
or UO_1831 (O_1831,N_14916,N_14972);
xnor UO_1832 (O_1832,N_14895,N_14799);
and UO_1833 (O_1833,N_14989,N_14807);
and UO_1834 (O_1834,N_14941,N_14887);
and UO_1835 (O_1835,N_14766,N_14984);
nor UO_1836 (O_1836,N_14890,N_14799);
nor UO_1837 (O_1837,N_14929,N_14975);
xor UO_1838 (O_1838,N_14799,N_14914);
nor UO_1839 (O_1839,N_14997,N_14899);
and UO_1840 (O_1840,N_14857,N_14958);
nor UO_1841 (O_1841,N_14975,N_14750);
or UO_1842 (O_1842,N_14794,N_14822);
or UO_1843 (O_1843,N_14797,N_14790);
xnor UO_1844 (O_1844,N_14980,N_14959);
nor UO_1845 (O_1845,N_14967,N_14996);
nand UO_1846 (O_1846,N_14777,N_14840);
or UO_1847 (O_1847,N_14761,N_14904);
and UO_1848 (O_1848,N_14794,N_14925);
xnor UO_1849 (O_1849,N_14800,N_14938);
nor UO_1850 (O_1850,N_14923,N_14809);
xor UO_1851 (O_1851,N_14774,N_14798);
or UO_1852 (O_1852,N_14957,N_14870);
nor UO_1853 (O_1853,N_14933,N_14909);
xnor UO_1854 (O_1854,N_14917,N_14773);
xor UO_1855 (O_1855,N_14815,N_14876);
and UO_1856 (O_1856,N_14887,N_14790);
or UO_1857 (O_1857,N_14918,N_14917);
xnor UO_1858 (O_1858,N_14835,N_14810);
nand UO_1859 (O_1859,N_14926,N_14816);
xnor UO_1860 (O_1860,N_14797,N_14774);
and UO_1861 (O_1861,N_14934,N_14797);
nor UO_1862 (O_1862,N_14927,N_14837);
or UO_1863 (O_1863,N_14864,N_14952);
nand UO_1864 (O_1864,N_14849,N_14941);
and UO_1865 (O_1865,N_14980,N_14768);
nor UO_1866 (O_1866,N_14767,N_14863);
and UO_1867 (O_1867,N_14872,N_14928);
nand UO_1868 (O_1868,N_14862,N_14812);
nand UO_1869 (O_1869,N_14839,N_14934);
xnor UO_1870 (O_1870,N_14825,N_14794);
nor UO_1871 (O_1871,N_14966,N_14978);
or UO_1872 (O_1872,N_14976,N_14928);
or UO_1873 (O_1873,N_14839,N_14961);
nand UO_1874 (O_1874,N_14977,N_14845);
nor UO_1875 (O_1875,N_14814,N_14813);
nand UO_1876 (O_1876,N_14960,N_14794);
nor UO_1877 (O_1877,N_14822,N_14790);
and UO_1878 (O_1878,N_14874,N_14945);
nand UO_1879 (O_1879,N_14922,N_14992);
and UO_1880 (O_1880,N_14823,N_14857);
and UO_1881 (O_1881,N_14899,N_14788);
xor UO_1882 (O_1882,N_14761,N_14850);
nand UO_1883 (O_1883,N_14987,N_14896);
nor UO_1884 (O_1884,N_14756,N_14963);
xnor UO_1885 (O_1885,N_14985,N_14859);
nand UO_1886 (O_1886,N_14768,N_14863);
nand UO_1887 (O_1887,N_14774,N_14848);
nand UO_1888 (O_1888,N_14788,N_14860);
or UO_1889 (O_1889,N_14893,N_14932);
nand UO_1890 (O_1890,N_14856,N_14916);
nor UO_1891 (O_1891,N_14936,N_14954);
nand UO_1892 (O_1892,N_14758,N_14754);
nand UO_1893 (O_1893,N_14767,N_14916);
or UO_1894 (O_1894,N_14854,N_14866);
and UO_1895 (O_1895,N_14863,N_14775);
nor UO_1896 (O_1896,N_14832,N_14891);
or UO_1897 (O_1897,N_14816,N_14849);
nand UO_1898 (O_1898,N_14857,N_14959);
nand UO_1899 (O_1899,N_14850,N_14913);
nor UO_1900 (O_1900,N_14826,N_14779);
or UO_1901 (O_1901,N_14880,N_14953);
nor UO_1902 (O_1902,N_14853,N_14833);
nand UO_1903 (O_1903,N_14951,N_14871);
and UO_1904 (O_1904,N_14970,N_14939);
or UO_1905 (O_1905,N_14881,N_14946);
nand UO_1906 (O_1906,N_14941,N_14792);
nand UO_1907 (O_1907,N_14917,N_14837);
nand UO_1908 (O_1908,N_14912,N_14967);
or UO_1909 (O_1909,N_14890,N_14778);
nor UO_1910 (O_1910,N_14815,N_14836);
nand UO_1911 (O_1911,N_14903,N_14884);
xor UO_1912 (O_1912,N_14905,N_14918);
xnor UO_1913 (O_1913,N_14801,N_14831);
and UO_1914 (O_1914,N_14776,N_14752);
or UO_1915 (O_1915,N_14916,N_14826);
and UO_1916 (O_1916,N_14797,N_14862);
nor UO_1917 (O_1917,N_14759,N_14868);
nand UO_1918 (O_1918,N_14802,N_14811);
or UO_1919 (O_1919,N_14759,N_14923);
and UO_1920 (O_1920,N_14998,N_14997);
nor UO_1921 (O_1921,N_14823,N_14983);
nor UO_1922 (O_1922,N_14830,N_14841);
xor UO_1923 (O_1923,N_14886,N_14941);
and UO_1924 (O_1924,N_14766,N_14781);
or UO_1925 (O_1925,N_14829,N_14796);
and UO_1926 (O_1926,N_14846,N_14959);
xor UO_1927 (O_1927,N_14823,N_14994);
xnor UO_1928 (O_1928,N_14946,N_14983);
nand UO_1929 (O_1929,N_14948,N_14983);
or UO_1930 (O_1930,N_14814,N_14961);
nand UO_1931 (O_1931,N_14882,N_14914);
nand UO_1932 (O_1932,N_14815,N_14805);
nand UO_1933 (O_1933,N_14973,N_14808);
and UO_1934 (O_1934,N_14901,N_14833);
and UO_1935 (O_1935,N_14756,N_14851);
and UO_1936 (O_1936,N_14971,N_14775);
nor UO_1937 (O_1937,N_14801,N_14913);
or UO_1938 (O_1938,N_14974,N_14785);
nor UO_1939 (O_1939,N_14882,N_14884);
and UO_1940 (O_1940,N_14885,N_14861);
nor UO_1941 (O_1941,N_14961,N_14882);
or UO_1942 (O_1942,N_14847,N_14926);
nand UO_1943 (O_1943,N_14855,N_14858);
and UO_1944 (O_1944,N_14795,N_14812);
nand UO_1945 (O_1945,N_14954,N_14919);
and UO_1946 (O_1946,N_14989,N_14924);
and UO_1947 (O_1947,N_14999,N_14915);
xor UO_1948 (O_1948,N_14936,N_14882);
nand UO_1949 (O_1949,N_14780,N_14968);
nand UO_1950 (O_1950,N_14822,N_14836);
xnor UO_1951 (O_1951,N_14856,N_14910);
and UO_1952 (O_1952,N_14981,N_14944);
and UO_1953 (O_1953,N_14976,N_14856);
and UO_1954 (O_1954,N_14876,N_14992);
or UO_1955 (O_1955,N_14804,N_14950);
xor UO_1956 (O_1956,N_14916,N_14762);
xnor UO_1957 (O_1957,N_14829,N_14803);
nand UO_1958 (O_1958,N_14940,N_14949);
nor UO_1959 (O_1959,N_14863,N_14945);
nor UO_1960 (O_1960,N_14850,N_14872);
and UO_1961 (O_1961,N_14959,N_14845);
nand UO_1962 (O_1962,N_14958,N_14767);
or UO_1963 (O_1963,N_14901,N_14874);
or UO_1964 (O_1964,N_14947,N_14848);
or UO_1965 (O_1965,N_14863,N_14941);
xor UO_1966 (O_1966,N_14969,N_14916);
nand UO_1967 (O_1967,N_14929,N_14901);
and UO_1968 (O_1968,N_14946,N_14893);
nand UO_1969 (O_1969,N_14962,N_14892);
xnor UO_1970 (O_1970,N_14863,N_14928);
nand UO_1971 (O_1971,N_14798,N_14782);
or UO_1972 (O_1972,N_14947,N_14961);
nand UO_1973 (O_1973,N_14855,N_14780);
nand UO_1974 (O_1974,N_14822,N_14948);
and UO_1975 (O_1975,N_14792,N_14934);
nor UO_1976 (O_1976,N_14990,N_14934);
xor UO_1977 (O_1977,N_14940,N_14841);
and UO_1978 (O_1978,N_14900,N_14970);
xor UO_1979 (O_1979,N_14948,N_14795);
nor UO_1980 (O_1980,N_14915,N_14768);
nor UO_1981 (O_1981,N_14884,N_14776);
nor UO_1982 (O_1982,N_14797,N_14800);
and UO_1983 (O_1983,N_14991,N_14931);
and UO_1984 (O_1984,N_14897,N_14790);
nand UO_1985 (O_1985,N_14981,N_14816);
and UO_1986 (O_1986,N_14847,N_14784);
nand UO_1987 (O_1987,N_14918,N_14885);
nand UO_1988 (O_1988,N_14918,N_14939);
nor UO_1989 (O_1989,N_14905,N_14935);
nor UO_1990 (O_1990,N_14907,N_14782);
or UO_1991 (O_1991,N_14874,N_14919);
nor UO_1992 (O_1992,N_14786,N_14754);
or UO_1993 (O_1993,N_14926,N_14952);
xnor UO_1994 (O_1994,N_14858,N_14851);
nand UO_1995 (O_1995,N_14791,N_14992);
and UO_1996 (O_1996,N_14833,N_14798);
nor UO_1997 (O_1997,N_14791,N_14868);
or UO_1998 (O_1998,N_14986,N_14774);
nand UO_1999 (O_1999,N_14791,N_14890);
endmodule