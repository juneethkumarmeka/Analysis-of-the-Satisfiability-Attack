module basic_1500_15000_2000_5_levels_2xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nor U0 (N_0,In_1195,In_1405);
or U1 (N_1,In_1,In_1110);
or U2 (N_2,In_1480,In_1228);
nor U3 (N_3,In_1011,In_981);
and U4 (N_4,In_622,In_793);
and U5 (N_5,In_1398,In_714);
nor U6 (N_6,In_781,In_1143);
nand U7 (N_7,In_1025,In_701);
or U8 (N_8,In_985,In_616);
and U9 (N_9,In_136,In_479);
or U10 (N_10,In_1274,In_1132);
and U11 (N_11,In_716,In_674);
nand U12 (N_12,In_1184,In_390);
nor U13 (N_13,In_445,In_1311);
or U14 (N_14,In_31,In_803);
and U15 (N_15,In_708,In_989);
nand U16 (N_16,In_9,In_417);
or U17 (N_17,In_867,In_896);
nor U18 (N_18,In_845,In_464);
or U19 (N_19,In_441,In_260);
or U20 (N_20,In_844,In_450);
nand U21 (N_21,In_1187,In_1083);
and U22 (N_22,In_1188,In_452);
nand U23 (N_23,In_94,In_992);
nor U24 (N_24,In_557,In_965);
or U25 (N_25,In_606,In_1355);
or U26 (N_26,In_864,In_402);
or U27 (N_27,In_405,In_952);
and U28 (N_28,In_1161,In_1384);
nor U29 (N_29,In_1352,In_1050);
or U30 (N_30,In_397,In_556);
nand U31 (N_31,In_843,In_69);
nor U32 (N_32,In_143,In_1285);
xor U33 (N_33,In_1014,In_1351);
and U34 (N_34,In_1030,In_185);
nor U35 (N_35,In_401,In_108);
nor U36 (N_36,In_384,In_1042);
and U37 (N_37,In_731,In_128);
or U38 (N_38,In_95,In_385);
nor U39 (N_39,In_500,In_539);
nor U40 (N_40,In_330,In_787);
nand U41 (N_41,In_1006,In_767);
nand U42 (N_42,In_635,In_795);
nor U43 (N_43,In_52,In_283);
or U44 (N_44,In_1099,In_532);
and U45 (N_45,In_1236,In_1058);
or U46 (N_46,In_518,In_407);
nand U47 (N_47,In_751,In_201);
or U48 (N_48,In_861,In_1107);
nor U49 (N_49,In_865,In_17);
or U50 (N_50,In_1339,In_866);
nand U51 (N_51,In_1012,In_756);
nand U52 (N_52,In_629,In_153);
nor U53 (N_53,In_618,In_1373);
nor U54 (N_54,In_770,In_361);
nor U55 (N_55,In_1466,In_683);
nor U56 (N_56,In_1139,In_416);
nor U57 (N_57,In_38,In_50);
and U58 (N_58,In_332,In_1381);
nand U59 (N_59,In_166,In_85);
nor U60 (N_60,In_1413,In_371);
nor U61 (N_61,In_1357,In_996);
nand U62 (N_62,In_1104,In_753);
nand U63 (N_63,In_1013,In_109);
or U64 (N_64,In_1377,In_1243);
or U65 (N_65,In_1002,In_901);
nor U66 (N_66,In_517,In_208);
and U67 (N_67,In_1437,In_316);
and U68 (N_68,In_451,In_575);
or U69 (N_69,In_192,In_605);
nand U70 (N_70,In_830,In_673);
and U71 (N_71,In_576,In_1036);
nor U72 (N_72,In_1237,In_839);
nor U73 (N_73,In_204,In_379);
or U74 (N_74,In_695,In_217);
or U75 (N_75,In_1231,In_463);
or U76 (N_76,In_394,In_1067);
and U77 (N_77,In_406,In_1476);
nand U78 (N_78,In_971,In_706);
or U79 (N_79,In_1094,In_720);
and U80 (N_80,In_317,In_596);
nand U81 (N_81,In_1296,In_587);
and U82 (N_82,In_363,In_1223);
xnor U83 (N_83,In_395,In_328);
nand U84 (N_84,In_988,In_804);
and U85 (N_85,In_376,In_722);
nand U86 (N_86,In_1475,In_24);
or U87 (N_87,In_216,In_1176);
and U88 (N_88,In_806,In_1166);
nand U89 (N_89,In_1305,In_476);
or U90 (N_90,In_1363,In_1368);
or U91 (N_91,In_1283,In_1290);
nand U92 (N_92,In_243,In_1164);
or U93 (N_93,In_917,In_1226);
or U94 (N_94,In_318,In_1263);
or U95 (N_95,In_1076,In_200);
nor U96 (N_96,In_598,In_885);
and U97 (N_97,In_1017,In_1273);
or U98 (N_98,In_297,In_1113);
nand U99 (N_99,In_1477,In_709);
or U100 (N_100,In_1111,In_287);
nor U101 (N_101,In_377,In_1252);
nand U102 (N_102,In_231,In_1383);
nand U103 (N_103,In_367,In_1314);
or U104 (N_104,In_1098,In_712);
xor U105 (N_105,In_1179,In_68);
and U106 (N_106,In_202,In_221);
xnor U107 (N_107,In_1335,In_951);
nand U108 (N_108,In_322,In_730);
nor U109 (N_109,In_1336,In_655);
nand U110 (N_110,In_595,In_940);
nor U111 (N_111,In_666,In_1136);
nor U112 (N_112,In_261,In_922);
or U113 (N_113,In_1287,In_87);
nor U114 (N_114,In_226,In_5);
and U115 (N_115,In_205,In_1016);
xor U116 (N_116,In_561,In_570);
or U117 (N_117,In_923,In_743);
or U118 (N_118,In_360,In_103);
nor U119 (N_119,In_638,In_579);
and U120 (N_120,In_636,In_1344);
nand U121 (N_121,In_1473,In_1400);
and U122 (N_122,In_926,In_617);
nand U123 (N_123,In_750,In_1007);
nor U124 (N_124,In_1376,In_121);
nand U125 (N_125,In_809,In_1434);
nor U126 (N_126,In_814,In_1337);
nor U127 (N_127,In_15,In_1169);
or U128 (N_128,In_776,In_620);
or U129 (N_129,In_664,In_1331);
nor U130 (N_130,In_1003,In_1464);
nor U131 (N_131,In_847,In_370);
nor U132 (N_132,In_490,In_560);
xor U133 (N_133,In_163,In_591);
nor U134 (N_134,In_534,In_1046);
nor U135 (N_135,In_1299,In_1061);
nor U136 (N_136,In_1436,In_6);
nand U137 (N_137,In_105,In_913);
nand U138 (N_138,In_883,In_1254);
nand U139 (N_139,In_232,In_67);
and U140 (N_140,In_1178,In_1279);
or U141 (N_141,In_1412,In_75);
and U142 (N_142,In_206,In_227);
xor U143 (N_143,In_1208,In_897);
or U144 (N_144,In_410,In_948);
nand U145 (N_145,In_29,In_1202);
and U146 (N_146,In_546,In_888);
or U147 (N_147,In_438,In_442);
nor U148 (N_148,In_822,In_25);
nor U149 (N_149,In_1211,In_149);
and U150 (N_150,In_969,In_1448);
and U151 (N_151,In_1418,In_626);
or U152 (N_152,In_1440,In_774);
and U153 (N_153,In_309,In_881);
nor U154 (N_154,In_1167,In_887);
or U155 (N_155,In_973,In_292);
nor U156 (N_156,In_1095,In_11);
or U157 (N_157,In_35,In_1186);
and U158 (N_158,In_439,In_1022);
nand U159 (N_159,In_977,In_443);
or U160 (N_160,In_1433,In_857);
nor U161 (N_161,In_53,In_909);
nor U162 (N_162,In_359,In_1115);
and U163 (N_163,In_207,In_979);
nor U164 (N_164,In_585,In_870);
and U165 (N_165,In_380,In_354);
nor U166 (N_166,In_78,In_190);
or U167 (N_167,In_412,In_1052);
and U168 (N_168,In_754,In_140);
and U169 (N_169,In_123,In_785);
nor U170 (N_170,In_22,In_1474);
or U171 (N_171,In_1389,In_1426);
xnor U172 (N_172,In_331,In_409);
and U173 (N_173,In_92,In_271);
nand U174 (N_174,In_241,In_1424);
or U175 (N_175,In_874,In_419);
and U176 (N_176,In_364,In_1453);
and U177 (N_177,In_1037,In_272);
nand U178 (N_178,In_1258,In_311);
or U179 (N_179,In_1342,In_1494);
or U180 (N_180,In_1492,In_39);
and U181 (N_181,In_1393,In_130);
and U182 (N_182,In_1347,In_939);
and U183 (N_183,In_122,In_389);
or U184 (N_184,In_295,In_1310);
nor U185 (N_185,In_900,In_193);
or U186 (N_186,In_1276,In_773);
nor U187 (N_187,In_453,In_552);
and U188 (N_188,In_1297,In_1268);
or U189 (N_189,In_448,In_1160);
and U190 (N_190,In_220,In_1271);
or U191 (N_191,In_251,In_928);
and U192 (N_192,In_538,In_877);
or U193 (N_193,In_1329,In_267);
nand U194 (N_194,In_1040,In_1218);
nand U195 (N_195,In_807,In_997);
nand U196 (N_196,In_1148,In_669);
nor U197 (N_197,In_194,In_1444);
nor U198 (N_198,In_593,In_171);
nor U199 (N_199,In_177,In_640);
and U200 (N_200,In_879,In_485);
or U201 (N_201,In_168,In_160);
or U202 (N_202,In_1253,In_1078);
or U203 (N_203,In_584,In_250);
nand U204 (N_204,In_280,In_404);
nor U205 (N_205,In_418,In_590);
nand U206 (N_206,In_119,In_215);
nand U207 (N_207,In_1032,In_600);
nor U208 (N_208,In_125,In_1275);
and U209 (N_209,In_902,In_1308);
nor U210 (N_210,In_599,In_508);
and U211 (N_211,In_1251,In_429);
nand U212 (N_212,In_930,In_1374);
nor U213 (N_213,In_447,In_621);
nand U214 (N_214,In_972,In_631);
or U215 (N_215,In_424,In_863);
or U216 (N_216,In_833,In_1499);
xor U217 (N_217,In_1490,In_308);
or U218 (N_218,In_657,In_355);
xnor U219 (N_219,In_1146,In_872);
nor U220 (N_220,In_796,In_566);
nor U221 (N_221,In_1239,In_728);
and U222 (N_222,In_643,In_1375);
nor U223 (N_223,In_1322,In_1072);
or U224 (N_224,In_1266,In_515);
nor U225 (N_225,In_837,In_851);
and U226 (N_226,In_942,In_772);
nor U227 (N_227,In_26,In_333);
nand U228 (N_228,In_727,In_746);
nand U229 (N_229,In_775,In_741);
and U230 (N_230,In_838,In_735);
or U231 (N_231,In_848,In_408);
or U232 (N_232,In_1068,In_90);
nand U233 (N_233,In_1485,In_1242);
or U234 (N_234,In_1292,In_1216);
or U235 (N_235,In_274,In_522);
or U236 (N_236,In_134,In_1079);
and U237 (N_237,In_1105,In_196);
xor U238 (N_238,In_219,In_466);
nand U239 (N_239,In_736,In_525);
nand U240 (N_240,In_588,In_689);
nand U241 (N_241,In_107,In_1484);
nor U242 (N_242,In_248,In_1153);
nand U243 (N_243,In_502,In_920);
and U244 (N_244,In_372,In_265);
nand U245 (N_245,In_541,In_257);
and U246 (N_246,In_1108,In_662);
nand U247 (N_247,In_478,In_914);
nor U248 (N_248,In_1289,In_1138);
and U249 (N_249,In_1177,In_65);
nand U250 (N_250,In_339,In_1222);
or U251 (N_251,In_393,In_732);
nor U252 (N_252,In_32,In_762);
and U253 (N_253,In_950,In_273);
and U254 (N_254,In_93,In_777);
nand U255 (N_255,In_904,In_924);
nand U256 (N_256,In_176,In_890);
and U257 (N_257,In_469,In_1119);
nor U258 (N_258,In_1348,In_889);
or U259 (N_259,In_540,In_812);
xor U260 (N_260,In_1451,In_66);
and U261 (N_261,In_158,In_1323);
nand U262 (N_262,In_400,In_711);
xor U263 (N_263,In_497,In_704);
nor U264 (N_264,In_1262,In_1152);
nand U265 (N_265,In_483,In_744);
and U266 (N_266,In_572,In_1399);
or U267 (N_267,In_133,In_677);
or U268 (N_268,In_894,In_1049);
nor U269 (N_269,In_188,In_535);
nand U270 (N_270,In_299,In_101);
nand U271 (N_271,In_1282,In_276);
xnor U272 (N_272,In_1356,In_473);
nand U273 (N_273,In_1286,In_288);
nand U274 (N_274,In_1074,In_262);
and U275 (N_275,In_1388,In_423);
or U276 (N_276,In_1315,In_1341);
nor U277 (N_277,In_195,In_504);
nor U278 (N_278,In_1359,In_1259);
nand U279 (N_279,In_1387,In_1124);
and U280 (N_280,In_49,In_936);
nor U281 (N_281,In_1333,In_827);
nor U282 (N_282,In_456,In_1225);
nor U283 (N_283,In_625,In_1361);
nor U284 (N_284,In_986,In_420);
and U285 (N_285,In_183,In_1238);
xor U286 (N_286,In_784,In_649);
or U287 (N_287,In_564,In_797);
or U288 (N_288,In_337,In_23);
nor U289 (N_289,In_582,In_647);
nand U290 (N_290,In_1441,In_810);
nor U291 (N_291,In_619,In_1461);
or U292 (N_292,In_912,In_642);
nand U293 (N_293,In_1257,In_567);
nand U294 (N_294,In_239,In_1171);
nand U295 (N_295,In_1154,In_59);
and U296 (N_296,In_161,In_375);
and U297 (N_297,In_966,In_382);
and U298 (N_298,In_724,In_148);
or U299 (N_299,In_1245,In_338);
and U300 (N_300,In_975,In_58);
and U301 (N_301,In_826,In_368);
nor U302 (N_302,In_173,In_30);
xnor U303 (N_303,In_1181,In_1396);
nor U304 (N_304,In_1151,In_999);
nor U305 (N_305,In_831,In_681);
or U306 (N_306,In_854,In_118);
or U307 (N_307,In_362,In_1364);
nor U308 (N_308,In_726,In_224);
nand U309 (N_309,In_790,In_1033);
and U310 (N_310,In_10,In_433);
nand U311 (N_311,In_277,In_738);
and U312 (N_312,In_1149,In_578);
or U313 (N_313,In_873,In_1390);
nor U314 (N_314,In_1338,In_356);
and U315 (N_315,In_1198,In_801);
nand U316 (N_316,In_1420,In_1004);
and U317 (N_317,In_1446,In_336);
or U318 (N_318,In_852,In_1325);
and U319 (N_319,In_868,In_841);
and U320 (N_320,In_747,In_1059);
or U321 (N_321,In_855,In_884);
or U322 (N_322,In_880,In_794);
and U323 (N_323,In_1093,In_813);
nand U324 (N_324,In_944,In_46);
and U325 (N_325,In_455,In_1156);
nand U326 (N_326,In_691,In_256);
nand U327 (N_327,In_113,In_832);
nor U328 (N_328,In_154,In_1077);
and U329 (N_329,In_1317,In_713);
and U330 (N_330,In_835,In_305);
and U331 (N_331,In_151,In_1199);
and U332 (N_332,In_1248,In_1439);
or U333 (N_333,In_54,In_218);
nor U334 (N_334,In_1109,In_1358);
nor U335 (N_335,In_388,In_120);
or U336 (N_336,In_399,In_1027);
and U337 (N_337,In_238,In_1397);
or U338 (N_338,In_602,In_306);
and U339 (N_339,In_302,In_446);
and U340 (N_340,In_223,In_1288);
or U341 (N_341,In_987,In_1019);
xor U342 (N_342,In_301,In_1103);
and U343 (N_343,In_342,In_100);
and U344 (N_344,In_703,In_1326);
nand U345 (N_345,In_124,In_1120);
nor U346 (N_346,In_1128,In_477);
and U347 (N_347,In_658,In_97);
or U348 (N_348,In_1442,In_77);
nor U349 (N_349,In_791,In_978);
nor U350 (N_350,In_348,In_934);
nand U351 (N_351,In_315,In_1057);
nor U352 (N_352,In_228,In_853);
nor U353 (N_353,In_1071,In_1121);
nand U354 (N_354,In_1015,In_651);
nand U355 (N_355,In_733,In_700);
and U356 (N_356,In_1213,In_1214);
nand U357 (N_357,In_671,In_1227);
or U358 (N_358,In_1470,In_960);
and U359 (N_359,In_1024,In_764);
or U360 (N_360,In_320,In_786);
nand U361 (N_361,In_1346,In_179);
nand U362 (N_362,In_805,In_1423);
and U363 (N_363,In_1415,In_705);
or U364 (N_364,In_717,In_266);
and U365 (N_365,In_454,In_96);
or U366 (N_366,In_182,In_862);
nor U367 (N_367,In_268,In_1137);
nand U368 (N_368,In_817,In_432);
nand U369 (N_369,In_789,In_1295);
nor U370 (N_370,In_435,In_14);
or U371 (N_371,In_214,In_656);
nor U372 (N_372,In_899,In_1233);
and U373 (N_373,In_396,In_1081);
and U374 (N_374,In_1117,In_373);
and U375 (N_375,In_70,In_110);
xor U376 (N_376,In_353,In_491);
or U377 (N_377,In_1190,In_1130);
nand U378 (N_378,In_178,In_1018);
nor U379 (N_379,In_1255,In_836);
nand U380 (N_380,In_645,In_1493);
or U381 (N_381,In_967,In_235);
nor U382 (N_382,In_734,In_1455);
and U383 (N_383,In_307,In_929);
and U384 (N_384,In_468,In_269);
and U385 (N_385,In_281,In_1391);
nand U386 (N_386,In_882,In_721);
nand U387 (N_387,In_1129,In_1054);
nand U388 (N_388,In_990,In_1334);
nand U389 (N_389,In_8,In_1053);
and U390 (N_390,In_898,In_678);
and U391 (N_391,In_347,In_1365);
nand U392 (N_392,In_1089,In_765);
nor U393 (N_393,In_1209,In_156);
nand U394 (N_394,In_1483,In_869);
or U395 (N_395,In_1215,In_480);
nor U396 (N_396,In_919,In_528);
nand U397 (N_397,In_729,In_1182);
or U398 (N_398,In_1496,In_537);
nand U399 (N_399,In_1407,In_165);
nand U400 (N_400,In_427,In_488);
nand U401 (N_401,In_1096,In_428);
nor U402 (N_402,In_104,In_83);
and U403 (N_403,In_1086,In_88);
or U404 (N_404,In_875,In_580);
or U405 (N_405,In_946,In_34);
or U406 (N_406,In_761,In_964);
or U407 (N_407,In_653,In_859);
and U408 (N_408,In_1159,In_1106);
or U409 (N_409,In_1431,In_63);
nor U410 (N_410,In_86,In_694);
nor U411 (N_411,In_1460,In_905);
or U412 (N_412,In_1409,In_1312);
nand U413 (N_413,In_1234,In_961);
nand U414 (N_414,In_630,In_1125);
nor U415 (N_415,In_296,In_953);
or U416 (N_416,In_976,In_684);
and U417 (N_417,In_1284,In_234);
and U418 (N_418,In_326,In_131);
nor U419 (N_419,In_1371,In_1065);
nand U420 (N_420,In_1345,In_1354);
nand U421 (N_421,In_1126,In_530);
or U422 (N_422,In_931,In_661);
nor U423 (N_423,In_551,In_693);
nor U424 (N_424,In_563,In_245);
or U425 (N_425,In_1192,In_632);
nand U426 (N_426,In_752,In_1435);
and U427 (N_427,In_670,In_1183);
and U428 (N_428,In_461,In_1165);
and U429 (N_429,In_956,In_474);
or U430 (N_430,In_559,In_1332);
or U431 (N_431,In_365,In_1321);
and U432 (N_432,In_222,In_1023);
and U433 (N_433,In_1478,In_698);
nand U434 (N_434,In_589,In_974);
or U435 (N_435,In_1230,In_440);
or U436 (N_436,In_278,In_335);
nand U437 (N_437,In_55,In_411);
xor U438 (N_438,In_514,In_247);
or U439 (N_439,In_203,In_545);
nand U440 (N_440,In_1403,In_680);
nand U441 (N_441,In_60,In_1467);
and U442 (N_442,In_321,In_1353);
nand U443 (N_443,In_1232,In_1265);
or U444 (N_444,In_1080,In_41);
nand U445 (N_445,In_676,In_768);
nand U446 (N_446,In_1487,In_1118);
and U447 (N_447,In_1280,In_513);
or U448 (N_448,In_28,In_1135);
or U449 (N_449,In_138,In_135);
nor U450 (N_450,In_300,In_189);
or U451 (N_451,In_291,In_933);
nor U452 (N_452,In_568,In_164);
or U453 (N_453,In_1449,In_725);
or U454 (N_454,In_1495,In_1454);
nor U455 (N_455,In_99,In_449);
or U456 (N_456,In_1244,In_1291);
or U457 (N_457,In_414,In_608);
or U458 (N_458,In_470,In_139);
nor U459 (N_459,In_1462,In_818);
nand U460 (N_460,In_187,In_484);
nand U461 (N_461,In_1249,In_48);
nand U462 (N_462,In_858,In_253);
and U463 (N_463,In_895,In_782);
nor U464 (N_464,In_1194,In_1185);
nor U465 (N_465,In_1457,In_679);
nor U466 (N_466,In_828,In_82);
nand U467 (N_467,In_13,In_652);
nor U468 (N_468,In_506,In_1378);
nand U469 (N_469,In_159,In_627);
nand U470 (N_470,In_1001,In_56);
nor U471 (N_471,In_209,In_341);
nand U472 (N_472,In_1468,In_637);
nor U473 (N_473,In_1264,In_460);
and U474 (N_474,In_1055,In_723);
and U475 (N_475,In_799,In_511);
nor U476 (N_476,In_503,In_398);
nor U477 (N_477,In_494,In_840);
and U478 (N_478,In_849,In_1173);
or U479 (N_479,In_829,In_697);
or U480 (N_480,In_57,In_941);
and U481 (N_481,In_748,In_1028);
and U482 (N_482,In_1256,In_1043);
and U483 (N_483,In_760,In_16);
and U484 (N_484,In_1340,In_554);
nor U485 (N_485,In_18,In_230);
or U486 (N_486,In_79,In_20);
or U487 (N_487,In_1367,In_43);
or U488 (N_488,In_597,In_240);
or U489 (N_489,In_938,In_1319);
and U490 (N_490,In_565,In_1343);
or U491 (N_491,In_1206,In_327);
or U492 (N_492,In_945,In_529);
or U493 (N_493,In_808,In_1294);
nor U494 (N_494,In_592,In_259);
nand U495 (N_495,In_1328,In_687);
and U496 (N_496,In_246,In_467);
nand U497 (N_497,In_1281,In_472);
nand U498 (N_498,In_667,In_27);
nor U499 (N_499,In_871,In_1205);
or U500 (N_500,In_1031,In_1459);
nand U501 (N_501,In_170,In_391);
xnor U502 (N_502,In_71,In_850);
nor U503 (N_503,In_282,In_1419);
and U504 (N_504,In_1082,In_1366);
nand U505 (N_505,In_1141,In_61);
nor U506 (N_506,In_672,In_1048);
nor U507 (N_507,In_1051,In_644);
and U508 (N_508,In_1417,In_1303);
and U509 (N_509,In_304,In_1116);
nor U510 (N_510,In_132,In_1122);
or U511 (N_511,In_358,In_778);
and U512 (N_512,In_1421,In_648);
nor U513 (N_513,In_574,In_334);
nand U514 (N_514,In_255,In_114);
nand U515 (N_515,In_37,In_550);
nand U516 (N_516,In_403,In_611);
nand U517 (N_517,In_769,In_1293);
and U518 (N_518,In_1497,In_954);
nor U519 (N_519,In_1008,In_682);
nand U520 (N_520,In_471,In_910);
or U521 (N_521,In_1144,In_1100);
nand U522 (N_522,In_1219,In_1372);
nand U523 (N_523,In_823,In_1471);
and U524 (N_524,In_1133,In_1157);
nand U525 (N_525,In_609,In_654);
or U526 (N_526,In_702,In_1021);
or U527 (N_527,In_815,In_586);
nand U528 (N_528,In_431,In_1085);
or U529 (N_529,In_270,In_533);
or U530 (N_530,In_1406,In_665);
and U531 (N_531,In_1392,In_1044);
nor U532 (N_532,In_229,In_980);
and U533 (N_533,In_1197,In_324);
or U534 (N_534,In_1414,In_12);
and U535 (N_535,In_686,In_76);
nand U536 (N_536,In_345,In_1330);
or U537 (N_537,In_581,In_1456);
nand U538 (N_538,In_505,In_615);
or U539 (N_539,In_36,In_145);
or U540 (N_540,In_719,In_1170);
or U541 (N_541,In_1306,In_425);
and U542 (N_542,In_1422,In_983);
nand U543 (N_543,In_1056,In_422);
nor U544 (N_544,In_1070,In_444);
nor U545 (N_545,In_963,In_526);
or U546 (N_546,In_162,In_421);
or U547 (N_547,In_1463,In_1489);
and U548 (N_548,In_915,In_357);
or U549 (N_549,In_352,In_1369);
and U550 (N_550,In_558,In_675);
or U551 (N_551,In_548,In_181);
nand U552 (N_552,In_519,In_745);
or U553 (N_553,In_907,In_1438);
nor U554 (N_554,In_1408,In_137);
nand U555 (N_555,In_199,In_1091);
nor U556 (N_556,In_779,In_1313);
and U557 (N_557,In_157,In_555);
or U558 (N_558,In_51,In_1270);
nor U559 (N_559,In_198,In_816);
nand U560 (N_560,In_498,In_1432);
nand U561 (N_561,In_1318,In_1009);
and U562 (N_562,In_457,In_387);
nand U563 (N_563,In_458,In_935);
nor U564 (N_564,In_1155,In_577);
or U565 (N_565,In_112,In_0);
nor U566 (N_566,In_213,In_1324);
and U567 (N_567,In_544,In_481);
and U568 (N_568,In_62,In_509);
and U569 (N_569,In_72,In_1212);
nor U570 (N_570,In_413,In_610);
nor U571 (N_571,In_1020,In_258);
nor U572 (N_572,In_641,In_527);
and U573 (N_573,In_739,In_1240);
nand U574 (N_574,In_465,In_995);
nor U575 (N_575,In_487,In_1479);
nor U576 (N_576,In_1026,In_1491);
and U577 (N_577,In_1427,In_542);
or U578 (N_578,In_908,In_493);
nand U579 (N_579,In_126,In_346);
and U580 (N_580,In_1395,In_152);
nand U581 (N_581,In_236,In_102);
nand U582 (N_582,In_1486,In_381);
or U583 (N_583,In_783,In_1370);
nor U584 (N_584,In_1380,In_668);
nor U585 (N_585,In_957,In_1220);
nor U586 (N_586,In_612,In_1410);
nand U587 (N_587,In_740,In_116);
nor U588 (N_588,In_937,In_146);
nor U589 (N_589,In_290,In_1430);
or U590 (N_590,In_507,In_553);
or U591 (N_591,In_1145,In_1304);
xnor U592 (N_592,In_233,In_127);
nand U593 (N_593,In_1073,In_1062);
nor U594 (N_594,In_495,In_970);
nand U595 (N_595,In_1401,In_825);
nor U596 (N_596,In_343,In_172);
nor U597 (N_597,In_998,In_1360);
or U598 (N_598,In_603,In_824);
or U599 (N_599,In_891,In_45);
nand U600 (N_600,In_374,In_279);
and U601 (N_601,In_1147,In_523);
and U602 (N_602,In_142,In_520);
or U603 (N_603,In_492,In_1045);
or U604 (N_604,In_918,In_4);
or U605 (N_605,In_147,In_982);
and U606 (N_606,In_84,In_1272);
nand U607 (N_607,In_659,In_984);
or U608 (N_608,In_284,In_366);
or U609 (N_609,In_1064,In_1134);
and U610 (N_610,In_710,In_521);
nand U611 (N_611,In_562,In_1088);
or U612 (N_612,In_415,In_604);
nor U613 (N_613,In_73,In_685);
xnor U614 (N_614,In_916,In_1241);
or U615 (N_615,In_921,In_47);
or U616 (N_616,In_482,In_800);
and U617 (N_617,In_3,In_759);
nor U618 (N_618,In_1224,In_21);
nand U619 (N_619,In_117,In_155);
nand U620 (N_620,In_571,In_74);
nand U621 (N_621,In_1385,In_834);
or U622 (N_622,In_690,In_594);
or U623 (N_623,In_688,In_237);
and U624 (N_624,In_351,In_1047);
nand U625 (N_625,In_80,In_293);
nor U626 (N_626,In_1316,In_1246);
nor U627 (N_627,In_1092,In_1452);
nor U628 (N_628,In_601,In_111);
nor U629 (N_629,In_383,In_294);
and U630 (N_630,In_628,In_252);
and U631 (N_631,In_89,In_144);
nand U632 (N_632,In_459,In_169);
nor U633 (N_633,In_1250,In_1267);
nand U634 (N_634,In_344,In_893);
nand U635 (N_635,In_1450,In_737);
nand U636 (N_636,In_141,In_180);
and U637 (N_637,In_1349,In_1207);
and U638 (N_638,In_819,In_1472);
or U639 (N_639,In_792,In_319);
and U640 (N_640,In_1307,In_1201);
nand U641 (N_641,In_210,In_106);
or U642 (N_642,In_1039,In_33);
and U643 (N_643,In_1298,In_329);
xor U644 (N_644,In_386,In_634);
nand U645 (N_645,In_646,In_696);
nor U646 (N_646,In_434,In_314);
nor U647 (N_647,In_1309,In_524);
nand U648 (N_648,In_1131,In_1458);
and U649 (N_649,In_1362,In_1035);
nand U650 (N_650,In_1302,In_660);
and U651 (N_651,In_1158,In_1038);
and U652 (N_652,In_573,In_842);
and U653 (N_653,In_40,In_516);
or U654 (N_654,In_959,In_1269);
nor U655 (N_655,In_1278,In_663);
nor U656 (N_656,In_496,In_1210);
nand U657 (N_657,In_1034,In_1247);
or U658 (N_658,In_633,In_994);
nand U659 (N_659,In_1320,In_1428);
or U660 (N_660,In_263,In_350);
nor U661 (N_661,In_1123,In_771);
or U662 (N_662,In_1481,In_303);
or U663 (N_663,In_878,In_1350);
or U664 (N_664,In_186,In_426);
or U665 (N_665,In_369,In_1404);
nand U666 (N_666,In_623,In_392);
nand U667 (N_667,In_699,In_1482);
nor U668 (N_668,In_325,In_780);
and U669 (N_669,In_1075,In_310);
nor U670 (N_670,In_1425,In_1229);
or U671 (N_671,In_692,In_191);
nand U672 (N_672,In_613,In_766);
and U673 (N_673,In_1469,In_44);
nand U674 (N_674,In_821,In_903);
and U675 (N_675,In_718,In_927);
or U676 (N_676,In_1102,In_64);
or U677 (N_677,In_462,In_1142);
and U678 (N_678,In_436,In_860);
nand U679 (N_679,In_1127,In_349);
nor U680 (N_680,In_569,In_378);
nand U681 (N_681,In_1150,In_1382);
nor U682 (N_682,In_225,In_1416);
or U683 (N_683,In_1090,In_1191);
nand U684 (N_684,In_115,In_501);
and U685 (N_685,In_955,In_289);
or U686 (N_686,In_312,In_1193);
and U687 (N_687,In_607,In_1235);
and U688 (N_688,In_1060,In_174);
and U689 (N_689,In_547,In_1163);
and U690 (N_690,In_925,In_313);
and U691 (N_691,In_1172,In_340);
nand U692 (N_692,In_1010,In_1063);
and U693 (N_693,In_244,In_249);
nor U694 (N_694,In_715,In_1386);
nor U695 (N_695,In_1498,In_211);
or U696 (N_696,In_820,In_531);
nor U697 (N_697,In_1069,In_42);
nand U698 (N_698,In_1175,In_1200);
and U699 (N_699,In_19,In_1301);
and U700 (N_700,In_1162,In_184);
or U701 (N_701,In_949,In_323);
or U702 (N_702,In_1445,In_129);
nand U703 (N_703,In_499,In_1217);
and U704 (N_704,In_1429,In_98);
and U705 (N_705,In_212,In_1174);
nand U706 (N_706,In_275,In_2);
nor U707 (N_707,In_1402,In_1114);
and U708 (N_708,In_430,In_650);
xnor U709 (N_709,In_911,In_958);
nand U710 (N_710,In_639,In_1261);
or U711 (N_711,In_1447,In_798);
nor U712 (N_712,In_707,In_624);
and U713 (N_713,In_175,In_1168);
and U714 (N_714,In_1379,In_549);
nor U715 (N_715,In_512,In_475);
and U716 (N_716,In_876,In_991);
or U717 (N_717,In_285,In_286);
and U718 (N_718,In_1180,In_1488);
nand U719 (N_719,In_1203,In_1327);
and U720 (N_720,In_91,In_614);
or U721 (N_721,In_962,In_742);
nand U722 (N_722,In_1411,In_1084);
nor U723 (N_723,In_1029,In_758);
nor U724 (N_724,In_242,In_1112);
nor U725 (N_725,In_150,In_856);
nand U726 (N_726,In_1101,In_763);
nor U727 (N_727,In_947,In_788);
nand U728 (N_728,In_1087,In_802);
nand U729 (N_729,In_1300,In_1000);
and U730 (N_730,In_1140,In_932);
nand U731 (N_731,In_536,In_486);
nor U732 (N_732,In_1041,In_1196);
nand U733 (N_733,In_1465,In_583);
nor U734 (N_734,In_993,In_437);
nor U735 (N_735,In_7,In_906);
or U736 (N_736,In_892,In_1277);
nor U737 (N_737,In_1005,In_755);
nand U738 (N_738,In_1097,In_489);
nand U739 (N_739,In_1394,In_264);
nand U740 (N_740,In_886,In_298);
nor U741 (N_741,In_510,In_846);
and U742 (N_742,In_1221,In_1260);
or U743 (N_743,In_1443,In_811);
or U744 (N_744,In_968,In_167);
or U745 (N_745,In_1189,In_749);
xnor U746 (N_746,In_81,In_1066);
and U747 (N_747,In_197,In_543);
nor U748 (N_748,In_943,In_1204);
or U749 (N_749,In_757,In_254);
nor U750 (N_750,In_83,In_932);
nand U751 (N_751,In_1413,In_182);
or U752 (N_752,In_636,In_65);
and U753 (N_753,In_1159,In_575);
and U754 (N_754,In_78,In_636);
or U755 (N_755,In_1149,In_521);
nand U756 (N_756,In_138,In_317);
nand U757 (N_757,In_1324,In_849);
nor U758 (N_758,In_1220,In_1209);
nand U759 (N_759,In_942,In_601);
or U760 (N_760,In_584,In_1426);
or U761 (N_761,In_781,In_979);
nor U762 (N_762,In_44,In_588);
nor U763 (N_763,In_1215,In_1008);
nor U764 (N_764,In_70,In_555);
nand U765 (N_765,In_1218,In_653);
and U766 (N_766,In_1338,In_887);
and U767 (N_767,In_190,In_922);
nand U768 (N_768,In_590,In_443);
nand U769 (N_769,In_350,In_792);
nand U770 (N_770,In_573,In_562);
nand U771 (N_771,In_44,In_469);
and U772 (N_772,In_319,In_544);
or U773 (N_773,In_1389,In_1206);
and U774 (N_774,In_643,In_539);
nor U775 (N_775,In_1314,In_835);
nor U776 (N_776,In_1166,In_1229);
nand U777 (N_777,In_258,In_1274);
and U778 (N_778,In_1038,In_817);
and U779 (N_779,In_30,In_723);
nor U780 (N_780,In_1247,In_267);
nand U781 (N_781,In_1005,In_1356);
xnor U782 (N_782,In_1013,In_417);
nor U783 (N_783,In_42,In_1064);
or U784 (N_784,In_1331,In_193);
nand U785 (N_785,In_977,In_1001);
nor U786 (N_786,In_355,In_617);
nor U787 (N_787,In_961,In_288);
nand U788 (N_788,In_777,In_54);
or U789 (N_789,In_941,In_1098);
nand U790 (N_790,In_1426,In_909);
and U791 (N_791,In_483,In_950);
nand U792 (N_792,In_508,In_1493);
nand U793 (N_793,In_1463,In_141);
and U794 (N_794,In_1414,In_444);
nand U795 (N_795,In_3,In_715);
nor U796 (N_796,In_167,In_1117);
nand U797 (N_797,In_751,In_86);
nor U798 (N_798,In_1077,In_356);
nor U799 (N_799,In_20,In_1197);
and U800 (N_800,In_1402,In_698);
xnor U801 (N_801,In_523,In_633);
nand U802 (N_802,In_801,In_25);
xor U803 (N_803,In_1297,In_944);
nand U804 (N_804,In_382,In_1290);
and U805 (N_805,In_993,In_173);
nor U806 (N_806,In_107,In_1039);
nand U807 (N_807,In_152,In_1361);
and U808 (N_808,In_414,In_1242);
and U809 (N_809,In_330,In_919);
nor U810 (N_810,In_161,In_754);
and U811 (N_811,In_1403,In_340);
nand U812 (N_812,In_1476,In_757);
nor U813 (N_813,In_1376,In_1002);
nand U814 (N_814,In_1186,In_1336);
and U815 (N_815,In_857,In_727);
nand U816 (N_816,In_817,In_462);
nand U817 (N_817,In_168,In_312);
or U818 (N_818,In_666,In_335);
or U819 (N_819,In_1279,In_1272);
and U820 (N_820,In_1068,In_610);
nand U821 (N_821,In_1029,In_724);
xnor U822 (N_822,In_1429,In_825);
nand U823 (N_823,In_231,In_57);
or U824 (N_824,In_849,In_1346);
and U825 (N_825,In_746,In_93);
or U826 (N_826,In_1232,In_945);
nand U827 (N_827,In_258,In_1355);
and U828 (N_828,In_1286,In_1463);
or U829 (N_829,In_272,In_485);
nor U830 (N_830,In_856,In_197);
nor U831 (N_831,In_611,In_165);
nor U832 (N_832,In_309,In_439);
and U833 (N_833,In_1025,In_1018);
or U834 (N_834,In_1114,In_679);
nand U835 (N_835,In_465,In_576);
and U836 (N_836,In_785,In_1360);
nand U837 (N_837,In_432,In_945);
nand U838 (N_838,In_1403,In_1226);
or U839 (N_839,In_654,In_1084);
and U840 (N_840,In_115,In_493);
and U841 (N_841,In_1125,In_178);
nand U842 (N_842,In_1334,In_646);
nor U843 (N_843,In_785,In_443);
nor U844 (N_844,In_860,In_1203);
nand U845 (N_845,In_405,In_967);
or U846 (N_846,In_223,In_1409);
or U847 (N_847,In_616,In_519);
nand U848 (N_848,In_35,In_394);
and U849 (N_849,In_236,In_1455);
nand U850 (N_850,In_299,In_1169);
and U851 (N_851,In_36,In_415);
or U852 (N_852,In_925,In_198);
and U853 (N_853,In_1039,In_779);
nand U854 (N_854,In_1071,In_634);
or U855 (N_855,In_514,In_488);
or U856 (N_856,In_153,In_753);
and U857 (N_857,In_1244,In_994);
and U858 (N_858,In_16,In_1173);
nand U859 (N_859,In_411,In_1112);
or U860 (N_860,In_154,In_714);
or U861 (N_861,In_1211,In_1247);
nor U862 (N_862,In_618,In_70);
nand U863 (N_863,In_1128,In_732);
xnor U864 (N_864,In_1316,In_831);
nand U865 (N_865,In_1481,In_1363);
or U866 (N_866,In_748,In_131);
nor U867 (N_867,In_1027,In_1291);
nand U868 (N_868,In_1311,In_1428);
xnor U869 (N_869,In_436,In_46);
nand U870 (N_870,In_485,In_948);
nor U871 (N_871,In_1294,In_1439);
nor U872 (N_872,In_720,In_1316);
nand U873 (N_873,In_269,In_453);
nor U874 (N_874,In_1310,In_890);
or U875 (N_875,In_1082,In_1069);
and U876 (N_876,In_96,In_1490);
and U877 (N_877,In_315,In_659);
nand U878 (N_878,In_1124,In_838);
nand U879 (N_879,In_36,In_579);
and U880 (N_880,In_113,In_657);
or U881 (N_881,In_587,In_38);
nand U882 (N_882,In_221,In_833);
nor U883 (N_883,In_1188,In_1019);
nand U884 (N_884,In_918,In_882);
and U885 (N_885,In_721,In_1332);
or U886 (N_886,In_878,In_1345);
nor U887 (N_887,In_734,In_1100);
and U888 (N_888,In_137,In_1168);
nor U889 (N_889,In_953,In_1459);
and U890 (N_890,In_1182,In_933);
nand U891 (N_891,In_1194,In_742);
and U892 (N_892,In_1490,In_120);
or U893 (N_893,In_1214,In_408);
and U894 (N_894,In_122,In_1227);
or U895 (N_895,In_87,In_265);
nor U896 (N_896,In_602,In_1090);
or U897 (N_897,In_597,In_865);
or U898 (N_898,In_811,In_1102);
nand U899 (N_899,In_115,In_213);
nand U900 (N_900,In_1092,In_904);
xnor U901 (N_901,In_489,In_1369);
nor U902 (N_902,In_122,In_8);
or U903 (N_903,In_1495,In_1216);
or U904 (N_904,In_1050,In_974);
xnor U905 (N_905,In_1034,In_1020);
and U906 (N_906,In_1477,In_1201);
or U907 (N_907,In_386,In_198);
xor U908 (N_908,In_1362,In_77);
xnor U909 (N_909,In_403,In_1440);
nor U910 (N_910,In_1186,In_772);
nor U911 (N_911,In_562,In_606);
and U912 (N_912,In_692,In_705);
nor U913 (N_913,In_1212,In_184);
nand U914 (N_914,In_1408,In_392);
and U915 (N_915,In_537,In_208);
and U916 (N_916,In_535,In_1231);
or U917 (N_917,In_1459,In_294);
or U918 (N_918,In_1256,In_1400);
and U919 (N_919,In_397,In_23);
nand U920 (N_920,In_1477,In_1070);
or U921 (N_921,In_537,In_575);
or U922 (N_922,In_41,In_128);
nand U923 (N_923,In_1426,In_1351);
nand U924 (N_924,In_149,In_1377);
nor U925 (N_925,In_236,In_265);
and U926 (N_926,In_1237,In_1160);
or U927 (N_927,In_72,In_1250);
nor U928 (N_928,In_1087,In_1107);
nand U929 (N_929,In_540,In_349);
or U930 (N_930,In_386,In_792);
or U931 (N_931,In_442,In_1182);
and U932 (N_932,In_947,In_488);
or U933 (N_933,In_980,In_567);
nand U934 (N_934,In_172,In_232);
xnor U935 (N_935,In_419,In_534);
nor U936 (N_936,In_32,In_800);
nand U937 (N_937,In_317,In_294);
and U938 (N_938,In_199,In_1493);
nand U939 (N_939,In_1000,In_660);
or U940 (N_940,In_227,In_417);
xor U941 (N_941,In_199,In_1030);
and U942 (N_942,In_1475,In_1403);
and U943 (N_943,In_277,In_430);
nand U944 (N_944,In_869,In_101);
nand U945 (N_945,In_838,In_94);
xnor U946 (N_946,In_376,In_1181);
and U947 (N_947,In_1338,In_470);
and U948 (N_948,In_774,In_739);
and U949 (N_949,In_1261,In_1071);
or U950 (N_950,In_435,In_395);
or U951 (N_951,In_824,In_1057);
and U952 (N_952,In_1183,In_1225);
and U953 (N_953,In_748,In_825);
nor U954 (N_954,In_1088,In_1107);
or U955 (N_955,In_434,In_1383);
nor U956 (N_956,In_900,In_1320);
and U957 (N_957,In_1189,In_732);
or U958 (N_958,In_81,In_1419);
and U959 (N_959,In_1207,In_415);
nand U960 (N_960,In_1414,In_461);
nand U961 (N_961,In_1387,In_528);
and U962 (N_962,In_666,In_480);
nor U963 (N_963,In_465,In_311);
nor U964 (N_964,In_1001,In_1162);
nand U965 (N_965,In_400,In_81);
nor U966 (N_966,In_896,In_289);
or U967 (N_967,In_1085,In_1076);
nor U968 (N_968,In_183,In_290);
nor U969 (N_969,In_424,In_703);
or U970 (N_970,In_491,In_754);
or U971 (N_971,In_160,In_347);
and U972 (N_972,In_1434,In_1229);
or U973 (N_973,In_779,In_982);
nor U974 (N_974,In_648,In_559);
nor U975 (N_975,In_712,In_846);
or U976 (N_976,In_88,In_767);
and U977 (N_977,In_338,In_853);
and U978 (N_978,In_157,In_254);
and U979 (N_979,In_53,In_1080);
or U980 (N_980,In_1442,In_1011);
or U981 (N_981,In_1204,In_1150);
and U982 (N_982,In_943,In_1090);
nor U983 (N_983,In_1106,In_1257);
or U984 (N_984,In_280,In_985);
or U985 (N_985,In_1326,In_944);
xnor U986 (N_986,In_1457,In_1292);
and U987 (N_987,In_159,In_307);
nor U988 (N_988,In_961,In_1232);
and U989 (N_989,In_1434,In_518);
nor U990 (N_990,In_556,In_634);
nand U991 (N_991,In_916,In_562);
and U992 (N_992,In_1303,In_1123);
nor U993 (N_993,In_507,In_1093);
and U994 (N_994,In_576,In_596);
nor U995 (N_995,In_1020,In_921);
and U996 (N_996,In_249,In_276);
and U997 (N_997,In_1424,In_1392);
nand U998 (N_998,In_971,In_1040);
nor U999 (N_999,In_940,In_1171);
nand U1000 (N_1000,In_892,In_1327);
nor U1001 (N_1001,In_302,In_828);
and U1002 (N_1002,In_1417,In_356);
nor U1003 (N_1003,In_1066,In_1148);
and U1004 (N_1004,In_507,In_945);
and U1005 (N_1005,In_847,In_1101);
or U1006 (N_1006,In_650,In_864);
and U1007 (N_1007,In_1131,In_406);
and U1008 (N_1008,In_372,In_433);
nand U1009 (N_1009,In_1102,In_1168);
or U1010 (N_1010,In_1280,In_755);
or U1011 (N_1011,In_1494,In_188);
and U1012 (N_1012,In_93,In_152);
and U1013 (N_1013,In_1330,In_1257);
nor U1014 (N_1014,In_951,In_1337);
xor U1015 (N_1015,In_1346,In_1252);
nor U1016 (N_1016,In_1210,In_471);
nand U1017 (N_1017,In_238,In_997);
or U1018 (N_1018,In_216,In_1351);
and U1019 (N_1019,In_1397,In_474);
nor U1020 (N_1020,In_1385,In_380);
nor U1021 (N_1021,In_192,In_1487);
nor U1022 (N_1022,In_501,In_874);
or U1023 (N_1023,In_1158,In_950);
nand U1024 (N_1024,In_788,In_551);
and U1025 (N_1025,In_1029,In_1255);
and U1026 (N_1026,In_410,In_364);
or U1027 (N_1027,In_377,In_252);
and U1028 (N_1028,In_992,In_311);
and U1029 (N_1029,In_470,In_1073);
and U1030 (N_1030,In_357,In_185);
or U1031 (N_1031,In_314,In_374);
nand U1032 (N_1032,In_872,In_1404);
nor U1033 (N_1033,In_183,In_644);
nor U1034 (N_1034,In_320,In_576);
and U1035 (N_1035,In_554,In_1297);
or U1036 (N_1036,In_1197,In_363);
nor U1037 (N_1037,In_1285,In_1174);
and U1038 (N_1038,In_396,In_1246);
and U1039 (N_1039,In_1261,In_257);
nor U1040 (N_1040,In_1365,In_512);
nand U1041 (N_1041,In_41,In_48);
xnor U1042 (N_1042,In_644,In_1134);
nor U1043 (N_1043,In_1250,In_809);
or U1044 (N_1044,In_65,In_1448);
and U1045 (N_1045,In_619,In_1168);
nand U1046 (N_1046,In_1304,In_1387);
or U1047 (N_1047,In_1374,In_7);
and U1048 (N_1048,In_743,In_843);
and U1049 (N_1049,In_674,In_633);
or U1050 (N_1050,In_1205,In_196);
nor U1051 (N_1051,In_1146,In_214);
and U1052 (N_1052,In_733,In_592);
nor U1053 (N_1053,In_721,In_1383);
or U1054 (N_1054,In_111,In_176);
nor U1055 (N_1055,In_1174,In_934);
nand U1056 (N_1056,In_590,In_1374);
nor U1057 (N_1057,In_718,In_596);
nor U1058 (N_1058,In_772,In_976);
nand U1059 (N_1059,In_1458,In_1438);
or U1060 (N_1060,In_859,In_598);
nand U1061 (N_1061,In_1147,In_234);
nor U1062 (N_1062,In_256,In_948);
nor U1063 (N_1063,In_1351,In_1319);
and U1064 (N_1064,In_308,In_693);
or U1065 (N_1065,In_441,In_1166);
and U1066 (N_1066,In_296,In_1029);
or U1067 (N_1067,In_729,In_923);
or U1068 (N_1068,In_145,In_712);
nor U1069 (N_1069,In_608,In_251);
nand U1070 (N_1070,In_827,In_738);
xnor U1071 (N_1071,In_1047,In_509);
or U1072 (N_1072,In_231,In_268);
and U1073 (N_1073,In_595,In_441);
nor U1074 (N_1074,In_1123,In_1063);
or U1075 (N_1075,In_1427,In_779);
or U1076 (N_1076,In_350,In_959);
nand U1077 (N_1077,In_1204,In_1318);
or U1078 (N_1078,In_1108,In_216);
nor U1079 (N_1079,In_419,In_1377);
nor U1080 (N_1080,In_1368,In_547);
nand U1081 (N_1081,In_1079,In_1245);
nor U1082 (N_1082,In_294,In_336);
nor U1083 (N_1083,In_1317,In_1055);
nand U1084 (N_1084,In_674,In_469);
and U1085 (N_1085,In_1166,In_55);
nand U1086 (N_1086,In_444,In_884);
nor U1087 (N_1087,In_212,In_1425);
nor U1088 (N_1088,In_1418,In_329);
nand U1089 (N_1089,In_1398,In_1358);
nand U1090 (N_1090,In_42,In_627);
nand U1091 (N_1091,In_910,In_65);
and U1092 (N_1092,In_1081,In_1080);
nor U1093 (N_1093,In_831,In_1269);
and U1094 (N_1094,In_995,In_872);
xor U1095 (N_1095,In_1496,In_768);
nor U1096 (N_1096,In_803,In_650);
or U1097 (N_1097,In_1063,In_504);
and U1098 (N_1098,In_1115,In_275);
nand U1099 (N_1099,In_855,In_1293);
nand U1100 (N_1100,In_996,In_378);
or U1101 (N_1101,In_309,In_1303);
nand U1102 (N_1102,In_627,In_318);
nand U1103 (N_1103,In_1353,In_535);
nor U1104 (N_1104,In_1287,In_148);
xnor U1105 (N_1105,In_87,In_1276);
and U1106 (N_1106,In_585,In_14);
and U1107 (N_1107,In_682,In_12);
and U1108 (N_1108,In_827,In_1006);
and U1109 (N_1109,In_59,In_533);
and U1110 (N_1110,In_709,In_233);
nand U1111 (N_1111,In_1221,In_560);
nor U1112 (N_1112,In_463,In_1109);
nor U1113 (N_1113,In_18,In_888);
or U1114 (N_1114,In_163,In_764);
or U1115 (N_1115,In_889,In_644);
or U1116 (N_1116,In_635,In_1258);
and U1117 (N_1117,In_730,In_820);
or U1118 (N_1118,In_1032,In_1490);
or U1119 (N_1119,In_555,In_521);
or U1120 (N_1120,In_1392,In_93);
nand U1121 (N_1121,In_1250,In_810);
and U1122 (N_1122,In_1081,In_423);
nand U1123 (N_1123,In_386,In_281);
nand U1124 (N_1124,In_784,In_1310);
nor U1125 (N_1125,In_1320,In_1365);
or U1126 (N_1126,In_1273,In_1351);
or U1127 (N_1127,In_675,In_228);
and U1128 (N_1128,In_198,In_1235);
or U1129 (N_1129,In_101,In_250);
nand U1130 (N_1130,In_627,In_918);
nor U1131 (N_1131,In_205,In_415);
and U1132 (N_1132,In_748,In_620);
nor U1133 (N_1133,In_50,In_514);
and U1134 (N_1134,In_321,In_1100);
nand U1135 (N_1135,In_787,In_142);
nand U1136 (N_1136,In_1147,In_1375);
nor U1137 (N_1137,In_716,In_1131);
nand U1138 (N_1138,In_1151,In_373);
and U1139 (N_1139,In_625,In_881);
and U1140 (N_1140,In_854,In_955);
nand U1141 (N_1141,In_702,In_493);
nor U1142 (N_1142,In_652,In_389);
nor U1143 (N_1143,In_192,In_306);
and U1144 (N_1144,In_738,In_945);
or U1145 (N_1145,In_1111,In_1272);
or U1146 (N_1146,In_1159,In_674);
nand U1147 (N_1147,In_1376,In_1305);
nor U1148 (N_1148,In_1361,In_1332);
and U1149 (N_1149,In_1009,In_143);
or U1150 (N_1150,In_1191,In_908);
or U1151 (N_1151,In_367,In_1039);
and U1152 (N_1152,In_84,In_64);
nor U1153 (N_1153,In_724,In_1126);
nand U1154 (N_1154,In_1256,In_1166);
and U1155 (N_1155,In_777,In_304);
nor U1156 (N_1156,In_748,In_784);
nand U1157 (N_1157,In_538,In_991);
and U1158 (N_1158,In_910,In_220);
nand U1159 (N_1159,In_25,In_24);
nor U1160 (N_1160,In_11,In_760);
and U1161 (N_1161,In_430,In_571);
nor U1162 (N_1162,In_954,In_926);
nand U1163 (N_1163,In_1054,In_96);
and U1164 (N_1164,In_1498,In_848);
and U1165 (N_1165,In_822,In_500);
nand U1166 (N_1166,In_1337,In_867);
or U1167 (N_1167,In_52,In_1069);
nor U1168 (N_1168,In_200,In_584);
nor U1169 (N_1169,In_866,In_1038);
nand U1170 (N_1170,In_528,In_847);
xor U1171 (N_1171,In_303,In_388);
and U1172 (N_1172,In_937,In_1383);
and U1173 (N_1173,In_549,In_632);
nand U1174 (N_1174,In_358,In_660);
or U1175 (N_1175,In_743,In_898);
or U1176 (N_1176,In_693,In_1479);
nand U1177 (N_1177,In_278,In_1292);
nor U1178 (N_1178,In_517,In_398);
nand U1179 (N_1179,In_423,In_191);
or U1180 (N_1180,In_384,In_147);
nand U1181 (N_1181,In_798,In_34);
or U1182 (N_1182,In_617,In_839);
nor U1183 (N_1183,In_1105,In_567);
nor U1184 (N_1184,In_1103,In_771);
nor U1185 (N_1185,In_1447,In_244);
or U1186 (N_1186,In_988,In_1180);
and U1187 (N_1187,In_839,In_1371);
nor U1188 (N_1188,In_1482,In_1417);
or U1189 (N_1189,In_874,In_336);
nor U1190 (N_1190,In_110,In_84);
xnor U1191 (N_1191,In_783,In_812);
nor U1192 (N_1192,In_917,In_429);
xnor U1193 (N_1193,In_946,In_726);
nor U1194 (N_1194,In_98,In_75);
or U1195 (N_1195,In_105,In_154);
nand U1196 (N_1196,In_919,In_1097);
or U1197 (N_1197,In_363,In_325);
nand U1198 (N_1198,In_1431,In_14);
and U1199 (N_1199,In_1331,In_728);
or U1200 (N_1200,In_1408,In_1118);
nor U1201 (N_1201,In_1374,In_132);
nand U1202 (N_1202,In_850,In_504);
or U1203 (N_1203,In_351,In_1201);
or U1204 (N_1204,In_54,In_56);
nor U1205 (N_1205,In_1165,In_353);
or U1206 (N_1206,In_270,In_360);
nor U1207 (N_1207,In_1310,In_1477);
nand U1208 (N_1208,In_330,In_1072);
nand U1209 (N_1209,In_1439,In_80);
or U1210 (N_1210,In_992,In_1271);
nand U1211 (N_1211,In_222,In_370);
nor U1212 (N_1212,In_477,In_172);
and U1213 (N_1213,In_162,In_429);
or U1214 (N_1214,In_557,In_468);
nor U1215 (N_1215,In_1292,In_1230);
and U1216 (N_1216,In_1001,In_1317);
and U1217 (N_1217,In_1088,In_1094);
and U1218 (N_1218,In_1381,In_164);
or U1219 (N_1219,In_137,In_802);
nand U1220 (N_1220,In_74,In_436);
nor U1221 (N_1221,In_950,In_1210);
or U1222 (N_1222,In_465,In_750);
and U1223 (N_1223,In_1243,In_134);
or U1224 (N_1224,In_902,In_903);
or U1225 (N_1225,In_1299,In_53);
and U1226 (N_1226,In_450,In_579);
or U1227 (N_1227,In_823,In_1126);
nor U1228 (N_1228,In_966,In_1168);
nand U1229 (N_1229,In_637,In_649);
nor U1230 (N_1230,In_263,In_1324);
nand U1231 (N_1231,In_1000,In_461);
nand U1232 (N_1232,In_443,In_769);
nand U1233 (N_1233,In_753,In_962);
nor U1234 (N_1234,In_509,In_1358);
nand U1235 (N_1235,In_283,In_890);
and U1236 (N_1236,In_1347,In_44);
and U1237 (N_1237,In_222,In_502);
nor U1238 (N_1238,In_1301,In_335);
and U1239 (N_1239,In_79,In_232);
and U1240 (N_1240,In_1116,In_180);
nor U1241 (N_1241,In_772,In_138);
nand U1242 (N_1242,In_948,In_460);
xnor U1243 (N_1243,In_158,In_1335);
or U1244 (N_1244,In_921,In_1379);
nand U1245 (N_1245,In_1155,In_54);
and U1246 (N_1246,In_1248,In_142);
nand U1247 (N_1247,In_1316,In_368);
nor U1248 (N_1248,In_474,In_504);
and U1249 (N_1249,In_884,In_396);
nand U1250 (N_1250,In_566,In_358);
nand U1251 (N_1251,In_409,In_184);
and U1252 (N_1252,In_130,In_118);
nor U1253 (N_1253,In_260,In_604);
nor U1254 (N_1254,In_954,In_107);
nor U1255 (N_1255,In_261,In_1363);
nor U1256 (N_1256,In_821,In_528);
nand U1257 (N_1257,In_1308,In_1042);
or U1258 (N_1258,In_1010,In_1300);
nor U1259 (N_1259,In_24,In_982);
nand U1260 (N_1260,In_229,In_1284);
nand U1261 (N_1261,In_1217,In_1158);
and U1262 (N_1262,In_988,In_143);
nand U1263 (N_1263,In_884,In_1235);
nor U1264 (N_1264,In_83,In_550);
xnor U1265 (N_1265,In_719,In_327);
and U1266 (N_1266,In_1271,In_51);
nand U1267 (N_1267,In_1404,In_1368);
nand U1268 (N_1268,In_571,In_460);
xor U1269 (N_1269,In_156,In_1013);
nor U1270 (N_1270,In_663,In_1364);
and U1271 (N_1271,In_1065,In_471);
nand U1272 (N_1272,In_461,In_514);
or U1273 (N_1273,In_209,In_490);
nand U1274 (N_1274,In_79,In_725);
nor U1275 (N_1275,In_1193,In_1440);
or U1276 (N_1276,In_547,In_1413);
or U1277 (N_1277,In_1055,In_621);
or U1278 (N_1278,In_1362,In_1259);
and U1279 (N_1279,In_2,In_334);
or U1280 (N_1280,In_280,In_781);
and U1281 (N_1281,In_1371,In_392);
nor U1282 (N_1282,In_47,In_923);
and U1283 (N_1283,In_1289,In_420);
nor U1284 (N_1284,In_971,In_118);
or U1285 (N_1285,In_1489,In_244);
or U1286 (N_1286,In_716,In_268);
nor U1287 (N_1287,In_1377,In_95);
nor U1288 (N_1288,In_1417,In_1387);
xnor U1289 (N_1289,In_91,In_628);
nand U1290 (N_1290,In_1358,In_349);
and U1291 (N_1291,In_897,In_1178);
nor U1292 (N_1292,In_642,In_221);
and U1293 (N_1293,In_988,In_734);
and U1294 (N_1294,In_809,In_1015);
nor U1295 (N_1295,In_781,In_562);
and U1296 (N_1296,In_413,In_622);
nand U1297 (N_1297,In_275,In_1228);
and U1298 (N_1298,In_19,In_652);
or U1299 (N_1299,In_951,In_787);
and U1300 (N_1300,In_1105,In_2);
nor U1301 (N_1301,In_1129,In_674);
and U1302 (N_1302,In_815,In_1);
nor U1303 (N_1303,In_818,In_1199);
nor U1304 (N_1304,In_708,In_962);
nand U1305 (N_1305,In_234,In_64);
nand U1306 (N_1306,In_369,In_96);
or U1307 (N_1307,In_484,In_864);
xor U1308 (N_1308,In_470,In_1314);
nand U1309 (N_1309,In_1204,In_70);
and U1310 (N_1310,In_170,In_164);
and U1311 (N_1311,In_1308,In_1481);
and U1312 (N_1312,In_666,In_1163);
nand U1313 (N_1313,In_847,In_716);
nor U1314 (N_1314,In_376,In_1017);
nor U1315 (N_1315,In_33,In_1499);
or U1316 (N_1316,In_1457,In_703);
nand U1317 (N_1317,In_272,In_946);
or U1318 (N_1318,In_852,In_1054);
nor U1319 (N_1319,In_591,In_1345);
and U1320 (N_1320,In_1238,In_1145);
nor U1321 (N_1321,In_937,In_1247);
and U1322 (N_1322,In_93,In_835);
xor U1323 (N_1323,In_640,In_970);
or U1324 (N_1324,In_897,In_689);
and U1325 (N_1325,In_777,In_318);
nor U1326 (N_1326,In_949,In_1235);
nand U1327 (N_1327,In_694,In_544);
nand U1328 (N_1328,In_250,In_1401);
and U1329 (N_1329,In_1386,In_493);
and U1330 (N_1330,In_1057,In_436);
and U1331 (N_1331,In_1212,In_1204);
and U1332 (N_1332,In_124,In_849);
or U1333 (N_1333,In_540,In_288);
nor U1334 (N_1334,In_276,In_1285);
nor U1335 (N_1335,In_507,In_229);
nand U1336 (N_1336,In_972,In_611);
and U1337 (N_1337,In_687,In_1289);
nor U1338 (N_1338,In_1001,In_267);
nand U1339 (N_1339,In_102,In_144);
and U1340 (N_1340,In_1436,In_126);
or U1341 (N_1341,In_1383,In_614);
or U1342 (N_1342,In_1404,In_256);
nor U1343 (N_1343,In_1349,In_1358);
or U1344 (N_1344,In_671,In_793);
and U1345 (N_1345,In_1420,In_336);
and U1346 (N_1346,In_1191,In_989);
and U1347 (N_1347,In_1448,In_1463);
and U1348 (N_1348,In_280,In_416);
or U1349 (N_1349,In_550,In_931);
and U1350 (N_1350,In_381,In_1420);
nand U1351 (N_1351,In_775,In_1343);
nor U1352 (N_1352,In_326,In_670);
xnor U1353 (N_1353,In_435,In_490);
nor U1354 (N_1354,In_544,In_1336);
or U1355 (N_1355,In_177,In_378);
nand U1356 (N_1356,In_238,In_484);
and U1357 (N_1357,In_389,In_128);
nor U1358 (N_1358,In_727,In_1161);
nor U1359 (N_1359,In_659,In_304);
or U1360 (N_1360,In_494,In_235);
and U1361 (N_1361,In_7,In_1459);
and U1362 (N_1362,In_854,In_626);
or U1363 (N_1363,In_1396,In_82);
nor U1364 (N_1364,In_696,In_283);
nand U1365 (N_1365,In_150,In_1471);
nor U1366 (N_1366,In_1048,In_1187);
nor U1367 (N_1367,In_835,In_969);
or U1368 (N_1368,In_1469,In_485);
or U1369 (N_1369,In_293,In_492);
nand U1370 (N_1370,In_1267,In_1455);
nand U1371 (N_1371,In_1228,In_793);
nor U1372 (N_1372,In_515,In_1195);
and U1373 (N_1373,In_1042,In_958);
nand U1374 (N_1374,In_573,In_519);
or U1375 (N_1375,In_66,In_1066);
nand U1376 (N_1376,In_103,In_347);
or U1377 (N_1377,In_127,In_317);
or U1378 (N_1378,In_768,In_1211);
nor U1379 (N_1379,In_255,In_1139);
or U1380 (N_1380,In_902,In_146);
nand U1381 (N_1381,In_110,In_960);
or U1382 (N_1382,In_1460,In_1313);
nand U1383 (N_1383,In_24,In_628);
nor U1384 (N_1384,In_1481,In_400);
and U1385 (N_1385,In_285,In_1184);
and U1386 (N_1386,In_377,In_69);
nand U1387 (N_1387,In_597,In_1460);
or U1388 (N_1388,In_484,In_347);
or U1389 (N_1389,In_779,In_211);
nand U1390 (N_1390,In_1132,In_78);
nand U1391 (N_1391,In_301,In_1228);
and U1392 (N_1392,In_727,In_1253);
and U1393 (N_1393,In_1307,In_395);
nor U1394 (N_1394,In_1220,In_106);
nand U1395 (N_1395,In_854,In_1136);
or U1396 (N_1396,In_1458,In_1066);
or U1397 (N_1397,In_1469,In_562);
and U1398 (N_1398,In_327,In_271);
nand U1399 (N_1399,In_575,In_705);
nand U1400 (N_1400,In_222,In_996);
nand U1401 (N_1401,In_1295,In_1464);
and U1402 (N_1402,In_669,In_1187);
nor U1403 (N_1403,In_538,In_563);
nor U1404 (N_1404,In_476,In_1365);
nor U1405 (N_1405,In_1299,In_975);
nand U1406 (N_1406,In_562,In_1249);
nor U1407 (N_1407,In_1058,In_1174);
and U1408 (N_1408,In_438,In_1332);
nand U1409 (N_1409,In_90,In_753);
and U1410 (N_1410,In_1307,In_384);
and U1411 (N_1411,In_246,In_38);
and U1412 (N_1412,In_952,In_99);
or U1413 (N_1413,In_225,In_904);
or U1414 (N_1414,In_1350,In_408);
nor U1415 (N_1415,In_38,In_784);
nor U1416 (N_1416,In_243,In_884);
nand U1417 (N_1417,In_1400,In_771);
nor U1418 (N_1418,In_621,In_566);
and U1419 (N_1419,In_1373,In_257);
or U1420 (N_1420,In_223,In_308);
and U1421 (N_1421,In_740,In_672);
nor U1422 (N_1422,In_113,In_1061);
xor U1423 (N_1423,In_1168,In_621);
nand U1424 (N_1424,In_75,In_1067);
nor U1425 (N_1425,In_225,In_1412);
and U1426 (N_1426,In_650,In_585);
nand U1427 (N_1427,In_1453,In_575);
or U1428 (N_1428,In_648,In_24);
nor U1429 (N_1429,In_932,In_851);
nor U1430 (N_1430,In_1470,In_800);
nor U1431 (N_1431,In_715,In_1189);
nand U1432 (N_1432,In_88,In_8);
or U1433 (N_1433,In_1053,In_1433);
or U1434 (N_1434,In_580,In_387);
and U1435 (N_1435,In_145,In_168);
nand U1436 (N_1436,In_1032,In_1383);
nand U1437 (N_1437,In_1215,In_596);
nand U1438 (N_1438,In_1213,In_1078);
nor U1439 (N_1439,In_382,In_378);
nand U1440 (N_1440,In_1355,In_1202);
nor U1441 (N_1441,In_841,In_1170);
nor U1442 (N_1442,In_589,In_553);
xnor U1443 (N_1443,In_1101,In_14);
or U1444 (N_1444,In_734,In_888);
nor U1445 (N_1445,In_879,In_1427);
or U1446 (N_1446,In_796,In_1102);
and U1447 (N_1447,In_928,In_1240);
nand U1448 (N_1448,In_196,In_1002);
and U1449 (N_1449,In_50,In_1402);
nor U1450 (N_1450,In_690,In_1358);
nor U1451 (N_1451,In_304,In_1089);
nand U1452 (N_1452,In_1281,In_496);
or U1453 (N_1453,In_882,In_3);
and U1454 (N_1454,In_183,In_946);
and U1455 (N_1455,In_1306,In_278);
nand U1456 (N_1456,In_408,In_880);
nor U1457 (N_1457,In_953,In_950);
nand U1458 (N_1458,In_759,In_1009);
and U1459 (N_1459,In_1025,In_230);
and U1460 (N_1460,In_311,In_251);
nor U1461 (N_1461,In_359,In_524);
nand U1462 (N_1462,In_782,In_1306);
nor U1463 (N_1463,In_778,In_772);
or U1464 (N_1464,In_459,In_442);
nand U1465 (N_1465,In_1254,In_356);
nor U1466 (N_1466,In_382,In_370);
xnor U1467 (N_1467,In_391,In_1063);
nand U1468 (N_1468,In_137,In_664);
nor U1469 (N_1469,In_688,In_207);
nand U1470 (N_1470,In_920,In_786);
nor U1471 (N_1471,In_1059,In_193);
nand U1472 (N_1472,In_780,In_458);
nor U1473 (N_1473,In_570,In_1328);
nand U1474 (N_1474,In_310,In_1027);
nor U1475 (N_1475,In_844,In_61);
or U1476 (N_1476,In_1210,In_1286);
nand U1477 (N_1477,In_1313,In_1222);
and U1478 (N_1478,In_378,In_433);
and U1479 (N_1479,In_1358,In_608);
and U1480 (N_1480,In_833,In_1086);
and U1481 (N_1481,In_721,In_1400);
and U1482 (N_1482,In_791,In_1311);
and U1483 (N_1483,In_1378,In_223);
and U1484 (N_1484,In_1393,In_137);
nand U1485 (N_1485,In_7,In_788);
or U1486 (N_1486,In_707,In_42);
nor U1487 (N_1487,In_901,In_476);
and U1488 (N_1488,In_1461,In_1057);
and U1489 (N_1489,In_1197,In_1403);
nand U1490 (N_1490,In_431,In_1322);
nand U1491 (N_1491,In_698,In_868);
and U1492 (N_1492,In_474,In_588);
nand U1493 (N_1493,In_397,In_339);
or U1494 (N_1494,In_902,In_413);
and U1495 (N_1495,In_450,In_466);
or U1496 (N_1496,In_24,In_10);
and U1497 (N_1497,In_420,In_329);
nor U1498 (N_1498,In_582,In_399);
nor U1499 (N_1499,In_346,In_181);
nor U1500 (N_1500,In_801,In_648);
and U1501 (N_1501,In_230,In_321);
nor U1502 (N_1502,In_661,In_1101);
or U1503 (N_1503,In_231,In_1368);
nand U1504 (N_1504,In_840,In_1427);
or U1505 (N_1505,In_1443,In_202);
or U1506 (N_1506,In_1393,In_281);
nand U1507 (N_1507,In_703,In_130);
or U1508 (N_1508,In_58,In_447);
or U1509 (N_1509,In_1028,In_428);
and U1510 (N_1510,In_1090,In_895);
nor U1511 (N_1511,In_1300,In_60);
nand U1512 (N_1512,In_1389,In_342);
or U1513 (N_1513,In_524,In_1271);
and U1514 (N_1514,In_763,In_263);
or U1515 (N_1515,In_974,In_611);
or U1516 (N_1516,In_1417,In_1167);
and U1517 (N_1517,In_545,In_1037);
nand U1518 (N_1518,In_824,In_601);
or U1519 (N_1519,In_1256,In_335);
nor U1520 (N_1520,In_211,In_1145);
nand U1521 (N_1521,In_461,In_715);
nor U1522 (N_1522,In_770,In_137);
or U1523 (N_1523,In_1306,In_1029);
nor U1524 (N_1524,In_534,In_528);
and U1525 (N_1525,In_405,In_923);
nand U1526 (N_1526,In_842,In_1435);
nor U1527 (N_1527,In_1325,In_164);
nor U1528 (N_1528,In_1293,In_300);
or U1529 (N_1529,In_586,In_444);
nand U1530 (N_1530,In_1144,In_259);
or U1531 (N_1531,In_0,In_1363);
nand U1532 (N_1532,In_1184,In_41);
or U1533 (N_1533,In_1125,In_1397);
and U1534 (N_1534,In_415,In_99);
or U1535 (N_1535,In_636,In_225);
nand U1536 (N_1536,In_1441,In_821);
nand U1537 (N_1537,In_659,In_1401);
and U1538 (N_1538,In_411,In_877);
or U1539 (N_1539,In_77,In_445);
nand U1540 (N_1540,In_1477,In_1249);
xor U1541 (N_1541,In_1358,In_1494);
nor U1542 (N_1542,In_1402,In_1042);
and U1543 (N_1543,In_1449,In_121);
or U1544 (N_1544,In_567,In_914);
or U1545 (N_1545,In_279,In_514);
nand U1546 (N_1546,In_540,In_1116);
nand U1547 (N_1547,In_271,In_808);
nand U1548 (N_1548,In_610,In_536);
and U1549 (N_1549,In_83,In_533);
xnor U1550 (N_1550,In_1487,In_1258);
or U1551 (N_1551,In_1488,In_1120);
nand U1552 (N_1552,In_17,In_1466);
nor U1553 (N_1553,In_576,In_703);
or U1554 (N_1554,In_614,In_1424);
nand U1555 (N_1555,In_925,In_219);
or U1556 (N_1556,In_585,In_1113);
and U1557 (N_1557,In_547,In_1247);
nand U1558 (N_1558,In_519,In_163);
or U1559 (N_1559,In_1262,In_565);
and U1560 (N_1560,In_729,In_444);
or U1561 (N_1561,In_370,In_1107);
and U1562 (N_1562,In_278,In_329);
and U1563 (N_1563,In_1144,In_1440);
or U1564 (N_1564,In_538,In_503);
and U1565 (N_1565,In_661,In_1494);
or U1566 (N_1566,In_1430,In_912);
nor U1567 (N_1567,In_60,In_1133);
nor U1568 (N_1568,In_1162,In_103);
nand U1569 (N_1569,In_1085,In_1440);
nor U1570 (N_1570,In_1283,In_64);
or U1571 (N_1571,In_964,In_452);
and U1572 (N_1572,In_1141,In_1025);
or U1573 (N_1573,In_1271,In_168);
and U1574 (N_1574,In_482,In_670);
nand U1575 (N_1575,In_548,In_763);
and U1576 (N_1576,In_385,In_221);
xnor U1577 (N_1577,In_940,In_957);
and U1578 (N_1578,In_944,In_889);
and U1579 (N_1579,In_586,In_353);
xnor U1580 (N_1580,In_847,In_871);
and U1581 (N_1581,In_41,In_920);
or U1582 (N_1582,In_1114,In_38);
nand U1583 (N_1583,In_408,In_102);
or U1584 (N_1584,In_490,In_579);
nand U1585 (N_1585,In_1160,In_850);
or U1586 (N_1586,In_1182,In_730);
nor U1587 (N_1587,In_1042,In_755);
and U1588 (N_1588,In_250,In_1210);
and U1589 (N_1589,In_365,In_209);
nor U1590 (N_1590,In_1474,In_923);
or U1591 (N_1591,In_1128,In_30);
nor U1592 (N_1592,In_381,In_353);
or U1593 (N_1593,In_579,In_665);
nand U1594 (N_1594,In_747,In_1340);
or U1595 (N_1595,In_1328,In_675);
nor U1596 (N_1596,In_482,In_424);
nor U1597 (N_1597,In_798,In_911);
and U1598 (N_1598,In_359,In_283);
nor U1599 (N_1599,In_855,In_1403);
or U1600 (N_1600,In_155,In_1361);
or U1601 (N_1601,In_860,In_525);
or U1602 (N_1602,In_1121,In_663);
nand U1603 (N_1603,In_341,In_775);
or U1604 (N_1604,In_462,In_102);
and U1605 (N_1605,In_203,In_138);
or U1606 (N_1606,In_460,In_1112);
or U1607 (N_1607,In_1246,In_30);
and U1608 (N_1608,In_709,In_628);
or U1609 (N_1609,In_1380,In_862);
nor U1610 (N_1610,In_161,In_872);
or U1611 (N_1611,In_1237,In_408);
or U1612 (N_1612,In_62,In_1205);
or U1613 (N_1613,In_1136,In_690);
and U1614 (N_1614,In_768,In_582);
nor U1615 (N_1615,In_1307,In_901);
nand U1616 (N_1616,In_666,In_43);
or U1617 (N_1617,In_561,In_962);
nor U1618 (N_1618,In_410,In_1418);
and U1619 (N_1619,In_28,In_1441);
nor U1620 (N_1620,In_1296,In_475);
nor U1621 (N_1621,In_629,In_1364);
or U1622 (N_1622,In_697,In_263);
and U1623 (N_1623,In_525,In_267);
or U1624 (N_1624,In_1462,In_725);
nand U1625 (N_1625,In_840,In_0);
and U1626 (N_1626,In_637,In_290);
nand U1627 (N_1627,In_1201,In_85);
nor U1628 (N_1628,In_1043,In_367);
nand U1629 (N_1629,In_756,In_493);
nand U1630 (N_1630,In_272,In_172);
nand U1631 (N_1631,In_667,In_688);
nor U1632 (N_1632,In_843,In_63);
or U1633 (N_1633,In_807,In_69);
nand U1634 (N_1634,In_983,In_1348);
and U1635 (N_1635,In_1093,In_119);
or U1636 (N_1636,In_1070,In_889);
xor U1637 (N_1637,In_44,In_888);
or U1638 (N_1638,In_6,In_55);
nand U1639 (N_1639,In_164,In_256);
and U1640 (N_1640,In_558,In_1084);
nand U1641 (N_1641,In_1033,In_981);
xnor U1642 (N_1642,In_163,In_521);
and U1643 (N_1643,In_10,In_119);
nand U1644 (N_1644,In_498,In_841);
and U1645 (N_1645,In_494,In_176);
nand U1646 (N_1646,In_648,In_500);
nor U1647 (N_1647,In_748,In_533);
nor U1648 (N_1648,In_200,In_156);
or U1649 (N_1649,In_383,In_477);
and U1650 (N_1650,In_1492,In_630);
and U1651 (N_1651,In_33,In_599);
and U1652 (N_1652,In_176,In_1141);
nand U1653 (N_1653,In_134,In_684);
and U1654 (N_1654,In_899,In_210);
and U1655 (N_1655,In_438,In_1053);
and U1656 (N_1656,In_1277,In_1471);
xnor U1657 (N_1657,In_1111,In_1458);
nor U1658 (N_1658,In_1324,In_891);
nand U1659 (N_1659,In_1090,In_817);
nand U1660 (N_1660,In_711,In_456);
and U1661 (N_1661,In_802,In_470);
nor U1662 (N_1662,In_1113,In_708);
nor U1663 (N_1663,In_173,In_250);
nand U1664 (N_1664,In_1457,In_132);
or U1665 (N_1665,In_256,In_674);
nor U1666 (N_1666,In_50,In_501);
nand U1667 (N_1667,In_1095,In_486);
nor U1668 (N_1668,In_894,In_842);
and U1669 (N_1669,In_968,In_173);
nor U1670 (N_1670,In_110,In_733);
nand U1671 (N_1671,In_384,In_772);
xnor U1672 (N_1672,In_325,In_345);
nand U1673 (N_1673,In_878,In_1176);
nand U1674 (N_1674,In_871,In_631);
nor U1675 (N_1675,In_176,In_1095);
nor U1676 (N_1676,In_6,In_127);
nand U1677 (N_1677,In_136,In_811);
xor U1678 (N_1678,In_1236,In_1192);
or U1679 (N_1679,In_646,In_1036);
xor U1680 (N_1680,In_738,In_626);
nand U1681 (N_1681,In_0,In_1452);
nor U1682 (N_1682,In_1044,In_906);
xnor U1683 (N_1683,In_1101,In_1111);
nand U1684 (N_1684,In_740,In_660);
nand U1685 (N_1685,In_739,In_533);
nand U1686 (N_1686,In_1,In_401);
nand U1687 (N_1687,In_217,In_10);
nor U1688 (N_1688,In_554,In_994);
nor U1689 (N_1689,In_1134,In_39);
or U1690 (N_1690,In_1019,In_477);
and U1691 (N_1691,In_194,In_1407);
and U1692 (N_1692,In_1432,In_1433);
nand U1693 (N_1693,In_256,In_229);
nand U1694 (N_1694,In_484,In_169);
nor U1695 (N_1695,In_1086,In_54);
or U1696 (N_1696,In_1468,In_1434);
nand U1697 (N_1697,In_573,In_939);
nor U1698 (N_1698,In_1260,In_1381);
nor U1699 (N_1699,In_845,In_51);
nand U1700 (N_1700,In_629,In_1418);
or U1701 (N_1701,In_1412,In_736);
and U1702 (N_1702,In_634,In_908);
and U1703 (N_1703,In_578,In_891);
nand U1704 (N_1704,In_29,In_516);
and U1705 (N_1705,In_1379,In_42);
and U1706 (N_1706,In_949,In_1216);
or U1707 (N_1707,In_513,In_1088);
or U1708 (N_1708,In_1471,In_796);
or U1709 (N_1709,In_1198,In_754);
nor U1710 (N_1710,In_269,In_580);
nand U1711 (N_1711,In_1087,In_1049);
nor U1712 (N_1712,In_430,In_878);
or U1713 (N_1713,In_715,In_891);
or U1714 (N_1714,In_1235,In_688);
nand U1715 (N_1715,In_473,In_204);
nor U1716 (N_1716,In_1243,In_1135);
and U1717 (N_1717,In_635,In_516);
nand U1718 (N_1718,In_864,In_345);
or U1719 (N_1719,In_1341,In_825);
nand U1720 (N_1720,In_783,In_1059);
nor U1721 (N_1721,In_126,In_1075);
nand U1722 (N_1722,In_858,In_842);
nand U1723 (N_1723,In_447,In_1191);
and U1724 (N_1724,In_244,In_896);
xor U1725 (N_1725,In_720,In_808);
or U1726 (N_1726,In_94,In_476);
nand U1727 (N_1727,In_989,In_413);
nand U1728 (N_1728,In_1095,In_598);
nand U1729 (N_1729,In_1353,In_1151);
or U1730 (N_1730,In_99,In_1365);
nand U1731 (N_1731,In_26,In_461);
nand U1732 (N_1732,In_826,In_146);
and U1733 (N_1733,In_496,In_106);
nor U1734 (N_1734,In_1246,In_1209);
nand U1735 (N_1735,In_1099,In_38);
and U1736 (N_1736,In_1307,In_1136);
or U1737 (N_1737,In_469,In_924);
xnor U1738 (N_1738,In_1377,In_1417);
or U1739 (N_1739,In_1444,In_413);
nand U1740 (N_1740,In_357,In_423);
and U1741 (N_1741,In_1297,In_1217);
nand U1742 (N_1742,In_1024,In_218);
or U1743 (N_1743,In_783,In_271);
nand U1744 (N_1744,In_588,In_7);
or U1745 (N_1745,In_1053,In_120);
or U1746 (N_1746,In_97,In_863);
and U1747 (N_1747,In_259,In_330);
or U1748 (N_1748,In_1085,In_527);
nor U1749 (N_1749,In_496,In_1052);
nor U1750 (N_1750,In_637,In_377);
nand U1751 (N_1751,In_1061,In_1322);
or U1752 (N_1752,In_61,In_1053);
nor U1753 (N_1753,In_448,In_412);
or U1754 (N_1754,In_1055,In_382);
nand U1755 (N_1755,In_851,In_283);
and U1756 (N_1756,In_958,In_1404);
and U1757 (N_1757,In_1016,In_329);
nor U1758 (N_1758,In_409,In_1244);
and U1759 (N_1759,In_197,In_592);
nand U1760 (N_1760,In_369,In_1095);
nor U1761 (N_1761,In_177,In_1159);
and U1762 (N_1762,In_1280,In_384);
nor U1763 (N_1763,In_822,In_705);
nor U1764 (N_1764,In_193,In_145);
and U1765 (N_1765,In_1470,In_1331);
nor U1766 (N_1766,In_1182,In_1099);
or U1767 (N_1767,In_1423,In_698);
nor U1768 (N_1768,In_676,In_785);
nand U1769 (N_1769,In_1094,In_742);
nand U1770 (N_1770,In_1140,In_497);
and U1771 (N_1771,In_1445,In_659);
nor U1772 (N_1772,In_377,In_842);
or U1773 (N_1773,In_11,In_1338);
nand U1774 (N_1774,In_1424,In_487);
nor U1775 (N_1775,In_1420,In_1157);
and U1776 (N_1776,In_1325,In_686);
nand U1777 (N_1777,In_791,In_1217);
and U1778 (N_1778,In_6,In_374);
and U1779 (N_1779,In_1198,In_875);
and U1780 (N_1780,In_640,In_1320);
nand U1781 (N_1781,In_1006,In_1258);
nor U1782 (N_1782,In_453,In_197);
nand U1783 (N_1783,In_1235,In_727);
nor U1784 (N_1784,In_169,In_428);
and U1785 (N_1785,In_1076,In_819);
and U1786 (N_1786,In_434,In_381);
or U1787 (N_1787,In_1220,In_348);
or U1788 (N_1788,In_357,In_1206);
xor U1789 (N_1789,In_45,In_443);
or U1790 (N_1790,In_277,In_655);
nor U1791 (N_1791,In_687,In_995);
nand U1792 (N_1792,In_478,In_489);
nand U1793 (N_1793,In_293,In_245);
nand U1794 (N_1794,In_157,In_1360);
and U1795 (N_1795,In_1473,In_146);
nor U1796 (N_1796,In_19,In_317);
and U1797 (N_1797,In_1264,In_501);
nor U1798 (N_1798,In_1292,In_511);
and U1799 (N_1799,In_310,In_807);
nand U1800 (N_1800,In_418,In_754);
xor U1801 (N_1801,In_146,In_1056);
nor U1802 (N_1802,In_534,In_661);
nor U1803 (N_1803,In_1162,In_952);
or U1804 (N_1804,In_747,In_0);
or U1805 (N_1805,In_561,In_392);
nor U1806 (N_1806,In_233,In_527);
nor U1807 (N_1807,In_138,In_1220);
and U1808 (N_1808,In_354,In_454);
or U1809 (N_1809,In_147,In_1241);
nand U1810 (N_1810,In_99,In_1147);
nand U1811 (N_1811,In_1266,In_87);
nand U1812 (N_1812,In_598,In_177);
and U1813 (N_1813,In_151,In_557);
and U1814 (N_1814,In_1262,In_206);
and U1815 (N_1815,In_1276,In_789);
nand U1816 (N_1816,In_1391,In_198);
and U1817 (N_1817,In_63,In_468);
nor U1818 (N_1818,In_245,In_883);
and U1819 (N_1819,In_1481,In_735);
and U1820 (N_1820,In_729,In_377);
or U1821 (N_1821,In_397,In_1354);
and U1822 (N_1822,In_384,In_1284);
and U1823 (N_1823,In_689,In_818);
and U1824 (N_1824,In_67,In_1235);
and U1825 (N_1825,In_188,In_671);
or U1826 (N_1826,In_1484,In_212);
nor U1827 (N_1827,In_930,In_1455);
or U1828 (N_1828,In_296,In_1456);
and U1829 (N_1829,In_449,In_367);
or U1830 (N_1830,In_1156,In_110);
nor U1831 (N_1831,In_1456,In_1294);
nor U1832 (N_1832,In_532,In_547);
nand U1833 (N_1833,In_392,In_17);
nor U1834 (N_1834,In_560,In_816);
nand U1835 (N_1835,In_112,In_92);
and U1836 (N_1836,In_97,In_1413);
nand U1837 (N_1837,In_204,In_96);
and U1838 (N_1838,In_196,In_629);
and U1839 (N_1839,In_1398,In_760);
nor U1840 (N_1840,In_962,In_681);
and U1841 (N_1841,In_554,In_868);
or U1842 (N_1842,In_525,In_1042);
or U1843 (N_1843,In_79,In_651);
nor U1844 (N_1844,In_472,In_775);
and U1845 (N_1845,In_157,In_357);
nor U1846 (N_1846,In_904,In_1380);
and U1847 (N_1847,In_1392,In_1105);
or U1848 (N_1848,In_1012,In_214);
nor U1849 (N_1849,In_1401,In_191);
nor U1850 (N_1850,In_1324,In_490);
nor U1851 (N_1851,In_1191,In_815);
nor U1852 (N_1852,In_103,In_614);
nand U1853 (N_1853,In_459,In_1332);
nor U1854 (N_1854,In_593,In_843);
and U1855 (N_1855,In_1166,In_412);
nand U1856 (N_1856,In_523,In_1103);
nor U1857 (N_1857,In_11,In_1151);
nor U1858 (N_1858,In_1059,In_465);
or U1859 (N_1859,In_977,In_1230);
and U1860 (N_1860,In_1055,In_342);
and U1861 (N_1861,In_1187,In_263);
or U1862 (N_1862,In_900,In_643);
or U1863 (N_1863,In_380,In_697);
nor U1864 (N_1864,In_858,In_1428);
or U1865 (N_1865,In_835,In_418);
and U1866 (N_1866,In_424,In_1124);
nand U1867 (N_1867,In_843,In_1456);
or U1868 (N_1868,In_776,In_231);
and U1869 (N_1869,In_451,In_20);
nand U1870 (N_1870,In_347,In_546);
and U1871 (N_1871,In_274,In_519);
nand U1872 (N_1872,In_895,In_833);
xnor U1873 (N_1873,In_581,In_1404);
nand U1874 (N_1874,In_33,In_439);
and U1875 (N_1875,In_1329,In_775);
nand U1876 (N_1876,In_1293,In_536);
nor U1877 (N_1877,In_783,In_709);
and U1878 (N_1878,In_1108,In_601);
or U1879 (N_1879,In_1401,In_41);
or U1880 (N_1880,In_223,In_466);
nor U1881 (N_1881,In_715,In_1346);
nor U1882 (N_1882,In_1063,In_513);
and U1883 (N_1883,In_215,In_719);
or U1884 (N_1884,In_853,In_565);
xor U1885 (N_1885,In_649,In_1189);
nor U1886 (N_1886,In_517,In_1449);
and U1887 (N_1887,In_910,In_849);
or U1888 (N_1888,In_862,In_409);
or U1889 (N_1889,In_803,In_1167);
nand U1890 (N_1890,In_1499,In_1485);
xor U1891 (N_1891,In_357,In_414);
or U1892 (N_1892,In_97,In_1257);
nand U1893 (N_1893,In_419,In_158);
nand U1894 (N_1894,In_1378,In_466);
and U1895 (N_1895,In_1203,In_1422);
or U1896 (N_1896,In_179,In_941);
and U1897 (N_1897,In_795,In_292);
nor U1898 (N_1898,In_908,In_1189);
nor U1899 (N_1899,In_1404,In_680);
or U1900 (N_1900,In_879,In_520);
nor U1901 (N_1901,In_427,In_351);
nand U1902 (N_1902,In_1120,In_1345);
and U1903 (N_1903,In_986,In_1118);
nor U1904 (N_1904,In_1382,In_1200);
or U1905 (N_1905,In_1437,In_1471);
nor U1906 (N_1906,In_1125,In_216);
nand U1907 (N_1907,In_1250,In_884);
nand U1908 (N_1908,In_336,In_321);
nor U1909 (N_1909,In_833,In_993);
nand U1910 (N_1910,In_649,In_691);
nand U1911 (N_1911,In_1396,In_901);
nand U1912 (N_1912,In_779,In_637);
nor U1913 (N_1913,In_320,In_266);
nor U1914 (N_1914,In_1433,In_1350);
nand U1915 (N_1915,In_571,In_438);
and U1916 (N_1916,In_892,In_1332);
and U1917 (N_1917,In_297,In_509);
or U1918 (N_1918,In_242,In_1472);
or U1919 (N_1919,In_576,In_387);
and U1920 (N_1920,In_313,In_967);
or U1921 (N_1921,In_75,In_1003);
and U1922 (N_1922,In_1092,In_402);
nand U1923 (N_1923,In_535,In_724);
and U1924 (N_1924,In_480,In_299);
or U1925 (N_1925,In_439,In_1172);
nand U1926 (N_1926,In_1156,In_201);
nand U1927 (N_1927,In_904,In_1144);
or U1928 (N_1928,In_68,In_114);
and U1929 (N_1929,In_989,In_515);
and U1930 (N_1930,In_686,In_327);
or U1931 (N_1931,In_957,In_199);
nor U1932 (N_1932,In_531,In_981);
nor U1933 (N_1933,In_685,In_1310);
and U1934 (N_1934,In_546,In_128);
nand U1935 (N_1935,In_141,In_344);
or U1936 (N_1936,In_618,In_858);
nand U1937 (N_1937,In_1130,In_1105);
or U1938 (N_1938,In_1021,In_30);
or U1939 (N_1939,In_1009,In_200);
nand U1940 (N_1940,In_1269,In_1051);
or U1941 (N_1941,In_397,In_514);
nor U1942 (N_1942,In_1143,In_1100);
nor U1943 (N_1943,In_97,In_487);
nor U1944 (N_1944,In_746,In_683);
and U1945 (N_1945,In_319,In_307);
nor U1946 (N_1946,In_293,In_447);
nand U1947 (N_1947,In_325,In_522);
and U1948 (N_1948,In_309,In_661);
or U1949 (N_1949,In_1406,In_1453);
nand U1950 (N_1950,In_109,In_1203);
and U1951 (N_1951,In_829,In_1274);
or U1952 (N_1952,In_527,In_526);
nand U1953 (N_1953,In_924,In_1101);
and U1954 (N_1954,In_404,In_1379);
and U1955 (N_1955,In_1158,In_801);
or U1956 (N_1956,In_414,In_421);
nor U1957 (N_1957,In_274,In_346);
nand U1958 (N_1958,In_1359,In_769);
and U1959 (N_1959,In_515,In_398);
and U1960 (N_1960,In_173,In_1287);
nand U1961 (N_1961,In_713,In_1345);
nand U1962 (N_1962,In_965,In_274);
nand U1963 (N_1963,In_400,In_407);
nor U1964 (N_1964,In_302,In_606);
nor U1965 (N_1965,In_204,In_182);
nor U1966 (N_1966,In_1105,In_769);
nand U1967 (N_1967,In_864,In_1309);
nor U1968 (N_1968,In_1484,In_305);
or U1969 (N_1969,In_1143,In_1121);
and U1970 (N_1970,In_493,In_404);
or U1971 (N_1971,In_1313,In_804);
xnor U1972 (N_1972,In_1220,In_951);
nor U1973 (N_1973,In_844,In_396);
nor U1974 (N_1974,In_768,In_218);
nor U1975 (N_1975,In_590,In_318);
and U1976 (N_1976,In_810,In_838);
and U1977 (N_1977,In_462,In_1069);
or U1978 (N_1978,In_567,In_802);
or U1979 (N_1979,In_998,In_986);
or U1980 (N_1980,In_782,In_257);
and U1981 (N_1981,In_1326,In_1201);
and U1982 (N_1982,In_715,In_1208);
nand U1983 (N_1983,In_184,In_1447);
and U1984 (N_1984,In_569,In_1426);
nand U1985 (N_1985,In_529,In_1367);
nor U1986 (N_1986,In_1198,In_991);
and U1987 (N_1987,In_180,In_961);
or U1988 (N_1988,In_821,In_171);
or U1989 (N_1989,In_983,In_780);
and U1990 (N_1990,In_418,In_1167);
nand U1991 (N_1991,In_448,In_911);
nor U1992 (N_1992,In_1343,In_664);
nor U1993 (N_1993,In_346,In_853);
nor U1994 (N_1994,In_864,In_1363);
and U1995 (N_1995,In_51,In_63);
and U1996 (N_1996,In_458,In_326);
and U1997 (N_1997,In_111,In_1442);
or U1998 (N_1998,In_93,In_1397);
or U1999 (N_1999,In_715,In_773);
and U2000 (N_2000,In_996,In_258);
nand U2001 (N_2001,In_749,In_425);
nor U2002 (N_2002,In_629,In_551);
nand U2003 (N_2003,In_1139,In_1208);
or U2004 (N_2004,In_337,In_784);
or U2005 (N_2005,In_933,In_653);
nand U2006 (N_2006,In_403,In_68);
nor U2007 (N_2007,In_1404,In_391);
nor U2008 (N_2008,In_12,In_643);
and U2009 (N_2009,In_320,In_800);
nor U2010 (N_2010,In_174,In_546);
and U2011 (N_2011,In_522,In_637);
nor U2012 (N_2012,In_1154,In_429);
nand U2013 (N_2013,In_40,In_835);
nand U2014 (N_2014,In_604,In_933);
and U2015 (N_2015,In_1113,In_503);
nand U2016 (N_2016,In_468,In_65);
or U2017 (N_2017,In_354,In_675);
and U2018 (N_2018,In_323,In_375);
nor U2019 (N_2019,In_535,In_1162);
and U2020 (N_2020,In_1233,In_1419);
xnor U2021 (N_2021,In_599,In_1113);
and U2022 (N_2022,In_1499,In_788);
or U2023 (N_2023,In_1491,In_73);
nand U2024 (N_2024,In_1478,In_827);
and U2025 (N_2025,In_556,In_1094);
nor U2026 (N_2026,In_739,In_1227);
nor U2027 (N_2027,In_1273,In_462);
xor U2028 (N_2028,In_509,In_433);
nor U2029 (N_2029,In_410,In_518);
nor U2030 (N_2030,In_679,In_1293);
and U2031 (N_2031,In_1030,In_1197);
nand U2032 (N_2032,In_889,In_1107);
and U2033 (N_2033,In_1342,In_832);
nor U2034 (N_2034,In_223,In_36);
nand U2035 (N_2035,In_204,In_1293);
nor U2036 (N_2036,In_1432,In_1390);
or U2037 (N_2037,In_20,In_1062);
or U2038 (N_2038,In_281,In_304);
nor U2039 (N_2039,In_1087,In_795);
or U2040 (N_2040,In_245,In_212);
nand U2041 (N_2041,In_920,In_649);
or U2042 (N_2042,In_1325,In_431);
nor U2043 (N_2043,In_987,In_1330);
nand U2044 (N_2044,In_1481,In_1073);
nand U2045 (N_2045,In_93,In_869);
nor U2046 (N_2046,In_391,In_629);
or U2047 (N_2047,In_703,In_1155);
nor U2048 (N_2048,In_1225,In_743);
nand U2049 (N_2049,In_1226,In_385);
nor U2050 (N_2050,In_1393,In_985);
nand U2051 (N_2051,In_338,In_246);
nor U2052 (N_2052,In_271,In_1030);
nor U2053 (N_2053,In_43,In_1407);
and U2054 (N_2054,In_1338,In_1365);
or U2055 (N_2055,In_1427,In_192);
and U2056 (N_2056,In_1147,In_1264);
nor U2057 (N_2057,In_1475,In_827);
and U2058 (N_2058,In_641,In_57);
nor U2059 (N_2059,In_1423,In_1029);
or U2060 (N_2060,In_1083,In_214);
nand U2061 (N_2061,In_1480,In_1303);
nor U2062 (N_2062,In_1062,In_187);
nand U2063 (N_2063,In_178,In_968);
and U2064 (N_2064,In_91,In_954);
nor U2065 (N_2065,In_769,In_720);
or U2066 (N_2066,In_1110,In_904);
and U2067 (N_2067,In_951,In_625);
or U2068 (N_2068,In_29,In_457);
nor U2069 (N_2069,In_590,In_1280);
or U2070 (N_2070,In_430,In_399);
nor U2071 (N_2071,In_1081,In_290);
nor U2072 (N_2072,In_270,In_1206);
nor U2073 (N_2073,In_176,In_368);
or U2074 (N_2074,In_420,In_1412);
nand U2075 (N_2075,In_100,In_607);
or U2076 (N_2076,In_38,In_561);
nor U2077 (N_2077,In_612,In_1169);
nand U2078 (N_2078,In_918,In_853);
nor U2079 (N_2079,In_709,In_998);
and U2080 (N_2080,In_824,In_151);
and U2081 (N_2081,In_1121,In_697);
or U2082 (N_2082,In_258,In_662);
nor U2083 (N_2083,In_23,In_940);
nand U2084 (N_2084,In_83,In_138);
and U2085 (N_2085,In_794,In_725);
or U2086 (N_2086,In_511,In_622);
and U2087 (N_2087,In_932,In_124);
nor U2088 (N_2088,In_1217,In_481);
nand U2089 (N_2089,In_96,In_501);
nor U2090 (N_2090,In_737,In_812);
nor U2091 (N_2091,In_321,In_784);
nor U2092 (N_2092,In_1265,In_566);
xnor U2093 (N_2093,In_1279,In_412);
nand U2094 (N_2094,In_868,In_1232);
nand U2095 (N_2095,In_56,In_810);
nand U2096 (N_2096,In_249,In_301);
nor U2097 (N_2097,In_387,In_110);
nand U2098 (N_2098,In_433,In_522);
and U2099 (N_2099,In_877,In_1363);
nand U2100 (N_2100,In_1406,In_736);
nor U2101 (N_2101,In_1403,In_964);
nand U2102 (N_2102,In_1330,In_464);
and U2103 (N_2103,In_699,In_140);
nor U2104 (N_2104,In_1268,In_812);
nor U2105 (N_2105,In_665,In_331);
nand U2106 (N_2106,In_838,In_218);
or U2107 (N_2107,In_856,In_548);
nand U2108 (N_2108,In_554,In_514);
xnor U2109 (N_2109,In_845,In_752);
and U2110 (N_2110,In_712,In_1488);
nor U2111 (N_2111,In_356,In_561);
or U2112 (N_2112,In_832,In_372);
xor U2113 (N_2113,In_270,In_937);
nand U2114 (N_2114,In_661,In_1138);
nand U2115 (N_2115,In_74,In_1473);
nor U2116 (N_2116,In_403,In_1150);
or U2117 (N_2117,In_1065,In_1470);
nor U2118 (N_2118,In_1102,In_1260);
or U2119 (N_2119,In_1339,In_1370);
or U2120 (N_2120,In_764,In_1101);
or U2121 (N_2121,In_28,In_485);
and U2122 (N_2122,In_1103,In_296);
or U2123 (N_2123,In_533,In_1413);
nand U2124 (N_2124,In_1119,In_17);
nor U2125 (N_2125,In_161,In_232);
nor U2126 (N_2126,In_881,In_538);
nor U2127 (N_2127,In_136,In_933);
or U2128 (N_2128,In_1276,In_1285);
nand U2129 (N_2129,In_1311,In_256);
nand U2130 (N_2130,In_580,In_755);
and U2131 (N_2131,In_348,In_474);
nor U2132 (N_2132,In_82,In_746);
nor U2133 (N_2133,In_753,In_1384);
nand U2134 (N_2134,In_996,In_384);
or U2135 (N_2135,In_1291,In_1467);
nor U2136 (N_2136,In_1027,In_1261);
nand U2137 (N_2137,In_1147,In_448);
and U2138 (N_2138,In_1113,In_268);
nor U2139 (N_2139,In_244,In_1375);
nand U2140 (N_2140,In_1150,In_1440);
and U2141 (N_2141,In_437,In_907);
and U2142 (N_2142,In_342,In_716);
or U2143 (N_2143,In_977,In_516);
or U2144 (N_2144,In_1044,In_26);
nand U2145 (N_2145,In_671,In_1076);
or U2146 (N_2146,In_583,In_469);
xor U2147 (N_2147,In_1170,In_25);
nand U2148 (N_2148,In_650,In_1294);
nor U2149 (N_2149,In_360,In_1273);
or U2150 (N_2150,In_390,In_506);
nand U2151 (N_2151,In_874,In_384);
nand U2152 (N_2152,In_1186,In_438);
nand U2153 (N_2153,In_1445,In_1486);
or U2154 (N_2154,In_502,In_1477);
and U2155 (N_2155,In_143,In_1195);
and U2156 (N_2156,In_1418,In_1373);
and U2157 (N_2157,In_394,In_167);
or U2158 (N_2158,In_939,In_458);
or U2159 (N_2159,In_1414,In_191);
nor U2160 (N_2160,In_1487,In_753);
nand U2161 (N_2161,In_742,In_568);
and U2162 (N_2162,In_262,In_477);
nand U2163 (N_2163,In_619,In_28);
or U2164 (N_2164,In_287,In_704);
or U2165 (N_2165,In_284,In_22);
and U2166 (N_2166,In_545,In_18);
nand U2167 (N_2167,In_1256,In_64);
nand U2168 (N_2168,In_612,In_1389);
nor U2169 (N_2169,In_1058,In_1477);
or U2170 (N_2170,In_837,In_990);
or U2171 (N_2171,In_1021,In_1197);
or U2172 (N_2172,In_394,In_935);
xor U2173 (N_2173,In_848,In_1005);
or U2174 (N_2174,In_370,In_393);
nand U2175 (N_2175,In_1487,In_705);
nor U2176 (N_2176,In_48,In_604);
nand U2177 (N_2177,In_516,In_427);
xnor U2178 (N_2178,In_424,In_1250);
and U2179 (N_2179,In_526,In_1123);
nand U2180 (N_2180,In_471,In_53);
nand U2181 (N_2181,In_98,In_889);
and U2182 (N_2182,In_1286,In_111);
and U2183 (N_2183,In_804,In_27);
nand U2184 (N_2184,In_291,In_748);
or U2185 (N_2185,In_1354,In_1411);
or U2186 (N_2186,In_1300,In_1405);
nand U2187 (N_2187,In_1071,In_1465);
xor U2188 (N_2188,In_284,In_550);
xnor U2189 (N_2189,In_62,In_1303);
or U2190 (N_2190,In_94,In_1116);
nand U2191 (N_2191,In_684,In_1480);
or U2192 (N_2192,In_601,In_774);
and U2193 (N_2193,In_954,In_973);
or U2194 (N_2194,In_457,In_540);
nor U2195 (N_2195,In_1089,In_370);
nor U2196 (N_2196,In_709,In_428);
nand U2197 (N_2197,In_852,In_209);
nand U2198 (N_2198,In_12,In_716);
nor U2199 (N_2199,In_1088,In_252);
nand U2200 (N_2200,In_1128,In_314);
or U2201 (N_2201,In_989,In_612);
or U2202 (N_2202,In_136,In_332);
or U2203 (N_2203,In_573,In_33);
and U2204 (N_2204,In_134,In_1306);
or U2205 (N_2205,In_989,In_1108);
or U2206 (N_2206,In_815,In_1275);
or U2207 (N_2207,In_322,In_548);
and U2208 (N_2208,In_1151,In_177);
and U2209 (N_2209,In_55,In_1381);
nor U2210 (N_2210,In_145,In_1237);
nor U2211 (N_2211,In_1151,In_777);
nor U2212 (N_2212,In_1479,In_797);
and U2213 (N_2213,In_1044,In_341);
or U2214 (N_2214,In_155,In_1191);
and U2215 (N_2215,In_487,In_1476);
nand U2216 (N_2216,In_779,In_906);
and U2217 (N_2217,In_1006,In_1039);
nor U2218 (N_2218,In_839,In_695);
nor U2219 (N_2219,In_570,In_238);
or U2220 (N_2220,In_1286,In_202);
nand U2221 (N_2221,In_145,In_1105);
and U2222 (N_2222,In_45,In_700);
nand U2223 (N_2223,In_1220,In_641);
xnor U2224 (N_2224,In_544,In_114);
nand U2225 (N_2225,In_631,In_262);
or U2226 (N_2226,In_1456,In_415);
and U2227 (N_2227,In_1472,In_1355);
and U2228 (N_2228,In_233,In_748);
and U2229 (N_2229,In_460,In_109);
and U2230 (N_2230,In_1490,In_919);
nand U2231 (N_2231,In_1253,In_480);
nand U2232 (N_2232,In_264,In_206);
and U2233 (N_2233,In_1498,In_482);
or U2234 (N_2234,In_761,In_421);
and U2235 (N_2235,In_233,In_1110);
nor U2236 (N_2236,In_591,In_191);
or U2237 (N_2237,In_289,In_391);
nor U2238 (N_2238,In_245,In_213);
nand U2239 (N_2239,In_1230,In_33);
or U2240 (N_2240,In_1047,In_1256);
xor U2241 (N_2241,In_1259,In_174);
or U2242 (N_2242,In_1320,In_1364);
or U2243 (N_2243,In_305,In_1245);
and U2244 (N_2244,In_1085,In_346);
and U2245 (N_2245,In_1192,In_747);
nand U2246 (N_2246,In_722,In_659);
nor U2247 (N_2247,In_714,In_432);
nor U2248 (N_2248,In_1142,In_583);
or U2249 (N_2249,In_883,In_191);
or U2250 (N_2250,In_109,In_121);
or U2251 (N_2251,In_585,In_128);
xnor U2252 (N_2252,In_1036,In_741);
and U2253 (N_2253,In_876,In_996);
nand U2254 (N_2254,In_839,In_96);
or U2255 (N_2255,In_307,In_1102);
and U2256 (N_2256,In_309,In_252);
and U2257 (N_2257,In_210,In_793);
or U2258 (N_2258,In_192,In_322);
or U2259 (N_2259,In_573,In_680);
and U2260 (N_2260,In_636,In_631);
or U2261 (N_2261,In_783,In_1241);
or U2262 (N_2262,In_279,In_923);
and U2263 (N_2263,In_1330,In_870);
or U2264 (N_2264,In_49,In_1164);
nor U2265 (N_2265,In_615,In_987);
nand U2266 (N_2266,In_999,In_1198);
nor U2267 (N_2267,In_460,In_1236);
or U2268 (N_2268,In_563,In_1126);
nand U2269 (N_2269,In_1481,In_474);
nor U2270 (N_2270,In_739,In_204);
nand U2271 (N_2271,In_583,In_41);
or U2272 (N_2272,In_876,In_1172);
and U2273 (N_2273,In_970,In_513);
or U2274 (N_2274,In_48,In_1379);
or U2275 (N_2275,In_1455,In_153);
or U2276 (N_2276,In_1326,In_1399);
nor U2277 (N_2277,In_1471,In_716);
and U2278 (N_2278,In_954,In_1250);
or U2279 (N_2279,In_1253,In_172);
nand U2280 (N_2280,In_450,In_349);
and U2281 (N_2281,In_984,In_710);
or U2282 (N_2282,In_209,In_607);
nand U2283 (N_2283,In_249,In_70);
and U2284 (N_2284,In_384,In_1490);
and U2285 (N_2285,In_1413,In_58);
or U2286 (N_2286,In_1427,In_506);
nand U2287 (N_2287,In_366,In_1455);
or U2288 (N_2288,In_665,In_854);
nor U2289 (N_2289,In_295,In_1232);
nand U2290 (N_2290,In_906,In_182);
and U2291 (N_2291,In_1414,In_1036);
or U2292 (N_2292,In_399,In_1205);
and U2293 (N_2293,In_784,In_1127);
nor U2294 (N_2294,In_175,In_1152);
or U2295 (N_2295,In_248,In_177);
or U2296 (N_2296,In_726,In_737);
and U2297 (N_2297,In_97,In_892);
and U2298 (N_2298,In_5,In_1044);
nand U2299 (N_2299,In_1229,In_680);
or U2300 (N_2300,In_757,In_577);
nand U2301 (N_2301,In_1042,In_1320);
nand U2302 (N_2302,In_721,In_212);
and U2303 (N_2303,In_912,In_507);
nor U2304 (N_2304,In_1465,In_885);
nor U2305 (N_2305,In_1088,In_390);
nor U2306 (N_2306,In_989,In_368);
xnor U2307 (N_2307,In_710,In_826);
nand U2308 (N_2308,In_1099,In_1235);
nand U2309 (N_2309,In_779,In_630);
and U2310 (N_2310,In_1071,In_1120);
nand U2311 (N_2311,In_102,In_1237);
or U2312 (N_2312,In_434,In_855);
or U2313 (N_2313,In_286,In_1230);
nor U2314 (N_2314,In_24,In_694);
nand U2315 (N_2315,In_124,In_650);
and U2316 (N_2316,In_454,In_743);
or U2317 (N_2317,In_595,In_119);
or U2318 (N_2318,In_899,In_917);
and U2319 (N_2319,In_572,In_305);
nor U2320 (N_2320,In_152,In_1321);
and U2321 (N_2321,In_351,In_1295);
nand U2322 (N_2322,In_332,In_129);
nor U2323 (N_2323,In_186,In_509);
or U2324 (N_2324,In_1395,In_135);
nand U2325 (N_2325,In_898,In_1405);
nor U2326 (N_2326,In_684,In_373);
xnor U2327 (N_2327,In_680,In_707);
nand U2328 (N_2328,In_264,In_566);
or U2329 (N_2329,In_930,In_346);
or U2330 (N_2330,In_1130,In_998);
nor U2331 (N_2331,In_262,In_197);
nand U2332 (N_2332,In_1357,In_655);
or U2333 (N_2333,In_756,In_777);
nor U2334 (N_2334,In_1197,In_1320);
or U2335 (N_2335,In_131,In_733);
or U2336 (N_2336,In_1346,In_1010);
and U2337 (N_2337,In_470,In_603);
and U2338 (N_2338,In_551,In_470);
and U2339 (N_2339,In_177,In_467);
nand U2340 (N_2340,In_964,In_56);
and U2341 (N_2341,In_1000,In_1298);
nand U2342 (N_2342,In_597,In_642);
nand U2343 (N_2343,In_1433,In_1079);
nor U2344 (N_2344,In_431,In_1245);
nand U2345 (N_2345,In_788,In_34);
and U2346 (N_2346,In_923,In_1214);
or U2347 (N_2347,In_964,In_1115);
nor U2348 (N_2348,In_324,In_927);
or U2349 (N_2349,In_987,In_1028);
nand U2350 (N_2350,In_1020,In_220);
and U2351 (N_2351,In_356,In_152);
nand U2352 (N_2352,In_1027,In_340);
nor U2353 (N_2353,In_10,In_125);
xor U2354 (N_2354,In_730,In_1159);
nor U2355 (N_2355,In_1372,In_115);
or U2356 (N_2356,In_630,In_1359);
nand U2357 (N_2357,In_66,In_945);
nor U2358 (N_2358,In_1027,In_659);
or U2359 (N_2359,In_555,In_663);
nor U2360 (N_2360,In_158,In_127);
nor U2361 (N_2361,In_802,In_228);
or U2362 (N_2362,In_612,In_2);
or U2363 (N_2363,In_1232,In_1247);
and U2364 (N_2364,In_550,In_696);
and U2365 (N_2365,In_280,In_165);
nor U2366 (N_2366,In_861,In_724);
and U2367 (N_2367,In_18,In_458);
nand U2368 (N_2368,In_416,In_1065);
xor U2369 (N_2369,In_772,In_1037);
and U2370 (N_2370,In_943,In_882);
nor U2371 (N_2371,In_266,In_1385);
or U2372 (N_2372,In_1314,In_1185);
and U2373 (N_2373,In_1338,In_368);
nand U2374 (N_2374,In_523,In_409);
nand U2375 (N_2375,In_124,In_1316);
nor U2376 (N_2376,In_1386,In_53);
nor U2377 (N_2377,In_1404,In_732);
or U2378 (N_2378,In_723,In_681);
or U2379 (N_2379,In_554,In_7);
xnor U2380 (N_2380,In_1124,In_762);
nor U2381 (N_2381,In_777,In_322);
nor U2382 (N_2382,In_250,In_1067);
xor U2383 (N_2383,In_920,In_1185);
and U2384 (N_2384,In_793,In_1373);
xnor U2385 (N_2385,In_962,In_780);
or U2386 (N_2386,In_1083,In_1263);
nor U2387 (N_2387,In_384,In_1092);
nand U2388 (N_2388,In_286,In_1335);
and U2389 (N_2389,In_331,In_1341);
or U2390 (N_2390,In_897,In_347);
xor U2391 (N_2391,In_947,In_688);
nand U2392 (N_2392,In_1065,In_1007);
nand U2393 (N_2393,In_1148,In_1291);
or U2394 (N_2394,In_688,In_1176);
and U2395 (N_2395,In_673,In_770);
and U2396 (N_2396,In_1086,In_1185);
and U2397 (N_2397,In_719,In_6);
or U2398 (N_2398,In_760,In_21);
nand U2399 (N_2399,In_1168,In_564);
and U2400 (N_2400,In_257,In_1218);
nor U2401 (N_2401,In_857,In_883);
or U2402 (N_2402,In_1238,In_221);
or U2403 (N_2403,In_244,In_1321);
nor U2404 (N_2404,In_54,In_503);
nor U2405 (N_2405,In_1324,In_563);
xor U2406 (N_2406,In_556,In_450);
or U2407 (N_2407,In_460,In_1280);
and U2408 (N_2408,In_880,In_1441);
or U2409 (N_2409,In_735,In_111);
or U2410 (N_2410,In_1317,In_1226);
or U2411 (N_2411,In_1091,In_765);
nor U2412 (N_2412,In_667,In_1336);
and U2413 (N_2413,In_1162,In_274);
or U2414 (N_2414,In_1205,In_51);
nor U2415 (N_2415,In_274,In_75);
and U2416 (N_2416,In_1230,In_184);
nand U2417 (N_2417,In_1062,In_810);
or U2418 (N_2418,In_887,In_62);
or U2419 (N_2419,In_496,In_586);
and U2420 (N_2420,In_197,In_156);
nor U2421 (N_2421,In_301,In_1147);
or U2422 (N_2422,In_137,In_547);
nor U2423 (N_2423,In_1157,In_1027);
nor U2424 (N_2424,In_128,In_647);
or U2425 (N_2425,In_803,In_624);
and U2426 (N_2426,In_1383,In_1178);
and U2427 (N_2427,In_756,In_1124);
and U2428 (N_2428,In_862,In_1174);
nand U2429 (N_2429,In_1113,In_1240);
and U2430 (N_2430,In_153,In_675);
and U2431 (N_2431,In_352,In_897);
and U2432 (N_2432,In_1209,In_1225);
nand U2433 (N_2433,In_1362,In_736);
and U2434 (N_2434,In_1481,In_1054);
or U2435 (N_2435,In_5,In_1092);
nand U2436 (N_2436,In_149,In_832);
or U2437 (N_2437,In_403,In_468);
or U2438 (N_2438,In_1319,In_664);
nand U2439 (N_2439,In_235,In_780);
and U2440 (N_2440,In_971,In_845);
nand U2441 (N_2441,In_203,In_1262);
or U2442 (N_2442,In_655,In_764);
or U2443 (N_2443,In_1470,In_1245);
nor U2444 (N_2444,In_247,In_10);
nand U2445 (N_2445,In_1025,In_248);
or U2446 (N_2446,In_295,In_370);
nand U2447 (N_2447,In_474,In_1330);
or U2448 (N_2448,In_291,In_556);
or U2449 (N_2449,In_627,In_22);
or U2450 (N_2450,In_1196,In_1032);
nand U2451 (N_2451,In_649,In_642);
nand U2452 (N_2452,In_1064,In_1079);
or U2453 (N_2453,In_768,In_1136);
nand U2454 (N_2454,In_368,In_746);
and U2455 (N_2455,In_716,In_1367);
and U2456 (N_2456,In_1296,In_651);
nand U2457 (N_2457,In_865,In_993);
and U2458 (N_2458,In_289,In_380);
and U2459 (N_2459,In_787,In_1484);
or U2460 (N_2460,In_58,In_1071);
and U2461 (N_2461,In_712,In_854);
and U2462 (N_2462,In_201,In_1099);
nand U2463 (N_2463,In_617,In_310);
and U2464 (N_2464,In_989,In_629);
or U2465 (N_2465,In_234,In_398);
nand U2466 (N_2466,In_1457,In_1135);
nand U2467 (N_2467,In_86,In_328);
and U2468 (N_2468,In_120,In_1484);
and U2469 (N_2469,In_53,In_989);
nor U2470 (N_2470,In_543,In_481);
nand U2471 (N_2471,In_367,In_1482);
or U2472 (N_2472,In_280,In_647);
nand U2473 (N_2473,In_1027,In_851);
or U2474 (N_2474,In_292,In_157);
nor U2475 (N_2475,In_65,In_835);
nor U2476 (N_2476,In_449,In_724);
nand U2477 (N_2477,In_726,In_170);
nand U2478 (N_2478,In_388,In_1158);
and U2479 (N_2479,In_1250,In_852);
nand U2480 (N_2480,In_1426,In_861);
nand U2481 (N_2481,In_1251,In_1438);
nor U2482 (N_2482,In_1240,In_863);
or U2483 (N_2483,In_189,In_1144);
nand U2484 (N_2484,In_1237,In_473);
nor U2485 (N_2485,In_1073,In_78);
nor U2486 (N_2486,In_859,In_567);
nor U2487 (N_2487,In_1238,In_890);
nor U2488 (N_2488,In_1392,In_1398);
xnor U2489 (N_2489,In_699,In_266);
nand U2490 (N_2490,In_1133,In_1254);
and U2491 (N_2491,In_633,In_150);
nor U2492 (N_2492,In_1342,In_1157);
nor U2493 (N_2493,In_951,In_773);
nor U2494 (N_2494,In_860,In_351);
or U2495 (N_2495,In_805,In_787);
nor U2496 (N_2496,In_64,In_663);
or U2497 (N_2497,In_199,In_432);
or U2498 (N_2498,In_271,In_194);
nor U2499 (N_2499,In_229,In_624);
nor U2500 (N_2500,In_943,In_296);
and U2501 (N_2501,In_1314,In_1041);
nand U2502 (N_2502,In_440,In_341);
nor U2503 (N_2503,In_250,In_946);
nand U2504 (N_2504,In_1009,In_1179);
nor U2505 (N_2505,In_337,In_1290);
and U2506 (N_2506,In_1196,In_1473);
and U2507 (N_2507,In_1317,In_836);
nand U2508 (N_2508,In_1206,In_855);
nand U2509 (N_2509,In_90,In_790);
and U2510 (N_2510,In_1371,In_437);
nor U2511 (N_2511,In_1184,In_18);
nor U2512 (N_2512,In_330,In_322);
or U2513 (N_2513,In_17,In_578);
or U2514 (N_2514,In_1122,In_493);
nand U2515 (N_2515,In_588,In_1249);
and U2516 (N_2516,In_1468,In_552);
and U2517 (N_2517,In_470,In_1092);
or U2518 (N_2518,In_964,In_280);
and U2519 (N_2519,In_1074,In_730);
or U2520 (N_2520,In_161,In_1289);
or U2521 (N_2521,In_1364,In_686);
or U2522 (N_2522,In_272,In_1290);
and U2523 (N_2523,In_40,In_1431);
and U2524 (N_2524,In_1248,In_208);
nor U2525 (N_2525,In_1029,In_1121);
nand U2526 (N_2526,In_1057,In_1052);
nor U2527 (N_2527,In_1214,In_156);
nor U2528 (N_2528,In_589,In_1421);
nor U2529 (N_2529,In_332,In_214);
or U2530 (N_2530,In_881,In_1397);
nor U2531 (N_2531,In_719,In_71);
or U2532 (N_2532,In_923,In_374);
nand U2533 (N_2533,In_1490,In_879);
or U2534 (N_2534,In_1435,In_266);
or U2535 (N_2535,In_960,In_736);
and U2536 (N_2536,In_957,In_628);
nor U2537 (N_2537,In_1320,In_991);
and U2538 (N_2538,In_99,In_454);
nor U2539 (N_2539,In_968,In_49);
nor U2540 (N_2540,In_722,In_753);
nor U2541 (N_2541,In_611,In_678);
and U2542 (N_2542,In_991,In_559);
nand U2543 (N_2543,In_1096,In_1302);
nor U2544 (N_2544,In_783,In_562);
nor U2545 (N_2545,In_113,In_704);
or U2546 (N_2546,In_1257,In_249);
and U2547 (N_2547,In_127,In_1293);
nor U2548 (N_2548,In_14,In_216);
nor U2549 (N_2549,In_1072,In_213);
and U2550 (N_2550,In_612,In_1426);
and U2551 (N_2551,In_1245,In_68);
or U2552 (N_2552,In_276,In_558);
or U2553 (N_2553,In_640,In_576);
nor U2554 (N_2554,In_796,In_1048);
and U2555 (N_2555,In_1485,In_1436);
nor U2556 (N_2556,In_634,In_272);
xor U2557 (N_2557,In_877,In_847);
nor U2558 (N_2558,In_619,In_430);
nand U2559 (N_2559,In_1076,In_752);
or U2560 (N_2560,In_815,In_226);
and U2561 (N_2561,In_862,In_800);
nand U2562 (N_2562,In_14,In_450);
or U2563 (N_2563,In_691,In_198);
or U2564 (N_2564,In_1044,In_1279);
nor U2565 (N_2565,In_1330,In_81);
nor U2566 (N_2566,In_475,In_1035);
and U2567 (N_2567,In_1409,In_535);
nor U2568 (N_2568,In_73,In_1473);
or U2569 (N_2569,In_999,In_1391);
and U2570 (N_2570,In_559,In_1439);
and U2571 (N_2571,In_990,In_341);
or U2572 (N_2572,In_270,In_1240);
nand U2573 (N_2573,In_809,In_1018);
nand U2574 (N_2574,In_1466,In_1162);
nand U2575 (N_2575,In_1022,In_1427);
or U2576 (N_2576,In_357,In_1275);
and U2577 (N_2577,In_373,In_883);
nor U2578 (N_2578,In_503,In_1265);
nor U2579 (N_2579,In_787,In_989);
or U2580 (N_2580,In_904,In_148);
and U2581 (N_2581,In_617,In_892);
or U2582 (N_2582,In_639,In_1070);
or U2583 (N_2583,In_717,In_1158);
and U2584 (N_2584,In_236,In_872);
or U2585 (N_2585,In_368,In_15);
nand U2586 (N_2586,In_45,In_26);
or U2587 (N_2587,In_440,In_234);
or U2588 (N_2588,In_1444,In_1023);
nand U2589 (N_2589,In_1100,In_519);
nor U2590 (N_2590,In_264,In_1404);
nand U2591 (N_2591,In_434,In_323);
or U2592 (N_2592,In_907,In_352);
nand U2593 (N_2593,In_496,In_296);
nand U2594 (N_2594,In_868,In_1376);
or U2595 (N_2595,In_13,In_888);
or U2596 (N_2596,In_801,In_144);
or U2597 (N_2597,In_1026,In_364);
nor U2598 (N_2598,In_817,In_1060);
and U2599 (N_2599,In_902,In_701);
or U2600 (N_2600,In_918,In_1270);
or U2601 (N_2601,In_1256,In_928);
xor U2602 (N_2602,In_364,In_604);
or U2603 (N_2603,In_708,In_1362);
and U2604 (N_2604,In_463,In_1056);
nor U2605 (N_2605,In_26,In_978);
and U2606 (N_2606,In_1200,In_301);
and U2607 (N_2607,In_1112,In_141);
and U2608 (N_2608,In_908,In_950);
nor U2609 (N_2609,In_21,In_574);
or U2610 (N_2610,In_1404,In_1144);
nor U2611 (N_2611,In_878,In_1150);
nor U2612 (N_2612,In_1080,In_621);
and U2613 (N_2613,In_135,In_970);
nand U2614 (N_2614,In_970,In_341);
and U2615 (N_2615,In_83,In_1045);
nand U2616 (N_2616,In_634,In_664);
nor U2617 (N_2617,In_724,In_238);
and U2618 (N_2618,In_384,In_334);
nand U2619 (N_2619,In_1181,In_480);
and U2620 (N_2620,In_773,In_341);
nand U2621 (N_2621,In_534,In_1302);
and U2622 (N_2622,In_913,In_1056);
nor U2623 (N_2623,In_781,In_1441);
or U2624 (N_2624,In_1372,In_711);
nor U2625 (N_2625,In_754,In_123);
or U2626 (N_2626,In_56,In_451);
nor U2627 (N_2627,In_193,In_1298);
nor U2628 (N_2628,In_1413,In_611);
or U2629 (N_2629,In_920,In_1008);
nor U2630 (N_2630,In_944,In_907);
nor U2631 (N_2631,In_1349,In_945);
and U2632 (N_2632,In_1260,In_1127);
or U2633 (N_2633,In_1109,In_1111);
nand U2634 (N_2634,In_1481,In_411);
nor U2635 (N_2635,In_132,In_1352);
xor U2636 (N_2636,In_872,In_271);
and U2637 (N_2637,In_318,In_496);
or U2638 (N_2638,In_1066,In_1050);
nor U2639 (N_2639,In_928,In_425);
nor U2640 (N_2640,In_323,In_1498);
nor U2641 (N_2641,In_599,In_687);
nor U2642 (N_2642,In_317,In_833);
nand U2643 (N_2643,In_728,In_918);
and U2644 (N_2644,In_548,In_1398);
nand U2645 (N_2645,In_277,In_37);
and U2646 (N_2646,In_1372,In_1271);
and U2647 (N_2647,In_772,In_1191);
and U2648 (N_2648,In_1340,In_909);
and U2649 (N_2649,In_286,In_1215);
or U2650 (N_2650,In_21,In_1481);
or U2651 (N_2651,In_374,In_821);
nor U2652 (N_2652,In_742,In_769);
and U2653 (N_2653,In_875,In_1206);
and U2654 (N_2654,In_2,In_1014);
and U2655 (N_2655,In_863,In_240);
nand U2656 (N_2656,In_1008,In_1364);
or U2657 (N_2657,In_634,In_164);
nor U2658 (N_2658,In_429,In_262);
nand U2659 (N_2659,In_838,In_140);
nor U2660 (N_2660,In_1336,In_981);
and U2661 (N_2661,In_1316,In_646);
or U2662 (N_2662,In_1187,In_633);
or U2663 (N_2663,In_622,In_167);
or U2664 (N_2664,In_707,In_156);
nand U2665 (N_2665,In_470,In_1063);
nor U2666 (N_2666,In_383,In_879);
or U2667 (N_2667,In_696,In_15);
and U2668 (N_2668,In_1444,In_1419);
or U2669 (N_2669,In_1090,In_672);
and U2670 (N_2670,In_417,In_18);
nor U2671 (N_2671,In_222,In_1293);
or U2672 (N_2672,In_105,In_1381);
nand U2673 (N_2673,In_977,In_1004);
and U2674 (N_2674,In_1340,In_760);
and U2675 (N_2675,In_1134,In_13);
and U2676 (N_2676,In_1290,In_505);
and U2677 (N_2677,In_187,In_754);
or U2678 (N_2678,In_1302,In_172);
or U2679 (N_2679,In_795,In_1078);
and U2680 (N_2680,In_780,In_186);
nand U2681 (N_2681,In_668,In_1226);
and U2682 (N_2682,In_363,In_838);
and U2683 (N_2683,In_861,In_802);
and U2684 (N_2684,In_1260,In_1413);
nand U2685 (N_2685,In_700,In_398);
nor U2686 (N_2686,In_316,In_730);
or U2687 (N_2687,In_11,In_1494);
nand U2688 (N_2688,In_895,In_703);
nor U2689 (N_2689,In_964,In_423);
or U2690 (N_2690,In_425,In_1061);
nand U2691 (N_2691,In_476,In_906);
nor U2692 (N_2692,In_1149,In_224);
nor U2693 (N_2693,In_1462,In_1137);
nand U2694 (N_2694,In_486,In_583);
or U2695 (N_2695,In_267,In_1118);
nand U2696 (N_2696,In_1371,In_63);
nand U2697 (N_2697,In_1419,In_1250);
and U2698 (N_2698,In_1347,In_1439);
nand U2699 (N_2699,In_357,In_1189);
nand U2700 (N_2700,In_112,In_1469);
nor U2701 (N_2701,In_1210,In_1309);
and U2702 (N_2702,In_1359,In_940);
or U2703 (N_2703,In_549,In_132);
or U2704 (N_2704,In_1288,In_1371);
nor U2705 (N_2705,In_1345,In_1082);
or U2706 (N_2706,In_1222,In_1228);
nand U2707 (N_2707,In_1359,In_736);
nor U2708 (N_2708,In_902,In_941);
and U2709 (N_2709,In_1068,In_283);
nand U2710 (N_2710,In_947,In_191);
and U2711 (N_2711,In_194,In_717);
nor U2712 (N_2712,In_668,In_961);
and U2713 (N_2713,In_1045,In_614);
nor U2714 (N_2714,In_73,In_1063);
nor U2715 (N_2715,In_380,In_1321);
or U2716 (N_2716,In_1010,In_1143);
nand U2717 (N_2717,In_1406,In_766);
nor U2718 (N_2718,In_1258,In_284);
and U2719 (N_2719,In_893,In_736);
nand U2720 (N_2720,In_236,In_530);
and U2721 (N_2721,In_576,In_1378);
nor U2722 (N_2722,In_653,In_1322);
or U2723 (N_2723,In_663,In_39);
nand U2724 (N_2724,In_105,In_115);
nand U2725 (N_2725,In_704,In_1469);
nor U2726 (N_2726,In_1247,In_549);
nor U2727 (N_2727,In_1496,In_228);
nor U2728 (N_2728,In_98,In_697);
and U2729 (N_2729,In_775,In_1205);
nand U2730 (N_2730,In_502,In_35);
and U2731 (N_2731,In_1325,In_208);
and U2732 (N_2732,In_680,In_1352);
nand U2733 (N_2733,In_381,In_827);
nand U2734 (N_2734,In_1449,In_518);
or U2735 (N_2735,In_456,In_46);
xor U2736 (N_2736,In_245,In_17);
nand U2737 (N_2737,In_906,In_683);
and U2738 (N_2738,In_1337,In_63);
nor U2739 (N_2739,In_624,In_1169);
or U2740 (N_2740,In_719,In_1006);
xnor U2741 (N_2741,In_208,In_1182);
nor U2742 (N_2742,In_1161,In_544);
or U2743 (N_2743,In_145,In_1383);
and U2744 (N_2744,In_47,In_1297);
nor U2745 (N_2745,In_864,In_644);
and U2746 (N_2746,In_786,In_696);
nand U2747 (N_2747,In_1495,In_508);
and U2748 (N_2748,In_524,In_357);
and U2749 (N_2749,In_371,In_394);
and U2750 (N_2750,In_162,In_1283);
and U2751 (N_2751,In_1339,In_382);
nand U2752 (N_2752,In_460,In_901);
or U2753 (N_2753,In_388,In_823);
nand U2754 (N_2754,In_242,In_1225);
nand U2755 (N_2755,In_33,In_1276);
nor U2756 (N_2756,In_36,In_123);
nand U2757 (N_2757,In_934,In_1154);
nand U2758 (N_2758,In_409,In_740);
or U2759 (N_2759,In_100,In_36);
nor U2760 (N_2760,In_875,In_787);
xor U2761 (N_2761,In_696,In_602);
nand U2762 (N_2762,In_382,In_1249);
nand U2763 (N_2763,In_1434,In_210);
and U2764 (N_2764,In_395,In_587);
and U2765 (N_2765,In_676,In_627);
nand U2766 (N_2766,In_1260,In_769);
and U2767 (N_2767,In_129,In_749);
nor U2768 (N_2768,In_1308,In_228);
or U2769 (N_2769,In_599,In_211);
nor U2770 (N_2770,In_1332,In_284);
or U2771 (N_2771,In_658,In_743);
nand U2772 (N_2772,In_132,In_631);
or U2773 (N_2773,In_1303,In_293);
nor U2774 (N_2774,In_734,In_1412);
and U2775 (N_2775,In_872,In_1173);
or U2776 (N_2776,In_222,In_156);
nor U2777 (N_2777,In_832,In_133);
or U2778 (N_2778,In_812,In_1384);
and U2779 (N_2779,In_967,In_403);
nand U2780 (N_2780,In_1156,In_328);
or U2781 (N_2781,In_1058,In_917);
nand U2782 (N_2782,In_808,In_1190);
nand U2783 (N_2783,In_1333,In_536);
and U2784 (N_2784,In_865,In_414);
nor U2785 (N_2785,In_1256,In_334);
nor U2786 (N_2786,In_1172,In_1202);
nor U2787 (N_2787,In_272,In_1286);
nand U2788 (N_2788,In_64,In_1051);
nor U2789 (N_2789,In_1351,In_156);
nand U2790 (N_2790,In_1442,In_514);
nand U2791 (N_2791,In_66,In_529);
and U2792 (N_2792,In_589,In_301);
nand U2793 (N_2793,In_1006,In_75);
and U2794 (N_2794,In_475,In_1067);
or U2795 (N_2795,In_245,In_881);
nand U2796 (N_2796,In_1472,In_379);
nor U2797 (N_2797,In_1353,In_50);
and U2798 (N_2798,In_952,In_251);
or U2799 (N_2799,In_608,In_1245);
nand U2800 (N_2800,In_143,In_764);
nor U2801 (N_2801,In_550,In_133);
or U2802 (N_2802,In_1125,In_1365);
nand U2803 (N_2803,In_634,In_1212);
nor U2804 (N_2804,In_1300,In_1443);
and U2805 (N_2805,In_250,In_1315);
nand U2806 (N_2806,In_1072,In_473);
xor U2807 (N_2807,In_629,In_805);
and U2808 (N_2808,In_66,In_489);
and U2809 (N_2809,In_967,In_1345);
nor U2810 (N_2810,In_1455,In_57);
nand U2811 (N_2811,In_619,In_193);
nand U2812 (N_2812,In_1244,In_339);
nand U2813 (N_2813,In_816,In_1259);
nor U2814 (N_2814,In_678,In_928);
nand U2815 (N_2815,In_674,In_391);
or U2816 (N_2816,In_610,In_794);
nand U2817 (N_2817,In_1451,In_188);
or U2818 (N_2818,In_846,In_526);
or U2819 (N_2819,In_519,In_1257);
or U2820 (N_2820,In_446,In_1318);
nor U2821 (N_2821,In_474,In_1146);
nand U2822 (N_2822,In_482,In_290);
nor U2823 (N_2823,In_634,In_387);
nand U2824 (N_2824,In_680,In_491);
xor U2825 (N_2825,In_892,In_904);
or U2826 (N_2826,In_1155,In_64);
nor U2827 (N_2827,In_258,In_18);
or U2828 (N_2828,In_1138,In_440);
and U2829 (N_2829,In_258,In_922);
nor U2830 (N_2830,In_801,In_127);
nor U2831 (N_2831,In_1476,In_877);
nand U2832 (N_2832,In_1473,In_1008);
xor U2833 (N_2833,In_947,In_1389);
or U2834 (N_2834,In_465,In_791);
nand U2835 (N_2835,In_112,In_99);
or U2836 (N_2836,In_121,In_435);
nor U2837 (N_2837,In_1097,In_1316);
and U2838 (N_2838,In_180,In_1321);
and U2839 (N_2839,In_567,In_1117);
nor U2840 (N_2840,In_1384,In_632);
and U2841 (N_2841,In_716,In_477);
or U2842 (N_2842,In_791,In_624);
nand U2843 (N_2843,In_174,In_1046);
nor U2844 (N_2844,In_1324,In_1456);
or U2845 (N_2845,In_316,In_671);
nor U2846 (N_2846,In_219,In_961);
nor U2847 (N_2847,In_101,In_1322);
nor U2848 (N_2848,In_1432,In_718);
nand U2849 (N_2849,In_373,In_1428);
or U2850 (N_2850,In_682,In_744);
nor U2851 (N_2851,In_314,In_1371);
nor U2852 (N_2852,In_1487,In_1218);
or U2853 (N_2853,In_521,In_1067);
nor U2854 (N_2854,In_278,In_383);
nor U2855 (N_2855,In_1471,In_712);
or U2856 (N_2856,In_211,In_611);
and U2857 (N_2857,In_828,In_633);
and U2858 (N_2858,In_334,In_1029);
and U2859 (N_2859,In_1406,In_883);
nor U2860 (N_2860,In_200,In_1315);
or U2861 (N_2861,In_1199,In_89);
nor U2862 (N_2862,In_622,In_155);
xor U2863 (N_2863,In_1498,In_1017);
nor U2864 (N_2864,In_1067,In_1048);
or U2865 (N_2865,In_177,In_1497);
nand U2866 (N_2866,In_779,In_342);
and U2867 (N_2867,In_799,In_1329);
nand U2868 (N_2868,In_1138,In_238);
nand U2869 (N_2869,In_612,In_1236);
nor U2870 (N_2870,In_1325,In_616);
or U2871 (N_2871,In_552,In_78);
and U2872 (N_2872,In_929,In_37);
nor U2873 (N_2873,In_808,In_6);
or U2874 (N_2874,In_297,In_1262);
nand U2875 (N_2875,In_1358,In_669);
nand U2876 (N_2876,In_1383,In_802);
nor U2877 (N_2877,In_1065,In_413);
and U2878 (N_2878,In_1022,In_1479);
nor U2879 (N_2879,In_1031,In_506);
nand U2880 (N_2880,In_1112,In_1432);
nand U2881 (N_2881,In_703,In_1319);
nand U2882 (N_2882,In_1043,In_472);
nor U2883 (N_2883,In_1415,In_765);
or U2884 (N_2884,In_349,In_545);
nor U2885 (N_2885,In_1211,In_1200);
nand U2886 (N_2886,In_415,In_940);
or U2887 (N_2887,In_1008,In_460);
xnor U2888 (N_2888,In_1133,In_1358);
nor U2889 (N_2889,In_1207,In_446);
nor U2890 (N_2890,In_759,In_1363);
xnor U2891 (N_2891,In_504,In_841);
nor U2892 (N_2892,In_660,In_770);
or U2893 (N_2893,In_1423,In_908);
xor U2894 (N_2894,In_334,In_277);
nand U2895 (N_2895,In_1496,In_438);
or U2896 (N_2896,In_1261,In_741);
xnor U2897 (N_2897,In_576,In_651);
and U2898 (N_2898,In_1161,In_1402);
xor U2899 (N_2899,In_33,In_988);
nor U2900 (N_2900,In_52,In_474);
or U2901 (N_2901,In_801,In_894);
nand U2902 (N_2902,In_1026,In_341);
nand U2903 (N_2903,In_472,In_71);
or U2904 (N_2904,In_925,In_406);
nor U2905 (N_2905,In_1102,In_1029);
and U2906 (N_2906,In_288,In_721);
nand U2907 (N_2907,In_230,In_1331);
xor U2908 (N_2908,In_991,In_1319);
or U2909 (N_2909,In_353,In_1013);
nor U2910 (N_2910,In_1233,In_1364);
nor U2911 (N_2911,In_182,In_697);
xnor U2912 (N_2912,In_365,In_836);
nand U2913 (N_2913,In_1447,In_1290);
and U2914 (N_2914,In_541,In_167);
nor U2915 (N_2915,In_486,In_1050);
and U2916 (N_2916,In_1199,In_688);
or U2917 (N_2917,In_995,In_588);
nand U2918 (N_2918,In_801,In_1449);
or U2919 (N_2919,In_447,In_923);
and U2920 (N_2920,In_494,In_1021);
or U2921 (N_2921,In_683,In_536);
nor U2922 (N_2922,In_43,In_365);
nor U2923 (N_2923,In_1471,In_1392);
nor U2924 (N_2924,In_818,In_868);
and U2925 (N_2925,In_1106,In_991);
and U2926 (N_2926,In_511,In_711);
nor U2927 (N_2927,In_1061,In_820);
nor U2928 (N_2928,In_1493,In_518);
or U2929 (N_2929,In_1277,In_525);
nand U2930 (N_2930,In_655,In_1400);
or U2931 (N_2931,In_600,In_1017);
or U2932 (N_2932,In_984,In_535);
or U2933 (N_2933,In_1171,In_687);
and U2934 (N_2934,In_971,In_1245);
and U2935 (N_2935,In_75,In_114);
nor U2936 (N_2936,In_953,In_446);
nand U2937 (N_2937,In_255,In_1492);
nand U2938 (N_2938,In_560,In_1385);
and U2939 (N_2939,In_691,In_1411);
and U2940 (N_2940,In_257,In_618);
or U2941 (N_2941,In_705,In_759);
and U2942 (N_2942,In_946,In_1252);
and U2943 (N_2943,In_673,In_653);
and U2944 (N_2944,In_852,In_570);
nor U2945 (N_2945,In_30,In_484);
nor U2946 (N_2946,In_1024,In_864);
nor U2947 (N_2947,In_269,In_369);
or U2948 (N_2948,In_956,In_734);
nand U2949 (N_2949,In_573,In_721);
nand U2950 (N_2950,In_145,In_811);
nor U2951 (N_2951,In_93,In_1172);
and U2952 (N_2952,In_1369,In_101);
xnor U2953 (N_2953,In_456,In_86);
or U2954 (N_2954,In_1122,In_348);
xnor U2955 (N_2955,In_197,In_1124);
or U2956 (N_2956,In_1334,In_1206);
or U2957 (N_2957,In_982,In_548);
and U2958 (N_2958,In_346,In_362);
nand U2959 (N_2959,In_1447,In_976);
nor U2960 (N_2960,In_200,In_450);
or U2961 (N_2961,In_1270,In_987);
or U2962 (N_2962,In_576,In_124);
and U2963 (N_2963,In_717,In_1088);
or U2964 (N_2964,In_1240,In_728);
nor U2965 (N_2965,In_662,In_1387);
and U2966 (N_2966,In_333,In_317);
nand U2967 (N_2967,In_1293,In_1352);
and U2968 (N_2968,In_1202,In_798);
xnor U2969 (N_2969,In_338,In_876);
nand U2970 (N_2970,In_197,In_1409);
nand U2971 (N_2971,In_875,In_1405);
nor U2972 (N_2972,In_709,In_42);
and U2973 (N_2973,In_92,In_123);
nand U2974 (N_2974,In_1288,In_498);
nor U2975 (N_2975,In_197,In_330);
nor U2976 (N_2976,In_300,In_467);
and U2977 (N_2977,In_1285,In_1178);
and U2978 (N_2978,In_990,In_733);
nor U2979 (N_2979,In_1389,In_1381);
or U2980 (N_2980,In_480,In_398);
and U2981 (N_2981,In_1419,In_922);
nor U2982 (N_2982,In_434,In_107);
or U2983 (N_2983,In_454,In_1085);
and U2984 (N_2984,In_1408,In_1226);
nor U2985 (N_2985,In_1358,In_444);
nand U2986 (N_2986,In_1253,In_484);
nand U2987 (N_2987,In_239,In_829);
xnor U2988 (N_2988,In_521,In_1241);
or U2989 (N_2989,In_516,In_887);
nand U2990 (N_2990,In_497,In_1455);
nand U2991 (N_2991,In_830,In_1296);
and U2992 (N_2992,In_814,In_1287);
or U2993 (N_2993,In_504,In_1309);
or U2994 (N_2994,In_277,In_858);
and U2995 (N_2995,In_229,In_301);
nor U2996 (N_2996,In_843,In_941);
nor U2997 (N_2997,In_264,In_105);
nor U2998 (N_2998,In_1479,In_17);
nor U2999 (N_2999,In_118,In_422);
and U3000 (N_3000,N_1628,N_2254);
and U3001 (N_3001,N_155,N_1274);
and U3002 (N_3002,N_1434,N_2898);
and U3003 (N_3003,N_1523,N_584);
nor U3004 (N_3004,N_617,N_1698);
nor U3005 (N_3005,N_1531,N_871);
and U3006 (N_3006,N_317,N_1684);
nand U3007 (N_3007,N_1233,N_866);
nand U3008 (N_3008,N_2496,N_934);
and U3009 (N_3009,N_2630,N_2750);
nor U3010 (N_3010,N_2946,N_1824);
nand U3011 (N_3011,N_2873,N_414);
nand U3012 (N_3012,N_327,N_873);
or U3013 (N_3013,N_1360,N_2222);
or U3014 (N_3014,N_861,N_2869);
or U3015 (N_3015,N_2766,N_1273);
and U3016 (N_3016,N_1305,N_1849);
nor U3017 (N_3017,N_1891,N_1419);
and U3018 (N_3018,N_769,N_1497);
nor U3019 (N_3019,N_2552,N_2439);
or U3020 (N_3020,N_969,N_1045);
and U3021 (N_3021,N_252,N_2374);
and U3022 (N_3022,N_1030,N_2690);
nor U3023 (N_3023,N_185,N_994);
or U3024 (N_3024,N_716,N_87);
or U3025 (N_3025,N_1676,N_876);
and U3026 (N_3026,N_1143,N_825);
nand U3027 (N_3027,N_1620,N_1644);
nor U3028 (N_3028,N_2595,N_1812);
or U3029 (N_3029,N_2246,N_1744);
nor U3030 (N_3030,N_1998,N_482);
nand U3031 (N_3031,N_2981,N_804);
and U3032 (N_3032,N_157,N_791);
and U3033 (N_3033,N_2270,N_2015);
or U3034 (N_3034,N_1560,N_2559);
nor U3035 (N_3035,N_1976,N_667);
or U3036 (N_3036,N_776,N_1321);
or U3037 (N_3037,N_2033,N_595);
or U3038 (N_3038,N_1788,N_536);
nand U3039 (N_3039,N_2112,N_2648);
nand U3040 (N_3040,N_2892,N_1734);
nor U3041 (N_3041,N_1974,N_402);
nand U3042 (N_3042,N_950,N_2206);
nand U3043 (N_3043,N_51,N_1341);
nand U3044 (N_3044,N_2776,N_451);
or U3045 (N_3045,N_2834,N_2515);
or U3046 (N_3046,N_2262,N_1185);
or U3047 (N_3047,N_212,N_2263);
or U3048 (N_3048,N_2364,N_1847);
nand U3049 (N_3049,N_1611,N_15);
or U3050 (N_3050,N_892,N_2797);
nand U3051 (N_3051,N_9,N_384);
and U3052 (N_3052,N_405,N_1906);
nor U3053 (N_3053,N_2914,N_2391);
or U3054 (N_3054,N_2907,N_1265);
and U3055 (N_3055,N_683,N_2144);
nand U3056 (N_3056,N_1845,N_160);
nand U3057 (N_3057,N_633,N_465);
nor U3058 (N_3058,N_2772,N_135);
nand U3059 (N_3059,N_189,N_489);
or U3060 (N_3060,N_1390,N_166);
and U3061 (N_3061,N_167,N_256);
xor U3062 (N_3062,N_455,N_365);
nand U3063 (N_3063,N_1863,N_2445);
and U3064 (N_3064,N_314,N_2302);
and U3065 (N_3065,N_250,N_1940);
and U3066 (N_3066,N_448,N_2700);
or U3067 (N_3067,N_2028,N_1899);
xor U3068 (N_3068,N_799,N_2352);
or U3069 (N_3069,N_968,N_26);
and U3070 (N_3070,N_2163,N_1603);
nand U3071 (N_3071,N_980,N_193);
nand U3072 (N_3072,N_2945,N_88);
nand U3073 (N_3073,N_2232,N_2444);
and U3074 (N_3074,N_2782,N_1078);
or U3075 (N_3075,N_294,N_2920);
and U3076 (N_3076,N_509,N_1748);
or U3077 (N_3077,N_1358,N_1890);
nor U3078 (N_3078,N_2878,N_2458);
or U3079 (N_3079,N_2737,N_715);
xor U3080 (N_3080,N_757,N_534);
nor U3081 (N_3081,N_1039,N_94);
and U3082 (N_3082,N_1289,N_2937);
nor U3083 (N_3083,N_2716,N_1941);
and U3084 (N_3084,N_608,N_920);
nor U3085 (N_3085,N_1414,N_349);
nor U3086 (N_3086,N_180,N_2377);
and U3087 (N_3087,N_2058,N_1756);
or U3088 (N_3088,N_1510,N_601);
nor U3089 (N_3089,N_1993,N_1687);
and U3090 (N_3090,N_1569,N_880);
and U3091 (N_3091,N_1095,N_1671);
xnor U3092 (N_3092,N_1908,N_1726);
and U3093 (N_3093,N_1913,N_2698);
nand U3094 (N_3094,N_850,N_2047);
nand U3095 (N_3095,N_1140,N_1666);
nor U3096 (N_3096,N_1715,N_2646);
and U3097 (N_3097,N_1134,N_1178);
and U3098 (N_3098,N_2727,N_2528);
and U3099 (N_3099,N_2061,N_1837);
nor U3100 (N_3100,N_1148,N_1464);
or U3101 (N_3101,N_8,N_1429);
and U3102 (N_3102,N_1945,N_2751);
and U3103 (N_3103,N_182,N_2579);
nor U3104 (N_3104,N_293,N_624);
nor U3105 (N_3105,N_471,N_2482);
and U3106 (N_3106,N_1068,N_772);
nor U3107 (N_3107,N_2862,N_792);
or U3108 (N_3108,N_1807,N_2516);
or U3109 (N_3109,N_253,N_2031);
nand U3110 (N_3110,N_100,N_1482);
nor U3111 (N_3111,N_1522,N_918);
nor U3112 (N_3112,N_2647,N_411);
nand U3113 (N_3113,N_756,N_1935);
nor U3114 (N_3114,N_2298,N_267);
or U3115 (N_3115,N_1081,N_1982);
nand U3116 (N_3116,N_1658,N_226);
and U3117 (N_3117,N_1480,N_425);
nand U3118 (N_3118,N_680,N_917);
nand U3119 (N_3119,N_1840,N_266);
xnor U3120 (N_3120,N_1714,N_1761);
or U3121 (N_3121,N_2423,N_2718);
or U3122 (N_3122,N_574,N_2904);
nor U3123 (N_3123,N_1617,N_712);
or U3124 (N_3124,N_2662,N_532);
nand U3125 (N_3125,N_1947,N_2483);
or U3126 (N_3126,N_2651,N_1584);
nand U3127 (N_3127,N_2196,N_2083);
and U3128 (N_3128,N_1448,N_1255);
nand U3129 (N_3129,N_718,N_93);
nor U3130 (N_3130,N_629,N_2027);
or U3131 (N_3131,N_810,N_2756);
nand U3132 (N_3132,N_36,N_2664);
nand U3133 (N_3133,N_2450,N_2717);
nor U3134 (N_3134,N_922,N_1736);
nor U3135 (N_3135,N_1023,N_921);
nand U3136 (N_3136,N_2051,N_909);
nand U3137 (N_3137,N_340,N_819);
or U3138 (N_3138,N_2174,N_1970);
xnor U3139 (N_3139,N_773,N_1354);
nor U3140 (N_3140,N_995,N_2612);
nand U3141 (N_3141,N_985,N_2130);
nand U3142 (N_3142,N_1461,N_285);
nor U3143 (N_3143,N_775,N_2135);
nand U3144 (N_3144,N_1477,N_474);
and U3145 (N_3145,N_2609,N_1020);
nand U3146 (N_3146,N_816,N_1443);
or U3147 (N_3147,N_1880,N_199);
and U3148 (N_3148,N_2712,N_919);
nand U3149 (N_3149,N_906,N_1174);
nor U3150 (N_3150,N_2799,N_1680);
nand U3151 (N_3151,N_1168,N_277);
and U3152 (N_3152,N_1339,N_1115);
and U3153 (N_3153,N_1019,N_2673);
or U3154 (N_3154,N_2703,N_2069);
nor U3155 (N_3155,N_750,N_2906);
or U3156 (N_3156,N_2514,N_329);
nand U3157 (N_3157,N_1991,N_297);
or U3158 (N_3158,N_2831,N_1145);
or U3159 (N_3159,N_923,N_282);
and U3160 (N_3160,N_2913,N_1088);
nand U3161 (N_3161,N_2755,N_2437);
nor U3162 (N_3162,N_1428,N_345);
nand U3163 (N_3163,N_206,N_993);
and U3164 (N_3164,N_1241,N_1504);
and U3165 (N_3165,N_2415,N_1122);
nand U3166 (N_3166,N_2495,N_143);
nand U3167 (N_3167,N_1280,N_2507);
nand U3168 (N_3168,N_2004,N_2477);
or U3169 (N_3169,N_882,N_2639);
or U3170 (N_3170,N_1730,N_1905);
nand U3171 (N_3171,N_1879,N_2052);
or U3172 (N_3172,N_1746,N_2443);
nor U3173 (N_3173,N_326,N_2422);
nand U3174 (N_3174,N_2855,N_140);
nor U3175 (N_3175,N_1541,N_2247);
or U3176 (N_3176,N_477,N_2753);
nand U3177 (N_3177,N_2654,N_2317);
nand U3178 (N_3178,N_2104,N_1636);
and U3179 (N_3179,N_1312,N_2223);
and U3180 (N_3180,N_659,N_124);
nor U3181 (N_3181,N_2728,N_2017);
or U3182 (N_3182,N_2592,N_867);
nand U3183 (N_3183,N_2999,N_2320);
or U3184 (N_3184,N_237,N_1985);
nand U3185 (N_3185,N_1641,N_358);
xor U3186 (N_3186,N_2375,N_518);
or U3187 (N_3187,N_1096,N_832);
nor U3188 (N_3188,N_2494,N_2952);
nand U3189 (N_3189,N_2412,N_447);
nor U3190 (N_3190,N_1110,N_869);
nor U3191 (N_3191,N_1745,N_394);
nand U3192 (N_3192,N_2838,N_1773);
nor U3193 (N_3193,N_615,N_2082);
nand U3194 (N_3194,N_2519,N_44);
nand U3195 (N_3195,N_2171,N_1085);
and U3196 (N_3196,N_1713,N_436);
or U3197 (N_3197,N_1892,N_1413);
and U3198 (N_3198,N_2471,N_2250);
or U3199 (N_3199,N_236,N_417);
and U3200 (N_3200,N_766,N_1979);
or U3201 (N_3201,N_2956,N_2793);
or U3202 (N_3202,N_1253,N_652);
nor U3203 (N_3203,N_796,N_1402);
or U3204 (N_3204,N_1723,N_2576);
or U3205 (N_3205,N_1415,N_815);
nand U3206 (N_3206,N_2820,N_801);
and U3207 (N_3207,N_1476,N_679);
and U3208 (N_3208,N_1240,N_732);
and U3209 (N_3209,N_1992,N_978);
nor U3210 (N_3210,N_105,N_1951);
nand U3211 (N_3211,N_1127,N_966);
nand U3212 (N_3212,N_530,N_884);
or U3213 (N_3213,N_486,N_400);
nor U3214 (N_3214,N_350,N_2784);
or U3215 (N_3215,N_1227,N_2113);
and U3216 (N_3216,N_2239,N_928);
nand U3217 (N_3217,N_2866,N_717);
nor U3218 (N_3218,N_854,N_2989);
nand U3219 (N_3219,N_1862,N_27);
or U3220 (N_3220,N_2996,N_2745);
nand U3221 (N_3221,N_211,N_472);
and U3222 (N_3222,N_2310,N_541);
nand U3223 (N_3223,N_2729,N_1798);
nand U3224 (N_3224,N_1685,N_586);
and U3225 (N_3225,N_2583,N_1931);
nor U3226 (N_3226,N_227,N_1138);
or U3227 (N_3227,N_2560,N_1380);
nand U3228 (N_3228,N_1490,N_713);
and U3229 (N_3229,N_1069,N_755);
nand U3230 (N_3230,N_2280,N_445);
nor U3231 (N_3231,N_175,N_2562);
or U3232 (N_3232,N_343,N_1961);
nand U3233 (N_3233,N_1614,N_834);
or U3234 (N_3234,N_930,N_2522);
nor U3235 (N_3235,N_458,N_2541);
or U3236 (N_3236,N_2986,N_2456);
or U3237 (N_3237,N_2199,N_1693);
and U3238 (N_3238,N_493,N_2466);
nor U3239 (N_3239,N_625,N_2710);
and U3240 (N_3240,N_1231,N_697);
and U3241 (N_3241,N_539,N_782);
nor U3242 (N_3242,N_1405,N_1692);
and U3243 (N_3243,N_542,N_2558);
or U3244 (N_3244,N_1200,N_2965);
and U3245 (N_3245,N_2304,N_2988);
and U3246 (N_3246,N_60,N_1883);
or U3247 (N_3247,N_2449,N_1747);
or U3248 (N_3248,N_552,N_2057);
or U3249 (N_3249,N_2119,N_115);
nor U3250 (N_3250,N_2365,N_1757);
and U3251 (N_3251,N_2441,N_2801);
or U3252 (N_3252,N_381,N_658);
or U3253 (N_3253,N_28,N_644);
nand U3254 (N_3254,N_341,N_2186);
and U3255 (N_3255,N_2888,N_262);
nor U3256 (N_3256,N_2532,N_2935);
nor U3257 (N_3257,N_2960,N_1234);
or U3258 (N_3258,N_2059,N_19);
nand U3259 (N_3259,N_1886,N_569);
nand U3260 (N_3260,N_2207,N_1889);
and U3261 (N_3261,N_2012,N_1086);
nor U3262 (N_3262,N_1842,N_1859);
and U3263 (N_3263,N_944,N_2297);
or U3264 (N_3264,N_2658,N_281);
or U3265 (N_3265,N_1832,N_434);
nand U3266 (N_3266,N_2676,N_1462);
and U3267 (N_3267,N_2337,N_2968);
nand U3268 (N_3268,N_1387,N_668);
nand U3269 (N_3269,N_1455,N_2887);
nor U3270 (N_3270,N_748,N_38);
nor U3271 (N_3271,N_1003,N_2764);
nand U3272 (N_3272,N_2770,N_1440);
nand U3273 (N_3273,N_2026,N_456);
nand U3274 (N_3274,N_1625,N_1806);
or U3275 (N_3275,N_690,N_550);
or U3276 (N_3276,N_557,N_1914);
nor U3277 (N_3277,N_1850,N_420);
nand U3278 (N_3278,N_1682,N_2627);
or U3279 (N_3279,N_2813,N_2889);
and U3280 (N_3280,N_2107,N_1416);
nor U3281 (N_3281,N_2021,N_2032);
nor U3282 (N_3282,N_1660,N_406);
nand U3283 (N_3283,N_176,N_591);
nor U3284 (N_3284,N_80,N_764);
nor U3285 (N_3285,N_225,N_383);
nor U3286 (N_3286,N_2355,N_1260);
or U3287 (N_3287,N_2569,N_741);
nor U3288 (N_3288,N_2931,N_767);
nor U3289 (N_3289,N_2667,N_362);
and U3290 (N_3290,N_1766,N_2752);
and U3291 (N_3291,N_259,N_2681);
nor U3292 (N_3292,N_2465,N_2068);
xnor U3293 (N_3293,N_1725,N_2732);
nand U3294 (N_3294,N_548,N_2497);
nand U3295 (N_3295,N_2553,N_354);
and U3296 (N_3296,N_676,N_1518);
or U3297 (N_3297,N_1437,N_2102);
nand U3298 (N_3298,N_809,N_2961);
xnor U3299 (N_3299,N_2255,N_2563);
or U3300 (N_3300,N_418,N_1808);
and U3301 (N_3301,N_1933,N_2932);
nand U3302 (N_3302,N_1348,N_1398);
xor U3303 (N_3303,N_2306,N_2918);
nor U3304 (N_3304,N_2598,N_941);
nor U3305 (N_3305,N_2565,N_1699);
nand U3306 (N_3306,N_2379,N_1749);
and U3307 (N_3307,N_583,N_355);
or U3308 (N_3308,N_172,N_2084);
nor U3309 (N_3309,N_1778,N_812);
nand U3310 (N_3310,N_240,N_311);
nor U3311 (N_3311,N_759,N_2435);
nand U3312 (N_3312,N_2279,N_1579);
and U3313 (N_3313,N_2679,N_1297);
nor U3314 (N_3314,N_2819,N_1025);
and U3315 (N_3315,N_1183,N_352);
or U3316 (N_3316,N_2479,N_2324);
or U3317 (N_3317,N_2396,N_1135);
nand U3318 (N_3318,N_2861,N_1681);
nor U3319 (N_3319,N_1008,N_1943);
and U3320 (N_3320,N_1018,N_2743);
nand U3321 (N_3321,N_551,N_1588);
and U3322 (N_3322,N_2603,N_2499);
nor U3323 (N_3323,N_1860,N_2001);
or U3324 (N_3324,N_2845,N_560);
nor U3325 (N_3325,N_2897,N_924);
or U3326 (N_3326,N_2318,N_1813);
or U3327 (N_3327,N_1417,N_2132);
nor U3328 (N_3328,N_2613,N_1703);
and U3329 (N_3329,N_173,N_1898);
and U3330 (N_3330,N_1270,N_2476);
or U3331 (N_3331,N_961,N_2959);
nor U3332 (N_3332,N_1539,N_646);
or U3333 (N_3333,N_200,N_846);
or U3334 (N_3334,N_1421,N_255);
or U3335 (N_3335,N_1787,N_806);
and U3336 (N_3336,N_239,N_2719);
nor U3337 (N_3337,N_1820,N_1498);
nor U3338 (N_3338,N_2393,N_1098);
and U3339 (N_3339,N_229,N_2674);
nand U3340 (N_3340,N_2886,N_2257);
and U3341 (N_3341,N_1279,N_2384);
or U3342 (N_3342,N_1281,N_1022);
nand U3343 (N_3343,N_1760,N_2075);
nand U3344 (N_3344,N_931,N_1169);
and U3345 (N_3345,N_1938,N_494);
nor U3346 (N_3346,N_130,N_324);
nor U3347 (N_3347,N_195,N_1500);
and U3348 (N_3348,N_466,N_2726);
nor U3349 (N_3349,N_1000,N_506);
or U3350 (N_3350,N_1332,N_1742);
or U3351 (N_3351,N_2475,N_2323);
or U3352 (N_3352,N_1975,N_339);
nand U3353 (N_3353,N_765,N_2909);
and U3354 (N_3354,N_2243,N_818);
and U3355 (N_3355,N_503,N_1156);
nand U3356 (N_3356,N_2418,N_2319);
nor U3357 (N_3357,N_555,N_2584);
and U3358 (N_3358,N_2036,N_887);
and U3359 (N_3359,N_1268,N_1491);
nor U3360 (N_3360,N_2636,N_2062);
nand U3361 (N_3361,N_396,N_2041);
nor U3362 (N_3362,N_1929,N_2330);
or U3363 (N_3363,N_1459,N_859);
or U3364 (N_3364,N_2709,N_144);
nor U3365 (N_3365,N_2594,N_330);
or U3366 (N_3366,N_544,N_170);
xor U3367 (N_3367,N_2749,N_2118);
and U3368 (N_3368,N_1131,N_2357);
and U3369 (N_3369,N_1894,N_1729);
nor U3370 (N_3370,N_2191,N_1229);
nor U3371 (N_3371,N_594,N_1800);
nor U3372 (N_3372,N_682,N_837);
or U3373 (N_3373,N_752,N_2166);
and U3374 (N_3374,N_1774,N_581);
or U3375 (N_3375,N_1014,N_2115);
and U3376 (N_3376,N_647,N_2721);
nand U3377 (N_3377,N_390,N_1483);
or U3378 (N_3378,N_2124,N_1343);
and U3379 (N_3379,N_2546,N_2350);
and U3380 (N_3380,N_2125,N_1410);
or U3381 (N_3381,N_556,N_320);
nor U3382 (N_3382,N_2212,N_2244);
nand U3383 (N_3383,N_929,N_1662);
and U3384 (N_3384,N_2521,N_2184);
nand U3385 (N_3385,N_2675,N_2977);
and U3386 (N_3386,N_1973,N_137);
nor U3387 (N_3387,N_1599,N_2484);
and U3388 (N_3388,N_1776,N_1221);
and U3389 (N_3389,N_2524,N_761);
or U3390 (N_3390,N_1656,N_942);
and U3391 (N_3391,N_2851,N_1154);
nor U3392 (N_3392,N_1118,N_1851);
or U3393 (N_3393,N_1206,N_2233);
nor U3394 (N_3394,N_1784,N_1566);
or U3395 (N_3395,N_2291,N_2140);
or U3396 (N_3396,N_1637,N_1338);
or U3397 (N_3397,N_1595,N_2172);
and U3398 (N_3398,N_1619,N_2329);
and U3399 (N_3399,N_90,N_899);
or U3400 (N_3400,N_824,N_1151);
and U3401 (N_3401,N_2505,N_2123);
nor U3402 (N_3402,N_813,N_2386);
and U3403 (N_3403,N_1137,N_1180);
nor U3404 (N_3404,N_1418,N_1374);
and U3405 (N_3405,N_20,N_1505);
nor U3406 (N_3406,N_2970,N_2669);
nand U3407 (N_3407,N_1853,N_45);
nand U3408 (N_3408,N_269,N_2373);
nand U3409 (N_3409,N_1921,N_2419);
and U3410 (N_3410,N_2202,N_1167);
or U3411 (N_3411,N_957,N_1564);
nor U3412 (N_3412,N_1953,N_2811);
or U3413 (N_3413,N_566,N_501);
xor U3414 (N_3414,N_1204,N_2401);
nor U3415 (N_3415,N_1647,N_18);
or U3416 (N_3416,N_2146,N_631);
and U3417 (N_3417,N_526,N_790);
or U3418 (N_3418,N_1283,N_69);
and U3419 (N_3419,N_1347,N_123);
and U3420 (N_3420,N_1422,N_2087);
and U3421 (N_3421,N_224,N_1456);
and U3422 (N_3422,N_1304,N_1865);
nor U3423 (N_3423,N_2485,N_1432);
nand U3424 (N_3424,N_2366,N_244);
and U3425 (N_3425,N_2659,N_2980);
nand U3426 (N_3426,N_1923,N_2953);
or U3427 (N_3427,N_1804,N_939);
and U3428 (N_3428,N_2067,N_645);
and U3429 (N_3429,N_1471,N_1769);
and U3430 (N_3430,N_1097,N_2705);
nand U3431 (N_3431,N_483,N_220);
nand U3432 (N_3432,N_228,N_2821);
nor U3433 (N_3433,N_222,N_1634);
nor U3434 (N_3434,N_1646,N_2597);
or U3435 (N_3435,N_700,N_1626);
nor U3436 (N_3436,N_1708,N_1399);
nand U3437 (N_3437,N_821,N_2336);
or U3438 (N_3438,N_579,N_1190);
nor U3439 (N_3439,N_2462,N_305);
nand U3440 (N_3440,N_1683,N_395);
nor U3441 (N_3441,N_962,N_1046);
and U3442 (N_3442,N_360,N_2915);
or U3443 (N_3443,N_1779,N_2641);
xnor U3444 (N_3444,N_747,N_714);
nor U3445 (N_3445,N_2704,N_1814);
or U3446 (N_3446,N_525,N_179);
and U3447 (N_3447,N_2226,N_2817);
nand U3448 (N_3448,N_1223,N_841);
and U3449 (N_3449,N_2005,N_947);
and U3450 (N_3450,N_213,N_2020);
and U3451 (N_3451,N_1246,N_2634);
nand U3452 (N_3452,N_2150,N_2814);
or U3453 (N_3453,N_2536,N_1430);
or U3454 (N_3454,N_2876,N_2734);
nand U3455 (N_3455,N_361,N_1142);
and U3456 (N_3456,N_2259,N_1763);
xnor U3457 (N_3457,N_1717,N_1084);
nand U3458 (N_3458,N_1986,N_901);
nor U3459 (N_3459,N_1802,N_877);
and U3460 (N_3460,N_408,N_2397);
and U3461 (N_3461,N_1770,N_2498);
nor U3462 (N_3462,N_2189,N_1344);
or U3463 (N_3463,N_2684,N_2545);
nor U3464 (N_3464,N_496,N_2686);
nand U3465 (N_3465,N_1288,N_2470);
and U3466 (N_3466,N_627,N_1616);
nand U3467 (N_3467,N_2929,N_2468);
or U3468 (N_3468,N_1805,N_2875);
and U3469 (N_3469,N_2106,N_1102);
or U3470 (N_3470,N_1479,N_2768);
and U3471 (N_3471,N_1365,N_1596);
and U3472 (N_3472,N_1112,N_1309);
xor U3473 (N_3473,N_925,N_142);
nor U3474 (N_3474,N_261,N_430);
nand U3475 (N_3475,N_77,N_705);
and U3476 (N_3476,N_1489,N_344);
or U3477 (N_3477,N_1968,N_1352);
nand U3478 (N_3478,N_1574,N_1205);
and U3479 (N_3479,N_2376,N_116);
nand U3480 (N_3480,N_2902,N_2582);
nor U3481 (N_3481,N_2618,N_1108);
or U3482 (N_3482,N_1694,N_154);
nor U3483 (N_3483,N_2905,N_848);
nand U3484 (N_3484,N_427,N_2794);
and U3485 (N_3485,N_953,N_890);
or U3486 (N_3486,N_450,N_2249);
or U3487 (N_3487,N_1932,N_2264);
nor U3488 (N_3488,N_1589,N_1907);
xnor U3489 (N_3489,N_1126,N_977);
nor U3490 (N_3490,N_2503,N_975);
xnor U3491 (N_3491,N_491,N_711);
nand U3492 (N_3492,N_1158,N_2587);
nor U3493 (N_3493,N_271,N_588);
or U3494 (N_3494,N_2370,N_117);
and U3495 (N_3495,N_2911,N_1409);
nand U3496 (N_3496,N_904,N_2155);
or U3497 (N_3497,N_2187,N_2637);
nand U3498 (N_3498,N_2478,N_2358);
nand U3499 (N_3499,N_865,N_1395);
nor U3500 (N_3500,N_2387,N_1882);
and U3501 (N_3501,N_1501,N_777);
and U3502 (N_3502,N_443,N_684);
nor U3503 (N_3503,N_2615,N_2551);
nand U3504 (N_3504,N_2241,N_1727);
or U3505 (N_3505,N_1495,N_1065);
and U3506 (N_3506,N_2850,N_1355);
nor U3507 (N_3507,N_1117,N_1600);
or U3508 (N_3508,N_1195,N_1606);
and U3509 (N_3509,N_798,N_986);
or U3510 (N_3510,N_2938,N_636);
nor U3511 (N_3511,N_270,N_580);
or U3512 (N_3512,N_2779,N_470);
or U3513 (N_3513,N_2735,N_246);
and U3514 (N_3514,N_2480,N_2413);
nor U3515 (N_3515,N_2327,N_1502);
nand U3516 (N_3516,N_2269,N_523);
and U3517 (N_3517,N_2837,N_1576);
and U3518 (N_3518,N_1711,N_204);
nor U3519 (N_3519,N_2808,N_1215);
or U3520 (N_3520,N_40,N_342);
nor U3521 (N_3521,N_2473,N_879);
or U3522 (N_3522,N_1678,N_1330);
nand U3523 (N_3523,N_2571,N_316);
nand U3524 (N_3524,N_2954,N_1060);
xor U3525 (N_3525,N_1176,N_499);
and U3526 (N_3526,N_1076,N_2823);
nand U3527 (N_3527,N_637,N_102);
nand U3528 (N_3528,N_2985,N_161);
nor U3529 (N_3529,N_2265,N_1264);
or U3530 (N_3530,N_446,N_1219);
and U3531 (N_3531,N_1189,N_2321);
nand U3532 (N_3532,N_1627,N_2701);
nor U3533 (N_3533,N_58,N_468);
nor U3534 (N_3534,N_231,N_2844);
nor U3535 (N_3535,N_2882,N_666);
or U3536 (N_3536,N_2805,N_1562);
and U3537 (N_3537,N_2169,N_2198);
nand U3538 (N_3538,N_1277,N_254);
nand U3539 (N_3539,N_1857,N_1591);
or U3540 (N_3540,N_1527,N_2871);
or U3541 (N_3541,N_1435,N_2029);
nand U3542 (N_3542,N_1967,N_1058);
or U3543 (N_3543,N_1055,N_1013);
or U3544 (N_3544,N_174,N_242);
and U3545 (N_3545,N_914,N_171);
nor U3546 (N_3546,N_363,N_1331);
nor U3547 (N_3547,N_1101,N_2500);
nor U3548 (N_3548,N_2235,N_1833);
and U3549 (N_3549,N_1400,N_565);
nand U3550 (N_3550,N_1450,N_1179);
nand U3551 (N_3551,N_2872,N_1296);
nor U3552 (N_3552,N_731,N_1593);
nand U3553 (N_3553,N_998,N_2767);
nand U3554 (N_3554,N_1538,N_710);
or U3555 (N_3555,N_1578,N_612);
nand U3556 (N_3556,N_1244,N_2141);
and U3557 (N_3557,N_2227,N_2190);
and U3558 (N_3558,N_2042,N_287);
nor U3559 (N_3559,N_1753,N_1827);
or U3560 (N_3560,N_1999,N_426);
nor U3561 (N_3561,N_1377,N_379);
or U3562 (N_3562,N_78,N_2835);
or U3563 (N_3563,N_233,N_2526);
nand U3564 (N_3564,N_521,N_43);
or U3565 (N_3565,N_1235,N_2007);
or U3566 (N_3566,N_2780,N_842);
nand U3567 (N_3567,N_1198,N_2620);
nand U3568 (N_3568,N_2486,N_2818);
nor U3569 (N_3569,N_720,N_725);
and U3570 (N_3570,N_1092,N_1216);
or U3571 (N_3571,N_181,N_597);
nor U3572 (N_3572,N_1393,N_951);
or U3573 (N_3573,N_2604,N_2188);
or U3574 (N_3574,N_1768,N_1737);
nand U3575 (N_3575,N_2816,N_399);
nor U3576 (N_3576,N_1981,N_2725);
nand U3577 (N_3577,N_2275,N_2847);
and U3578 (N_3578,N_371,N_260);
xor U3579 (N_3579,N_943,N_2848);
nor U3580 (N_3580,N_1972,N_2461);
or U3581 (N_3581,N_454,N_2213);
nand U3582 (N_3582,N_2665,N_1545);
or U3583 (N_3583,N_1006,N_2783);
and U3584 (N_3584,N_276,N_110);
and U3585 (N_3585,N_392,N_2955);
and U3586 (N_3586,N_31,N_1664);
nor U3587 (N_3587,N_2788,N_2660);
nand U3588 (N_3588,N_1622,N_2775);
and U3589 (N_3589,N_152,N_564);
or U3590 (N_3590,N_431,N_1962);
and U3591 (N_3591,N_2289,N_207);
and U3592 (N_3592,N_41,N_54);
and U3593 (N_3593,N_2707,N_1441);
or U3594 (N_3594,N_742,N_1696);
nor U3595 (N_3595,N_2997,N_150);
and U3596 (N_3596,N_562,N_1266);
nor U3597 (N_3597,N_415,N_2900);
nor U3598 (N_3598,N_2543,N_1881);
nor U3599 (N_3599,N_2930,N_670);
nand U3600 (N_3600,N_2237,N_527);
nor U3601 (N_3601,N_2746,N_1359);
nor U3602 (N_3602,N_299,N_695);
nor U3603 (N_3603,N_1944,N_2722);
or U3604 (N_3604,N_1426,N_2574);
nor U3605 (N_3605,N_2713,N_1533);
nor U3606 (N_3606,N_1555,N_441);
and U3607 (N_3607,N_1320,N_656);
xor U3608 (N_3608,N_2378,N_1577);
xnor U3609 (N_3609,N_1040,N_2969);
nand U3610 (N_3610,N_2180,N_440);
and U3611 (N_3611,N_423,N_490);
or U3612 (N_3612,N_484,N_1775);
nor U3613 (N_3613,N_2353,N_2408);
nand U3614 (N_3614,N_2683,N_2152);
and U3615 (N_3615,N_151,N_582);
or U3616 (N_3616,N_1444,N_2447);
or U3617 (N_3617,N_554,N_1299);
or U3618 (N_3618,N_1335,N_1655);
nor U3619 (N_3619,N_2607,N_2151);
nor U3620 (N_3620,N_760,N_784);
or U3621 (N_3621,N_64,N_1830);
nand U3622 (N_3622,N_2631,N_1648);
or U3623 (N_3623,N_85,N_2078);
nor U3624 (N_3624,N_467,N_1408);
nor U3625 (N_3625,N_602,N_1278);
nand U3626 (N_3626,N_1741,N_208);
nor U3627 (N_3627,N_232,N_2296);
or U3628 (N_3628,N_2539,N_2841);
and U3629 (N_3629,N_2940,N_1718);
nand U3630 (N_3630,N_2696,N_2910);
or U3631 (N_3631,N_2281,N_852);
nor U3632 (N_3632,N_1630,N_1217);
xnor U3633 (N_3633,N_952,N_1559);
xor U3634 (N_3634,N_258,N_2635);
nor U3635 (N_3635,N_1446,N_643);
nand U3636 (N_3636,N_2129,N_507);
nand U3637 (N_3637,N_678,N_2699);
nor U3638 (N_3638,N_896,N_2110);
or U3639 (N_3639,N_1199,N_2773);
and U3640 (N_3640,N_2697,N_1050);
and U3641 (N_3641,N_187,N_2185);
nor U3642 (N_3642,N_2272,N_1601);
or U3643 (N_3643,N_1751,N_2436);
or U3644 (N_3644,N_13,N_21);
or U3645 (N_3645,N_1568,N_1071);
nor U3646 (N_3646,N_621,N_2072);
nor U3647 (N_3647,N_2292,N_2846);
or U3648 (N_3648,N_639,N_2810);
and U3649 (N_3649,N_348,N_2738);
nand U3650 (N_3650,N_76,N_2139);
nand U3651 (N_3651,N_1353,N_1392);
or U3652 (N_3652,N_164,N_2984);
nand U3653 (N_3653,N_688,N_1783);
nand U3654 (N_3654,N_2013,N_111);
xor U3655 (N_3655,N_2944,N_2839);
nand U3656 (N_3656,N_2216,N_39);
and U3657 (N_3657,N_1243,N_444);
and U3658 (N_3658,N_2286,N_779);
nand U3659 (N_3659,N_531,N_1653);
and U3660 (N_3660,N_217,N_407);
and U3661 (N_3661,N_571,N_1258);
and U3662 (N_3662,N_2804,N_817);
nor U3663 (N_3663,N_2116,N_1212);
or U3664 (N_3664,N_1554,N_1866);
and U3665 (N_3665,N_910,N_337);
or U3666 (N_3666,N_1350,N_1150);
and U3667 (N_3667,N_1192,N_2464);
nor U3668 (N_3668,N_1275,N_1042);
or U3669 (N_3669,N_2400,N_1317);
nand U3670 (N_3670,N_1836,N_382);
nand U3671 (N_3671,N_1363,N_1074);
or U3672 (N_3672,N_1116,N_1079);
nand U3673 (N_3673,N_524,N_856);
and U3674 (N_3674,N_1997,N_2070);
nor U3675 (N_3675,N_1412,N_1230);
xnor U3676 (N_3676,N_1303,N_2548);
nor U3677 (N_3677,N_2702,N_72);
nand U3678 (N_3678,N_2050,N_1702);
and U3679 (N_3679,N_2715,N_438);
and U3680 (N_3680,N_2778,N_675);
xor U3681 (N_3681,N_203,N_2008);
or U3682 (N_3682,N_1984,N_2388);
and U3683 (N_3683,N_1287,N_2504);
nand U3684 (N_3684,N_1295,N_128);
nor U3685 (N_3685,N_719,N_2809);
or U3686 (N_3686,N_479,N_307);
nor U3687 (N_3687,N_2383,N_1994);
xnor U3688 (N_3688,N_1926,N_2867);
or U3689 (N_3689,N_1308,N_2142);
or U3690 (N_3690,N_1575,N_2638);
and U3691 (N_3691,N_2802,N_849);
xor U3692 (N_3692,N_42,N_10);
nor U3693 (N_3693,N_1870,N_1439);
nor U3694 (N_3694,N_2170,N_2972);
or U3695 (N_3695,N_1872,N_938);
or U3696 (N_3696,N_517,N_22);
nor U3697 (N_3697,N_1937,N_1856);
nand U3698 (N_3698,N_1404,N_1759);
nor U3699 (N_3699,N_2951,N_972);
or U3700 (N_3700,N_937,N_915);
or U3701 (N_3701,N_903,N_788);
nand U3702 (N_3702,N_2994,N_265);
or U3703 (N_3703,N_475,N_540);
and U3704 (N_3704,N_322,N_1996);
or U3705 (N_3705,N_17,N_2097);
and U3706 (N_3706,N_1147,N_1721);
or U3707 (N_3707,N_2824,N_131);
and U3708 (N_3708,N_2421,N_1608);
nand U3709 (N_3709,N_894,N_592);
and U3710 (N_3710,N_2209,N_963);
or U3711 (N_3711,N_1059,N_99);
or U3712 (N_3712,N_1781,N_2164);
nand U3713 (N_3713,N_2621,N_452);
nor U3714 (N_3714,N_874,N_1722);
or U3715 (N_3715,N_205,N_2833);
nor U3716 (N_3716,N_981,N_613);
nand U3717 (N_3717,N_437,N_1534);
nor U3718 (N_3718,N_2126,N_1224);
and U3719 (N_3719,N_1376,N_2936);
or U3720 (N_3720,N_1561,N_2081);
and U3721 (N_3721,N_2195,N_397);
and U3722 (N_3722,N_2547,N_2939);
nand U3723 (N_3723,N_2739,N_1475);
and U3724 (N_3724,N_638,N_1166);
nand U3725 (N_3725,N_886,N_2407);
nand U3726 (N_3726,N_701,N_1613);
nand U3727 (N_3727,N_247,N_984);
and U3728 (N_3728,N_2744,N_1823);
nor U3729 (N_3729,N_2459,N_1269);
and U3730 (N_3730,N_2640,N_2555);
or U3731 (N_3731,N_1910,N_1397);
xnor U3732 (N_3732,N_651,N_413);
or U3733 (N_3733,N_2276,N_724);
nand U3734 (N_3734,N_2175,N_2258);
and U3735 (N_3735,N_2274,N_57);
or U3736 (N_3736,N_1799,N_567);
and U3737 (N_3737,N_1438,N_332);
and U3738 (N_3738,N_2593,N_268);
nor U3739 (N_3739,N_2065,N_2998);
nand U3740 (N_3740,N_858,N_1043);
or U3741 (N_3741,N_2176,N_2857);
or U3742 (N_3742,N_1005,N_2245);
or U3743 (N_3743,N_1739,N_433);
nand U3744 (N_3744,N_2978,N_1165);
nor U3745 (N_3745,N_1184,N_1334);
nand U3746 (N_3746,N_1103,N_2742);
nor U3747 (N_3747,N_1752,N_686);
nor U3748 (N_3748,N_2035,N_672);
and U3749 (N_3749,N_1885,N_1928);
or U3750 (N_3750,N_2894,N_1838);
and U3751 (N_3751,N_1496,N_1407);
or U3752 (N_3752,N_664,N_235);
xor U3753 (N_3753,N_1871,N_1191);
nor U3754 (N_3754,N_1367,N_1011);
or U3755 (N_3755,N_572,N_1663);
or U3756 (N_3756,N_1091,N_634);
and U3757 (N_3757,N_1302,N_847);
nor U3758 (N_3758,N_1897,N_109);
nor U3759 (N_3759,N_1843,N_1669);
nand U3760 (N_3760,N_2220,N_318);
nor U3761 (N_3761,N_2619,N_2520);
nand U3762 (N_3762,N_1811,N_2644);
nand U3763 (N_3763,N_1027,N_1794);
xnor U3764 (N_3764,N_2305,N_1329);
nand U3765 (N_3765,N_146,N_288);
nor U3766 (N_3766,N_2363,N_1492);
nand U3767 (N_3767,N_662,N_2356);
nor U3768 (N_3768,N_2828,N_2409);
and U3769 (N_3769,N_1451,N_822);
nand U3770 (N_3770,N_2018,N_457);
nand U3771 (N_3771,N_1969,N_2463);
or U3772 (N_3772,N_1958,N_1712);
or U3773 (N_3773,N_1639,N_263);
xnor U3774 (N_3774,N_2852,N_296);
nor U3775 (N_3775,N_1623,N_2351);
nand U3776 (N_3776,N_888,N_1345);
or U3777 (N_3777,N_306,N_1083);
and U3778 (N_3778,N_1487,N_1316);
nand U3779 (N_3779,N_25,N_485);
and U3780 (N_3780,N_2643,N_2076);
nor U3781 (N_3781,N_398,N_376);
nand U3782 (N_3782,N_2016,N_2099);
or U3783 (N_3783,N_190,N_1181);
nor U3784 (N_3784,N_1754,N_2723);
nor U3785 (N_3785,N_113,N_1272);
and U3786 (N_3786,N_1672,N_52);
nand U3787 (N_3787,N_1313,N_696);
and U3788 (N_3788,N_156,N_2633);
nand U3789 (N_3789,N_1378,N_1732);
and U3790 (N_3790,N_1549,N_2114);
nor U3791 (N_3791,N_2933,N_606);
or U3792 (N_3792,N_2137,N_1196);
or U3793 (N_3793,N_2385,N_65);
nand U3794 (N_3794,N_1136,N_2577);
or U3795 (N_3795,N_2995,N_34);
or U3796 (N_3796,N_1532,N_2322);
nor U3797 (N_3797,N_1858,N_694);
nand U3798 (N_3798,N_954,N_2089);
and U3799 (N_3799,N_932,N_1835);
and U3800 (N_3800,N_279,N_1077);
or U3801 (N_3801,N_2979,N_2399);
or U3802 (N_3802,N_1093,N_1988);
or U3803 (N_3803,N_1900,N_119);
nand U3804 (N_3804,N_1323,N_378);
or U3805 (N_3805,N_545,N_1878);
or U3806 (N_3806,N_55,N_661);
nor U3807 (N_3807,N_35,N_1520);
and U3808 (N_3808,N_2096,N_2653);
and U3809 (N_3809,N_1594,N_1815);
and U3810 (N_3810,N_2,N_1731);
xnor U3811 (N_3811,N_2518,N_449);
or U3812 (N_3812,N_2748,N_912);
nor U3813 (N_3813,N_514,N_1689);
nand U3814 (N_3814,N_2045,N_2891);
nor U3815 (N_3815,N_2925,N_753);
and U3816 (N_3816,N_480,N_1743);
nor U3817 (N_3817,N_1016,N_14);
and U3818 (N_3818,N_66,N_1822);
xnor U3819 (N_3819,N_735,N_657);
nor U3820 (N_3820,N_2481,N_2865);
and U3821 (N_3821,N_1740,N_1916);
and U3822 (N_3822,N_488,N_380);
and U3823 (N_3823,N_1797,N_1346);
and U3824 (N_3824,N_1259,N_838);
or U3825 (N_3825,N_1010,N_2080);
nor U3826 (N_3826,N_1553,N_1955);
nor U3827 (N_3827,N_249,N_476);
nor U3828 (N_3828,N_771,N_1791);
or U3829 (N_3829,N_1173,N_2361);
nor U3830 (N_3830,N_68,N_1542);
or U3831 (N_3831,N_1481,N_346);
and U3832 (N_3832,N_2203,N_463);
and U3833 (N_3833,N_2856,N_570);
nand U3834 (N_3834,N_607,N_2508);
nand U3835 (N_3835,N_1582,N_1659);
or U3836 (N_3836,N_2411,N_870);
nand U3837 (N_3837,N_1638,N_2590);
and U3838 (N_3838,N_797,N_620);
or U3839 (N_3839,N_2253,N_1528);
nor U3840 (N_3840,N_192,N_1256);
or U3841 (N_3841,N_1139,N_1433);
and U3842 (N_3842,N_2611,N_2650);
nand U3843 (N_3843,N_1445,N_827);
and U3844 (N_3844,N_2371,N_2825);
and U3845 (N_3845,N_2687,N_1980);
or U3846 (N_3846,N_1846,N_2566);
or U3847 (N_3847,N_1113,N_83);
nor U3848 (N_3848,N_2215,N_1194);
nand U3849 (N_3849,N_875,N_734);
and U3850 (N_3850,N_2942,N_241);
or U3851 (N_3851,N_1704,N_1667);
nand U3852 (N_3852,N_687,N_603);
or U3853 (N_3853,N_2284,N_63);
or U3854 (N_3854,N_1765,N_783);
nand U3855 (N_3855,N_186,N_129);
nand U3856 (N_3856,N_2885,N_744);
and U3857 (N_3857,N_62,N_1826);
xnor U3858 (N_3858,N_1821,N_2428);
or U3859 (N_3859,N_422,N_1114);
or U3860 (N_3860,N_1855,N_1271);
and U3861 (N_3861,N_1133,N_74);
nor U3862 (N_3862,N_2714,N_2807);
nand U3863 (N_3863,N_495,N_2525);
and U3864 (N_3864,N_289,N_2883);
nor U3865 (N_3865,N_2754,N_2896);
and U3866 (N_3866,N_2927,N_1657);
xnor U3867 (N_3867,N_2093,N_723);
nor U3868 (N_3868,N_898,N_84);
nand U3869 (N_3869,N_729,N_333);
xor U3870 (N_3870,N_2055,N_1987);
or U3871 (N_3871,N_148,N_2348);
or U3872 (N_3872,N_2605,N_2670);
or U3873 (N_3873,N_964,N_1379);
and U3874 (N_3874,N_1051,N_1552);
nand U3875 (N_3875,N_1170,N_2785);
nor U3876 (N_3876,N_2843,N_1120);
or U3877 (N_3877,N_641,N_2431);
and U3878 (N_3878,N_1057,N_1563);
nand U3879 (N_3879,N_585,N_2109);
nand U3880 (N_3880,N_1550,N_215);
nor U3881 (N_3881,N_2975,N_2091);
and U3882 (N_3882,N_1458,N_2916);
or U3883 (N_3883,N_2086,N_1104);
or U3884 (N_3884,N_2800,N_1884);
nor U3885 (N_3885,N_1888,N_1469);
nand U3886 (N_3886,N_302,N_2368);
nor U3887 (N_3887,N_1790,N_2006);
nand U3888 (N_3888,N_1673,N_2806);
nor U3889 (N_3889,N_201,N_2389);
and U3890 (N_3890,N_803,N_2120);
nand U3891 (N_3891,N_1052,N_1915);
nand U3892 (N_3892,N_2622,N_1854);
and U3893 (N_3893,N_2832,N_2864);
nand U3894 (N_3894,N_2685,N_2433);
and U3895 (N_3895,N_1473,N_1072);
and U3896 (N_3896,N_610,N_2840);
or U3897 (N_3897,N_2493,N_1922);
or U3898 (N_3898,N_464,N_626);
nor U3899 (N_3899,N_1649,N_1971);
or U3900 (N_3900,N_2787,N_290);
or U3901 (N_3901,N_2299,N_1381);
and U3902 (N_3902,N_469,N_515);
xor U3903 (N_3903,N_1285,N_478);
or U3904 (N_3904,N_1570,N_1581);
nand U3905 (N_3905,N_2453,N_194);
and U3906 (N_3906,N_1089,N_2792);
nor U3907 (N_3907,N_1153,N_2095);
nor U3908 (N_3908,N_1701,N_1220);
and U3909 (N_3909,N_1161,N_33);
or U3910 (N_3910,N_2472,N_2432);
nand U3911 (N_3911,N_502,N_347);
or U3912 (N_3912,N_691,N_1061);
nor U3913 (N_3913,N_251,N_1391);
xor U3914 (N_3914,N_2947,N_648);
nor U3915 (N_3915,N_1758,N_1130);
nand U3916 (N_3916,N_2053,N_2448);
xor U3917 (N_3917,N_1252,N_71);
or U3918 (N_3918,N_739,N_1087);
nor U3919 (N_3919,N_1282,N_671);
or U3920 (N_3920,N_1066,N_2127);
nor U3921 (N_3921,N_2617,N_863);
nor U3922 (N_3922,N_2757,N_2899);
nand U3923 (N_3923,N_2706,N_1690);
nand U3924 (N_3924,N_338,N_1454);
and U3925 (N_3925,N_2103,N_1803);
or U3926 (N_3926,N_1571,N_1478);
nor U3927 (N_3927,N_926,N_23);
nor U3928 (N_3928,N_1525,N_2430);
and U3929 (N_3929,N_2666,N_1090);
and U3930 (N_3930,N_1100,N_935);
xnor U3931 (N_3931,N_1795,N_1427);
xnor U3932 (N_3932,N_1670,N_1201);
or U3933 (N_3933,N_1580,N_2283);
nand U3934 (N_3934,N_820,N_2066);
and U3935 (N_3935,N_2219,N_1128);
or U3936 (N_3936,N_598,N_1232);
nor U3937 (N_3937,N_1917,N_2672);
nand U3938 (N_3938,N_933,N_2402);
and U3939 (N_3939,N_508,N_653);
and U3940 (N_3940,N_2307,N_2315);
nand U3941 (N_3941,N_461,N_2829);
and U3942 (N_3942,N_1848,N_389);
nand U3943 (N_3943,N_300,N_2973);
or U3944 (N_3944,N_2517,N_2204);
nor U3945 (N_3945,N_1514,N_987);
nor U3946 (N_3946,N_1004,N_2655);
nor U3947 (N_3947,N_745,N_2214);
nand U3948 (N_3948,N_1119,N_1261);
nor U3949 (N_3949,N_622,N_2596);
nand U3950 (N_3950,N_1809,N_2108);
or U3951 (N_3951,N_2585,N_1144);
nand U3952 (N_3952,N_1474,N_628);
or U3953 (N_3953,N_1431,N_1152);
nand U3954 (N_3954,N_979,N_1155);
or U3955 (N_3955,N_1300,N_2781);
nand U3956 (N_3956,N_2599,N_487);
or U3957 (N_3957,N_59,N_2533);
nor U3958 (N_3958,N_1551,N_138);
nor U3959 (N_3959,N_1524,N_1592);
xor U3960 (N_3960,N_1590,N_1511);
nand U3961 (N_3961,N_1,N_2331);
nand U3962 (N_3962,N_1314,N_321);
nor U3963 (N_3963,N_1315,N_2157);
or U3964 (N_3964,N_1203,N_2711);
nand U3965 (N_3965,N_2455,N_955);
nor U3966 (N_3966,N_2879,N_2589);
and U3967 (N_3967,N_2903,N_1075);
nor U3968 (N_3968,N_2708,N_2287);
nor U3969 (N_3969,N_2758,N_1420);
nor U3970 (N_3970,N_2534,N_2308);
nand U3971 (N_3971,N_743,N_1290);
nor U3972 (N_3972,N_1688,N_835);
or U3973 (N_3973,N_364,N_1182);
nor U3974 (N_3974,N_844,N_2554);
and U3975 (N_3975,N_836,N_1604);
and U3976 (N_3976,N_1810,N_2343);
xor U3977 (N_3977,N_2009,N_1306);
nor U3978 (N_3978,N_2085,N_1911);
xor U3979 (N_3979,N_1328,N_1436);
or U3980 (N_3980,N_2210,N_2544);
nor U3981 (N_3981,N_2529,N_2424);
or U3982 (N_3982,N_1293,N_1109);
nand U3983 (N_3983,N_500,N_2268);
or U3984 (N_3984,N_609,N_1733);
nor U3985 (N_3985,N_1499,N_2868);
and U3986 (N_3986,N_1209,N_2616);
and U3987 (N_3987,N_970,N_2762);
nand U3988 (N_3988,N_1159,N_973);
nor U3989 (N_3989,N_2798,N_1977);
and U3990 (N_3990,N_1106,N_210);
nand U3991 (N_3991,N_1372,N_1319);
or U3992 (N_3992,N_2601,N_2535);
nand U3993 (N_3993,N_1948,N_1485);
or U3994 (N_3994,N_404,N_214);
and U3995 (N_3995,N_2300,N_2260);
nor U3996 (N_3996,N_726,N_278);
and U3997 (N_3997,N_1056,N_86);
nor U3998 (N_3998,N_309,N_768);
nand U3999 (N_3999,N_529,N_2335);
or U4000 (N_4000,N_2312,N_1044);
and U4001 (N_4001,N_1652,N_248);
and U4002 (N_4002,N_2691,N_2294);
nand U4003 (N_4003,N_1401,N_1442);
nor U4004 (N_4004,N_2231,N_1357);
and U4005 (N_4005,N_1724,N_1383);
or U4006 (N_4006,N_2311,N_1073);
nand U4007 (N_4007,N_900,N_2815);
nor U4008 (N_4008,N_178,N_2094);
nor U4009 (N_4009,N_2218,N_2971);
nor U4010 (N_4010,N_2789,N_2156);
nor U4011 (N_4011,N_1537,N_1047);
xnor U4012 (N_4012,N_721,N_945);
nand U4013 (N_4013,N_1516,N_2786);
nand U4014 (N_4014,N_291,N_2487);
and U4015 (N_4015,N_274,N_703);
nand U4016 (N_4016,N_2211,N_1728);
nand U4017 (N_4017,N_292,N_2588);
nor U4018 (N_4018,N_1336,N_2740);
xnor U4019 (N_4019,N_2614,N_1094);
or U4020 (N_4020,N_2987,N_1111);
or U4021 (N_4021,N_916,N_1033);
nand U4022 (N_4022,N_1460,N_2884);
or U4023 (N_4023,N_800,N_2842);
nor U4024 (N_4024,N_1547,N_1844);
or U4025 (N_4025,N_2438,N_2024);
nand U4026 (N_4026,N_2880,N_2372);
nand U4027 (N_4027,N_95,N_79);
nand U4028 (N_4028,N_948,N_1573);
nand U4029 (N_4029,N_221,N_1503);
nor U4030 (N_4030,N_120,N_432);
nand U4031 (N_4031,N_2063,N_673);
nor U4032 (N_4032,N_336,N_2677);
nand U4033 (N_4033,N_2288,N_2325);
or U4034 (N_4034,N_2147,N_845);
nor U4035 (N_4035,N_1002,N_577);
nand U4036 (N_4036,N_1236,N_2425);
nor U4037 (N_4037,N_839,N_2642);
nor U4038 (N_4038,N_1877,N_1535);
nor U4039 (N_4039,N_2168,N_2347);
nand U4040 (N_4040,N_2626,N_1565);
or U4041 (N_4041,N_2074,N_642);
nor U4042 (N_4042,N_2736,N_2181);
nand U4043 (N_4043,N_2488,N_29);
or U4044 (N_4044,N_283,N_2957);
or U4045 (N_4045,N_428,N_47);
or U4046 (N_4046,N_122,N_1318);
xor U4047 (N_4047,N_1370,N_751);
or U4048 (N_4048,N_1508,N_1558);
xor U4049 (N_4049,N_2092,N_587);
nor U4050 (N_4050,N_2277,N_2333);
or U4051 (N_4051,N_2564,N_2949);
or U4052 (N_4052,N_50,N_67);
nor U4053 (N_4053,N_1640,N_965);
and U4054 (N_4054,N_1767,N_2530);
or U4055 (N_4055,N_127,N_1772);
and U4056 (N_4056,N_2309,N_1949);
nand U4057 (N_4057,N_2192,N_1267);
or U4058 (N_4058,N_763,N_2966);
or U4059 (N_4059,N_2238,N_1394);
nand U4060 (N_4060,N_2440,N_596);
nand U4061 (N_4061,N_2967,N_619);
nor U4062 (N_4062,N_12,N_1598);
or U4063 (N_4063,N_1735,N_2452);
nor U4064 (N_4064,N_2454,N_325);
or U4065 (N_4065,N_136,N_1629);
and U4066 (N_4066,N_563,N_1543);
or U4067 (N_4067,N_412,N_2962);
nor U4068 (N_4068,N_749,N_618);
xnor U4069 (N_4069,N_1817,N_264);
nand U4070 (N_4070,N_737,N_2145);
and U4071 (N_4071,N_1661,N_125);
nand U4072 (N_4072,N_2870,N_2720);
xor U4073 (N_4073,N_1536,N_2334);
nor U4074 (N_4074,N_1896,N_2039);
or U4075 (N_4075,N_528,N_1612);
nor U4076 (N_4076,N_1163,N_2133);
nor U4077 (N_4077,N_2625,N_2165);
or U4078 (N_4078,N_2248,N_851);
and U4079 (N_4079,N_1602,N_1124);
nor U4080 (N_4080,N_702,N_2434);
and U4081 (N_4081,N_368,N_372);
or U4082 (N_4082,N_2632,N_1493);
and U4083 (N_4083,N_196,N_387);
nor U4084 (N_4084,N_1251,N_1311);
nand U4085 (N_4085,N_2282,N_112);
or U4086 (N_4086,N_2344,N_2557);
or U4087 (N_4087,N_787,N_2567);
nor U4088 (N_4088,N_1867,N_1700);
or U4089 (N_4089,N_81,N_2580);
or U4090 (N_4090,N_2490,N_2261);
and U4091 (N_4091,N_936,N_2763);
nand U4092 (N_4092,N_1609,N_2230);
and U4093 (N_4093,N_1037,N_537);
and U4094 (N_4094,N_1632,N_1946);
and U4095 (N_4095,N_2457,N_1710);
nor U4096 (N_4096,N_831,N_2056);
xnor U4097 (N_4097,N_2197,N_1007);
and U4098 (N_4098,N_1029,N_2759);
nand U4099 (N_4099,N_308,N_1294);
or U4100 (N_4100,N_1366,N_733);
or U4101 (N_4101,N_419,N_1895);
nand U4102 (N_4102,N_543,N_1466);
nor U4103 (N_4103,N_990,N_409);
nand U4104 (N_4104,N_1924,N_1793);
nand U4105 (N_4105,N_2941,N_2100);
and U4106 (N_4106,N_786,N_2692);
xor U4107 (N_4107,N_2730,N_1633);
nand U4108 (N_4108,N_5,N_473);
and U4109 (N_4109,N_974,N_1132);
or U4110 (N_4110,N_2071,N_2167);
nor U4111 (N_4111,N_2934,N_2943);
and U4112 (N_4112,N_1978,N_391);
nor U4113 (N_4113,N_1425,N_1512);
nor U4114 (N_4114,N_940,N_2578);
nor U4115 (N_4115,N_92,N_1572);
and U4116 (N_4116,N_2326,N_410);
nor U4117 (N_4117,N_992,N_1966);
and U4118 (N_4118,N_1406,N_2628);
or U4119 (N_4119,N_2090,N_2863);
nand U4120 (N_4120,N_1995,N_1337);
nor U4121 (N_4121,N_758,N_1864);
or U4122 (N_4122,N_2610,N_1925);
nand U4123 (N_4123,N_498,N_1371);
nor U4124 (N_4124,N_1515,N_2890);
or U4125 (N_4125,N_1868,N_762);
or U4126 (N_4126,N_1720,N_1918);
and U4127 (N_4127,N_1250,N_535);
or U4128 (N_4128,N_1841,N_7);
or U4129 (N_4129,N_2229,N_245);
nor U4130 (N_4130,N_2073,N_781);
or U4131 (N_4131,N_2153,N_2149);
nand U4132 (N_4132,N_2060,N_1284);
and U4133 (N_4133,N_2591,N_2624);
or U4134 (N_4134,N_575,N_334);
and U4135 (N_4135,N_1654,N_1567);
and U4136 (N_4136,N_2414,N_1876);
or U4137 (N_4137,N_2992,N_1674);
and U4138 (N_4138,N_1063,N_2346);
nor U4139 (N_4139,N_891,N_1009);
and U4140 (N_4140,N_826,N_2922);
nor U4141 (N_4141,N_2537,N_356);
nand U4142 (N_4142,N_2313,N_2406);
nand U4143 (N_4143,N_2853,N_91);
or U4144 (N_4144,N_1762,N_1172);
and U4145 (N_4145,N_2410,N_2830);
nor U4146 (N_4146,N_1544,N_2527);
nor U4147 (N_4147,N_868,N_106);
or U4148 (N_4148,N_2011,N_1960);
nand U4149 (N_4149,N_785,N_1322);
nor U4150 (N_4150,N_600,N_1818);
xor U4151 (N_4151,N_3,N_1675);
nand U4152 (N_4152,N_147,N_1587);
nand U4153 (N_4153,N_1356,N_2179);
or U4154 (N_4154,N_1771,N_1207);
nor U4155 (N_4155,N_2043,N_1327);
or U4156 (N_4156,N_2079,N_1146);
or U4157 (N_4157,N_1164,N_559);
and U4158 (N_4158,N_2836,N_1024);
and U4159 (N_4159,N_1129,N_669);
or U4160 (N_4160,N_198,N_2540);
nor U4161 (N_4161,N_2912,N_830);
nor U4162 (N_4162,N_927,N_385);
nand U4163 (N_4163,N_275,N_2228);
nor U4164 (N_4164,N_1388,N_2777);
or U4165 (N_4165,N_795,N_2162);
or U4166 (N_4166,N_1839,N_273);
nor U4167 (N_4167,N_2561,N_649);
nand U4168 (N_4168,N_605,N_1411);
and U4169 (N_4169,N_1829,N_1665);
or U4170 (N_4170,N_1540,N_864);
or U4171 (N_4171,N_883,N_1939);
nor U4172 (N_4172,N_243,N_1064);
or U4173 (N_4173,N_497,N_1942);
or U4174 (N_4174,N_335,N_2182);
nand U4175 (N_4175,N_1874,N_197);
nor U4176 (N_4176,N_2919,N_533);
nand U4177 (N_4177,N_462,N_740);
nand U4178 (N_4178,N_2608,N_315);
nand U4179 (N_4179,N_640,N_590);
or U4180 (N_4180,N_2769,N_331);
or U4181 (N_4181,N_1340,N_2048);
nand U4182 (N_4182,N_2208,N_2148);
or U4183 (N_4183,N_1028,N_2049);
or U4184 (N_4184,N_424,N_2200);
nor U4185 (N_4185,N_794,N_1750);
nand U4186 (N_4186,N_2881,N_2367);
nand U4187 (N_4187,N_2581,N_133);
nand U4188 (N_4188,N_2895,N_2731);
and U4189 (N_4189,N_516,N_1472);
and U4190 (N_4190,N_2240,N_2143);
or U4191 (N_4191,N_401,N_2030);
and U4192 (N_4192,N_2469,N_374);
nand U4193 (N_4193,N_1382,N_1697);
nand U4194 (N_4194,N_971,N_632);
and U4195 (N_4195,N_1403,N_2034);
nand U4196 (N_4196,N_833,N_1298);
and U4197 (N_4197,N_897,N_1226);
nand U4198 (N_4198,N_298,N_2390);
or U4199 (N_4199,N_660,N_857);
nand U4200 (N_4200,N_1369,N_893);
or U4201 (N_4201,N_2492,N_2338);
nor U4202 (N_4202,N_2225,N_2682);
nor U4203 (N_4203,N_370,N_1585);
and U4204 (N_4204,N_2193,N_37);
nand U4205 (N_4205,N_1162,N_2088);
nor U4206 (N_4206,N_1904,N_2467);
nand U4207 (N_4207,N_1519,N_604);
nor U4208 (N_4208,N_2963,N_1362);
nor U4209 (N_4209,N_2252,N_2694);
nor U4210 (N_4210,N_429,N_1952);
nand U4211 (N_4211,N_2022,N_860);
or U4212 (N_4212,N_11,N_2874);
nor U4213 (N_4213,N_82,N_2791);
nand U4214 (N_4214,N_481,N_2908);
or U4215 (N_4215,N_393,N_1187);
nor U4216 (N_4216,N_1755,N_1463);
and U4217 (N_4217,N_24,N_2138);
nand U4218 (N_4218,N_2812,N_2993);
nand U4219 (N_4219,N_2689,N_2741);
or U4220 (N_4220,N_511,N_1171);
or U4221 (N_4221,N_1001,N_1887);
nor U4222 (N_4222,N_823,N_578);
nand U4223 (N_4223,N_2111,N_2695);
xnor U4224 (N_4224,N_2570,N_114);
nor U4225 (N_4225,N_1286,N_1965);
or U4226 (N_4226,N_2183,N_1384);
nand U4227 (N_4227,N_1557,N_1307);
nor U4228 (N_4228,N_1828,N_1239);
and U4229 (N_4229,N_1361,N_1615);
nor U4230 (N_4230,N_2098,N_2267);
nor U4231 (N_4231,N_2760,N_104);
or U4232 (N_4232,N_359,N_1424);
nand U4233 (N_4233,N_1610,N_1691);
and U4234 (N_4234,N_2556,N_386);
nor U4235 (N_4235,N_1342,N_665);
or U4236 (N_4236,N_1927,N_2382);
and U4237 (N_4237,N_1368,N_2657);
and U4238 (N_4238,N_1107,N_49);
nor U4239 (N_4239,N_983,N_1213);
nor U4240 (N_4240,N_1834,N_2340);
nand U4241 (N_4241,N_2568,N_1214);
or U4242 (N_4242,N_949,N_677);
nor U4243 (N_4243,N_2924,N_2369);
nor U4244 (N_4244,N_727,N_2427);
nand U4245 (N_4245,N_1465,N_1292);
or U4246 (N_4246,N_855,N_2859);
nor U4247 (N_4247,N_1249,N_1053);
nor U4248 (N_4248,N_872,N_75);
or U4249 (N_4249,N_357,N_70);
nand U4250 (N_4250,N_323,N_492);
and U4251 (N_4251,N_1642,N_1486);
nand U4252 (N_4252,N_2990,N_685);
and U4253 (N_4253,N_1852,N_2513);
and U4254 (N_4254,N_519,N_616);
and U4255 (N_4255,N_223,N_808);
nor U4256 (N_4256,N_286,N_2077);
or U4257 (N_4257,N_2429,N_2293);
nor U4258 (N_4258,N_353,N_2295);
nand U4259 (N_4259,N_988,N_2177);
and U4260 (N_4260,N_2054,N_388);
and U4261 (N_4261,N_1506,N_2796);
nand U4262 (N_4262,N_862,N_153);
or U4263 (N_4263,N_2854,N_1324);
or U4264 (N_4264,N_2128,N_2661);
nand U4265 (N_4265,N_611,N_709);
nor U4266 (N_4266,N_2549,N_149);
and U4267 (N_4267,N_141,N_73);
nor U4268 (N_4268,N_1631,N_2649);
and U4269 (N_4269,N_2511,N_1351);
nand U4270 (N_4270,N_2003,N_2575);
nand U4271 (N_4271,N_16,N_145);
nand U4272 (N_4272,N_2774,N_53);
or U4273 (N_4273,N_1605,N_793);
nor U4274 (N_4274,N_2285,N_2044);
nand U4275 (N_4275,N_1225,N_238);
nand U4276 (N_4276,N_513,N_840);
and U4277 (N_4277,N_1254,N_689);
nor U4278 (N_4278,N_1597,N_312);
and U4279 (N_4279,N_1247,N_1651);
nand U4280 (N_4280,N_2550,N_1310);
and U4281 (N_4281,N_1237,N_2795);
and U4282 (N_4282,N_2019,N_1067);
nor U4283 (N_4283,N_2656,N_1621);
and U4284 (N_4284,N_2822,N_183);
nor U4285 (N_4285,N_158,N_1364);
nor U4286 (N_4286,N_1831,N_2460);
nor U4287 (N_4287,N_2671,N_162);
and U4288 (N_4288,N_881,N_1893);
and U4289 (N_4289,N_2359,N_2771);
nand U4290 (N_4290,N_2950,N_2826);
nand U4291 (N_4291,N_184,N_635);
and U4292 (N_4292,N_1188,N_2803);
or U4293 (N_4293,N_2398,N_1526);
or U4294 (N_4294,N_284,N_310);
and U4295 (N_4295,N_2290,N_1036);
and U4296 (N_4296,N_2572,N_1105);
nor U4297 (N_4297,N_504,N_2159);
nand U4298 (N_4298,N_2234,N_889);
nor U4299 (N_4299,N_905,N_1546);
or U4300 (N_4300,N_576,N_1034);
nor U4301 (N_4301,N_2040,N_1257);
nand U4302 (N_4302,N_97,N_1934);
nor U4303 (N_4303,N_538,N_814);
and U4304 (N_4304,N_2328,N_257);
nor U4305 (N_4305,N_2023,N_2154);
nor U4306 (N_4306,N_778,N_1989);
nand U4307 (N_4307,N_216,N_982);
and U4308 (N_4308,N_959,N_1963);
or U4309 (N_4309,N_1785,N_416);
nor U4310 (N_4310,N_1643,N_2523);
or U4311 (N_4311,N_2678,N_2134);
nor U4312 (N_4312,N_2747,N_328);
and U4313 (N_4313,N_1070,N_1447);
or U4314 (N_4314,N_1021,N_2693);
nand U4315 (N_4315,N_853,N_693);
or U4316 (N_4316,N_623,N_2849);
and U4317 (N_4317,N_630,N_774);
or U4318 (N_4318,N_913,N_2512);
and U4319 (N_4319,N_654,N_1583);
and U4320 (N_4320,N_1819,N_2303);
and U4321 (N_4321,N_1707,N_1738);
nor U4322 (N_4322,N_1792,N_2420);
and U4323 (N_4323,N_1764,N_738);
and U4324 (N_4324,N_1936,N_1333);
and U4325 (N_4325,N_1375,N_1719);
and U4326 (N_4326,N_1099,N_1618);
nor U4327 (N_4327,N_1920,N_165);
nand U4328 (N_4328,N_1026,N_1556);
and U4329 (N_4329,N_2733,N_460);
or U4330 (N_4330,N_2976,N_805);
and U4331 (N_4331,N_280,N_780);
nand U4332 (N_4332,N_435,N_1957);
nor U4333 (N_4333,N_2251,N_1048);
and U4334 (N_4334,N_2064,N_1903);
nand U4335 (N_4335,N_802,N_2392);
and U4336 (N_4336,N_169,N_754);
nand U4337 (N_4337,N_2194,N_1263);
nor U4338 (N_4338,N_1121,N_2991);
or U4339 (N_4339,N_2506,N_1177);
nand U4340 (N_4340,N_650,N_599);
nand U4341 (N_4341,N_1509,N_1245);
xnor U4342 (N_4342,N_2394,N_1015);
nand U4343 (N_4343,N_2510,N_807);
nand U4344 (N_4344,N_2790,N_2341);
nand U4345 (N_4345,N_2893,N_98);
nand U4346 (N_4346,N_1635,N_1801);
nor U4347 (N_4347,N_1262,N_2381);
nand U4348 (N_4348,N_2271,N_2339);
and U4349 (N_4349,N_2489,N_828);
or U4350 (N_4350,N_304,N_1517);
and U4351 (N_4351,N_2442,N_2380);
nand U4352 (N_4352,N_188,N_272);
and U4353 (N_4353,N_2101,N_442);
nor U4354 (N_4354,N_614,N_366);
or U4355 (N_4355,N_2278,N_1082);
nor U4356 (N_4356,N_1873,N_218);
or U4357 (N_4357,N_1218,N_1909);
nor U4358 (N_4358,N_301,N_976);
or U4359 (N_4359,N_4,N_1038);
or U4360 (N_4360,N_375,N_1291);
nor U4361 (N_4361,N_1325,N_1186);
nor U4362 (N_4362,N_1396,N_2417);
or U4363 (N_4363,N_1705,N_139);
and U4364 (N_4364,N_1869,N_1326);
or U4365 (N_4365,N_6,N_2948);
or U4366 (N_4366,N_126,N_997);
nor U4367 (N_4367,N_46,N_589);
nor U4368 (N_4368,N_549,N_61);
and U4369 (N_4369,N_908,N_553);
nand U4370 (N_4370,N_351,N_593);
xnor U4371 (N_4371,N_2958,N_2405);
or U4372 (N_4372,N_2014,N_1301);
and U4373 (N_4373,N_108,N_1777);
nand U4374 (N_4374,N_2502,N_1990);
and U4375 (N_4375,N_1054,N_1789);
nor U4376 (N_4376,N_2600,N_295);
and U4377 (N_4377,N_1389,N_1686);
or U4378 (N_4378,N_1507,N_1238);
or U4379 (N_4379,N_2025,N_1468);
nand U4380 (N_4380,N_2724,N_1062);
or U4381 (N_4381,N_2046,N_2160);
or U4382 (N_4382,N_698,N_107);
and U4383 (N_4383,N_1202,N_989);
or U4384 (N_4384,N_2491,N_996);
and U4385 (N_4385,N_895,N_1228);
nor U4386 (N_4386,N_2827,N_1386);
and U4387 (N_4387,N_843,N_96);
and U4388 (N_4388,N_1423,N_2983);
nand U4389 (N_4389,N_2256,N_999);
or U4390 (N_4390,N_2136,N_1650);
nand U4391 (N_4391,N_2217,N_736);
nand U4392 (N_4392,N_2606,N_377);
or U4393 (N_4393,N_510,N_0);
nor U4394 (N_4394,N_911,N_2416);
nand U4395 (N_4395,N_2663,N_1208);
nand U4396 (N_4396,N_1529,N_2860);
nor U4397 (N_4397,N_2964,N_2354);
or U4398 (N_4398,N_2451,N_902);
and U4399 (N_4399,N_2000,N_946);
or U4400 (N_4400,N_558,N_2117);
nor U4401 (N_4401,N_1679,N_234);
and U4402 (N_4402,N_1494,N_2236);
nor U4403 (N_4403,N_2501,N_373);
or U4404 (N_4404,N_101,N_1930);
nor U4405 (N_4405,N_2010,N_168);
nand U4406 (N_4406,N_2342,N_2761);
or U4407 (N_4407,N_707,N_1954);
and U4408 (N_4408,N_30,N_2038);
nand U4409 (N_4409,N_1349,N_369);
and U4410 (N_4410,N_2273,N_1901);
nor U4411 (N_4411,N_159,N_2652);
nor U4412 (N_4412,N_2349,N_2404);
and U4413 (N_4413,N_2161,N_681);
nand U4414 (N_4414,N_219,N_1786);
nand U4415 (N_4415,N_1175,N_2509);
or U4416 (N_4416,N_1276,N_1548);
and U4417 (N_4417,N_967,N_1049);
nand U4418 (N_4418,N_699,N_2205);
nand U4419 (N_4419,N_1041,N_960);
nor U4420 (N_4420,N_706,N_1956);
or U4421 (N_4421,N_2602,N_163);
nand U4422 (N_4422,N_1017,N_2474);
nor U4423 (N_4423,N_568,N_303);
and U4424 (N_4424,N_1919,N_421);
nand U4425 (N_4425,N_121,N_459);
and U4426 (N_4426,N_2002,N_2901);
xnor U4427 (N_4427,N_1248,N_2668);
and U4428 (N_4428,N_1983,N_991);
nand U4429 (N_4429,N_1157,N_2877);
nor U4430 (N_4430,N_1080,N_2531);
and U4431 (N_4431,N_1457,N_2680);
or U4432 (N_4432,N_1467,N_1453);
nor U4433 (N_4433,N_1032,N_1012);
and U4434 (N_4434,N_958,N_2395);
nand U4435 (N_4435,N_439,N_2629);
nor U4436 (N_4436,N_1902,N_1373);
nand U4437 (N_4437,N_202,N_2224);
and U4438 (N_4438,N_829,N_1521);
nor U4439 (N_4439,N_1875,N_2688);
and U4440 (N_4440,N_103,N_811);
nor U4441 (N_4441,N_2105,N_1796);
nor U4442 (N_4442,N_209,N_573);
nor U4443 (N_4443,N_2362,N_367);
nor U4444 (N_4444,N_708,N_1484);
and U4445 (N_4445,N_1470,N_1125);
nand U4446 (N_4446,N_1385,N_89);
or U4447 (N_4447,N_2917,N_1695);
and U4448 (N_4448,N_2332,N_522);
and U4449 (N_4449,N_505,N_2921);
and U4450 (N_4450,N_1222,N_2158);
nand U4451 (N_4451,N_730,N_2586);
nand U4452 (N_4452,N_1709,N_2178);
or U4453 (N_4453,N_1530,N_1624);
or U4454 (N_4454,N_2266,N_2623);
and U4455 (N_4455,N_520,N_56);
or U4456 (N_4456,N_878,N_546);
and U4457 (N_4457,N_728,N_2201);
or U4458 (N_4458,N_2926,N_2242);
nor U4459 (N_4459,N_2923,N_1513);
nor U4460 (N_4460,N_746,N_722);
xnor U4461 (N_4461,N_1668,N_2301);
nand U4462 (N_4462,N_2131,N_1149);
nand U4463 (N_4463,N_2037,N_1716);
and U4464 (N_4464,N_1586,N_1035);
or U4465 (N_4465,N_704,N_1607);
nand U4466 (N_4466,N_1645,N_2316);
or U4467 (N_4467,N_2982,N_770);
or U4468 (N_4468,N_2858,N_2974);
nor U4469 (N_4469,N_2122,N_1242);
and U4470 (N_4470,N_2173,N_313);
xnor U4471 (N_4471,N_1706,N_2538);
nor U4472 (N_4472,N_1031,N_1449);
or U4473 (N_4473,N_2314,N_1950);
or U4474 (N_4474,N_132,N_692);
nor U4475 (N_4475,N_1488,N_2345);
nor U4476 (N_4476,N_1816,N_1677);
xnor U4477 (N_4477,N_2360,N_1193);
nor U4478 (N_4478,N_1912,N_2446);
nand U4479 (N_4479,N_2542,N_1141);
xor U4480 (N_4480,N_2573,N_319);
nand U4481 (N_4481,N_1452,N_956);
nor U4482 (N_4482,N_663,N_177);
nand U4483 (N_4483,N_547,N_1210);
nand U4484 (N_4484,N_118,N_1825);
nand U4485 (N_4485,N_453,N_789);
or U4486 (N_4486,N_674,N_1197);
or U4487 (N_4487,N_2928,N_1861);
and U4488 (N_4488,N_885,N_2645);
or U4489 (N_4489,N_2221,N_512);
nor U4490 (N_4490,N_230,N_1964);
nor U4491 (N_4491,N_32,N_2121);
nand U4492 (N_4492,N_134,N_403);
nand U4493 (N_4493,N_1160,N_907);
nand U4494 (N_4494,N_2426,N_1782);
nand U4495 (N_4495,N_2403,N_191);
nor U4496 (N_4496,N_561,N_2765);
nand U4497 (N_4497,N_1780,N_1211);
nor U4498 (N_4498,N_48,N_1959);
and U4499 (N_4499,N_655,N_1123);
or U4500 (N_4500,N_407,N_2358);
and U4501 (N_4501,N_498,N_157);
and U4502 (N_4502,N_2265,N_2816);
and U4503 (N_4503,N_540,N_383);
or U4504 (N_4504,N_2732,N_1272);
nand U4505 (N_4505,N_2727,N_1655);
and U4506 (N_4506,N_2971,N_1357);
or U4507 (N_4507,N_2249,N_2705);
nand U4508 (N_4508,N_857,N_2898);
or U4509 (N_4509,N_2776,N_950);
nor U4510 (N_4510,N_1699,N_1074);
or U4511 (N_4511,N_950,N_617);
or U4512 (N_4512,N_957,N_1240);
nand U4513 (N_4513,N_880,N_613);
nor U4514 (N_4514,N_1898,N_2202);
or U4515 (N_4515,N_1566,N_1922);
and U4516 (N_4516,N_1971,N_2880);
or U4517 (N_4517,N_2737,N_462);
nor U4518 (N_4518,N_1876,N_1172);
nand U4519 (N_4519,N_737,N_1814);
nor U4520 (N_4520,N_2361,N_151);
or U4521 (N_4521,N_786,N_1379);
nand U4522 (N_4522,N_270,N_2106);
or U4523 (N_4523,N_2178,N_1050);
and U4524 (N_4524,N_807,N_2726);
or U4525 (N_4525,N_1789,N_1180);
nand U4526 (N_4526,N_1858,N_2740);
nor U4527 (N_4527,N_45,N_2423);
and U4528 (N_4528,N_1863,N_2835);
nand U4529 (N_4529,N_615,N_350);
nand U4530 (N_4530,N_1274,N_9);
and U4531 (N_4531,N_1542,N_1909);
nor U4532 (N_4532,N_1905,N_300);
and U4533 (N_4533,N_2977,N_1879);
or U4534 (N_4534,N_519,N_2682);
nor U4535 (N_4535,N_193,N_1411);
and U4536 (N_4536,N_147,N_1942);
nand U4537 (N_4537,N_2474,N_366);
or U4538 (N_4538,N_2110,N_2155);
xnor U4539 (N_4539,N_1763,N_1087);
or U4540 (N_4540,N_260,N_1238);
or U4541 (N_4541,N_2426,N_660);
and U4542 (N_4542,N_2578,N_2357);
nand U4543 (N_4543,N_191,N_1759);
nand U4544 (N_4544,N_2152,N_1483);
and U4545 (N_4545,N_938,N_1336);
nand U4546 (N_4546,N_2150,N_2757);
or U4547 (N_4547,N_2956,N_1258);
nand U4548 (N_4548,N_263,N_2645);
nor U4549 (N_4549,N_481,N_2955);
nor U4550 (N_4550,N_872,N_346);
and U4551 (N_4551,N_1706,N_2002);
or U4552 (N_4552,N_2990,N_1991);
nor U4553 (N_4553,N_2979,N_2961);
nor U4554 (N_4554,N_431,N_2634);
and U4555 (N_4555,N_1590,N_2359);
nor U4556 (N_4556,N_2209,N_2745);
nand U4557 (N_4557,N_1236,N_2683);
and U4558 (N_4558,N_470,N_294);
nor U4559 (N_4559,N_1550,N_903);
or U4560 (N_4560,N_495,N_2902);
nor U4561 (N_4561,N_1171,N_2763);
nand U4562 (N_4562,N_1066,N_2433);
nor U4563 (N_4563,N_226,N_1732);
xor U4564 (N_4564,N_2058,N_2095);
or U4565 (N_4565,N_2593,N_2839);
nor U4566 (N_4566,N_101,N_311);
nand U4567 (N_4567,N_739,N_810);
and U4568 (N_4568,N_1260,N_2647);
or U4569 (N_4569,N_543,N_1345);
or U4570 (N_4570,N_2746,N_1295);
or U4571 (N_4571,N_160,N_592);
nor U4572 (N_4572,N_750,N_704);
nand U4573 (N_4573,N_1743,N_1194);
nor U4574 (N_4574,N_214,N_2396);
or U4575 (N_4575,N_2749,N_526);
nand U4576 (N_4576,N_1336,N_830);
nor U4577 (N_4577,N_1352,N_877);
or U4578 (N_4578,N_2412,N_2858);
nor U4579 (N_4579,N_687,N_2778);
or U4580 (N_4580,N_2465,N_1198);
and U4581 (N_4581,N_1648,N_794);
and U4582 (N_4582,N_2019,N_1017);
or U4583 (N_4583,N_2384,N_1606);
or U4584 (N_4584,N_1500,N_2316);
nor U4585 (N_4585,N_2055,N_2103);
xor U4586 (N_4586,N_1742,N_2236);
nand U4587 (N_4587,N_1240,N_2753);
or U4588 (N_4588,N_1976,N_1390);
nor U4589 (N_4589,N_2252,N_1541);
and U4590 (N_4590,N_75,N_2504);
nor U4591 (N_4591,N_959,N_820);
nand U4592 (N_4592,N_181,N_1810);
nor U4593 (N_4593,N_2869,N_2185);
nand U4594 (N_4594,N_1479,N_1925);
and U4595 (N_4595,N_1331,N_1028);
and U4596 (N_4596,N_67,N_1349);
nand U4597 (N_4597,N_2644,N_465);
nand U4598 (N_4598,N_1141,N_1654);
nor U4599 (N_4599,N_295,N_1385);
and U4600 (N_4600,N_514,N_1202);
nand U4601 (N_4601,N_590,N_2106);
nand U4602 (N_4602,N_2212,N_1792);
nand U4603 (N_4603,N_84,N_2526);
or U4604 (N_4604,N_2620,N_289);
or U4605 (N_4605,N_865,N_1605);
and U4606 (N_4606,N_1783,N_1132);
and U4607 (N_4607,N_1348,N_1359);
and U4608 (N_4608,N_997,N_2432);
nor U4609 (N_4609,N_1016,N_947);
nor U4610 (N_4610,N_106,N_1983);
or U4611 (N_4611,N_2489,N_598);
nor U4612 (N_4612,N_1654,N_2596);
nor U4613 (N_4613,N_43,N_1665);
and U4614 (N_4614,N_168,N_1853);
nand U4615 (N_4615,N_2436,N_1436);
and U4616 (N_4616,N_621,N_2917);
nand U4617 (N_4617,N_2796,N_1557);
nor U4618 (N_4618,N_1412,N_2423);
or U4619 (N_4619,N_214,N_1515);
and U4620 (N_4620,N_70,N_244);
or U4621 (N_4621,N_1156,N_1658);
nand U4622 (N_4622,N_388,N_1295);
and U4623 (N_4623,N_1179,N_2654);
or U4624 (N_4624,N_2004,N_2646);
nor U4625 (N_4625,N_2481,N_887);
and U4626 (N_4626,N_815,N_2839);
nor U4627 (N_4627,N_2326,N_859);
nand U4628 (N_4628,N_2983,N_1715);
or U4629 (N_4629,N_980,N_1780);
nor U4630 (N_4630,N_873,N_988);
nand U4631 (N_4631,N_2280,N_485);
nor U4632 (N_4632,N_2537,N_1477);
or U4633 (N_4633,N_10,N_780);
nor U4634 (N_4634,N_735,N_2958);
nand U4635 (N_4635,N_1568,N_965);
nand U4636 (N_4636,N_1511,N_2196);
and U4637 (N_4637,N_2197,N_2606);
nand U4638 (N_4638,N_298,N_761);
nor U4639 (N_4639,N_2597,N_856);
and U4640 (N_4640,N_1196,N_1159);
nand U4641 (N_4641,N_380,N_515);
and U4642 (N_4642,N_2631,N_1066);
nor U4643 (N_4643,N_1448,N_2945);
nor U4644 (N_4644,N_2415,N_552);
nand U4645 (N_4645,N_534,N_1853);
and U4646 (N_4646,N_1701,N_2421);
and U4647 (N_4647,N_1972,N_1669);
or U4648 (N_4648,N_360,N_2674);
or U4649 (N_4649,N_476,N_2490);
or U4650 (N_4650,N_2210,N_2470);
xnor U4651 (N_4651,N_1968,N_1007);
or U4652 (N_4652,N_88,N_2164);
nand U4653 (N_4653,N_2614,N_228);
nor U4654 (N_4654,N_1305,N_2098);
or U4655 (N_4655,N_1002,N_2070);
nand U4656 (N_4656,N_2919,N_2258);
and U4657 (N_4657,N_2701,N_1451);
xor U4658 (N_4658,N_63,N_1952);
nor U4659 (N_4659,N_1659,N_2874);
and U4660 (N_4660,N_1979,N_1804);
nor U4661 (N_4661,N_1527,N_1323);
or U4662 (N_4662,N_663,N_1708);
or U4663 (N_4663,N_415,N_2152);
nand U4664 (N_4664,N_543,N_492);
and U4665 (N_4665,N_810,N_1265);
and U4666 (N_4666,N_1946,N_2467);
or U4667 (N_4667,N_2083,N_2197);
nor U4668 (N_4668,N_176,N_815);
and U4669 (N_4669,N_2514,N_232);
and U4670 (N_4670,N_565,N_431);
and U4671 (N_4671,N_577,N_1365);
nand U4672 (N_4672,N_1120,N_125);
nand U4673 (N_4673,N_1395,N_1279);
nor U4674 (N_4674,N_386,N_2229);
and U4675 (N_4675,N_2409,N_82);
or U4676 (N_4676,N_2215,N_1379);
and U4677 (N_4677,N_2220,N_1209);
nand U4678 (N_4678,N_746,N_1523);
and U4679 (N_4679,N_424,N_922);
or U4680 (N_4680,N_1682,N_605);
nor U4681 (N_4681,N_223,N_755);
and U4682 (N_4682,N_2992,N_2440);
nand U4683 (N_4683,N_1834,N_815);
or U4684 (N_4684,N_574,N_1524);
and U4685 (N_4685,N_1874,N_2194);
nor U4686 (N_4686,N_501,N_1300);
or U4687 (N_4687,N_2190,N_5);
nand U4688 (N_4688,N_2876,N_2229);
nor U4689 (N_4689,N_1210,N_1549);
nor U4690 (N_4690,N_1051,N_896);
nor U4691 (N_4691,N_365,N_663);
nand U4692 (N_4692,N_1582,N_535);
nor U4693 (N_4693,N_421,N_816);
and U4694 (N_4694,N_1206,N_1876);
nand U4695 (N_4695,N_938,N_1010);
nand U4696 (N_4696,N_2347,N_1699);
nand U4697 (N_4697,N_2091,N_2436);
nand U4698 (N_4698,N_2875,N_1180);
nand U4699 (N_4699,N_1246,N_873);
nand U4700 (N_4700,N_250,N_1984);
or U4701 (N_4701,N_696,N_1969);
and U4702 (N_4702,N_1955,N_2306);
and U4703 (N_4703,N_838,N_221);
nand U4704 (N_4704,N_1105,N_782);
or U4705 (N_4705,N_1108,N_1572);
or U4706 (N_4706,N_1618,N_535);
and U4707 (N_4707,N_225,N_2107);
or U4708 (N_4708,N_1235,N_248);
nand U4709 (N_4709,N_194,N_2571);
nand U4710 (N_4710,N_565,N_1488);
nor U4711 (N_4711,N_995,N_1799);
nor U4712 (N_4712,N_341,N_1514);
or U4713 (N_4713,N_1669,N_1546);
and U4714 (N_4714,N_2153,N_577);
nor U4715 (N_4715,N_82,N_2882);
nor U4716 (N_4716,N_1091,N_1127);
and U4717 (N_4717,N_1081,N_1890);
nor U4718 (N_4718,N_2251,N_2780);
and U4719 (N_4719,N_1807,N_1520);
nor U4720 (N_4720,N_1346,N_2016);
or U4721 (N_4721,N_1185,N_1355);
and U4722 (N_4722,N_1636,N_484);
nor U4723 (N_4723,N_2665,N_1164);
and U4724 (N_4724,N_2559,N_1800);
nor U4725 (N_4725,N_1003,N_399);
nand U4726 (N_4726,N_2309,N_71);
nand U4727 (N_4727,N_478,N_1138);
nor U4728 (N_4728,N_2319,N_366);
nor U4729 (N_4729,N_1501,N_1402);
nor U4730 (N_4730,N_504,N_1838);
nand U4731 (N_4731,N_300,N_742);
xor U4732 (N_4732,N_963,N_11);
nand U4733 (N_4733,N_1140,N_1252);
nor U4734 (N_4734,N_247,N_661);
nand U4735 (N_4735,N_891,N_416);
and U4736 (N_4736,N_578,N_780);
or U4737 (N_4737,N_1479,N_1797);
xor U4738 (N_4738,N_2238,N_1093);
and U4739 (N_4739,N_2971,N_1959);
xor U4740 (N_4740,N_1520,N_2949);
or U4741 (N_4741,N_2578,N_2404);
nor U4742 (N_4742,N_1652,N_294);
nand U4743 (N_4743,N_2021,N_1175);
xor U4744 (N_4744,N_693,N_602);
or U4745 (N_4745,N_2418,N_518);
xor U4746 (N_4746,N_10,N_1571);
xor U4747 (N_4747,N_1044,N_496);
or U4748 (N_4748,N_1651,N_12);
nor U4749 (N_4749,N_1021,N_821);
or U4750 (N_4750,N_121,N_76);
or U4751 (N_4751,N_986,N_1319);
or U4752 (N_4752,N_694,N_1064);
or U4753 (N_4753,N_1259,N_2929);
nor U4754 (N_4754,N_525,N_1811);
or U4755 (N_4755,N_2114,N_2247);
nand U4756 (N_4756,N_2769,N_556);
or U4757 (N_4757,N_2948,N_2268);
nor U4758 (N_4758,N_895,N_1840);
and U4759 (N_4759,N_991,N_212);
and U4760 (N_4760,N_378,N_1793);
nor U4761 (N_4761,N_740,N_36);
and U4762 (N_4762,N_1517,N_1007);
nor U4763 (N_4763,N_1030,N_2309);
and U4764 (N_4764,N_854,N_1958);
nand U4765 (N_4765,N_376,N_557);
nand U4766 (N_4766,N_215,N_2438);
nor U4767 (N_4767,N_868,N_644);
nor U4768 (N_4768,N_881,N_2494);
nand U4769 (N_4769,N_41,N_1116);
nor U4770 (N_4770,N_2691,N_2156);
and U4771 (N_4771,N_1516,N_1445);
xor U4772 (N_4772,N_2172,N_1363);
nand U4773 (N_4773,N_1268,N_365);
nand U4774 (N_4774,N_2114,N_2735);
or U4775 (N_4775,N_2276,N_2592);
xor U4776 (N_4776,N_1818,N_394);
and U4777 (N_4777,N_754,N_1866);
nor U4778 (N_4778,N_571,N_1589);
nor U4779 (N_4779,N_513,N_1999);
or U4780 (N_4780,N_792,N_1142);
and U4781 (N_4781,N_244,N_1055);
nand U4782 (N_4782,N_1596,N_1660);
and U4783 (N_4783,N_589,N_195);
and U4784 (N_4784,N_934,N_71);
nor U4785 (N_4785,N_2279,N_1407);
nand U4786 (N_4786,N_1771,N_1633);
and U4787 (N_4787,N_2782,N_2128);
nor U4788 (N_4788,N_2680,N_364);
or U4789 (N_4789,N_2878,N_88);
nand U4790 (N_4790,N_2302,N_892);
nor U4791 (N_4791,N_1556,N_2678);
or U4792 (N_4792,N_206,N_142);
or U4793 (N_4793,N_2771,N_33);
or U4794 (N_4794,N_724,N_2302);
nor U4795 (N_4795,N_620,N_2707);
nand U4796 (N_4796,N_251,N_1142);
or U4797 (N_4797,N_1795,N_2935);
and U4798 (N_4798,N_2802,N_1209);
nand U4799 (N_4799,N_192,N_1997);
or U4800 (N_4800,N_1498,N_2703);
and U4801 (N_4801,N_1659,N_2597);
xor U4802 (N_4802,N_511,N_397);
or U4803 (N_4803,N_1075,N_2428);
nor U4804 (N_4804,N_141,N_602);
nor U4805 (N_4805,N_236,N_2396);
nor U4806 (N_4806,N_1633,N_198);
and U4807 (N_4807,N_105,N_2268);
nor U4808 (N_4808,N_2284,N_1684);
nor U4809 (N_4809,N_1045,N_828);
or U4810 (N_4810,N_1134,N_2143);
nand U4811 (N_4811,N_1416,N_867);
or U4812 (N_4812,N_530,N_2699);
nand U4813 (N_4813,N_1385,N_587);
nor U4814 (N_4814,N_2975,N_233);
nor U4815 (N_4815,N_1234,N_293);
nor U4816 (N_4816,N_583,N_657);
nand U4817 (N_4817,N_1525,N_2350);
nor U4818 (N_4818,N_692,N_2422);
nor U4819 (N_4819,N_2476,N_1141);
and U4820 (N_4820,N_2720,N_54);
nand U4821 (N_4821,N_454,N_2668);
nand U4822 (N_4822,N_1898,N_2628);
or U4823 (N_4823,N_345,N_2316);
or U4824 (N_4824,N_2401,N_1854);
nor U4825 (N_4825,N_578,N_1273);
xor U4826 (N_4826,N_1,N_1652);
nand U4827 (N_4827,N_2812,N_2557);
nand U4828 (N_4828,N_513,N_1323);
or U4829 (N_4829,N_548,N_2363);
nor U4830 (N_4830,N_951,N_2514);
nand U4831 (N_4831,N_2610,N_2933);
or U4832 (N_4832,N_793,N_977);
and U4833 (N_4833,N_828,N_206);
nand U4834 (N_4834,N_1415,N_2394);
nor U4835 (N_4835,N_614,N_2775);
nor U4836 (N_4836,N_1951,N_550);
nor U4837 (N_4837,N_255,N_665);
nand U4838 (N_4838,N_1591,N_1961);
and U4839 (N_4839,N_254,N_2783);
and U4840 (N_4840,N_919,N_2581);
and U4841 (N_4841,N_2922,N_1418);
nor U4842 (N_4842,N_1865,N_2244);
xnor U4843 (N_4843,N_1116,N_2431);
and U4844 (N_4844,N_1285,N_2513);
or U4845 (N_4845,N_1019,N_577);
or U4846 (N_4846,N_2399,N_164);
or U4847 (N_4847,N_2096,N_58);
nand U4848 (N_4848,N_340,N_2406);
nand U4849 (N_4849,N_2187,N_2325);
or U4850 (N_4850,N_2916,N_2441);
or U4851 (N_4851,N_2968,N_2231);
and U4852 (N_4852,N_1379,N_1592);
or U4853 (N_4853,N_629,N_2087);
and U4854 (N_4854,N_125,N_1772);
nand U4855 (N_4855,N_323,N_667);
nor U4856 (N_4856,N_234,N_663);
nor U4857 (N_4857,N_1306,N_3);
nand U4858 (N_4858,N_839,N_1834);
nor U4859 (N_4859,N_899,N_740);
or U4860 (N_4860,N_172,N_525);
or U4861 (N_4861,N_1888,N_843);
nor U4862 (N_4862,N_224,N_1640);
nand U4863 (N_4863,N_865,N_971);
and U4864 (N_4864,N_658,N_911);
or U4865 (N_4865,N_1960,N_994);
and U4866 (N_4866,N_475,N_1900);
or U4867 (N_4867,N_2599,N_851);
nor U4868 (N_4868,N_1622,N_403);
nand U4869 (N_4869,N_893,N_423);
nor U4870 (N_4870,N_764,N_1788);
nand U4871 (N_4871,N_406,N_2655);
nand U4872 (N_4872,N_55,N_2708);
nor U4873 (N_4873,N_1110,N_1861);
and U4874 (N_4874,N_2101,N_262);
and U4875 (N_4875,N_245,N_1485);
or U4876 (N_4876,N_811,N_27);
or U4877 (N_4877,N_2876,N_898);
nand U4878 (N_4878,N_2018,N_1729);
nor U4879 (N_4879,N_2309,N_1773);
or U4880 (N_4880,N_574,N_1236);
nand U4881 (N_4881,N_495,N_1215);
nand U4882 (N_4882,N_1155,N_940);
or U4883 (N_4883,N_442,N_1714);
and U4884 (N_4884,N_1306,N_1179);
or U4885 (N_4885,N_1996,N_956);
or U4886 (N_4886,N_1359,N_1667);
and U4887 (N_4887,N_2531,N_2330);
xnor U4888 (N_4888,N_1424,N_479);
and U4889 (N_4889,N_1417,N_2514);
or U4890 (N_4890,N_200,N_1344);
nor U4891 (N_4891,N_1993,N_320);
and U4892 (N_4892,N_640,N_1793);
nor U4893 (N_4893,N_663,N_927);
nor U4894 (N_4894,N_1646,N_152);
nor U4895 (N_4895,N_1820,N_2660);
nand U4896 (N_4896,N_1572,N_2109);
or U4897 (N_4897,N_1614,N_2083);
nor U4898 (N_4898,N_2494,N_2774);
nand U4899 (N_4899,N_1307,N_2439);
or U4900 (N_4900,N_289,N_598);
nor U4901 (N_4901,N_2725,N_1149);
nor U4902 (N_4902,N_1312,N_2169);
or U4903 (N_4903,N_540,N_2606);
or U4904 (N_4904,N_641,N_269);
nor U4905 (N_4905,N_2063,N_2814);
xnor U4906 (N_4906,N_2630,N_365);
nand U4907 (N_4907,N_1432,N_1631);
nor U4908 (N_4908,N_1995,N_891);
and U4909 (N_4909,N_753,N_1834);
xnor U4910 (N_4910,N_2742,N_121);
nor U4911 (N_4911,N_2414,N_2083);
and U4912 (N_4912,N_1188,N_1471);
and U4913 (N_4913,N_2420,N_290);
and U4914 (N_4914,N_1523,N_1641);
or U4915 (N_4915,N_1129,N_2151);
nand U4916 (N_4916,N_2334,N_185);
nand U4917 (N_4917,N_299,N_2182);
or U4918 (N_4918,N_670,N_1234);
nor U4919 (N_4919,N_2303,N_2519);
nor U4920 (N_4920,N_2256,N_2692);
and U4921 (N_4921,N_579,N_650);
nand U4922 (N_4922,N_678,N_442);
or U4923 (N_4923,N_1488,N_1697);
nand U4924 (N_4924,N_2763,N_2473);
or U4925 (N_4925,N_759,N_479);
and U4926 (N_4926,N_2455,N_1939);
nor U4927 (N_4927,N_1876,N_1313);
and U4928 (N_4928,N_697,N_2665);
or U4929 (N_4929,N_1286,N_2231);
nor U4930 (N_4930,N_44,N_1068);
and U4931 (N_4931,N_1833,N_1086);
nand U4932 (N_4932,N_1020,N_2575);
nand U4933 (N_4933,N_2189,N_12);
or U4934 (N_4934,N_2773,N_2598);
nor U4935 (N_4935,N_1371,N_2473);
nand U4936 (N_4936,N_1033,N_732);
nor U4937 (N_4937,N_2704,N_2714);
or U4938 (N_4938,N_2022,N_5);
nor U4939 (N_4939,N_2861,N_870);
and U4940 (N_4940,N_2063,N_2470);
or U4941 (N_4941,N_375,N_925);
nand U4942 (N_4942,N_579,N_1160);
or U4943 (N_4943,N_2526,N_2);
nand U4944 (N_4944,N_1631,N_2272);
nor U4945 (N_4945,N_295,N_2690);
nand U4946 (N_4946,N_73,N_2882);
nand U4947 (N_4947,N_1119,N_1760);
nand U4948 (N_4948,N_150,N_2094);
or U4949 (N_4949,N_2932,N_227);
nand U4950 (N_4950,N_1821,N_227);
nand U4951 (N_4951,N_1310,N_757);
nand U4952 (N_4952,N_419,N_2076);
nor U4953 (N_4953,N_284,N_1565);
nor U4954 (N_4954,N_436,N_832);
and U4955 (N_4955,N_379,N_1541);
or U4956 (N_4956,N_2119,N_1233);
nor U4957 (N_4957,N_882,N_805);
nand U4958 (N_4958,N_2125,N_1207);
nand U4959 (N_4959,N_1607,N_135);
nor U4960 (N_4960,N_523,N_2859);
or U4961 (N_4961,N_2352,N_1033);
nor U4962 (N_4962,N_2174,N_2649);
and U4963 (N_4963,N_364,N_1708);
nor U4964 (N_4964,N_2566,N_2948);
nand U4965 (N_4965,N_2120,N_229);
nor U4966 (N_4966,N_2393,N_991);
and U4967 (N_4967,N_2273,N_2593);
nor U4968 (N_4968,N_2843,N_352);
or U4969 (N_4969,N_2885,N_2949);
or U4970 (N_4970,N_2627,N_2303);
nand U4971 (N_4971,N_2107,N_89);
nor U4972 (N_4972,N_475,N_1608);
nand U4973 (N_4973,N_1373,N_1917);
nand U4974 (N_4974,N_1895,N_2632);
and U4975 (N_4975,N_1140,N_933);
nand U4976 (N_4976,N_2590,N_2656);
nand U4977 (N_4977,N_2822,N_2544);
and U4978 (N_4978,N_545,N_1658);
or U4979 (N_4979,N_1056,N_274);
nor U4980 (N_4980,N_52,N_1468);
and U4981 (N_4981,N_476,N_1633);
nand U4982 (N_4982,N_1684,N_983);
nor U4983 (N_4983,N_2312,N_2927);
nand U4984 (N_4984,N_448,N_1422);
and U4985 (N_4985,N_2283,N_633);
nand U4986 (N_4986,N_106,N_2782);
or U4987 (N_4987,N_1760,N_1703);
nand U4988 (N_4988,N_2516,N_1845);
or U4989 (N_4989,N_2302,N_2727);
nor U4990 (N_4990,N_2745,N_1070);
nor U4991 (N_4991,N_2133,N_1950);
nand U4992 (N_4992,N_541,N_618);
nand U4993 (N_4993,N_486,N_2681);
nand U4994 (N_4994,N_2523,N_1013);
or U4995 (N_4995,N_1371,N_2750);
nor U4996 (N_4996,N_1108,N_488);
or U4997 (N_4997,N_210,N_0);
or U4998 (N_4998,N_1218,N_2672);
and U4999 (N_4999,N_1917,N_2988);
or U5000 (N_5000,N_2020,N_2268);
nor U5001 (N_5001,N_1489,N_1695);
or U5002 (N_5002,N_2636,N_134);
or U5003 (N_5003,N_1727,N_20);
nor U5004 (N_5004,N_2223,N_1626);
or U5005 (N_5005,N_1246,N_667);
and U5006 (N_5006,N_2209,N_778);
or U5007 (N_5007,N_125,N_209);
xor U5008 (N_5008,N_23,N_414);
nand U5009 (N_5009,N_109,N_822);
nand U5010 (N_5010,N_322,N_1210);
and U5011 (N_5011,N_1273,N_1202);
nand U5012 (N_5012,N_2916,N_820);
and U5013 (N_5013,N_2625,N_1580);
nor U5014 (N_5014,N_1619,N_2388);
nor U5015 (N_5015,N_1504,N_236);
nor U5016 (N_5016,N_358,N_1086);
nor U5017 (N_5017,N_1429,N_648);
or U5018 (N_5018,N_2391,N_574);
nor U5019 (N_5019,N_1204,N_1663);
and U5020 (N_5020,N_2905,N_1826);
and U5021 (N_5021,N_2415,N_1022);
or U5022 (N_5022,N_1500,N_572);
nor U5023 (N_5023,N_1139,N_2358);
nand U5024 (N_5024,N_1771,N_465);
or U5025 (N_5025,N_641,N_2580);
and U5026 (N_5026,N_66,N_698);
and U5027 (N_5027,N_2162,N_313);
and U5028 (N_5028,N_511,N_2974);
xor U5029 (N_5029,N_1807,N_1020);
or U5030 (N_5030,N_547,N_1095);
nor U5031 (N_5031,N_2718,N_2277);
nand U5032 (N_5032,N_2482,N_35);
nor U5033 (N_5033,N_624,N_2307);
or U5034 (N_5034,N_2278,N_1002);
nor U5035 (N_5035,N_340,N_1305);
and U5036 (N_5036,N_1841,N_980);
or U5037 (N_5037,N_2524,N_1803);
and U5038 (N_5038,N_2679,N_2486);
or U5039 (N_5039,N_903,N_476);
or U5040 (N_5040,N_1622,N_1915);
nand U5041 (N_5041,N_1970,N_1175);
nand U5042 (N_5042,N_390,N_954);
and U5043 (N_5043,N_1307,N_2638);
and U5044 (N_5044,N_2095,N_1566);
nand U5045 (N_5045,N_981,N_1440);
nand U5046 (N_5046,N_2896,N_833);
xor U5047 (N_5047,N_1893,N_1077);
nand U5048 (N_5048,N_1903,N_1554);
and U5049 (N_5049,N_1473,N_2362);
and U5050 (N_5050,N_2815,N_2920);
nor U5051 (N_5051,N_1841,N_1446);
nor U5052 (N_5052,N_1387,N_1928);
or U5053 (N_5053,N_761,N_491);
nand U5054 (N_5054,N_69,N_1268);
and U5055 (N_5055,N_2850,N_1863);
nand U5056 (N_5056,N_2033,N_1863);
or U5057 (N_5057,N_2827,N_2303);
or U5058 (N_5058,N_1686,N_761);
nor U5059 (N_5059,N_2272,N_1164);
nor U5060 (N_5060,N_2370,N_2235);
nand U5061 (N_5061,N_1171,N_2017);
nand U5062 (N_5062,N_554,N_1434);
nand U5063 (N_5063,N_1338,N_2896);
and U5064 (N_5064,N_655,N_181);
nand U5065 (N_5065,N_2977,N_2012);
nand U5066 (N_5066,N_522,N_1890);
and U5067 (N_5067,N_1055,N_2371);
and U5068 (N_5068,N_2001,N_1174);
nor U5069 (N_5069,N_2989,N_2605);
and U5070 (N_5070,N_2768,N_1791);
nand U5071 (N_5071,N_2052,N_1056);
and U5072 (N_5072,N_1579,N_1086);
or U5073 (N_5073,N_166,N_363);
xnor U5074 (N_5074,N_2101,N_2673);
nand U5075 (N_5075,N_2107,N_2476);
or U5076 (N_5076,N_1414,N_1469);
or U5077 (N_5077,N_2479,N_2533);
nor U5078 (N_5078,N_2127,N_1979);
xnor U5079 (N_5079,N_315,N_1822);
nor U5080 (N_5080,N_2600,N_1491);
nor U5081 (N_5081,N_2028,N_1777);
or U5082 (N_5082,N_1062,N_2793);
and U5083 (N_5083,N_865,N_1687);
nor U5084 (N_5084,N_1809,N_2060);
or U5085 (N_5085,N_300,N_1614);
and U5086 (N_5086,N_326,N_1852);
and U5087 (N_5087,N_2150,N_2453);
nor U5088 (N_5088,N_9,N_1855);
nor U5089 (N_5089,N_2441,N_1664);
nor U5090 (N_5090,N_1259,N_1659);
nor U5091 (N_5091,N_1508,N_402);
or U5092 (N_5092,N_2307,N_1119);
or U5093 (N_5093,N_2398,N_292);
and U5094 (N_5094,N_1170,N_1631);
nand U5095 (N_5095,N_261,N_797);
and U5096 (N_5096,N_576,N_2030);
or U5097 (N_5097,N_2346,N_1006);
nor U5098 (N_5098,N_2567,N_279);
nand U5099 (N_5099,N_2945,N_887);
nor U5100 (N_5100,N_2224,N_1161);
and U5101 (N_5101,N_351,N_1078);
nand U5102 (N_5102,N_2815,N_1638);
or U5103 (N_5103,N_2643,N_2060);
and U5104 (N_5104,N_999,N_2339);
nand U5105 (N_5105,N_2711,N_2568);
and U5106 (N_5106,N_787,N_194);
or U5107 (N_5107,N_502,N_200);
or U5108 (N_5108,N_2644,N_2563);
nor U5109 (N_5109,N_1877,N_2306);
nor U5110 (N_5110,N_349,N_1843);
or U5111 (N_5111,N_999,N_1685);
and U5112 (N_5112,N_1216,N_1206);
nand U5113 (N_5113,N_725,N_2410);
or U5114 (N_5114,N_1009,N_2259);
or U5115 (N_5115,N_1008,N_2590);
nor U5116 (N_5116,N_2733,N_784);
and U5117 (N_5117,N_1333,N_2192);
or U5118 (N_5118,N_677,N_178);
nand U5119 (N_5119,N_2553,N_2658);
or U5120 (N_5120,N_929,N_985);
nand U5121 (N_5121,N_38,N_2477);
and U5122 (N_5122,N_1278,N_1098);
or U5123 (N_5123,N_2019,N_1818);
and U5124 (N_5124,N_961,N_313);
or U5125 (N_5125,N_474,N_2166);
or U5126 (N_5126,N_2403,N_142);
and U5127 (N_5127,N_754,N_422);
nor U5128 (N_5128,N_870,N_482);
nor U5129 (N_5129,N_2571,N_1149);
and U5130 (N_5130,N_2971,N_2532);
nand U5131 (N_5131,N_10,N_1936);
nor U5132 (N_5132,N_2024,N_2425);
nand U5133 (N_5133,N_875,N_520);
nand U5134 (N_5134,N_489,N_1131);
nand U5135 (N_5135,N_2153,N_2067);
and U5136 (N_5136,N_2022,N_1785);
and U5137 (N_5137,N_2589,N_627);
or U5138 (N_5138,N_1773,N_982);
nand U5139 (N_5139,N_1513,N_2244);
or U5140 (N_5140,N_1579,N_1447);
or U5141 (N_5141,N_208,N_1146);
nor U5142 (N_5142,N_2757,N_2111);
or U5143 (N_5143,N_1113,N_1650);
or U5144 (N_5144,N_2913,N_985);
or U5145 (N_5145,N_2046,N_44);
and U5146 (N_5146,N_2005,N_31);
nand U5147 (N_5147,N_2589,N_763);
or U5148 (N_5148,N_784,N_1145);
and U5149 (N_5149,N_1999,N_566);
nand U5150 (N_5150,N_2096,N_710);
nor U5151 (N_5151,N_1630,N_1277);
and U5152 (N_5152,N_804,N_2042);
and U5153 (N_5153,N_2030,N_522);
or U5154 (N_5154,N_2668,N_2002);
nor U5155 (N_5155,N_1702,N_1807);
nand U5156 (N_5156,N_1945,N_92);
xnor U5157 (N_5157,N_1431,N_2197);
or U5158 (N_5158,N_861,N_977);
nor U5159 (N_5159,N_769,N_297);
nand U5160 (N_5160,N_2862,N_1930);
and U5161 (N_5161,N_624,N_1370);
nor U5162 (N_5162,N_1979,N_58);
xnor U5163 (N_5163,N_759,N_1186);
and U5164 (N_5164,N_344,N_409);
or U5165 (N_5165,N_830,N_13);
nor U5166 (N_5166,N_1033,N_913);
nand U5167 (N_5167,N_2787,N_1754);
nand U5168 (N_5168,N_1337,N_1063);
and U5169 (N_5169,N_2853,N_1447);
and U5170 (N_5170,N_1215,N_736);
nor U5171 (N_5171,N_67,N_2715);
nor U5172 (N_5172,N_2613,N_2506);
or U5173 (N_5173,N_913,N_1162);
nor U5174 (N_5174,N_2722,N_1767);
or U5175 (N_5175,N_1735,N_1663);
and U5176 (N_5176,N_1028,N_385);
nor U5177 (N_5177,N_277,N_453);
nand U5178 (N_5178,N_1661,N_1340);
or U5179 (N_5179,N_2833,N_2287);
or U5180 (N_5180,N_2652,N_1791);
nor U5181 (N_5181,N_318,N_457);
and U5182 (N_5182,N_1248,N_2414);
or U5183 (N_5183,N_1158,N_770);
nand U5184 (N_5184,N_158,N_1705);
nor U5185 (N_5185,N_272,N_1859);
or U5186 (N_5186,N_1679,N_487);
nand U5187 (N_5187,N_1278,N_2863);
or U5188 (N_5188,N_1202,N_2190);
nor U5189 (N_5189,N_2368,N_1607);
nand U5190 (N_5190,N_2,N_646);
nor U5191 (N_5191,N_2810,N_2742);
nor U5192 (N_5192,N_2090,N_2261);
and U5193 (N_5193,N_2284,N_2103);
and U5194 (N_5194,N_2726,N_484);
and U5195 (N_5195,N_2862,N_1501);
or U5196 (N_5196,N_304,N_2913);
nor U5197 (N_5197,N_899,N_2982);
xnor U5198 (N_5198,N_243,N_877);
nand U5199 (N_5199,N_995,N_2826);
and U5200 (N_5200,N_698,N_360);
or U5201 (N_5201,N_2983,N_905);
or U5202 (N_5202,N_1020,N_716);
nor U5203 (N_5203,N_2457,N_2188);
nand U5204 (N_5204,N_362,N_1429);
nand U5205 (N_5205,N_1115,N_798);
or U5206 (N_5206,N_879,N_1063);
nor U5207 (N_5207,N_1561,N_31);
and U5208 (N_5208,N_2869,N_102);
or U5209 (N_5209,N_679,N_1763);
nand U5210 (N_5210,N_2215,N_290);
nor U5211 (N_5211,N_821,N_2773);
nand U5212 (N_5212,N_2010,N_2791);
and U5213 (N_5213,N_2817,N_74);
nand U5214 (N_5214,N_1597,N_1645);
nand U5215 (N_5215,N_2060,N_1342);
nor U5216 (N_5216,N_2261,N_1529);
and U5217 (N_5217,N_2191,N_2513);
nor U5218 (N_5218,N_1474,N_834);
and U5219 (N_5219,N_2420,N_479);
and U5220 (N_5220,N_2049,N_2048);
or U5221 (N_5221,N_2244,N_199);
nand U5222 (N_5222,N_1282,N_2680);
nand U5223 (N_5223,N_240,N_2367);
nor U5224 (N_5224,N_2607,N_573);
or U5225 (N_5225,N_666,N_2969);
nor U5226 (N_5226,N_1216,N_1847);
nor U5227 (N_5227,N_2624,N_91);
nand U5228 (N_5228,N_2203,N_1262);
or U5229 (N_5229,N_1830,N_2758);
and U5230 (N_5230,N_2124,N_2415);
nand U5231 (N_5231,N_1480,N_765);
nor U5232 (N_5232,N_2540,N_2554);
nand U5233 (N_5233,N_2015,N_2407);
nand U5234 (N_5234,N_2265,N_49);
nor U5235 (N_5235,N_2896,N_1215);
or U5236 (N_5236,N_482,N_504);
nor U5237 (N_5237,N_1942,N_1174);
nor U5238 (N_5238,N_1689,N_547);
or U5239 (N_5239,N_122,N_2309);
and U5240 (N_5240,N_1868,N_1078);
or U5241 (N_5241,N_1630,N_2404);
and U5242 (N_5242,N_1347,N_1557);
and U5243 (N_5243,N_1841,N_658);
nand U5244 (N_5244,N_2674,N_979);
and U5245 (N_5245,N_502,N_333);
or U5246 (N_5246,N_2838,N_757);
or U5247 (N_5247,N_215,N_2345);
and U5248 (N_5248,N_2524,N_2540);
or U5249 (N_5249,N_1364,N_1148);
nand U5250 (N_5250,N_2806,N_1239);
and U5251 (N_5251,N_1024,N_1941);
or U5252 (N_5252,N_2894,N_2826);
and U5253 (N_5253,N_1620,N_588);
and U5254 (N_5254,N_1882,N_2269);
nor U5255 (N_5255,N_366,N_1364);
nand U5256 (N_5256,N_2461,N_1240);
or U5257 (N_5257,N_2092,N_488);
nor U5258 (N_5258,N_2062,N_2031);
xor U5259 (N_5259,N_1356,N_334);
or U5260 (N_5260,N_1571,N_1812);
or U5261 (N_5261,N_781,N_594);
and U5262 (N_5262,N_692,N_2766);
or U5263 (N_5263,N_1950,N_2191);
nand U5264 (N_5264,N_2839,N_2463);
or U5265 (N_5265,N_117,N_2453);
nand U5266 (N_5266,N_446,N_1889);
or U5267 (N_5267,N_2484,N_614);
nor U5268 (N_5268,N_2750,N_2823);
or U5269 (N_5269,N_2400,N_2669);
nor U5270 (N_5270,N_2455,N_396);
nor U5271 (N_5271,N_11,N_412);
and U5272 (N_5272,N_2017,N_2582);
and U5273 (N_5273,N_2589,N_79);
nand U5274 (N_5274,N_252,N_1457);
nand U5275 (N_5275,N_360,N_2472);
nor U5276 (N_5276,N_2099,N_627);
or U5277 (N_5277,N_1220,N_1969);
and U5278 (N_5278,N_196,N_1050);
nor U5279 (N_5279,N_2481,N_1930);
and U5280 (N_5280,N_2998,N_2309);
nand U5281 (N_5281,N_312,N_2616);
nor U5282 (N_5282,N_2307,N_2427);
nor U5283 (N_5283,N_2306,N_2747);
or U5284 (N_5284,N_1117,N_240);
or U5285 (N_5285,N_2222,N_1010);
and U5286 (N_5286,N_2020,N_2924);
nor U5287 (N_5287,N_2860,N_203);
or U5288 (N_5288,N_1656,N_872);
xnor U5289 (N_5289,N_2257,N_1816);
nor U5290 (N_5290,N_85,N_2102);
or U5291 (N_5291,N_1167,N_2135);
nand U5292 (N_5292,N_1323,N_1992);
nor U5293 (N_5293,N_397,N_2822);
or U5294 (N_5294,N_208,N_2091);
or U5295 (N_5295,N_2852,N_1401);
or U5296 (N_5296,N_2775,N_2371);
or U5297 (N_5297,N_291,N_1440);
or U5298 (N_5298,N_2956,N_2317);
or U5299 (N_5299,N_1682,N_1403);
or U5300 (N_5300,N_2715,N_43);
nand U5301 (N_5301,N_2749,N_243);
nor U5302 (N_5302,N_21,N_936);
nor U5303 (N_5303,N_531,N_1479);
or U5304 (N_5304,N_1672,N_1139);
nand U5305 (N_5305,N_549,N_1482);
and U5306 (N_5306,N_2432,N_928);
nor U5307 (N_5307,N_2178,N_2801);
and U5308 (N_5308,N_1288,N_1403);
nor U5309 (N_5309,N_2417,N_1591);
or U5310 (N_5310,N_1640,N_2653);
nand U5311 (N_5311,N_10,N_389);
or U5312 (N_5312,N_2681,N_2694);
xnor U5313 (N_5313,N_1870,N_1532);
xnor U5314 (N_5314,N_1937,N_404);
nor U5315 (N_5315,N_718,N_213);
nor U5316 (N_5316,N_1355,N_2543);
nor U5317 (N_5317,N_2515,N_2694);
nor U5318 (N_5318,N_1124,N_341);
nand U5319 (N_5319,N_2580,N_2246);
nor U5320 (N_5320,N_2523,N_2595);
or U5321 (N_5321,N_625,N_999);
or U5322 (N_5322,N_2013,N_918);
and U5323 (N_5323,N_2007,N_2543);
or U5324 (N_5324,N_908,N_1453);
nand U5325 (N_5325,N_1619,N_2219);
or U5326 (N_5326,N_2792,N_909);
or U5327 (N_5327,N_2655,N_2329);
and U5328 (N_5328,N_1227,N_2701);
or U5329 (N_5329,N_2157,N_2543);
or U5330 (N_5330,N_1705,N_689);
nor U5331 (N_5331,N_2932,N_781);
or U5332 (N_5332,N_1585,N_2857);
and U5333 (N_5333,N_620,N_1997);
nand U5334 (N_5334,N_402,N_2297);
or U5335 (N_5335,N_1722,N_420);
nand U5336 (N_5336,N_201,N_2075);
nor U5337 (N_5337,N_2834,N_2604);
or U5338 (N_5338,N_1055,N_629);
nor U5339 (N_5339,N_726,N_1644);
nor U5340 (N_5340,N_2683,N_1616);
nand U5341 (N_5341,N_2733,N_393);
nand U5342 (N_5342,N_2270,N_999);
nand U5343 (N_5343,N_2057,N_2226);
nor U5344 (N_5344,N_1750,N_173);
nor U5345 (N_5345,N_324,N_2980);
and U5346 (N_5346,N_2654,N_205);
nor U5347 (N_5347,N_1139,N_1203);
xor U5348 (N_5348,N_1481,N_1139);
and U5349 (N_5349,N_1767,N_1318);
or U5350 (N_5350,N_1897,N_948);
nor U5351 (N_5351,N_1277,N_1739);
nor U5352 (N_5352,N_1528,N_2675);
nand U5353 (N_5353,N_1495,N_1880);
and U5354 (N_5354,N_1340,N_918);
or U5355 (N_5355,N_2970,N_53);
and U5356 (N_5356,N_518,N_1082);
nor U5357 (N_5357,N_2177,N_2475);
nor U5358 (N_5358,N_1430,N_2330);
nor U5359 (N_5359,N_1360,N_1724);
or U5360 (N_5360,N_481,N_2304);
or U5361 (N_5361,N_1352,N_1317);
or U5362 (N_5362,N_2981,N_1805);
and U5363 (N_5363,N_2295,N_867);
nand U5364 (N_5364,N_1384,N_121);
or U5365 (N_5365,N_2562,N_912);
or U5366 (N_5366,N_660,N_2640);
nand U5367 (N_5367,N_492,N_127);
nor U5368 (N_5368,N_936,N_986);
or U5369 (N_5369,N_1980,N_2049);
and U5370 (N_5370,N_497,N_398);
and U5371 (N_5371,N_1607,N_1294);
or U5372 (N_5372,N_2024,N_668);
nand U5373 (N_5373,N_1406,N_2035);
and U5374 (N_5374,N_292,N_1861);
or U5375 (N_5375,N_181,N_1645);
and U5376 (N_5376,N_811,N_2083);
or U5377 (N_5377,N_456,N_755);
and U5378 (N_5378,N_2399,N_2455);
or U5379 (N_5379,N_1960,N_2303);
nor U5380 (N_5380,N_272,N_1241);
or U5381 (N_5381,N_1093,N_1169);
xor U5382 (N_5382,N_1176,N_2630);
nand U5383 (N_5383,N_947,N_2083);
nand U5384 (N_5384,N_1363,N_1742);
or U5385 (N_5385,N_1789,N_1796);
xnor U5386 (N_5386,N_720,N_2257);
nand U5387 (N_5387,N_1152,N_365);
xor U5388 (N_5388,N_312,N_124);
nand U5389 (N_5389,N_2838,N_313);
nor U5390 (N_5390,N_800,N_2752);
xor U5391 (N_5391,N_2427,N_2989);
nor U5392 (N_5392,N_329,N_1084);
nor U5393 (N_5393,N_2702,N_1232);
xor U5394 (N_5394,N_60,N_2243);
nand U5395 (N_5395,N_1074,N_1894);
or U5396 (N_5396,N_2744,N_2002);
or U5397 (N_5397,N_2945,N_2230);
nand U5398 (N_5398,N_1996,N_2806);
or U5399 (N_5399,N_115,N_2978);
nor U5400 (N_5400,N_279,N_1451);
nand U5401 (N_5401,N_1230,N_2432);
nand U5402 (N_5402,N_1660,N_1730);
nor U5403 (N_5403,N_663,N_477);
nand U5404 (N_5404,N_2896,N_1648);
nand U5405 (N_5405,N_2149,N_935);
nand U5406 (N_5406,N_1809,N_1165);
nand U5407 (N_5407,N_2663,N_1232);
nand U5408 (N_5408,N_2683,N_784);
or U5409 (N_5409,N_31,N_1098);
or U5410 (N_5410,N_1,N_2134);
and U5411 (N_5411,N_641,N_1460);
nor U5412 (N_5412,N_2767,N_574);
nor U5413 (N_5413,N_880,N_1900);
or U5414 (N_5414,N_2681,N_1341);
nand U5415 (N_5415,N_2721,N_2129);
nor U5416 (N_5416,N_1040,N_675);
and U5417 (N_5417,N_2675,N_2904);
or U5418 (N_5418,N_158,N_468);
nor U5419 (N_5419,N_461,N_1028);
nor U5420 (N_5420,N_1868,N_118);
or U5421 (N_5421,N_729,N_1484);
and U5422 (N_5422,N_1303,N_733);
xor U5423 (N_5423,N_1496,N_2741);
nor U5424 (N_5424,N_1001,N_1469);
nand U5425 (N_5425,N_2937,N_158);
nor U5426 (N_5426,N_1761,N_1029);
or U5427 (N_5427,N_2027,N_1690);
and U5428 (N_5428,N_2164,N_1846);
or U5429 (N_5429,N_1728,N_1233);
nand U5430 (N_5430,N_713,N_2663);
nor U5431 (N_5431,N_870,N_2935);
or U5432 (N_5432,N_1915,N_1594);
xor U5433 (N_5433,N_2352,N_2527);
nand U5434 (N_5434,N_179,N_2304);
nor U5435 (N_5435,N_1116,N_1465);
nand U5436 (N_5436,N_2564,N_1229);
nor U5437 (N_5437,N_2028,N_1919);
and U5438 (N_5438,N_1397,N_168);
nand U5439 (N_5439,N_180,N_436);
and U5440 (N_5440,N_416,N_706);
nor U5441 (N_5441,N_309,N_32);
nor U5442 (N_5442,N_1243,N_2161);
or U5443 (N_5443,N_329,N_270);
or U5444 (N_5444,N_128,N_2990);
and U5445 (N_5445,N_1179,N_779);
and U5446 (N_5446,N_339,N_445);
nand U5447 (N_5447,N_557,N_1207);
and U5448 (N_5448,N_787,N_773);
and U5449 (N_5449,N_2668,N_2330);
nor U5450 (N_5450,N_1066,N_1389);
and U5451 (N_5451,N_424,N_2339);
or U5452 (N_5452,N_944,N_685);
or U5453 (N_5453,N_2661,N_1054);
nor U5454 (N_5454,N_381,N_1472);
nor U5455 (N_5455,N_2129,N_2670);
nor U5456 (N_5456,N_2964,N_1658);
nand U5457 (N_5457,N_2921,N_1598);
nand U5458 (N_5458,N_212,N_1912);
nor U5459 (N_5459,N_1426,N_2669);
or U5460 (N_5460,N_1235,N_2350);
and U5461 (N_5461,N_2836,N_1489);
nor U5462 (N_5462,N_1709,N_1739);
or U5463 (N_5463,N_433,N_1493);
or U5464 (N_5464,N_2257,N_2071);
or U5465 (N_5465,N_1521,N_176);
nand U5466 (N_5466,N_268,N_810);
or U5467 (N_5467,N_2398,N_2213);
or U5468 (N_5468,N_1992,N_1133);
and U5469 (N_5469,N_927,N_2320);
and U5470 (N_5470,N_1165,N_1381);
nand U5471 (N_5471,N_1396,N_1409);
or U5472 (N_5472,N_134,N_1584);
and U5473 (N_5473,N_2819,N_2832);
nand U5474 (N_5474,N_2223,N_1584);
nand U5475 (N_5475,N_2414,N_1390);
and U5476 (N_5476,N_2465,N_1805);
nor U5477 (N_5477,N_742,N_2968);
nand U5478 (N_5478,N_705,N_2931);
or U5479 (N_5479,N_2251,N_2120);
and U5480 (N_5480,N_2645,N_1916);
or U5481 (N_5481,N_62,N_949);
and U5482 (N_5482,N_1580,N_1707);
and U5483 (N_5483,N_1766,N_199);
or U5484 (N_5484,N_1694,N_1954);
and U5485 (N_5485,N_661,N_2939);
nor U5486 (N_5486,N_1347,N_929);
xnor U5487 (N_5487,N_2510,N_2233);
and U5488 (N_5488,N_2603,N_2037);
nor U5489 (N_5489,N_2298,N_79);
and U5490 (N_5490,N_2462,N_1681);
or U5491 (N_5491,N_509,N_1953);
nand U5492 (N_5492,N_1696,N_1717);
or U5493 (N_5493,N_2831,N_610);
and U5494 (N_5494,N_2392,N_536);
nand U5495 (N_5495,N_145,N_1830);
or U5496 (N_5496,N_680,N_2495);
or U5497 (N_5497,N_357,N_1974);
nor U5498 (N_5498,N_2352,N_263);
nand U5499 (N_5499,N_1601,N_1512);
nor U5500 (N_5500,N_2136,N_712);
or U5501 (N_5501,N_14,N_552);
and U5502 (N_5502,N_2407,N_919);
nor U5503 (N_5503,N_2267,N_1194);
and U5504 (N_5504,N_2835,N_1446);
nor U5505 (N_5505,N_21,N_1977);
or U5506 (N_5506,N_1604,N_2300);
nor U5507 (N_5507,N_890,N_1949);
nand U5508 (N_5508,N_2864,N_1978);
and U5509 (N_5509,N_2643,N_206);
or U5510 (N_5510,N_1041,N_983);
nand U5511 (N_5511,N_1893,N_2950);
nor U5512 (N_5512,N_2191,N_1604);
or U5513 (N_5513,N_1186,N_841);
nor U5514 (N_5514,N_2875,N_1671);
and U5515 (N_5515,N_2887,N_1195);
nand U5516 (N_5516,N_2160,N_2813);
nor U5517 (N_5517,N_1102,N_314);
nor U5518 (N_5518,N_1019,N_1212);
xor U5519 (N_5519,N_2123,N_51);
and U5520 (N_5520,N_1010,N_671);
nor U5521 (N_5521,N_468,N_1181);
or U5522 (N_5522,N_2205,N_2377);
nand U5523 (N_5523,N_2063,N_7);
and U5524 (N_5524,N_1917,N_1276);
nand U5525 (N_5525,N_1986,N_1116);
nor U5526 (N_5526,N_236,N_27);
and U5527 (N_5527,N_1364,N_2480);
nor U5528 (N_5528,N_37,N_1924);
nand U5529 (N_5529,N_2008,N_17);
nor U5530 (N_5530,N_2871,N_2279);
nor U5531 (N_5531,N_1816,N_2635);
nor U5532 (N_5532,N_2808,N_2144);
and U5533 (N_5533,N_2868,N_2809);
nor U5534 (N_5534,N_1505,N_1728);
nor U5535 (N_5535,N_2964,N_164);
xor U5536 (N_5536,N_1622,N_2549);
nand U5537 (N_5537,N_2242,N_2098);
nor U5538 (N_5538,N_284,N_2159);
nor U5539 (N_5539,N_2207,N_681);
and U5540 (N_5540,N_955,N_2065);
and U5541 (N_5541,N_1396,N_322);
and U5542 (N_5542,N_2615,N_1948);
nor U5543 (N_5543,N_1979,N_1136);
nor U5544 (N_5544,N_2549,N_2478);
and U5545 (N_5545,N_1003,N_1754);
nand U5546 (N_5546,N_961,N_1182);
and U5547 (N_5547,N_1679,N_364);
or U5548 (N_5548,N_116,N_474);
and U5549 (N_5549,N_667,N_2644);
nand U5550 (N_5550,N_2353,N_494);
nand U5551 (N_5551,N_1378,N_2596);
nand U5552 (N_5552,N_2300,N_2668);
nand U5553 (N_5553,N_972,N_579);
nand U5554 (N_5554,N_198,N_2825);
nor U5555 (N_5555,N_2548,N_2315);
and U5556 (N_5556,N_256,N_2622);
and U5557 (N_5557,N_678,N_2800);
and U5558 (N_5558,N_1831,N_1528);
or U5559 (N_5559,N_1231,N_2670);
or U5560 (N_5560,N_2216,N_2980);
nand U5561 (N_5561,N_649,N_658);
nor U5562 (N_5562,N_88,N_1649);
or U5563 (N_5563,N_1283,N_2387);
nor U5564 (N_5564,N_877,N_2311);
xor U5565 (N_5565,N_826,N_1124);
or U5566 (N_5566,N_2711,N_2940);
nor U5567 (N_5567,N_1066,N_2405);
nor U5568 (N_5568,N_2409,N_612);
or U5569 (N_5569,N_1785,N_541);
or U5570 (N_5570,N_657,N_129);
nor U5571 (N_5571,N_1590,N_122);
nor U5572 (N_5572,N_1890,N_2031);
or U5573 (N_5573,N_524,N_2602);
or U5574 (N_5574,N_153,N_70);
or U5575 (N_5575,N_2769,N_1520);
or U5576 (N_5576,N_1680,N_2244);
nand U5577 (N_5577,N_207,N_1744);
and U5578 (N_5578,N_2623,N_393);
or U5579 (N_5579,N_1599,N_2428);
nand U5580 (N_5580,N_2978,N_5);
nor U5581 (N_5581,N_1380,N_1038);
nor U5582 (N_5582,N_2268,N_2135);
and U5583 (N_5583,N_1741,N_684);
nand U5584 (N_5584,N_2162,N_2987);
or U5585 (N_5585,N_2260,N_2725);
and U5586 (N_5586,N_1454,N_1308);
and U5587 (N_5587,N_104,N_1654);
or U5588 (N_5588,N_128,N_1388);
or U5589 (N_5589,N_1624,N_1089);
nand U5590 (N_5590,N_1785,N_2488);
nor U5591 (N_5591,N_1132,N_2923);
nand U5592 (N_5592,N_112,N_526);
nor U5593 (N_5593,N_589,N_2771);
nor U5594 (N_5594,N_1519,N_116);
or U5595 (N_5595,N_1434,N_573);
nor U5596 (N_5596,N_1741,N_829);
nand U5597 (N_5597,N_1045,N_2219);
nor U5598 (N_5598,N_2510,N_299);
nor U5599 (N_5599,N_1500,N_1902);
or U5600 (N_5600,N_2210,N_2157);
nand U5601 (N_5601,N_76,N_1003);
or U5602 (N_5602,N_2922,N_172);
xnor U5603 (N_5603,N_2145,N_1657);
or U5604 (N_5604,N_1901,N_423);
or U5605 (N_5605,N_341,N_1469);
xnor U5606 (N_5606,N_2066,N_1403);
and U5607 (N_5607,N_1684,N_2220);
nor U5608 (N_5608,N_2085,N_363);
nor U5609 (N_5609,N_2687,N_695);
or U5610 (N_5610,N_907,N_879);
nor U5611 (N_5611,N_1430,N_1106);
nor U5612 (N_5612,N_605,N_1314);
and U5613 (N_5613,N_1026,N_2443);
nor U5614 (N_5614,N_940,N_2893);
nand U5615 (N_5615,N_54,N_1573);
nand U5616 (N_5616,N_1324,N_1535);
nand U5617 (N_5617,N_1128,N_601);
xor U5618 (N_5618,N_2866,N_2436);
or U5619 (N_5619,N_1984,N_2252);
nand U5620 (N_5620,N_1524,N_1422);
nand U5621 (N_5621,N_2891,N_2590);
and U5622 (N_5622,N_2904,N_452);
nand U5623 (N_5623,N_1602,N_1633);
or U5624 (N_5624,N_1472,N_1623);
and U5625 (N_5625,N_1850,N_2434);
nand U5626 (N_5626,N_1999,N_1381);
nor U5627 (N_5627,N_2695,N_757);
and U5628 (N_5628,N_30,N_1910);
and U5629 (N_5629,N_455,N_529);
and U5630 (N_5630,N_872,N_1467);
or U5631 (N_5631,N_1109,N_2835);
nor U5632 (N_5632,N_2325,N_1291);
and U5633 (N_5633,N_2131,N_1550);
nor U5634 (N_5634,N_1421,N_121);
nand U5635 (N_5635,N_1174,N_211);
or U5636 (N_5636,N_2674,N_228);
and U5637 (N_5637,N_2588,N_788);
nand U5638 (N_5638,N_570,N_1957);
and U5639 (N_5639,N_2090,N_1197);
nand U5640 (N_5640,N_527,N_678);
or U5641 (N_5641,N_1637,N_72);
nand U5642 (N_5642,N_216,N_2047);
nand U5643 (N_5643,N_426,N_1678);
and U5644 (N_5644,N_1992,N_1917);
or U5645 (N_5645,N_2738,N_319);
and U5646 (N_5646,N_761,N_2244);
nand U5647 (N_5647,N_1705,N_1190);
and U5648 (N_5648,N_1190,N_2065);
nand U5649 (N_5649,N_2167,N_2091);
nand U5650 (N_5650,N_2300,N_586);
and U5651 (N_5651,N_605,N_1304);
nor U5652 (N_5652,N_444,N_572);
or U5653 (N_5653,N_727,N_2533);
nand U5654 (N_5654,N_2938,N_361);
nor U5655 (N_5655,N_1321,N_2160);
or U5656 (N_5656,N_2079,N_268);
or U5657 (N_5657,N_1048,N_1322);
and U5658 (N_5658,N_2274,N_830);
and U5659 (N_5659,N_196,N_21);
nor U5660 (N_5660,N_154,N_1358);
or U5661 (N_5661,N_1576,N_2788);
and U5662 (N_5662,N_2756,N_292);
and U5663 (N_5663,N_34,N_1787);
and U5664 (N_5664,N_860,N_244);
or U5665 (N_5665,N_1531,N_2694);
and U5666 (N_5666,N_2489,N_1814);
or U5667 (N_5667,N_600,N_2887);
or U5668 (N_5668,N_1911,N_1480);
nor U5669 (N_5669,N_1676,N_49);
xnor U5670 (N_5670,N_1677,N_1907);
and U5671 (N_5671,N_1287,N_1035);
nor U5672 (N_5672,N_1582,N_2295);
or U5673 (N_5673,N_747,N_2466);
nand U5674 (N_5674,N_710,N_2831);
or U5675 (N_5675,N_479,N_1658);
or U5676 (N_5676,N_216,N_1677);
nor U5677 (N_5677,N_1182,N_1543);
and U5678 (N_5678,N_1797,N_604);
nand U5679 (N_5679,N_1543,N_2197);
and U5680 (N_5680,N_1449,N_1182);
nor U5681 (N_5681,N_1447,N_279);
nor U5682 (N_5682,N_2510,N_1461);
and U5683 (N_5683,N_216,N_1362);
or U5684 (N_5684,N_2296,N_2386);
xnor U5685 (N_5685,N_2001,N_2493);
nand U5686 (N_5686,N_2091,N_1659);
nor U5687 (N_5687,N_1798,N_1992);
or U5688 (N_5688,N_2399,N_156);
or U5689 (N_5689,N_452,N_2714);
nor U5690 (N_5690,N_2658,N_107);
nor U5691 (N_5691,N_693,N_2151);
and U5692 (N_5692,N_1317,N_867);
nand U5693 (N_5693,N_321,N_1942);
and U5694 (N_5694,N_2926,N_2762);
nor U5695 (N_5695,N_806,N_1202);
nor U5696 (N_5696,N_734,N_93);
and U5697 (N_5697,N_2397,N_196);
or U5698 (N_5698,N_635,N_2311);
nor U5699 (N_5699,N_2891,N_2484);
and U5700 (N_5700,N_1647,N_2930);
and U5701 (N_5701,N_1464,N_1793);
or U5702 (N_5702,N_857,N_2427);
and U5703 (N_5703,N_2727,N_1569);
nand U5704 (N_5704,N_2547,N_426);
or U5705 (N_5705,N_2262,N_554);
nor U5706 (N_5706,N_464,N_2411);
or U5707 (N_5707,N_253,N_1854);
or U5708 (N_5708,N_119,N_1380);
nor U5709 (N_5709,N_773,N_1057);
and U5710 (N_5710,N_458,N_1551);
or U5711 (N_5711,N_1203,N_1348);
or U5712 (N_5712,N_396,N_2157);
and U5713 (N_5713,N_399,N_1610);
and U5714 (N_5714,N_2421,N_2440);
xnor U5715 (N_5715,N_1383,N_615);
or U5716 (N_5716,N_1837,N_2040);
and U5717 (N_5717,N_181,N_1584);
and U5718 (N_5718,N_1926,N_2015);
nor U5719 (N_5719,N_2936,N_1245);
nor U5720 (N_5720,N_2458,N_357);
nor U5721 (N_5721,N_1202,N_834);
or U5722 (N_5722,N_2964,N_1742);
or U5723 (N_5723,N_837,N_1351);
nand U5724 (N_5724,N_2403,N_2877);
xor U5725 (N_5725,N_2873,N_1037);
nor U5726 (N_5726,N_2139,N_2738);
nor U5727 (N_5727,N_777,N_514);
nor U5728 (N_5728,N_974,N_108);
and U5729 (N_5729,N_879,N_1551);
xnor U5730 (N_5730,N_2881,N_627);
nor U5731 (N_5731,N_579,N_555);
nand U5732 (N_5732,N_2051,N_1661);
nand U5733 (N_5733,N_2288,N_2211);
nand U5734 (N_5734,N_1369,N_562);
nand U5735 (N_5735,N_1453,N_1786);
and U5736 (N_5736,N_1740,N_314);
or U5737 (N_5737,N_2922,N_563);
and U5738 (N_5738,N_2485,N_2772);
and U5739 (N_5739,N_2097,N_918);
and U5740 (N_5740,N_1851,N_375);
or U5741 (N_5741,N_1212,N_244);
nand U5742 (N_5742,N_1565,N_1139);
nand U5743 (N_5743,N_1766,N_2885);
nand U5744 (N_5744,N_1619,N_2715);
or U5745 (N_5745,N_2314,N_527);
or U5746 (N_5746,N_635,N_2248);
and U5747 (N_5747,N_1653,N_132);
and U5748 (N_5748,N_1168,N_2535);
or U5749 (N_5749,N_1406,N_856);
or U5750 (N_5750,N_2433,N_694);
or U5751 (N_5751,N_85,N_1326);
or U5752 (N_5752,N_1118,N_1789);
nor U5753 (N_5753,N_1919,N_437);
nand U5754 (N_5754,N_1824,N_262);
and U5755 (N_5755,N_301,N_190);
and U5756 (N_5756,N_987,N_1828);
and U5757 (N_5757,N_1697,N_1647);
nand U5758 (N_5758,N_749,N_2421);
or U5759 (N_5759,N_2310,N_333);
nand U5760 (N_5760,N_1743,N_1010);
nor U5761 (N_5761,N_1,N_465);
nor U5762 (N_5762,N_695,N_2627);
or U5763 (N_5763,N_1199,N_2234);
or U5764 (N_5764,N_1665,N_2957);
nand U5765 (N_5765,N_513,N_2513);
nor U5766 (N_5766,N_266,N_79);
and U5767 (N_5767,N_2176,N_133);
nor U5768 (N_5768,N_1098,N_2638);
and U5769 (N_5769,N_1797,N_782);
nand U5770 (N_5770,N_116,N_2318);
or U5771 (N_5771,N_1874,N_979);
nor U5772 (N_5772,N_2602,N_2869);
nand U5773 (N_5773,N_958,N_1178);
or U5774 (N_5774,N_1141,N_346);
nand U5775 (N_5775,N_432,N_681);
and U5776 (N_5776,N_628,N_949);
or U5777 (N_5777,N_2852,N_1723);
and U5778 (N_5778,N_2714,N_2175);
and U5779 (N_5779,N_2291,N_344);
nor U5780 (N_5780,N_276,N_2834);
and U5781 (N_5781,N_268,N_920);
or U5782 (N_5782,N_2156,N_2542);
nor U5783 (N_5783,N_1467,N_2170);
nand U5784 (N_5784,N_2175,N_1173);
nand U5785 (N_5785,N_2771,N_1598);
nor U5786 (N_5786,N_754,N_687);
or U5787 (N_5787,N_997,N_2887);
nand U5788 (N_5788,N_355,N_1843);
or U5789 (N_5789,N_2146,N_2429);
or U5790 (N_5790,N_1389,N_638);
nand U5791 (N_5791,N_272,N_2998);
and U5792 (N_5792,N_1649,N_1370);
nand U5793 (N_5793,N_223,N_2906);
or U5794 (N_5794,N_533,N_1903);
nor U5795 (N_5795,N_1164,N_332);
nor U5796 (N_5796,N_1709,N_92);
and U5797 (N_5797,N_1375,N_410);
and U5798 (N_5798,N_2603,N_340);
or U5799 (N_5799,N_2059,N_1194);
and U5800 (N_5800,N_1690,N_717);
nor U5801 (N_5801,N_1034,N_1452);
or U5802 (N_5802,N_2365,N_1681);
nor U5803 (N_5803,N_336,N_953);
nand U5804 (N_5804,N_1448,N_2270);
nand U5805 (N_5805,N_188,N_178);
nor U5806 (N_5806,N_2558,N_2970);
or U5807 (N_5807,N_1307,N_2399);
or U5808 (N_5808,N_2281,N_841);
nor U5809 (N_5809,N_2738,N_1127);
nor U5810 (N_5810,N_1936,N_1544);
and U5811 (N_5811,N_2361,N_1177);
nor U5812 (N_5812,N_1812,N_2692);
nand U5813 (N_5813,N_1594,N_1753);
nor U5814 (N_5814,N_153,N_851);
or U5815 (N_5815,N_1800,N_322);
or U5816 (N_5816,N_2738,N_2295);
nor U5817 (N_5817,N_1281,N_486);
nor U5818 (N_5818,N_1850,N_2582);
nor U5819 (N_5819,N_690,N_1831);
xor U5820 (N_5820,N_910,N_604);
and U5821 (N_5821,N_1400,N_2258);
and U5822 (N_5822,N_2774,N_2969);
and U5823 (N_5823,N_1289,N_1278);
nor U5824 (N_5824,N_1067,N_1788);
and U5825 (N_5825,N_2240,N_653);
and U5826 (N_5826,N_1004,N_1907);
or U5827 (N_5827,N_2946,N_2852);
or U5828 (N_5828,N_1085,N_1989);
nor U5829 (N_5829,N_910,N_2892);
nor U5830 (N_5830,N_772,N_2567);
and U5831 (N_5831,N_595,N_2788);
or U5832 (N_5832,N_1768,N_1504);
and U5833 (N_5833,N_1594,N_1917);
nor U5834 (N_5834,N_297,N_2746);
and U5835 (N_5835,N_350,N_2455);
nor U5836 (N_5836,N_611,N_2233);
nor U5837 (N_5837,N_2382,N_612);
nand U5838 (N_5838,N_663,N_770);
or U5839 (N_5839,N_424,N_281);
nor U5840 (N_5840,N_1602,N_733);
xnor U5841 (N_5841,N_578,N_2227);
nand U5842 (N_5842,N_198,N_1599);
or U5843 (N_5843,N_1854,N_660);
or U5844 (N_5844,N_51,N_2388);
and U5845 (N_5845,N_2945,N_782);
nand U5846 (N_5846,N_1921,N_883);
and U5847 (N_5847,N_733,N_2929);
nor U5848 (N_5848,N_1095,N_807);
or U5849 (N_5849,N_209,N_564);
and U5850 (N_5850,N_1901,N_1304);
or U5851 (N_5851,N_2077,N_2540);
nand U5852 (N_5852,N_761,N_136);
and U5853 (N_5853,N_1307,N_2820);
or U5854 (N_5854,N_1482,N_888);
nor U5855 (N_5855,N_2296,N_2314);
nor U5856 (N_5856,N_537,N_2638);
nand U5857 (N_5857,N_2072,N_1264);
or U5858 (N_5858,N_1702,N_1790);
nand U5859 (N_5859,N_1512,N_412);
or U5860 (N_5860,N_324,N_2204);
and U5861 (N_5861,N_1333,N_1302);
and U5862 (N_5862,N_960,N_271);
or U5863 (N_5863,N_1042,N_2402);
nand U5864 (N_5864,N_918,N_1300);
nor U5865 (N_5865,N_2871,N_2232);
nor U5866 (N_5866,N_2329,N_2735);
or U5867 (N_5867,N_616,N_1210);
nand U5868 (N_5868,N_2950,N_645);
and U5869 (N_5869,N_87,N_2873);
and U5870 (N_5870,N_2253,N_626);
or U5871 (N_5871,N_2059,N_2252);
or U5872 (N_5872,N_979,N_1015);
and U5873 (N_5873,N_2962,N_1978);
nor U5874 (N_5874,N_1138,N_1773);
nand U5875 (N_5875,N_682,N_1995);
nand U5876 (N_5876,N_725,N_430);
nand U5877 (N_5877,N_1571,N_2174);
or U5878 (N_5878,N_2578,N_2084);
nor U5879 (N_5879,N_1189,N_2318);
or U5880 (N_5880,N_2830,N_1409);
and U5881 (N_5881,N_2701,N_1271);
nor U5882 (N_5882,N_1918,N_359);
nand U5883 (N_5883,N_2497,N_1928);
xor U5884 (N_5884,N_1111,N_1214);
nor U5885 (N_5885,N_18,N_2866);
and U5886 (N_5886,N_1501,N_666);
nand U5887 (N_5887,N_508,N_916);
and U5888 (N_5888,N_1566,N_712);
nor U5889 (N_5889,N_2485,N_1774);
nand U5890 (N_5890,N_2197,N_741);
and U5891 (N_5891,N_2286,N_1163);
and U5892 (N_5892,N_1854,N_2610);
nor U5893 (N_5893,N_773,N_1084);
nand U5894 (N_5894,N_2802,N_1616);
or U5895 (N_5895,N_2905,N_2512);
and U5896 (N_5896,N_1245,N_2526);
nor U5897 (N_5897,N_2094,N_1930);
and U5898 (N_5898,N_2707,N_678);
nor U5899 (N_5899,N_2005,N_824);
nand U5900 (N_5900,N_1340,N_596);
and U5901 (N_5901,N_2435,N_2809);
and U5902 (N_5902,N_2806,N_1363);
nor U5903 (N_5903,N_1521,N_1057);
xor U5904 (N_5904,N_635,N_2255);
nor U5905 (N_5905,N_1607,N_1054);
nand U5906 (N_5906,N_2238,N_2158);
nand U5907 (N_5907,N_792,N_1575);
xnor U5908 (N_5908,N_1066,N_790);
or U5909 (N_5909,N_1396,N_783);
nand U5910 (N_5910,N_2756,N_1126);
or U5911 (N_5911,N_364,N_339);
nand U5912 (N_5912,N_428,N_2474);
or U5913 (N_5913,N_839,N_1504);
or U5914 (N_5914,N_2577,N_1492);
or U5915 (N_5915,N_433,N_2237);
nand U5916 (N_5916,N_1477,N_285);
or U5917 (N_5917,N_646,N_1596);
nand U5918 (N_5918,N_1354,N_1659);
nand U5919 (N_5919,N_2935,N_1574);
or U5920 (N_5920,N_328,N_458);
or U5921 (N_5921,N_1881,N_106);
nor U5922 (N_5922,N_2979,N_2392);
nor U5923 (N_5923,N_201,N_1138);
and U5924 (N_5924,N_1806,N_2897);
nor U5925 (N_5925,N_446,N_2177);
or U5926 (N_5926,N_2935,N_2326);
and U5927 (N_5927,N_2191,N_58);
nor U5928 (N_5928,N_2,N_1089);
and U5929 (N_5929,N_2203,N_2560);
nand U5930 (N_5930,N_747,N_928);
or U5931 (N_5931,N_1862,N_1263);
nor U5932 (N_5932,N_2116,N_2298);
and U5933 (N_5933,N_98,N_1428);
nand U5934 (N_5934,N_2743,N_2333);
nor U5935 (N_5935,N_1722,N_520);
and U5936 (N_5936,N_2061,N_617);
or U5937 (N_5937,N_597,N_972);
and U5938 (N_5938,N_1982,N_1899);
nor U5939 (N_5939,N_2675,N_1356);
and U5940 (N_5940,N_1496,N_2532);
nand U5941 (N_5941,N_1415,N_977);
or U5942 (N_5942,N_1817,N_1303);
nor U5943 (N_5943,N_2274,N_435);
nor U5944 (N_5944,N_1216,N_606);
or U5945 (N_5945,N_1397,N_1663);
nand U5946 (N_5946,N_619,N_2801);
nand U5947 (N_5947,N_2204,N_408);
nor U5948 (N_5948,N_2340,N_2152);
nor U5949 (N_5949,N_2768,N_863);
nand U5950 (N_5950,N_2728,N_271);
or U5951 (N_5951,N_85,N_2133);
or U5952 (N_5952,N_389,N_331);
nor U5953 (N_5953,N_1696,N_1038);
and U5954 (N_5954,N_2462,N_1516);
nand U5955 (N_5955,N_2503,N_593);
or U5956 (N_5956,N_2487,N_1945);
or U5957 (N_5957,N_481,N_303);
nand U5958 (N_5958,N_770,N_305);
and U5959 (N_5959,N_2318,N_1141);
nor U5960 (N_5960,N_45,N_723);
nor U5961 (N_5961,N_607,N_2377);
nand U5962 (N_5962,N_2132,N_2294);
or U5963 (N_5963,N_520,N_2002);
or U5964 (N_5964,N_138,N_894);
or U5965 (N_5965,N_1662,N_2181);
and U5966 (N_5966,N_1469,N_1733);
nand U5967 (N_5967,N_1428,N_1051);
nor U5968 (N_5968,N_1288,N_774);
and U5969 (N_5969,N_247,N_305);
nor U5970 (N_5970,N_1792,N_2857);
and U5971 (N_5971,N_2398,N_2528);
or U5972 (N_5972,N_7,N_1856);
nand U5973 (N_5973,N_2553,N_1068);
nor U5974 (N_5974,N_731,N_2810);
nor U5975 (N_5975,N_2412,N_986);
xor U5976 (N_5976,N_2362,N_1230);
or U5977 (N_5977,N_2164,N_1748);
xnor U5978 (N_5978,N_1020,N_1966);
or U5979 (N_5979,N_1836,N_447);
or U5980 (N_5980,N_1913,N_467);
and U5981 (N_5981,N_631,N_663);
nor U5982 (N_5982,N_1627,N_2599);
or U5983 (N_5983,N_2818,N_2965);
nor U5984 (N_5984,N_2474,N_765);
nand U5985 (N_5985,N_827,N_2365);
or U5986 (N_5986,N_2629,N_2258);
or U5987 (N_5987,N_2269,N_1438);
and U5988 (N_5988,N_478,N_2516);
or U5989 (N_5989,N_1209,N_2362);
or U5990 (N_5990,N_2428,N_296);
nor U5991 (N_5991,N_2759,N_579);
nand U5992 (N_5992,N_2212,N_2022);
or U5993 (N_5993,N_472,N_2596);
nor U5994 (N_5994,N_645,N_2193);
nor U5995 (N_5995,N_522,N_1041);
nor U5996 (N_5996,N_2787,N_2507);
or U5997 (N_5997,N_1605,N_34);
nor U5998 (N_5998,N_2801,N_1164);
nand U5999 (N_5999,N_2988,N_1781);
or U6000 (N_6000,N_4725,N_5641);
or U6001 (N_6001,N_5517,N_3347);
and U6002 (N_6002,N_4128,N_4139);
and U6003 (N_6003,N_4205,N_4608);
or U6004 (N_6004,N_3815,N_5779);
and U6005 (N_6005,N_4285,N_4635);
or U6006 (N_6006,N_3092,N_5362);
or U6007 (N_6007,N_3318,N_5745);
or U6008 (N_6008,N_4540,N_4632);
or U6009 (N_6009,N_3247,N_3584);
nand U6010 (N_6010,N_4743,N_4880);
or U6011 (N_6011,N_3337,N_3252);
nor U6012 (N_6012,N_5079,N_3180);
nand U6013 (N_6013,N_3805,N_5558);
and U6014 (N_6014,N_4012,N_5173);
or U6015 (N_6015,N_3690,N_3233);
nand U6016 (N_6016,N_4127,N_4685);
nand U6017 (N_6017,N_4583,N_5848);
nand U6018 (N_6018,N_3866,N_5029);
and U6019 (N_6019,N_4223,N_5816);
or U6020 (N_6020,N_5952,N_4078);
nor U6021 (N_6021,N_4652,N_3873);
nor U6022 (N_6022,N_3073,N_5014);
or U6023 (N_6023,N_3622,N_3679);
or U6024 (N_6024,N_5306,N_3406);
and U6025 (N_6025,N_4852,N_5936);
or U6026 (N_6026,N_3278,N_5752);
nand U6027 (N_6027,N_4301,N_3552);
nor U6028 (N_6028,N_5453,N_4544);
and U6029 (N_6029,N_4947,N_4516);
and U6030 (N_6030,N_4912,N_4911);
or U6031 (N_6031,N_5751,N_3658);
or U6032 (N_6032,N_3362,N_3245);
or U6033 (N_6033,N_4850,N_4614);
or U6034 (N_6034,N_3328,N_5750);
and U6035 (N_6035,N_3917,N_3508);
and U6036 (N_6036,N_4024,N_3382);
nand U6037 (N_6037,N_3042,N_4167);
and U6038 (N_6038,N_3141,N_4750);
or U6039 (N_6039,N_4797,N_4288);
nor U6040 (N_6040,N_4539,N_3413);
nor U6041 (N_6041,N_4392,N_4768);
or U6042 (N_6042,N_5591,N_5769);
and U6043 (N_6043,N_4791,N_5513);
nor U6044 (N_6044,N_3032,N_5922);
nor U6045 (N_6045,N_3848,N_5499);
nor U6046 (N_6046,N_5086,N_4792);
nor U6047 (N_6047,N_5676,N_3155);
or U6048 (N_6048,N_4184,N_5589);
and U6049 (N_6049,N_4869,N_3862);
and U6050 (N_6050,N_5077,N_5804);
nand U6051 (N_6051,N_4393,N_4469);
or U6052 (N_6052,N_3923,N_3545);
nor U6053 (N_6053,N_4551,N_5802);
or U6054 (N_6054,N_4359,N_4065);
or U6055 (N_6055,N_5340,N_4385);
or U6056 (N_6056,N_3230,N_3087);
nand U6057 (N_6057,N_4093,N_4588);
and U6058 (N_6058,N_3446,N_4915);
nand U6059 (N_6059,N_5342,N_3633);
nand U6060 (N_6060,N_4851,N_5935);
or U6061 (N_6061,N_4124,N_4038);
and U6062 (N_6062,N_4700,N_3320);
nand U6063 (N_6063,N_4709,N_3701);
nor U6064 (N_6064,N_3438,N_4194);
nor U6065 (N_6065,N_4620,N_5372);
or U6066 (N_6066,N_3225,N_3922);
or U6067 (N_6067,N_5934,N_3104);
nand U6068 (N_6068,N_5376,N_5593);
and U6069 (N_6069,N_5179,N_3309);
or U6070 (N_6070,N_4278,N_4962);
and U6071 (N_6071,N_5455,N_3525);
and U6072 (N_6072,N_5442,N_3392);
nand U6073 (N_6073,N_5711,N_3389);
and U6074 (N_6074,N_4819,N_5949);
and U6075 (N_6075,N_4906,N_5617);
or U6076 (N_6076,N_3015,N_5056);
xnor U6077 (N_6077,N_4363,N_3736);
nor U6078 (N_6078,N_4156,N_4858);
and U6079 (N_6079,N_5776,N_4818);
nor U6080 (N_6080,N_3538,N_5845);
and U6081 (N_6081,N_5681,N_4970);
or U6082 (N_6082,N_5326,N_5231);
and U6083 (N_6083,N_3174,N_3581);
and U6084 (N_6084,N_3031,N_4413);
or U6085 (N_6085,N_3644,N_3513);
and U6086 (N_6086,N_4997,N_3297);
nor U6087 (N_6087,N_3147,N_3807);
or U6088 (N_6088,N_3789,N_4802);
or U6089 (N_6089,N_5140,N_3900);
and U6090 (N_6090,N_4816,N_5904);
nor U6091 (N_6091,N_5467,N_5383);
and U6092 (N_6092,N_5397,N_5293);
or U6093 (N_6093,N_5002,N_5070);
nor U6094 (N_6094,N_5898,N_4905);
nand U6095 (N_6095,N_3181,N_3550);
nor U6096 (N_6096,N_3137,N_5803);
or U6097 (N_6097,N_3083,N_5206);
nand U6098 (N_6098,N_5956,N_5859);
and U6099 (N_6099,N_4414,N_4887);
nand U6100 (N_6100,N_5735,N_5118);
nand U6101 (N_6101,N_5006,N_4875);
and U6102 (N_6102,N_5434,N_3340);
nand U6103 (N_6103,N_4200,N_3070);
nand U6104 (N_6104,N_5043,N_4210);
or U6105 (N_6105,N_5401,N_5894);
and U6106 (N_6106,N_4129,N_4310);
and U6107 (N_6107,N_3030,N_3925);
nor U6108 (N_6108,N_4087,N_3836);
nand U6109 (N_6109,N_3416,N_4164);
and U6110 (N_6110,N_3840,N_5855);
nor U6111 (N_6111,N_3455,N_4737);
and U6112 (N_6112,N_4216,N_3645);
or U6113 (N_6113,N_4444,N_5095);
nand U6114 (N_6114,N_3270,N_4463);
xor U6115 (N_6115,N_3727,N_5198);
nand U6116 (N_6116,N_4581,N_4309);
nand U6117 (N_6117,N_3169,N_3852);
or U6118 (N_6118,N_4846,N_3440);
nand U6119 (N_6119,N_4121,N_4389);
or U6120 (N_6120,N_4396,N_4621);
nor U6121 (N_6121,N_4192,N_5984);
or U6122 (N_6122,N_4681,N_3891);
nor U6123 (N_6123,N_5626,N_3672);
or U6124 (N_6124,N_4215,N_5970);
nand U6125 (N_6125,N_4881,N_5102);
nor U6126 (N_6126,N_5169,N_4909);
and U6127 (N_6127,N_5396,N_3964);
nor U6128 (N_6128,N_5721,N_3966);
nand U6129 (N_6129,N_3706,N_4716);
nand U6130 (N_6130,N_3419,N_4021);
nor U6131 (N_6131,N_4094,N_5512);
and U6132 (N_6132,N_3534,N_4611);
nor U6133 (N_6133,N_3623,N_5780);
nand U6134 (N_6134,N_4370,N_5287);
or U6135 (N_6135,N_4160,N_4233);
nand U6136 (N_6136,N_3001,N_5562);
or U6137 (N_6137,N_4580,N_3609);
nor U6138 (N_6138,N_3681,N_3175);
nor U6139 (N_6139,N_3962,N_4415);
or U6140 (N_6140,N_5852,N_3612);
and U6141 (N_6141,N_3144,N_5618);
nor U6142 (N_6142,N_4193,N_3774);
or U6143 (N_6143,N_3604,N_5621);
or U6144 (N_6144,N_3729,N_5121);
or U6145 (N_6145,N_3956,N_4573);
and U6146 (N_6146,N_4361,N_4597);
nand U6147 (N_6147,N_3481,N_5725);
nand U6148 (N_6148,N_5682,N_4558);
or U6149 (N_6149,N_3259,N_5219);
and U6150 (N_6150,N_5565,N_3772);
and U6151 (N_6151,N_4933,N_4826);
or U6152 (N_6152,N_3102,N_4493);
or U6153 (N_6153,N_3049,N_5724);
and U6154 (N_6154,N_4943,N_4960);
and U6155 (N_6155,N_3152,N_5114);
nand U6156 (N_6156,N_3817,N_5472);
and U6157 (N_6157,N_5609,N_4062);
or U6158 (N_6158,N_4762,N_4648);
or U6159 (N_6159,N_5315,N_4830);
nor U6160 (N_6160,N_5851,N_3022);
nor U6161 (N_6161,N_4694,N_4232);
or U6162 (N_6162,N_4541,N_3091);
and U6163 (N_6163,N_4538,N_4372);
nor U6164 (N_6164,N_3076,N_4805);
and U6165 (N_6165,N_4060,N_5947);
and U6166 (N_6166,N_3506,N_3096);
nor U6167 (N_6167,N_3248,N_3546);
nand U6168 (N_6168,N_4290,N_3881);
nand U6169 (N_6169,N_5433,N_4394);
nor U6170 (N_6170,N_4458,N_3308);
nor U6171 (N_6171,N_5348,N_5263);
nand U6172 (N_6172,N_3920,N_5932);
nand U6173 (N_6173,N_5085,N_4665);
or U6174 (N_6174,N_3822,N_5792);
and U6175 (N_6175,N_5013,N_5036);
or U6176 (N_6176,N_4847,N_4522);
nand U6177 (N_6177,N_3627,N_3196);
nand U6178 (N_6178,N_5182,N_5388);
or U6179 (N_6179,N_3116,N_4923);
nor U6180 (N_6180,N_3423,N_5216);
nor U6181 (N_6181,N_4657,N_5252);
nand U6182 (N_6182,N_5463,N_5945);
or U6183 (N_6183,N_5475,N_4462);
xor U6184 (N_6184,N_5946,N_4170);
nor U6185 (N_6185,N_5394,N_4249);
or U6186 (N_6186,N_3950,N_3655);
or U6187 (N_6187,N_3268,N_3149);
or U6188 (N_6188,N_3357,N_5138);
or U6189 (N_6189,N_5008,N_3728);
nand U6190 (N_6190,N_5613,N_5921);
nand U6191 (N_6191,N_4322,N_5603);
and U6192 (N_6192,N_3113,N_4976);
nor U6193 (N_6193,N_3305,N_4910);
nor U6194 (N_6194,N_3947,N_4276);
or U6195 (N_6195,N_4701,N_3482);
nor U6196 (N_6196,N_4320,N_5088);
and U6197 (N_6197,N_5529,N_3496);
or U6198 (N_6198,N_4577,N_3847);
nor U6199 (N_6199,N_3686,N_4236);
and U6200 (N_6200,N_4147,N_5212);
nand U6201 (N_6201,N_4429,N_5518);
and U6202 (N_6202,N_4109,N_3710);
nand U6203 (N_6203,N_5624,N_4299);
and U6204 (N_6204,N_5683,N_5639);
xnor U6205 (N_6205,N_5010,N_4145);
or U6206 (N_6206,N_4587,N_5262);
xor U6207 (N_6207,N_4457,N_3187);
nand U6208 (N_6208,N_3965,N_4379);
and U6209 (N_6209,N_4863,N_3857);
nor U6210 (N_6210,N_4047,N_3702);
nand U6211 (N_6211,N_4639,N_5261);
nand U6212 (N_6212,N_3039,N_5057);
xnor U6213 (N_6213,N_5849,N_4119);
or U6214 (N_6214,N_4046,N_3541);
nand U6215 (N_6215,N_3026,N_5431);
nor U6216 (N_6216,N_3616,N_5700);
nor U6217 (N_6217,N_3237,N_4091);
and U6218 (N_6218,N_3786,N_4710);
or U6219 (N_6219,N_5053,N_3720);
nor U6220 (N_6220,N_5130,N_3458);
and U6221 (N_6221,N_4569,N_5236);
nand U6222 (N_6222,N_3475,N_4563);
or U6223 (N_6223,N_5555,N_4228);
or U6224 (N_6224,N_5411,N_5820);
xor U6225 (N_6225,N_5800,N_5580);
and U6226 (N_6226,N_3528,N_5577);
nand U6227 (N_6227,N_3078,N_4059);
and U6228 (N_6228,N_4677,N_5765);
nor U6229 (N_6229,N_3664,N_4026);
and U6230 (N_6230,N_5992,N_3631);
and U6231 (N_6231,N_3488,N_3176);
nand U6232 (N_6232,N_4111,N_3172);
or U6233 (N_6233,N_3937,N_5622);
or U6234 (N_6234,N_5390,N_5044);
or U6235 (N_6235,N_3164,N_3934);
nand U6236 (N_6236,N_3275,N_4346);
nor U6237 (N_6237,N_3165,N_4153);
or U6238 (N_6238,N_3704,N_3867);
nor U6239 (N_6239,N_5350,N_5590);
nor U6240 (N_6240,N_3865,N_4545);
and U6241 (N_6241,N_5920,N_5030);
nand U6242 (N_6242,N_4448,N_4894);
xor U6243 (N_6243,N_4023,N_4628);
nor U6244 (N_6244,N_4231,N_4130);
nand U6245 (N_6245,N_5727,N_3424);
nor U6246 (N_6246,N_4187,N_3468);
or U6247 (N_6247,N_4465,N_5719);
nor U6248 (N_6248,N_4422,N_4019);
and U6249 (N_6249,N_5135,N_5055);
nand U6250 (N_6250,N_5843,N_5502);
or U6251 (N_6251,N_3045,N_3918);
nor U6252 (N_6252,N_3837,N_4813);
nor U6253 (N_6253,N_5889,N_3454);
nor U6254 (N_6254,N_3855,N_3879);
or U6255 (N_6255,N_4572,N_5392);
or U6256 (N_6256,N_5019,N_5237);
nor U6257 (N_6257,N_5217,N_4785);
and U6258 (N_6258,N_3530,N_5979);
or U6259 (N_6259,N_4823,N_4533);
and U6260 (N_6260,N_5279,N_5993);
or U6261 (N_6261,N_5828,N_5854);
nand U6262 (N_6262,N_5597,N_3010);
and U6263 (N_6263,N_4799,N_5354);
and U6264 (N_6264,N_5958,N_5437);
or U6265 (N_6265,N_4421,N_4061);
nor U6266 (N_6266,N_5155,N_5552);
nand U6267 (N_6267,N_3294,N_5801);
or U6268 (N_6268,N_5199,N_4020);
or U6269 (N_6269,N_5406,N_4932);
nor U6270 (N_6270,N_5668,N_5585);
or U6271 (N_6271,N_4786,N_4935);
nand U6272 (N_6272,N_3839,N_5021);
nor U6273 (N_6273,N_3334,N_5402);
or U6274 (N_6274,N_4746,N_3586);
nor U6275 (N_6275,N_5451,N_5989);
or U6276 (N_6276,N_4636,N_3111);
nor U6277 (N_6277,N_4501,N_4084);
and U6278 (N_6278,N_4507,N_5810);
or U6279 (N_6279,N_4732,N_5887);
nor U6280 (N_6280,N_4376,N_4077);
or U6281 (N_6281,N_3628,N_5201);
or U6282 (N_6282,N_4579,N_5484);
and U6283 (N_6283,N_3249,N_5345);
nor U6284 (N_6284,N_4778,N_4264);
and U6285 (N_6285,N_3476,N_3620);
or U6286 (N_6286,N_3210,N_3053);
nand U6287 (N_6287,N_4296,N_3992);
or U6288 (N_6288,N_3601,N_5045);
nor U6289 (N_6289,N_5826,N_4692);
or U6290 (N_6290,N_5938,N_3444);
or U6291 (N_6291,N_3253,N_3089);
or U6292 (N_6292,N_5310,N_5302);
nand U6293 (N_6293,N_5159,N_3666);
nand U6294 (N_6294,N_5246,N_3740);
or U6295 (N_6295,N_4736,N_3222);
or U6296 (N_6296,N_4893,N_3944);
and U6297 (N_6297,N_3273,N_5571);
nand U6298 (N_6298,N_3461,N_5846);
and U6299 (N_6299,N_5062,N_3411);
or U6300 (N_6300,N_3596,N_3148);
or U6301 (N_6301,N_3012,N_5783);
and U6302 (N_6302,N_4637,N_4679);
nor U6303 (N_6303,N_4821,N_5663);
xnor U6304 (N_6304,N_4502,N_5823);
and U6305 (N_6305,N_3874,N_5426);
or U6306 (N_6306,N_3003,N_3484);
or U6307 (N_6307,N_4650,N_5551);
and U6308 (N_6308,N_4305,N_3281);
nor U6309 (N_6309,N_5838,N_5366);
or U6310 (N_6310,N_5353,N_3134);
nor U6311 (N_6311,N_3816,N_3778);
and U6312 (N_6312,N_4377,N_3898);
and U6313 (N_6313,N_3409,N_3159);
and U6314 (N_6314,N_4494,N_5146);
nand U6315 (N_6315,N_5523,N_4027);
and U6316 (N_6316,N_5895,N_5665);
nand U6317 (N_6317,N_3842,N_5243);
and U6318 (N_6318,N_4325,N_3415);
nand U6319 (N_6319,N_5098,N_4654);
and U6320 (N_6320,N_3689,N_4593);
or U6321 (N_6321,N_5772,N_4988);
or U6322 (N_6322,N_3629,N_5399);
and U6323 (N_6323,N_4779,N_3977);
and U6324 (N_6324,N_3041,N_3033);
xor U6325 (N_6325,N_5643,N_4327);
nor U6326 (N_6326,N_3283,N_3796);
and U6327 (N_6327,N_5535,N_3684);
nor U6328 (N_6328,N_4547,N_4162);
or U6329 (N_6329,N_3251,N_3452);
or U6330 (N_6330,N_3119,N_5951);
nand U6331 (N_6331,N_5297,N_4420);
nor U6332 (N_6332,N_4945,N_4693);
or U6333 (N_6333,N_5746,N_5209);
nor U6334 (N_6334,N_5532,N_3008);
and U6335 (N_6335,N_5228,N_3433);
nor U6336 (N_6336,N_4495,N_4841);
nor U6337 (N_6337,N_5988,N_4365);
or U6338 (N_6338,N_5793,N_3860);
and U6339 (N_6339,N_5900,N_3342);
or U6340 (N_6340,N_5975,N_3279);
and U6341 (N_6341,N_5123,N_4054);
or U6342 (N_6342,N_3395,N_3975);
nand U6343 (N_6343,N_4901,N_4401);
or U6344 (N_6344,N_4316,N_3761);
or U6345 (N_6345,N_4756,N_3106);
nor U6346 (N_6346,N_3126,N_4971);
nor U6347 (N_6347,N_5166,N_4536);
and U6348 (N_6348,N_5129,N_4795);
or U6349 (N_6349,N_3683,N_5117);
or U6350 (N_6350,N_4827,N_4029);
nor U6351 (N_6351,N_3005,N_4848);
nand U6352 (N_6352,N_4727,N_5807);
or U6353 (N_6353,N_3198,N_4279);
or U6354 (N_6354,N_4035,N_5505);
or U6355 (N_6355,N_5911,N_5456);
nor U6356 (N_6356,N_4644,N_5796);
or U6357 (N_6357,N_4284,N_3870);
nor U6358 (N_6358,N_3450,N_5701);
nor U6359 (N_6359,N_5497,N_4982);
or U6360 (N_6360,N_4803,N_3124);
and U6361 (N_6361,N_4515,N_4855);
nand U6362 (N_6362,N_4381,N_4102);
nand U6363 (N_6363,N_3613,N_5295);
nor U6364 (N_6364,N_4810,N_5332);
or U6365 (N_6365,N_5890,N_5501);
or U6366 (N_6366,N_3969,N_3863);
and U6367 (N_6367,N_4996,N_3678);
and U6368 (N_6368,N_3286,N_3561);
and U6369 (N_6369,N_3674,N_4482);
nand U6370 (N_6370,N_4386,N_5358);
or U6371 (N_6371,N_4036,N_4144);
nor U6372 (N_6372,N_3611,N_4721);
nand U6373 (N_6373,N_5825,N_5918);
nand U6374 (N_6374,N_3331,N_3858);
or U6375 (N_6375,N_4069,N_5128);
and U6376 (N_6376,N_5664,N_4828);
or U6377 (N_6377,N_5888,N_4926);
nand U6378 (N_6378,N_3034,N_5032);
or U6379 (N_6379,N_3722,N_3054);
nor U6380 (N_6380,N_3732,N_3735);
or U6381 (N_6381,N_5266,N_3202);
nand U6382 (N_6382,N_3341,N_5931);
nor U6383 (N_6383,N_3634,N_3765);
nor U6384 (N_6384,N_3539,N_3749);
or U6385 (N_6385,N_4978,N_5316);
and U6386 (N_6386,N_3442,N_3373);
and U6387 (N_6387,N_5730,N_5998);
and U6388 (N_6388,N_4856,N_4760);
and U6389 (N_6389,N_3698,N_5599);
xor U6390 (N_6390,N_3125,N_5413);
nand U6391 (N_6391,N_5506,N_5334);
and U6392 (N_6392,N_3290,N_5020);
nor U6393 (N_6393,N_3537,N_4566);
nand U6394 (N_6394,N_4142,N_4991);
nand U6395 (N_6395,N_5205,N_4936);
nand U6396 (N_6396,N_5432,N_5059);
nand U6397 (N_6397,N_3266,N_4297);
or U6398 (N_6398,N_4341,N_4719);
nand U6399 (N_6399,N_4949,N_3699);
or U6400 (N_6400,N_4002,N_3117);
nor U6401 (N_6401,N_3140,N_3793);
and U6402 (N_6402,N_5753,N_4340);
or U6403 (N_6403,N_3687,N_5879);
nor U6404 (N_6404,N_3560,N_4987);
nand U6405 (N_6405,N_3585,N_5317);
nand U6406 (N_6406,N_5759,N_3128);
or U6407 (N_6407,N_4983,N_3348);
and U6408 (N_6408,N_3303,N_4758);
nand U6409 (N_6409,N_3156,N_4067);
or U6410 (N_6410,N_4979,N_4470);
nand U6411 (N_6411,N_3067,N_5042);
and U6412 (N_6412,N_3650,N_4742);
and U6413 (N_6413,N_5874,N_5961);
or U6414 (N_6414,N_5156,N_5927);
and U6415 (N_6415,N_5351,N_5623);
and U6416 (N_6416,N_5011,N_4641);
or U6417 (N_6417,N_4706,N_3302);
and U6418 (N_6418,N_5344,N_4527);
or U6419 (N_6419,N_5997,N_4159);
nor U6420 (N_6420,N_4564,N_3453);
nand U6421 (N_6421,N_5809,N_4859);
nand U6422 (N_6422,N_3497,N_5758);
nor U6423 (N_6423,N_5028,N_5449);
xnor U6424 (N_6424,N_3833,N_5177);
nand U6425 (N_6425,N_5270,N_3547);
nor U6426 (N_6426,N_4559,N_3798);
nand U6427 (N_6427,N_4313,N_4968);
or U6428 (N_6428,N_4100,N_3715);
or U6429 (N_6429,N_5241,N_5487);
nor U6430 (N_6430,N_5582,N_3963);
or U6431 (N_6431,N_3094,N_3465);
nor U6432 (N_6432,N_4686,N_5136);
or U6433 (N_6433,N_3555,N_3353);
and U6434 (N_6434,N_4291,N_3460);
or U6435 (N_6435,N_3189,N_5857);
or U6436 (N_6436,N_4211,N_3499);
nor U6437 (N_6437,N_3770,N_4355);
nand U6438 (N_6438,N_4118,N_4348);
nand U6439 (N_6439,N_5737,N_5578);
nor U6440 (N_6440,N_4339,N_5880);
nor U6441 (N_6441,N_4043,N_3536);
nor U6442 (N_6442,N_5937,N_4584);
and U6443 (N_6443,N_4416,N_5052);
and U6444 (N_6444,N_5100,N_5969);
nor U6445 (N_6445,N_5507,N_3824);
or U6446 (N_6446,N_4082,N_4618);
or U6447 (N_6447,N_3746,N_3671);
and U6448 (N_6448,N_4051,N_5923);
nand U6449 (N_6449,N_5654,N_4884);
and U6450 (N_6450,N_4999,N_3051);
or U6451 (N_6451,N_3329,N_3647);
nand U6452 (N_6452,N_3921,N_5235);
and U6453 (N_6453,N_5728,N_4298);
or U6454 (N_6454,N_3669,N_4113);
nor U6455 (N_6455,N_5592,N_5500);
nor U6456 (N_6456,N_3818,N_5299);
and U6457 (N_6457,N_3976,N_5170);
and U6458 (N_6458,N_3058,N_5766);
nand U6459 (N_6459,N_5488,N_5048);
or U6460 (N_6460,N_3326,N_4304);
nor U6461 (N_6461,N_5026,N_5631);
and U6462 (N_6462,N_5515,N_5188);
and U6463 (N_6463,N_5187,N_4445);
nor U6464 (N_6464,N_4366,N_4504);
nand U6465 (N_6465,N_5761,N_5304);
nor U6466 (N_6466,N_5791,N_3459);
nor U6467 (N_6467,N_4549,N_4531);
xor U6468 (N_6468,N_4419,N_3907);
nand U6469 (N_6469,N_3845,N_3349);
and U6470 (N_6470,N_4479,N_4537);
or U6471 (N_6471,N_5991,N_5651);
nor U6472 (N_6472,N_3953,N_3121);
xor U6473 (N_6473,N_3274,N_3028);
nor U6474 (N_6474,N_5644,N_5151);
nand U6475 (N_6475,N_4168,N_3930);
nor U6476 (N_6476,N_5131,N_3263);
nor U6477 (N_6477,N_5331,N_4879);
nand U6478 (N_6478,N_5215,N_5091);
nand U6479 (N_6479,N_3851,N_4934);
nor U6480 (N_6480,N_4227,N_4399);
and U6481 (N_6481,N_5318,N_4446);
or U6482 (N_6482,N_5203,N_3295);
nor U6483 (N_6483,N_4695,N_3351);
nand U6484 (N_6484,N_5716,N_3378);
nand U6485 (N_6485,N_5642,N_5440);
or U6486 (N_6486,N_4992,N_3651);
nand U6487 (N_6487,N_4675,N_3742);
or U6488 (N_6488,N_5272,N_3142);
nand U6489 (N_6489,N_3705,N_4378);
or U6490 (N_6490,N_4519,N_4543);
and U6491 (N_6491,N_4072,N_4169);
nand U6492 (N_6492,N_4206,N_5105);
and U6493 (N_6493,N_3603,N_5714);
and U6494 (N_6494,N_4900,N_4831);
nor U6495 (N_6495,N_3422,N_4784);
nor U6496 (N_6496,N_5649,N_4990);
nor U6497 (N_6497,N_4518,N_5824);
and U6498 (N_6498,N_5398,N_5158);
and U6499 (N_6499,N_3810,N_3296);
nor U6500 (N_6500,N_5569,N_5275);
and U6501 (N_6501,N_5309,N_5625);
nor U6502 (N_6502,N_3792,N_4481);
or U6503 (N_6503,N_3470,N_4066);
xnor U6504 (N_6504,N_3945,N_4281);
and U6505 (N_6505,N_4181,N_3112);
nand U6506 (N_6506,N_4857,N_4674);
nor U6507 (N_6507,N_4050,N_4532);
or U6508 (N_6508,N_5972,N_5608);
nor U6509 (N_6509,N_3077,N_3246);
nand U6510 (N_6510,N_5533,N_5420);
or U6511 (N_6511,N_4007,N_3928);
nor U6512 (N_6512,N_3780,N_5811);
or U6513 (N_6513,N_4360,N_4653);
nand U6514 (N_6514,N_3949,N_4410);
nor U6515 (N_6515,N_5839,N_4808);
nor U6516 (N_6516,N_5818,N_3972);
nor U6517 (N_6517,N_5125,N_5944);
and U6518 (N_6518,N_5594,N_5202);
and U6519 (N_6519,N_5276,N_4993);
nor U6520 (N_6520,N_5210,N_4690);
nand U6521 (N_6521,N_3521,N_4649);
or U6522 (N_6522,N_4838,N_3261);
or U6523 (N_6523,N_5521,N_5570);
nor U6524 (N_6524,N_5324,N_4454);
nand U6525 (N_6525,N_3044,N_3402);
nand U6526 (N_6526,N_3725,N_3518);
nand U6527 (N_6527,N_3883,N_5576);
and U6528 (N_6528,N_4807,N_5168);
nand U6529 (N_6529,N_3061,N_3346);
and U6530 (N_6530,N_5003,N_5595);
or U6531 (N_6531,N_4877,N_5775);
xnor U6532 (N_6532,N_5035,N_5990);
nor U6533 (N_6533,N_5448,N_3800);
or U6534 (N_6534,N_4977,N_5646);
nand U6535 (N_6535,N_3489,N_3914);
and U6536 (N_6536,N_4049,N_5288);
nor U6537 (N_6537,N_5687,N_4487);
nor U6538 (N_6538,N_5339,N_5524);
and U6539 (N_6539,N_3363,N_5148);
nand U6540 (N_6540,N_4717,N_5183);
nand U6541 (N_6541,N_4865,N_4835);
nand U6542 (N_6542,N_4508,N_4268);
nor U6543 (N_6543,N_3178,N_5731);
and U6544 (N_6544,N_4398,N_5549);
and U6545 (N_6545,N_5435,N_4295);
nor U6546 (N_6546,N_5994,N_3434);
and U6547 (N_6547,N_4451,N_3575);
and U6548 (N_6548,N_3635,N_4280);
and U6549 (N_6549,N_4726,N_4619);
nand U6550 (N_6550,N_3208,N_5422);
or U6551 (N_6551,N_5080,N_5788);
nor U6552 (N_6552,N_5872,N_4384);
or U6553 (N_6553,N_5581,N_5903);
and U6554 (N_6554,N_3753,N_3335);
and U6555 (N_6555,N_5559,N_4234);
or U6556 (N_6556,N_5213,N_5610);
or U6557 (N_6557,N_5722,N_3764);
and U6558 (N_6558,N_4045,N_3370);
nor U6559 (N_6559,N_3659,N_5412);
nand U6560 (N_6560,N_4594,N_5416);
nand U6561 (N_6561,N_4520,N_4209);
and U6562 (N_6562,N_4552,N_5656);
nor U6563 (N_6563,N_4222,N_5691);
nand U6564 (N_6564,N_3957,N_5999);
and U6565 (N_6565,N_5531,N_3675);
nor U6566 (N_6566,N_3526,N_4001);
nor U6567 (N_6567,N_4702,N_5089);
and U6568 (N_6568,N_3615,N_4039);
and U6569 (N_6569,N_4447,N_3946);
and U6570 (N_6570,N_3052,N_3619);
nor U6571 (N_6571,N_3942,N_4018);
nor U6572 (N_6572,N_5167,N_3018);
nor U6573 (N_6573,N_4357,N_4418);
nor U6574 (N_6574,N_5389,N_4585);
and U6575 (N_6575,N_4524,N_3410);
nor U6576 (N_6576,N_4456,N_5616);
and U6577 (N_6577,N_5554,N_4964);
or U6578 (N_6578,N_4406,N_5365);
and U6579 (N_6579,N_3043,N_3379);
nand U6580 (N_6580,N_5335,N_5072);
nand U6581 (N_6581,N_3872,N_4453);
nor U6582 (N_6582,N_3826,N_3238);
xnor U6583 (N_6583,N_3979,N_3485);
and U6584 (N_6584,N_3564,N_5149);
and U6585 (N_6585,N_3280,N_5347);
nor U6586 (N_6586,N_5382,N_3777);
and U6587 (N_6587,N_3504,N_5878);
nand U6588 (N_6588,N_3955,N_4651);
nor U6589 (N_6589,N_3751,N_4120);
nor U6590 (N_6590,N_5066,N_4257);
nand U6591 (N_6591,N_3430,N_5224);
nor U6592 (N_6592,N_3075,N_4629);
and U6593 (N_6593,N_5104,N_5101);
nor U6594 (N_6594,N_3161,N_4950);
nor U6595 (N_6595,N_3663,N_3531);
and U6596 (N_6596,N_5457,N_3327);
nand U6597 (N_6597,N_4980,N_3062);
and U6598 (N_6598,N_5680,N_5473);
xnor U6599 (N_6599,N_4240,N_4088);
nor U6600 (N_6600,N_4178,N_3606);
nand U6601 (N_6601,N_5740,N_4275);
or U6602 (N_6602,N_5419,N_3048);
or U6603 (N_6603,N_5485,N_5983);
nand U6604 (N_6604,N_3890,N_5153);
xor U6605 (N_6605,N_5980,N_5611);
nor U6606 (N_6606,N_4262,N_4070);
or U6607 (N_6607,N_5004,N_5841);
nor U6608 (N_6608,N_4490,N_3624);
nand U6609 (N_6609,N_3726,N_5563);
nand U6610 (N_6610,N_4319,N_4343);
or U6611 (N_6611,N_5090,N_4899);
nand U6612 (N_6612,N_4505,N_3670);
or U6613 (N_6613,N_3400,N_5094);
or U6614 (N_6614,N_3183,N_5007);
nor U6615 (N_6615,N_5244,N_5959);
nand U6616 (N_6616,N_5278,N_5679);
nand U6617 (N_6617,N_3205,N_3213);
and U6618 (N_6618,N_3029,N_3594);
or U6619 (N_6619,N_5822,N_3897);
nand U6620 (N_6620,N_5892,N_5190);
xnor U6621 (N_6621,N_3692,N_5330);
nor U6622 (N_6622,N_4829,N_5560);
xnor U6623 (N_6623,N_3192,N_3657);
nor U6624 (N_6624,N_3162,N_5370);
or U6625 (N_6625,N_4172,N_5352);
nand U6626 (N_6626,N_4994,N_4781);
nand U6627 (N_6627,N_5885,N_5707);
nand U6628 (N_6628,N_5971,N_4161);
nor U6629 (N_6629,N_3548,N_4437);
and U6630 (N_6630,N_3998,N_4220);
and U6631 (N_6631,N_5954,N_3703);
nor U6632 (N_6632,N_5587,N_4426);
nor U6633 (N_6633,N_5251,N_3951);
nor U6634 (N_6634,N_4000,N_5865);
nand U6635 (N_6635,N_5414,N_5925);
or U6636 (N_6636,N_3024,N_4660);
or U6637 (N_6637,N_5756,N_4683);
nand U6638 (N_6638,N_3532,N_3677);
nor U6639 (N_6639,N_3020,N_3806);
or U6640 (N_6640,N_4705,N_4844);
nor U6641 (N_6641,N_5550,N_4391);
nor U6642 (N_6642,N_4432,N_5522);
nor U6643 (N_6643,N_5819,N_5060);
xnor U6644 (N_6644,N_4126,N_3399);
nand U6645 (N_6645,N_4350,N_3723);
nand U6646 (N_6646,N_3404,N_3101);
and U6647 (N_6647,N_4567,N_4624);
nand U6648 (N_6648,N_3838,N_5710);
nand U6649 (N_6649,N_4937,N_4796);
nand U6650 (N_6650,N_3566,N_3790);
nor U6651 (N_6651,N_4525,N_4764);
nor U6652 (N_6652,N_3931,N_4634);
and U6653 (N_6653,N_3724,N_3403);
nor U6654 (N_6654,N_3429,N_3355);
nor U6655 (N_6655,N_4259,N_5441);
nor U6656 (N_6656,N_3662,N_4946);
nand U6657 (N_6657,N_4497,N_3590);
xnor U6658 (N_6658,N_4954,N_3750);
nand U6659 (N_6659,N_4722,N_4833);
and U6660 (N_6660,N_5509,N_4907);
and U6661 (N_6661,N_5729,N_4148);
and U6662 (N_6662,N_3516,N_5797);
and U6663 (N_6663,N_3785,N_5410);
or U6664 (N_6664,N_3940,N_3551);
nand U6665 (N_6665,N_5815,N_3577);
nor U6666 (N_6666,N_4840,N_5447);
nand U6667 (N_6667,N_4655,N_4824);
nand U6668 (N_6668,N_5548,N_4308);
nand U6669 (N_6669,N_3088,N_4166);
or U6670 (N_6670,N_4740,N_5341);
and U6671 (N_6671,N_5133,N_5061);
or U6672 (N_6672,N_5914,N_4105);
nand U6673 (N_6673,N_5033,N_3477);
and U6674 (N_6674,N_5870,N_5322);
nand U6675 (N_6675,N_5527,N_4400);
nand U6676 (N_6676,N_3960,N_5242);
nor U6677 (N_6677,N_3559,N_3136);
nand U6678 (N_6678,N_4435,N_5939);
nand U6679 (N_6679,N_3876,N_5525);
or U6680 (N_6680,N_5160,N_4430);
nand U6681 (N_6681,N_3730,N_4057);
nor U6682 (N_6682,N_5038,N_5821);
nor U6683 (N_6683,N_4097,N_3843);
nor U6684 (N_6684,N_5553,N_5850);
nand U6685 (N_6685,N_3741,N_3697);
xor U6686 (N_6686,N_4870,N_4853);
xnor U6687 (N_6687,N_5039,N_5995);
or U6688 (N_6688,N_4472,N_4733);
nand U6689 (N_6689,N_5957,N_3595);
or U6690 (N_6690,N_5023,N_4330);
and U6691 (N_6691,N_5490,N_4436);
and U6692 (N_6692,N_5047,N_4599);
or U6693 (N_6693,N_5480,N_5063);
or U6694 (N_6694,N_5790,N_5734);
nand U6695 (N_6695,N_5225,N_4068);
nand U6696 (N_6696,N_3325,N_4009);
and U6697 (N_6697,N_5327,N_3204);
or U6698 (N_6698,N_3693,N_5386);
nand U6699 (N_6699,N_4226,N_3804);
and U6700 (N_6700,N_4441,N_4849);
or U6701 (N_6701,N_4277,N_5896);
and U6702 (N_6702,N_4595,N_3916);
or U6703 (N_6703,N_3129,N_4575);
and U6704 (N_6704,N_5657,N_4604);
or U6705 (N_6705,N_3243,N_3700);
nand U6706 (N_6706,N_3989,N_3573);
nor U6707 (N_6707,N_5429,N_3257);
and U6708 (N_6708,N_5054,N_4820);
and U6709 (N_6709,N_3652,N_4942);
nor U6710 (N_6710,N_3235,N_3894);
nor U6711 (N_6711,N_3338,N_5255);
or U6712 (N_6712,N_5071,N_3776);
and U6713 (N_6713,N_4741,N_4612);
and U6714 (N_6714,N_4478,N_3490);
xnor U6715 (N_6715,N_3823,N_4117);
and U6716 (N_6716,N_4591,N_3209);
and U6717 (N_6717,N_5690,N_5635);
and U6718 (N_6718,N_3574,N_3899);
nand U6719 (N_6719,N_5661,N_4969);
xor U6720 (N_6720,N_3260,N_5343);
nor U6721 (N_6721,N_4488,N_3797);
nand U6722 (N_6722,N_4245,N_5678);
or U6723 (N_6723,N_3242,N_4188);
nand U6724 (N_6724,N_4191,N_4042);
or U6725 (N_6725,N_3556,N_3637);
nor U6726 (N_6726,N_3709,N_5637);
nand U6727 (N_6727,N_4468,N_5284);
nand U6728 (N_6728,N_4659,N_3927);
nor U6729 (N_6729,N_5899,N_4010);
nor U6730 (N_6730,N_3011,N_3082);
and U6731 (N_6731,N_5605,N_5503);
or U6732 (N_6732,N_3641,N_4951);
and U6733 (N_6733,N_3171,N_3522);
nand U6734 (N_6734,N_3025,N_4955);
or U6735 (N_6735,N_4403,N_4283);
nand U6736 (N_6736,N_5789,N_3713);
and U6737 (N_6737,N_3759,N_4473);
or U6738 (N_6738,N_4380,N_3680);
and U6739 (N_6739,N_5520,N_4337);
and U6740 (N_6740,N_5798,N_5883);
and U6741 (N_6741,N_4048,N_4794);
nor U6742 (N_6742,N_5785,N_3775);
or U6743 (N_6743,N_3056,N_3908);
nor U6744 (N_6744,N_4938,N_3122);
nand U6745 (N_6745,N_3227,N_3074);
and U6746 (N_6746,N_5781,N_3769);
nor U6747 (N_6747,N_4872,N_4995);
nand U6748 (N_6748,N_4104,N_3361);
or U6749 (N_6749,N_3646,N_5670);
and U6750 (N_6750,N_5659,N_3610);
or U6751 (N_6751,N_4886,N_5606);
nand U6752 (N_6752,N_4952,N_5754);
and U6753 (N_6753,N_4959,N_5703);
or U6754 (N_6754,N_5282,N_5012);
or U6755 (N_6755,N_5688,N_3109);
xor U6756 (N_6756,N_3913,N_3428);
nand U6757 (N_6757,N_4777,N_4221);
or U6758 (N_6758,N_5704,N_3719);
nand U6759 (N_6759,N_3773,N_3027);
and U6760 (N_6760,N_4271,N_5705);
and U6761 (N_6761,N_4704,N_4202);
and U6762 (N_6762,N_5489,N_5645);
nor U6763 (N_6763,N_4058,N_5083);
or U6764 (N_6764,N_3160,N_3768);
nand U6765 (N_6765,N_3491,N_3691);
xnor U6766 (N_6766,N_5638,N_3794);
and U6767 (N_6767,N_3878,N_4203);
nand U6768 (N_6768,N_3756,N_3212);
and U6769 (N_6769,N_3987,N_3215);
nand U6770 (N_6770,N_4154,N_4423);
and U6771 (N_6771,N_3967,N_4506);
or U6772 (N_6772,N_5277,N_4196);
and U6773 (N_6773,N_3562,N_3177);
nor U6774 (N_6774,N_5702,N_4157);
or U6775 (N_6775,N_3549,N_3287);
or U6776 (N_6776,N_4697,N_4134);
nor U6777 (N_6777,N_5669,N_5771);
nand U6778 (N_6778,N_5672,N_3145);
nor U6779 (N_6779,N_3184,N_5770);
xor U6780 (N_6780,N_5373,N_3512);
xnor U6781 (N_6781,N_5511,N_4083);
and U6782 (N_6782,N_5955,N_4610);
nor U6783 (N_6783,N_3068,N_4546);
nand U6784 (N_6784,N_3599,N_5204);
nand U6785 (N_6785,N_3667,N_5357);
nor U6786 (N_6786,N_3214,N_4730);
nor U6787 (N_6787,N_3654,N_5446);
and U6788 (N_6788,N_4273,N_4122);
nand U6789 (N_6789,N_5508,N_4613);
xor U6790 (N_6790,N_4511,N_3451);
nor U6791 (N_6791,N_3108,N_3333);
or U6792 (N_6792,N_3783,N_3846);
or U6793 (N_6793,N_5543,N_5653);
or U6794 (N_6794,N_3059,N_3339);
and U6795 (N_6795,N_5866,N_4090);
and U6796 (N_6796,N_4956,N_5405);
nand U6797 (N_6797,N_5321,N_3618);
or U6798 (N_6798,N_5112,N_3046);
nor U6799 (N_6799,N_4438,N_4707);
and U6800 (N_6800,N_5040,N_3961);
or U6801 (N_6801,N_5720,N_5320);
nand U6802 (N_6802,N_3383,N_5108);
or U6803 (N_6803,N_4250,N_4534);
and U6804 (N_6804,N_4625,N_4931);
nor U6805 (N_6805,N_4904,N_3405);
or U6806 (N_6806,N_4013,N_3207);
or U6807 (N_6807,N_4387,N_3240);
nand U6808 (N_6808,N_4972,N_5583);
or U6809 (N_6809,N_5360,N_3304);
nor U6810 (N_6810,N_5075,N_3414);
or U6811 (N_6811,N_4008,N_4151);
and U6812 (N_6812,N_3217,N_3830);
nand U6813 (N_6813,N_3580,N_3038);
or U6814 (N_6814,N_5425,N_4266);
and U6815 (N_6815,N_3110,N_5915);
or U6816 (N_6816,N_5319,N_3995);
nor U6817 (N_6817,N_5930,N_3323);
nand U6818 (N_6818,N_3982,N_4440);
nand U6819 (N_6819,N_4351,N_5229);
nand U6820 (N_6820,N_4485,N_4914);
and U6821 (N_6821,N_3391,N_5391);
or U6822 (N_6822,N_3023,N_5636);
or U6823 (N_6823,N_3037,N_3582);
nor U6824 (N_6824,N_4606,N_5046);
nand U6825 (N_6825,N_3186,N_3332);
nor U6826 (N_6826,N_5541,N_4460);
and U6827 (N_6827,N_5214,N_4944);
nor U6828 (N_6828,N_3344,N_5162);
and U6829 (N_6829,N_3371,N_4219);
nand U6830 (N_6830,N_4455,N_5817);
nor U6831 (N_6831,N_3291,N_4177);
nor U6832 (N_6832,N_3903,N_5684);
nor U6833 (N_6833,N_3103,N_3540);
or U6834 (N_6834,N_3006,N_5692);
or U6835 (N_6835,N_3902,N_3236);
nor U6836 (N_6836,N_5808,N_5832);
nor U6837 (N_6837,N_5430,N_4925);
nand U6838 (N_6838,N_5181,N_5987);
or U6839 (N_6839,N_5257,N_4225);
nand U6840 (N_6840,N_3425,N_3151);
and U6841 (N_6841,N_5876,N_3385);
nor U6842 (N_6842,N_4044,N_5154);
nor U6843 (N_6843,N_5940,N_3387);
nand U6844 (N_6844,N_3587,N_3828);
or U6845 (N_6845,N_5813,N_4922);
nor U6846 (N_6846,N_5942,N_3201);
nor U6847 (N_6847,N_3386,N_5962);
nand U6848 (N_6848,N_5510,N_5666);
and U6849 (N_6849,N_3366,N_4592);
nor U6850 (N_6850,N_4115,N_5113);
or U6851 (N_6851,N_5726,N_4981);
and U6852 (N_6852,N_3494,N_3835);
nand U6853 (N_6853,N_5733,N_5504);
or U6854 (N_6854,N_4483,N_3936);
or U6855 (N_6855,N_5579,N_5069);
and U6856 (N_6856,N_4404,N_4425);
nor U6857 (N_6857,N_3986,N_3292);
or U6858 (N_6858,N_5782,N_4928);
nor U6859 (N_6859,N_3721,N_3597);
nand U6860 (N_6860,N_3120,N_4801);
nand U6861 (N_6861,N_5093,N_4347);
nor U6862 (N_6862,N_3621,N_4373);
xor U6863 (N_6863,N_3939,N_3206);
nand U6864 (N_6864,N_3276,N_4229);
or U6865 (N_6865,N_4103,N_5709);
and U6866 (N_6866,N_3600,N_4739);
and U6867 (N_6867,N_4270,N_5573);
nand U6868 (N_6868,N_4825,N_4260);
and U6869 (N_6869,N_3507,N_5627);
or U6870 (N_6870,N_5853,N_3665);
nor U6871 (N_6871,N_3271,N_3277);
or U6872 (N_6872,N_5650,N_5253);
nand U6873 (N_6873,N_3502,N_3529);
nand U6874 (N_6874,N_5840,N_5893);
or U6875 (N_6875,N_4712,N_5496);
nor U6876 (N_6876,N_4753,N_4086);
or U6877 (N_6877,N_5234,N_3885);
and U6878 (N_6878,N_3098,N_5407);
nand U6879 (N_6879,N_5546,N_3211);
or U6880 (N_6880,N_4961,N_5658);
or U6881 (N_6881,N_4289,N_3443);
or U6882 (N_6882,N_5403,N_5655);
or U6883 (N_6883,N_3267,N_5768);
nand U6884 (N_6884,N_4645,N_3009);
and U6885 (N_6885,N_3758,N_5185);
nand U6886 (N_6886,N_5584,N_4676);
nor U6887 (N_6887,N_4703,N_4646);
nand U6888 (N_6888,N_4135,N_4402);
nand U6889 (N_6889,N_4041,N_3282);
or U6890 (N_6890,N_5891,N_3754);
and U6891 (N_6891,N_4163,N_3752);
nand U6892 (N_6892,N_5557,N_5675);
and U6893 (N_6893,N_4586,N_5065);
or U6894 (N_6894,N_3421,N_5450);
xnor U6895 (N_6895,N_4658,N_5732);
or U6896 (N_6896,N_4673,N_3168);
nand U6897 (N_6897,N_3829,N_4056);
nand U6898 (N_6898,N_3888,N_5230);
or U6899 (N_6899,N_3814,N_5498);
nor U6900 (N_6900,N_3492,N_4965);
nor U6901 (N_6901,N_3869,N_3493);
nor U6902 (N_6902,N_4967,N_5191);
nor U6903 (N_6903,N_3457,N_3445);
or U6904 (N_6904,N_4724,N_4913);
nor U6905 (N_6905,N_4390,N_4876);
or U6906 (N_6906,N_3733,N_4336);
or U6907 (N_6907,N_5303,N_5837);
and U6908 (N_6908,N_5486,N_4958);
or U6909 (N_6909,N_4204,N_4123);
and U6910 (N_6910,N_3441,N_4682);
nor U6911 (N_6911,N_5226,N_3060);
xnor U6912 (N_6912,N_4861,N_4759);
xnor U6913 (N_6913,N_5178,N_3463);
nor U6914 (N_6914,N_5468,N_4556);
and U6915 (N_6915,N_3081,N_3467);
and U6916 (N_6916,N_4261,N_4542);
nand U6917 (N_6917,N_3973,N_5308);
and U6918 (N_6918,N_5881,N_5482);
or U6919 (N_6919,N_4582,N_4417);
nor U6920 (N_6920,N_4684,N_5926);
or U6921 (N_6921,N_4560,N_4333);
nor U6922 (N_6922,N_5864,N_3100);
and U6923 (N_6923,N_5256,N_3307);
or U6924 (N_6924,N_4315,N_5461);
nor U6925 (N_6925,N_5976,N_3398);
and U6926 (N_6926,N_3832,N_4099);
and U6927 (N_6927,N_5384,N_4755);
nand U6928 (N_6928,N_3974,N_3139);
or U6929 (N_6929,N_3397,N_3958);
or U6930 (N_6930,N_3004,N_4656);
nor U6931 (N_6931,N_3256,N_3194);
and U6932 (N_6932,N_4230,N_5271);
nand U6933 (N_6933,N_5424,N_4189);
nor U6934 (N_6934,N_4311,N_3643);
or U6935 (N_6935,N_4769,N_4512);
nand U6936 (N_6936,N_5152,N_5325);
and U6937 (N_6937,N_3352,N_4031);
nand U6938 (N_6938,N_5096,N_5909);
or U6939 (N_6939,N_3676,N_4173);
nor U6940 (N_6940,N_3384,N_3519);
or U6941 (N_6941,N_4411,N_5861);
nand U6942 (N_6942,N_5905,N_4037);
and U6943 (N_6943,N_4258,N_3234);
nor U6944 (N_6944,N_4642,N_4860);
and U6945 (N_6945,N_5001,N_5418);
nor U6946 (N_6946,N_5612,N_5280);
or U6947 (N_6947,N_5110,N_4186);
and U6948 (N_6948,N_3063,N_3047);
nor U6949 (N_6949,N_5027,N_3133);
nand U6950 (N_6950,N_5847,N_5743);
or U6951 (N_6951,N_3170,N_3583);
nor U6952 (N_6952,N_3834,N_5337);
nand U6953 (N_6953,N_4141,N_5897);
nor U6954 (N_6954,N_3892,N_3638);
nor U6955 (N_6955,N_5078,N_4486);
and U6956 (N_6956,N_4765,N_3199);
nand U6957 (N_6957,N_3298,N_3743);
or U6958 (N_6958,N_5977,N_4663);
nand U6959 (N_6959,N_4843,N_3854);
nand U6960 (N_6960,N_4878,N_5208);
and U6961 (N_6961,N_3367,N_5786);
and U6962 (N_6962,N_5671,N_3319);
nor U6963 (N_6963,N_3418,N_3002);
or U6964 (N_6964,N_4079,N_5860);
and U6965 (N_6965,N_4908,N_3182);
nand U6966 (N_6966,N_5106,N_4409);
and U6967 (N_6967,N_3132,N_5763);
nor U6968 (N_6968,N_5172,N_4150);
nor U6969 (N_6969,N_3831,N_4957);
or U6970 (N_6970,N_5239,N_5863);
nand U6971 (N_6971,N_3231,N_3464);
or U6972 (N_6972,N_3760,N_3040);
or U6973 (N_6973,N_5258,N_4535);
nand U6974 (N_6974,N_3801,N_4714);
or U6975 (N_6975,N_3368,N_3578);
nand U6976 (N_6976,N_5708,N_4948);
xor U6977 (N_6977,N_5596,N_3614);
nor U6978 (N_6978,N_5452,N_3322);
nand U6979 (N_6979,N_4318,N_4321);
nor U6980 (N_6980,N_5120,N_3163);
nor U6981 (N_6981,N_3381,N_4265);
or U6982 (N_6982,N_5836,N_4517);
and U6983 (N_6983,N_3107,N_5223);
nand U6984 (N_6984,N_4862,N_3593);
nor U6985 (N_6985,N_5134,N_4293);
or U6986 (N_6986,N_3781,N_4427);
nand U6987 (N_6987,N_4491,N_3498);
or U6988 (N_6988,N_3895,N_3408);
or U6989 (N_6989,N_3369,N_3431);
nand U6990 (N_6990,N_4666,N_4570);
or U6991 (N_6991,N_4845,N_4466);
and U6992 (N_6992,N_5760,N_5479);
nor U6993 (N_6993,N_3300,N_4680);
nand U6994 (N_6994,N_4731,N_3887);
nand U6995 (N_6995,N_3360,N_5757);
nor U6996 (N_6996,N_4197,N_3602);
nand U6997 (N_6997,N_4407,N_3694);
and U6998 (N_6998,N_4025,N_3695);
or U6999 (N_6999,N_3388,N_3153);
nand U7000 (N_7000,N_3803,N_5305);
or U7001 (N_7001,N_3880,N_5371);
nor U7002 (N_7002,N_3436,N_4252);
nor U7003 (N_7003,N_5677,N_5323);
or U7004 (N_7004,N_4405,N_3466);
and U7005 (N_7005,N_4885,N_4218);
or U7006 (N_7006,N_4688,N_3707);
or U7007 (N_7007,N_3808,N_3095);
nor U7008 (N_7008,N_5005,N_3118);
and U7009 (N_7009,N_3738,N_3336);
nor U7010 (N_7010,N_5494,N_4367);
nand U7011 (N_7011,N_5774,N_5674);
or U7012 (N_7012,N_3191,N_5377);
nand U7013 (N_7013,N_4329,N_4345);
nand U7014 (N_7014,N_3377,N_4095);
nor U7015 (N_7015,N_3625,N_3324);
and U7016 (N_7016,N_5157,N_5034);
or U7017 (N_7017,N_3988,N_3203);
and U7018 (N_7018,N_5787,N_5443);
nand U7019 (N_7019,N_3799,N_4898);
or U7020 (N_7020,N_4467,N_3682);
nor U7021 (N_7021,N_5265,N_4185);
nand U7022 (N_7022,N_5145,N_5886);
nor U7023 (N_7023,N_5119,N_4735);
and U7024 (N_7024,N_4775,N_4708);
nand U7025 (N_7025,N_4190,N_4116);
nand U7026 (N_7026,N_5696,N_4713);
or U7027 (N_7027,N_5474,N_3510);
nand U7028 (N_7028,N_3269,N_4397);
or U7029 (N_7029,N_3511,N_3605);
nand U7030 (N_7030,N_4015,N_3439);
nor U7031 (N_7031,N_4989,N_5948);
xor U7032 (N_7032,N_3289,N_4798);
or U7033 (N_7033,N_5736,N_4806);
nor U7034 (N_7034,N_5466,N_3563);
or U7035 (N_7035,N_3984,N_4578);
and U7036 (N_7036,N_5470,N_5254);
and U7037 (N_7037,N_5694,N_5260);
or U7038 (N_7038,N_3882,N_4063);
and U7039 (N_7039,N_5380,N_3093);
or U7040 (N_7040,N_5477,N_5015);
and U7041 (N_7041,N_4529,N_4328);
or U7042 (N_7042,N_5647,N_3819);
or U7043 (N_7043,N_3086,N_4555);
and U7044 (N_7044,N_3668,N_4307);
and U7045 (N_7045,N_5375,N_3938);
or U7046 (N_7046,N_5662,N_5249);
or U7047 (N_7047,N_3407,N_5068);
nor U7048 (N_7048,N_3910,N_5144);
and U7049 (N_7049,N_3221,N_4553);
and U7050 (N_7050,N_4312,N_5367);
nor U7051 (N_7051,N_4489,N_4269);
and U7052 (N_7052,N_3985,N_4179);
nand U7053 (N_7053,N_4353,N_5805);
nand U7054 (N_7054,N_4526,N_3514);
and U7055 (N_7055,N_4510,N_5107);
or U7056 (N_7056,N_5227,N_4664);
or U7057 (N_7057,N_4028,N_5084);
nand U7058 (N_7058,N_4459,N_4022);
nor U7059 (N_7059,N_3999,N_3782);
nand U7060 (N_7060,N_3158,N_3569);
or U7061 (N_7061,N_4975,N_4689);
nor U7062 (N_7062,N_4369,N_3306);
or U7063 (N_7063,N_3250,N_4075);
nand U7064 (N_7064,N_5834,N_3167);
or U7065 (N_7065,N_5454,N_4771);
nand U7066 (N_7066,N_4033,N_4892);
and U7067 (N_7067,N_4335,N_5022);
nand U7068 (N_7068,N_3471,N_4475);
and U7069 (N_7069,N_3896,N_3090);
or U7070 (N_7070,N_5197,N_3717);
xnor U7071 (N_7071,N_5281,N_3188);
nor U7072 (N_7072,N_5814,N_5189);
and U7073 (N_7073,N_4916,N_4484);
nor U7074 (N_7074,N_3688,N_4986);
nand U7075 (N_7075,N_3762,N_5614);
and U7076 (N_7076,N_3515,N_3166);
and U7077 (N_7077,N_4640,N_4749);
or U7078 (N_7078,N_5698,N_5115);
or U7079 (N_7079,N_3739,N_5718);
nor U7080 (N_7080,N_4358,N_5374);
or U7081 (N_7081,N_5196,N_4395);
nor U7082 (N_7082,N_4267,N_3877);
and U7083 (N_7083,N_4788,N_3941);
and U7084 (N_7084,N_4342,N_3143);
nand U7085 (N_7085,N_5495,N_5289);
nand U7086 (N_7086,N_4623,N_4032);
or U7087 (N_7087,N_4324,N_4643);
nand U7088 (N_7088,N_4303,N_3244);
nand U7089 (N_7089,N_4182,N_5767);
or U7090 (N_7090,N_4199,N_3708);
nand U7091 (N_7091,N_5996,N_4603);
nand U7092 (N_7092,N_5139,N_5176);
and U7093 (N_7093,N_5329,N_4412);
nor U7094 (N_7094,N_3264,N_4718);
nor U7095 (N_7095,N_3841,N_5492);
nor U7096 (N_7096,N_4554,N_4605);
or U7097 (N_7097,N_5965,N_3990);
nor U7098 (N_7098,N_4146,N_3853);
or U7099 (N_7099,N_5528,N_4548);
or U7100 (N_7100,N_3959,N_3884);
and U7101 (N_7101,N_3350,N_5967);
and U7102 (N_7102,N_3673,N_4136);
or U7103 (N_7103,N_5884,N_4183);
nand U7104 (N_7104,N_4837,N_4600);
and U7105 (N_7105,N_3146,N_4966);
and U7106 (N_7106,N_5739,N_3376);
or U7107 (N_7107,N_4253,N_5928);
nand U7108 (N_7108,N_4774,N_3013);
nor U7109 (N_7109,N_4433,N_4089);
nand U7110 (N_7110,N_5379,N_3288);
xnor U7111 (N_7111,N_4464,N_3737);
and U7112 (N_7112,N_3157,N_4375);
xor U7113 (N_7113,N_4248,N_4246);
or U7114 (N_7114,N_3401,N_5795);
nand U7115 (N_7115,N_5986,N_4609);
or U7116 (N_7116,N_5359,N_3131);
and U7117 (N_7117,N_3718,N_3653);
nor U7118 (N_7118,N_3420,N_5385);
nand U7119 (N_7119,N_3226,N_4576);
nor U7120 (N_7120,N_3071,N_3114);
and U7121 (N_7121,N_5273,N_4812);
nor U7122 (N_7122,N_5943,N_5908);
and U7123 (N_7123,N_3893,N_4744);
nand U7124 (N_7124,N_5349,N_4081);
xnor U7125 (N_7125,N_3080,N_3948);
nand U7126 (N_7126,N_4776,N_3997);
nand U7127 (N_7127,N_3315,N_5882);
or U7128 (N_7128,N_5749,N_4052);
nand U7129 (N_7129,N_3138,N_5141);
nor U7130 (N_7130,N_4214,N_5607);
or U7131 (N_7131,N_3813,N_4561);
nand U7132 (N_7132,N_5082,N_3520);
nor U7133 (N_7133,N_3390,N_3812);
and U7134 (N_7134,N_4477,N_5673);
nor U7135 (N_7135,N_3859,N_3889);
nor U7136 (N_7136,N_5933,N_3755);
xor U7137 (N_7137,N_4902,N_3968);
xnor U7138 (N_7138,N_4138,N_4096);
nor U7139 (N_7139,N_3123,N_4474);
and U7140 (N_7140,N_4424,N_3374);
and U7141 (N_7141,N_3784,N_4811);
nor U7142 (N_7142,N_3844,N_5620);
nand U7143 (N_7143,N_5290,N_4627);
nor U7144 (N_7144,N_4224,N_3448);
or U7145 (N_7145,N_4006,N_5264);
nor U7146 (N_7146,N_4004,N_5333);
or U7147 (N_7147,N_4763,N_4691);
and U7148 (N_7148,N_3150,N_5081);
nor U7149 (N_7149,N_5530,N_4897);
or U7150 (N_7150,N_4131,N_5369);
and U7151 (N_7151,N_3254,N_5738);
or U7152 (N_7152,N_3115,N_5124);
or U7153 (N_7153,N_4274,N_5537);
and U7154 (N_7154,N_5438,N_5628);
nor U7155 (N_7155,N_4809,N_4998);
or U7156 (N_7156,N_4678,N_3285);
nor U7157 (N_7157,N_4953,N_3919);
nor U7158 (N_7158,N_5566,N_3417);
or U7159 (N_7159,N_4053,N_5534);
nand U7160 (N_7160,N_4895,N_4671);
or U7161 (N_7161,N_5193,N_3079);
nand U7162 (N_7162,N_4571,N_3779);
nand U7163 (N_7163,N_5913,N_4930);
nor U7164 (N_7164,N_5147,N_3517);
nand U7165 (N_7165,N_4034,N_4668);
nand U7166 (N_7166,N_5539,N_3639);
nor U7167 (N_7167,N_3356,N_3007);
and U7168 (N_7168,N_5180,N_3200);
or U7169 (N_7169,N_5598,N_5164);
xnor U7170 (N_7170,N_4751,N_3954);
nand U7171 (N_7171,N_5542,N_3649);
and U7172 (N_7172,N_3648,N_5460);
and U7173 (N_7173,N_4630,N_5363);
nor U7174 (N_7174,N_4817,N_5116);
and U7175 (N_7175,N_3626,N_4344);
nor U7176 (N_7176,N_4235,N_5109);
and U7177 (N_7177,N_3316,N_5404);
nand U7178 (N_7178,N_5421,N_4924);
or U7179 (N_7179,N_5831,N_5686);
nand U7180 (N_7180,N_3630,N_5827);
nand U7181 (N_7181,N_4241,N_3055);
nor U7182 (N_7182,N_4371,N_4326);
and U7183 (N_7183,N_5916,N_4125);
nand U7184 (N_7184,N_4738,N_3744);
xnor U7185 (N_7185,N_5762,N_4207);
nor U7186 (N_7186,N_3632,N_3660);
and U7187 (N_7187,N_3097,N_4101);
nand U7188 (N_7188,N_5122,N_4452);
nand U7189 (N_7189,N_3661,N_4528);
and U7190 (N_7190,N_5778,N_5833);
and U7191 (N_7191,N_5964,N_5875);
nor U7192 (N_7192,N_3193,N_5963);
or U7193 (N_7193,N_5415,N_3449);
and U7194 (N_7194,N_5285,N_4638);
nand U7195 (N_7195,N_5126,N_3996);
nor U7196 (N_7196,N_5835,N_5291);
nor U7197 (N_7197,N_5283,N_5602);
and U7198 (N_7198,N_4752,N_4574);
nand U7199 (N_7199,N_3553,N_3952);
nor U7200 (N_7200,N_3802,N_3685);
and U7201 (N_7201,N_3358,N_5267);
or U7202 (N_7202,N_3084,N_4286);
nor U7203 (N_7203,N_5245,N_3788);
or U7204 (N_7204,N_5910,N_4017);
or U7205 (N_7205,N_5073,N_4772);
and U7206 (N_7206,N_5161,N_5462);
nor U7207 (N_7207,N_5192,N_5037);
or U7208 (N_7208,N_5667,N_5346);
nand U7209 (N_7209,N_5355,N_3570);
or U7210 (N_7210,N_5381,N_3313);
nand U7211 (N_7211,N_5469,N_4836);
nand U7212 (N_7212,N_3105,N_4854);
or U7213 (N_7213,N_4667,N_5269);
xor U7214 (N_7214,N_3312,N_3135);
nor U7215 (N_7215,N_3983,N_4711);
and U7216 (N_7216,N_5184,N_5695);
and U7217 (N_7217,N_4780,N_5715);
nor U7218 (N_7218,N_4530,N_3731);
and U7219 (N_7219,N_4237,N_5784);
nand U7220 (N_7220,N_5311,N_4030);
or U7221 (N_7221,N_5018,N_5378);
nand U7222 (N_7222,N_5356,N_4449);
and U7223 (N_7223,N_4767,N_5812);
and U7224 (N_7224,N_3864,N_5481);
and U7225 (N_7225,N_3219,N_4165);
nor U7226 (N_7226,N_5632,N_5877);
nor U7227 (N_7227,N_4670,N_4568);
and U7228 (N_7228,N_3265,N_3712);
nor U7229 (N_7229,N_4317,N_3099);
and U7230 (N_7230,N_3642,N_3608);
nand U7231 (N_7231,N_4562,N_3016);
nand U7232 (N_7232,N_5163,N_5723);
nor U7233 (N_7233,N_5294,N_3050);
nor U7234 (N_7234,N_4626,N_4471);
nor U7235 (N_7235,N_4919,N_3850);
xnor U7236 (N_7236,N_3926,N_4368);
nor U7237 (N_7237,N_3787,N_5049);
or U7238 (N_7238,N_3557,N_3255);
nor U7239 (N_7239,N_4255,N_5917);
nand U7240 (N_7240,N_4662,N_5697);
and U7241 (N_7241,N_5712,N_4868);
and U7242 (N_7242,N_4814,N_5871);
and U7243 (N_7243,N_3565,N_4239);
or U7244 (N_7244,N_4790,N_5137);
nand U7245 (N_7245,N_4720,N_3924);
nand U7246 (N_7246,N_4747,N_3875);
nor U7247 (N_7247,N_3427,N_4783);
nor U7248 (N_7248,N_5445,N_3228);
or U7249 (N_7249,N_3154,N_4891);
and U7250 (N_7250,N_4080,N_3435);
and U7251 (N_7251,N_5000,N_4770);
and U7252 (N_7252,N_5777,N_4287);
xnor U7253 (N_7253,N_5547,N_5601);
nand U7254 (N_7254,N_5744,N_5660);
nand U7255 (N_7255,N_3994,N_4208);
nor U7256 (N_7256,N_4064,N_5103);
nor U7257 (N_7257,N_5165,N_4598);
nand U7258 (N_7258,N_4804,N_5232);
nand U7259 (N_7259,N_3272,N_5143);
nor U7260 (N_7260,N_3827,N_4550);
or U7261 (N_7261,N_4171,N_4698);
or U7262 (N_7262,N_5973,N_4633);
nand U7263 (N_7263,N_3330,N_5259);
and U7264 (N_7264,N_4787,N_5799);
or U7265 (N_7265,N_3501,N_4842);
or U7266 (N_7266,N_5368,N_5540);
nor U7267 (N_7267,N_5907,N_3195);
or U7268 (N_7268,N_3321,N_5150);
nand U7269 (N_7269,N_5444,N_3127);
nor U7270 (N_7270,N_5194,N_4793);
or U7271 (N_7271,N_5806,N_4195);
nor U7272 (N_7272,N_4883,N_4110);
and U7273 (N_7273,N_5693,N_5142);
nand U7274 (N_7274,N_3757,N_3929);
and U7275 (N_7275,N_4696,N_3364);
nor U7276 (N_7276,N_3456,N_3576);
or U7277 (N_7277,N_3820,N_5575);
and U7278 (N_7278,N_3216,N_4773);
or U7279 (N_7279,N_4108,N_4616);
and U7280 (N_7280,N_3871,N_4354);
nor U7281 (N_7281,N_5862,N_4754);
and U7282 (N_7282,N_5829,N_4687);
nand U7283 (N_7283,N_5211,N_5706);
nor U7284 (N_7284,N_3886,N_5493);
nand U7285 (N_7285,N_3766,N_4866);
nor U7286 (N_7286,N_3554,N_5604);
nor U7287 (N_7287,N_4180,N_5400);
and U7288 (N_7288,N_4294,N_5950);
and U7289 (N_7289,N_3019,N_5648);
nor U7290 (N_7290,N_5458,N_3486);
nor U7291 (N_7291,N_4480,N_4198);
or U7292 (N_7292,N_4745,N_4631);
and U7293 (N_7293,N_5459,N_4323);
nor U7294 (N_7294,N_5968,N_4834);
nand U7295 (N_7295,N_3905,N_5250);
nand U7296 (N_7296,N_5953,N_3229);
nor U7297 (N_7297,N_4669,N_4011);
and U7298 (N_7298,N_5978,N_5218);
nand U7299 (N_7299,N_4985,N_4941);
and U7300 (N_7300,N_5314,N_4617);
or U7301 (N_7301,N_4917,N_3901);
xnor U7302 (N_7302,N_4114,N_5428);
and U7303 (N_7303,N_4974,N_4622);
or U7304 (N_7304,N_3607,N_5076);
and U7305 (N_7305,N_4513,N_3066);
and U7306 (N_7306,N_4349,N_3711);
or U7307 (N_7307,N_3462,N_3568);
or U7308 (N_7308,N_4434,N_4521);
and U7309 (N_7309,N_5087,N_5025);
and U7310 (N_7310,N_5393,N_5652);
nand U7311 (N_7311,N_4723,N_3714);
nand U7312 (N_7312,N_3474,N_5200);
or U7313 (N_7313,N_4761,N_4782);
and U7314 (N_7314,N_4408,N_3579);
or U7315 (N_7315,N_5248,N_4647);
nand U7316 (N_7316,N_4247,N_5545);
nand U7317 (N_7317,N_5713,N_3478);
or U7318 (N_7318,N_5640,N_4557);
nor U7319 (N_7319,N_3190,N_5041);
nand U7320 (N_7320,N_5941,N_3503);
and U7321 (N_7321,N_4428,N_3636);
or U7322 (N_7322,N_5919,N_3239);
nor U7323 (N_7323,N_5868,N_4514);
nor U7324 (N_7324,N_4137,N_4254);
or U7325 (N_7325,N_5491,N_5336);
nand U7326 (N_7326,N_4244,N_5536);
xor U7327 (N_7327,N_4661,N_3656);
or U7328 (N_7328,N_4498,N_5794);
or U7329 (N_7329,N_5464,N_5050);
nand U7330 (N_7330,N_4874,N_3791);
nand U7331 (N_7331,N_3000,N_3220);
nand U7332 (N_7332,N_3572,N_5220);
nor U7333 (N_7333,N_5906,N_3394);
xor U7334 (N_7334,N_3978,N_3185);
and U7335 (N_7335,N_4155,N_3057);
nand U7336 (N_7336,N_4314,N_5856);
nor U7337 (N_7337,N_5274,N_5561);
and U7338 (N_7338,N_3933,N_3915);
nor U7339 (N_7339,N_3473,N_3469);
nand U7340 (N_7340,N_5296,N_5981);
or U7341 (N_7341,N_3991,N_4867);
and U7342 (N_7342,N_4589,N_5268);
nor U7343 (N_7343,N_4362,N_5016);
nand U7344 (N_7344,N_3825,N_5312);
nor U7345 (N_7345,N_5417,N_4213);
or U7346 (N_7346,N_5051,N_5960);
or U7347 (N_7347,N_4499,N_3535);
and U7348 (N_7348,N_5514,N_3284);
nand U7349 (N_7349,N_3293,N_5764);
and U7350 (N_7350,N_3640,N_3821);
or U7351 (N_7351,N_5526,N_5568);
or U7352 (N_7352,N_3495,N_3224);
nor U7353 (N_7353,N_3432,N_4140);
or U7354 (N_7354,N_4903,N_3856);
nor U7355 (N_7355,N_4439,N_3064);
nor U7356 (N_7356,N_3017,N_5175);
or U7357 (N_7357,N_5633,N_4132);
and U7358 (N_7358,N_3849,N_3716);
or U7359 (N_7359,N_4040,N_5742);
nor U7360 (N_7360,N_4352,N_5328);
and U7361 (N_7361,N_3904,N_4092);
xnor U7362 (N_7362,N_3971,N_4699);
nor U7363 (N_7363,N_5024,N_5858);
nand U7364 (N_7364,N_4003,N_3912);
nand U7365 (N_7365,N_3365,N_5748);
or U7366 (N_7366,N_4864,N_5031);
nor U7367 (N_7367,N_5017,N_4302);
and U7368 (N_7368,N_4331,N_4728);
or U7369 (N_7369,N_3173,N_4085);
and U7370 (N_7370,N_5409,N_5629);
and U7371 (N_7371,N_4201,N_3359);
nor U7372 (N_7372,N_4334,N_3035);
or U7373 (N_7373,N_3343,N_5307);
and U7374 (N_7374,N_3747,N_5588);
nor U7375 (N_7375,N_4158,N_5476);
xor U7376 (N_7376,N_4174,N_3437);
or U7377 (N_7377,N_4839,N_3588);
or U7378 (N_7378,N_4300,N_4074);
or U7379 (N_7379,N_3412,N_3472);
nor U7380 (N_7380,N_4918,N_3232);
nor U7381 (N_7381,N_3533,N_4800);
and U7382 (N_7382,N_4496,N_4332);
nor U7383 (N_7383,N_4492,N_3375);
nand U7384 (N_7384,N_3696,N_4238);
and U7385 (N_7385,N_5395,N_5902);
or U7386 (N_7386,N_4014,N_5233);
nor U7387 (N_7387,N_3372,N_5929);
or U7388 (N_7388,N_3589,N_4242);
nor U7389 (N_7389,N_5221,N_5966);
nor U7390 (N_7390,N_4565,N_3085);
nor U7391 (N_7391,N_3487,N_3480);
nand U7392 (N_7392,N_3544,N_3771);
or U7393 (N_7393,N_4815,N_4356);
nand U7394 (N_7394,N_4106,N_5174);
and U7395 (N_7395,N_3980,N_3911);
and U7396 (N_7396,N_4112,N_4734);
nor U7397 (N_7397,N_3935,N_3909);
and U7398 (N_7398,N_4832,N_4450);
and U7399 (N_7399,N_5171,N_3591);
and U7400 (N_7400,N_3262,N_5699);
nand U7401 (N_7401,N_4602,N_5873);
nand U7402 (N_7402,N_5387,N_4500);
or U7403 (N_7403,N_3036,N_5478);
nand U7404 (N_7404,N_5519,N_3943);
nor U7405 (N_7405,N_3218,N_5619);
nor U7406 (N_7406,N_5567,N_4076);
and U7407 (N_7407,N_3396,N_4442);
nand U7408 (N_7408,N_3748,N_4055);
and U7409 (N_7409,N_4176,N_5689);
and U7410 (N_7410,N_3542,N_3393);
nand U7411 (N_7411,N_5222,N_5099);
nor U7412 (N_7412,N_5423,N_4282);
and U7413 (N_7413,N_3809,N_4509);
or U7414 (N_7414,N_5985,N_3571);
or U7415 (N_7415,N_5741,N_3981);
nand U7416 (N_7416,N_5186,N_3970);
and U7417 (N_7417,N_4963,N_4107);
or U7418 (N_7418,N_4590,N_4921);
or U7419 (N_7419,N_4757,N_5685);
nor U7420 (N_7420,N_3317,N_5338);
nor U7421 (N_7421,N_4920,N_5408);
or U7422 (N_7422,N_5092,N_4715);
nor U7423 (N_7423,N_5564,N_4748);
nand U7424 (N_7424,N_3509,N_5572);
or U7425 (N_7425,N_4073,N_4382);
nor U7426 (N_7426,N_5301,N_3745);
nand U7427 (N_7427,N_3932,N_3906);
and U7428 (N_7428,N_5127,N_3310);
nor U7429 (N_7429,N_5436,N_4217);
nor U7430 (N_7430,N_5912,N_3868);
xnor U7431 (N_7431,N_4251,N_4601);
nor U7432 (N_7432,N_3354,N_5067);
and U7433 (N_7433,N_3479,N_5483);
nor U7434 (N_7434,N_5364,N_4607);
and U7435 (N_7435,N_3598,N_5298);
nand U7436 (N_7436,N_5238,N_3505);
nand U7437 (N_7437,N_3558,N_5844);
or U7438 (N_7438,N_5538,N_4822);
nor U7439 (N_7439,N_4871,N_4292);
or U7440 (N_7440,N_3380,N_4306);
nand U7441 (N_7441,N_3811,N_5755);
or U7442 (N_7442,N_4896,N_4016);
nand U7443 (N_7443,N_3524,N_5747);
nor U7444 (N_7444,N_5869,N_3301);
or U7445 (N_7445,N_5361,N_4071);
nor U7446 (N_7446,N_3021,N_5556);
nor U7447 (N_7447,N_4729,N_3767);
nor U7448 (N_7448,N_4374,N_3795);
and U7449 (N_7449,N_3592,N_3993);
or U7450 (N_7450,N_4503,N_3543);
or U7451 (N_7451,N_5471,N_5544);
nand U7452 (N_7452,N_4596,N_4388);
nor U7453 (N_7453,N_5974,N_4431);
and U7454 (N_7454,N_4939,N_3311);
nand U7455 (N_7455,N_5286,N_3130);
and U7456 (N_7456,N_4364,N_4243);
and U7457 (N_7457,N_3065,N_4256);
nand U7458 (N_7458,N_4149,N_4890);
or U7459 (N_7459,N_3258,N_5465);
and U7460 (N_7460,N_4133,N_5074);
nor U7461 (N_7461,N_5097,N_3299);
nor U7462 (N_7462,N_4672,N_5717);
nand U7463 (N_7463,N_4338,N_4098);
nand U7464 (N_7464,N_3314,N_4263);
or U7465 (N_7465,N_5773,N_5313);
or U7466 (N_7466,N_5058,N_3523);
or U7467 (N_7467,N_4476,N_4882);
nor U7468 (N_7468,N_3179,N_3223);
nand U7469 (N_7469,N_5064,N_4443);
and U7470 (N_7470,N_4615,N_5207);
and U7471 (N_7471,N_5982,N_5574);
or U7472 (N_7472,N_3734,N_5867);
nor U7473 (N_7473,N_5292,N_3197);
nor U7474 (N_7474,N_4927,N_4940);
nand U7475 (N_7475,N_4005,N_3617);
nor U7476 (N_7476,N_3014,N_5600);
or U7477 (N_7477,N_5634,N_5830);
nand U7478 (N_7478,N_5247,N_5615);
or U7479 (N_7479,N_5516,N_4383);
and U7480 (N_7480,N_3426,N_4873);
and U7481 (N_7481,N_4272,N_5132);
nor U7482 (N_7482,N_3527,N_4152);
and U7483 (N_7483,N_5195,N_3241);
nand U7484 (N_7484,N_3345,N_4929);
xor U7485 (N_7485,N_4984,N_4888);
or U7486 (N_7486,N_5630,N_4973);
nor U7487 (N_7487,N_3483,N_5300);
nand U7488 (N_7488,N_3500,N_3447);
nor U7489 (N_7489,N_5111,N_4212);
nand U7490 (N_7490,N_4143,N_5924);
or U7491 (N_7491,N_4789,N_4889);
nor U7492 (N_7492,N_4766,N_5901);
nor U7493 (N_7493,N_3567,N_3069);
nor U7494 (N_7494,N_4175,N_4523);
nor U7495 (N_7495,N_3763,N_5842);
nand U7496 (N_7496,N_5009,N_5427);
and U7497 (N_7497,N_3861,N_4461);
nor U7498 (N_7498,N_5439,N_3072);
and U7499 (N_7499,N_5586,N_5240);
and U7500 (N_7500,N_4286,N_3248);
xnor U7501 (N_7501,N_3358,N_4288);
nand U7502 (N_7502,N_3869,N_5617);
or U7503 (N_7503,N_4862,N_4013);
nand U7504 (N_7504,N_5000,N_5265);
nor U7505 (N_7505,N_5052,N_4792);
and U7506 (N_7506,N_5521,N_4275);
nor U7507 (N_7507,N_3787,N_3140);
nand U7508 (N_7508,N_3815,N_4220);
nor U7509 (N_7509,N_4350,N_4517);
nand U7510 (N_7510,N_4399,N_5683);
nand U7511 (N_7511,N_4053,N_5709);
nand U7512 (N_7512,N_3614,N_5118);
or U7513 (N_7513,N_4376,N_4103);
xnor U7514 (N_7514,N_5627,N_5333);
and U7515 (N_7515,N_4719,N_4099);
and U7516 (N_7516,N_3779,N_5646);
or U7517 (N_7517,N_4373,N_4395);
and U7518 (N_7518,N_4557,N_4094);
xor U7519 (N_7519,N_4500,N_5317);
and U7520 (N_7520,N_5007,N_4448);
nor U7521 (N_7521,N_3814,N_4344);
nand U7522 (N_7522,N_4038,N_4364);
nor U7523 (N_7523,N_4866,N_3746);
nor U7524 (N_7524,N_4138,N_5570);
nor U7525 (N_7525,N_5481,N_5325);
nand U7526 (N_7526,N_3025,N_5239);
or U7527 (N_7527,N_5794,N_4790);
and U7528 (N_7528,N_4089,N_3400);
or U7529 (N_7529,N_4169,N_3601);
and U7530 (N_7530,N_3103,N_3242);
or U7531 (N_7531,N_4612,N_4734);
nand U7532 (N_7532,N_4211,N_5892);
nand U7533 (N_7533,N_4203,N_5960);
and U7534 (N_7534,N_4548,N_4998);
and U7535 (N_7535,N_4516,N_5985);
and U7536 (N_7536,N_5735,N_4824);
and U7537 (N_7537,N_4901,N_4948);
and U7538 (N_7538,N_3053,N_3467);
or U7539 (N_7539,N_3734,N_5940);
nor U7540 (N_7540,N_4654,N_4206);
nor U7541 (N_7541,N_4209,N_3800);
and U7542 (N_7542,N_3010,N_4553);
or U7543 (N_7543,N_5168,N_3298);
nand U7544 (N_7544,N_5518,N_4872);
and U7545 (N_7545,N_5705,N_4244);
xnor U7546 (N_7546,N_5119,N_4382);
nand U7547 (N_7547,N_4113,N_3601);
nand U7548 (N_7548,N_5240,N_3271);
and U7549 (N_7549,N_3314,N_5839);
or U7550 (N_7550,N_4553,N_4349);
nand U7551 (N_7551,N_4331,N_3086);
or U7552 (N_7552,N_3927,N_5282);
or U7553 (N_7553,N_5368,N_4876);
and U7554 (N_7554,N_5011,N_3232);
nor U7555 (N_7555,N_3417,N_4442);
and U7556 (N_7556,N_3004,N_3788);
or U7557 (N_7557,N_3308,N_4062);
nor U7558 (N_7558,N_4559,N_4581);
and U7559 (N_7559,N_3200,N_5682);
or U7560 (N_7560,N_4160,N_3943);
and U7561 (N_7561,N_4854,N_5498);
nand U7562 (N_7562,N_4202,N_4556);
nand U7563 (N_7563,N_5215,N_3029);
nand U7564 (N_7564,N_3090,N_5761);
nor U7565 (N_7565,N_3923,N_3896);
nand U7566 (N_7566,N_4786,N_3012);
nor U7567 (N_7567,N_5169,N_4975);
and U7568 (N_7568,N_4310,N_4854);
nand U7569 (N_7569,N_4623,N_3817);
nand U7570 (N_7570,N_5725,N_4733);
xor U7571 (N_7571,N_5610,N_4570);
and U7572 (N_7572,N_5091,N_5723);
xnor U7573 (N_7573,N_5983,N_5021);
and U7574 (N_7574,N_3813,N_5965);
nand U7575 (N_7575,N_4666,N_4267);
or U7576 (N_7576,N_5205,N_4402);
nor U7577 (N_7577,N_4167,N_5513);
nand U7578 (N_7578,N_4288,N_4394);
or U7579 (N_7579,N_3237,N_3229);
nor U7580 (N_7580,N_5963,N_3195);
or U7581 (N_7581,N_5293,N_4783);
nor U7582 (N_7582,N_3922,N_3387);
nor U7583 (N_7583,N_4601,N_5567);
nand U7584 (N_7584,N_4869,N_4348);
nor U7585 (N_7585,N_3970,N_3804);
nand U7586 (N_7586,N_4917,N_5434);
or U7587 (N_7587,N_3172,N_5737);
nor U7588 (N_7588,N_5427,N_4533);
nand U7589 (N_7589,N_3176,N_4460);
nand U7590 (N_7590,N_3797,N_5019);
nor U7591 (N_7591,N_3123,N_5639);
xor U7592 (N_7592,N_5730,N_3320);
or U7593 (N_7593,N_5134,N_4911);
nor U7594 (N_7594,N_4257,N_3739);
and U7595 (N_7595,N_4868,N_4568);
nor U7596 (N_7596,N_5725,N_5191);
or U7597 (N_7597,N_4091,N_4900);
nor U7598 (N_7598,N_5909,N_4094);
nor U7599 (N_7599,N_5128,N_5668);
nand U7600 (N_7600,N_3722,N_5677);
nand U7601 (N_7601,N_3444,N_4985);
or U7602 (N_7602,N_5174,N_4699);
and U7603 (N_7603,N_3135,N_3285);
and U7604 (N_7604,N_4841,N_3116);
xor U7605 (N_7605,N_3208,N_3876);
nand U7606 (N_7606,N_3193,N_5866);
nor U7607 (N_7607,N_3984,N_3964);
nor U7608 (N_7608,N_4782,N_3797);
xor U7609 (N_7609,N_5787,N_5745);
or U7610 (N_7610,N_4004,N_4349);
and U7611 (N_7611,N_5559,N_4373);
nand U7612 (N_7612,N_4872,N_4801);
nand U7613 (N_7613,N_5596,N_4983);
xnor U7614 (N_7614,N_3872,N_4805);
or U7615 (N_7615,N_5618,N_5721);
or U7616 (N_7616,N_5952,N_4072);
nor U7617 (N_7617,N_5042,N_3880);
nand U7618 (N_7618,N_5867,N_5780);
nand U7619 (N_7619,N_4148,N_4795);
nand U7620 (N_7620,N_4103,N_3535);
nor U7621 (N_7621,N_4355,N_5712);
nor U7622 (N_7622,N_5362,N_5374);
nor U7623 (N_7623,N_4612,N_5550);
and U7624 (N_7624,N_3219,N_4379);
or U7625 (N_7625,N_4712,N_5912);
nand U7626 (N_7626,N_4806,N_3952);
or U7627 (N_7627,N_5089,N_3183);
or U7628 (N_7628,N_3949,N_3449);
nand U7629 (N_7629,N_4834,N_3484);
nand U7630 (N_7630,N_5472,N_5652);
nand U7631 (N_7631,N_3207,N_3216);
nor U7632 (N_7632,N_5027,N_3524);
or U7633 (N_7633,N_3449,N_4850);
nor U7634 (N_7634,N_4803,N_3922);
nand U7635 (N_7635,N_4680,N_5840);
nor U7636 (N_7636,N_4998,N_3353);
or U7637 (N_7637,N_5323,N_4260);
nand U7638 (N_7638,N_4993,N_3454);
or U7639 (N_7639,N_5686,N_5132);
and U7640 (N_7640,N_4804,N_5857);
or U7641 (N_7641,N_5213,N_3355);
nand U7642 (N_7642,N_4241,N_5036);
and U7643 (N_7643,N_4014,N_3414);
xor U7644 (N_7644,N_3088,N_4558);
and U7645 (N_7645,N_5891,N_5934);
nand U7646 (N_7646,N_3722,N_3183);
nand U7647 (N_7647,N_5408,N_3740);
and U7648 (N_7648,N_4593,N_3086);
nor U7649 (N_7649,N_4249,N_4821);
nor U7650 (N_7650,N_4877,N_4129);
nand U7651 (N_7651,N_3023,N_3668);
nand U7652 (N_7652,N_3033,N_5141);
nand U7653 (N_7653,N_3907,N_4163);
and U7654 (N_7654,N_5825,N_5916);
nor U7655 (N_7655,N_3488,N_3259);
nor U7656 (N_7656,N_3965,N_4688);
or U7657 (N_7657,N_3008,N_3960);
or U7658 (N_7658,N_5424,N_4960);
or U7659 (N_7659,N_3387,N_4543);
and U7660 (N_7660,N_3445,N_5122);
nand U7661 (N_7661,N_5971,N_5250);
or U7662 (N_7662,N_3457,N_3285);
nand U7663 (N_7663,N_3274,N_5406);
and U7664 (N_7664,N_5043,N_4695);
or U7665 (N_7665,N_4164,N_4217);
nor U7666 (N_7666,N_5031,N_5134);
nor U7667 (N_7667,N_4610,N_3565);
nor U7668 (N_7668,N_4206,N_4377);
nor U7669 (N_7669,N_5424,N_5396);
nor U7670 (N_7670,N_3220,N_4216);
nand U7671 (N_7671,N_4047,N_5374);
or U7672 (N_7672,N_3014,N_5039);
or U7673 (N_7673,N_5995,N_3802);
xnor U7674 (N_7674,N_3655,N_4325);
nand U7675 (N_7675,N_5100,N_5647);
and U7676 (N_7676,N_3995,N_3856);
and U7677 (N_7677,N_4692,N_4506);
or U7678 (N_7678,N_5954,N_5385);
or U7679 (N_7679,N_3835,N_5684);
and U7680 (N_7680,N_5456,N_3168);
xnor U7681 (N_7681,N_5996,N_4693);
and U7682 (N_7682,N_4812,N_5974);
or U7683 (N_7683,N_4654,N_4281);
nand U7684 (N_7684,N_5037,N_4607);
nand U7685 (N_7685,N_4490,N_4552);
nand U7686 (N_7686,N_4404,N_4468);
and U7687 (N_7687,N_3920,N_3686);
and U7688 (N_7688,N_4210,N_4115);
and U7689 (N_7689,N_5285,N_5748);
and U7690 (N_7690,N_3557,N_3964);
nand U7691 (N_7691,N_3547,N_5778);
and U7692 (N_7692,N_4029,N_3249);
or U7693 (N_7693,N_3183,N_3800);
or U7694 (N_7694,N_5040,N_3278);
and U7695 (N_7695,N_5844,N_5428);
nand U7696 (N_7696,N_5191,N_4846);
nand U7697 (N_7697,N_4989,N_4355);
and U7698 (N_7698,N_5321,N_4290);
nand U7699 (N_7699,N_5146,N_4280);
or U7700 (N_7700,N_4035,N_4536);
and U7701 (N_7701,N_5712,N_5005);
nor U7702 (N_7702,N_5547,N_4618);
nand U7703 (N_7703,N_5899,N_4410);
and U7704 (N_7704,N_3438,N_4197);
and U7705 (N_7705,N_3328,N_3122);
nor U7706 (N_7706,N_4188,N_5701);
or U7707 (N_7707,N_4279,N_3264);
or U7708 (N_7708,N_4003,N_4341);
or U7709 (N_7709,N_5015,N_5643);
or U7710 (N_7710,N_3897,N_5197);
and U7711 (N_7711,N_5221,N_3234);
or U7712 (N_7712,N_5782,N_3137);
nor U7713 (N_7713,N_3326,N_3075);
or U7714 (N_7714,N_3182,N_4122);
xnor U7715 (N_7715,N_3965,N_4659);
nand U7716 (N_7716,N_3619,N_5941);
or U7717 (N_7717,N_3082,N_3832);
nor U7718 (N_7718,N_5353,N_3759);
xor U7719 (N_7719,N_3614,N_4358);
and U7720 (N_7720,N_5035,N_3944);
nand U7721 (N_7721,N_5446,N_3361);
nor U7722 (N_7722,N_5490,N_5569);
or U7723 (N_7723,N_4756,N_4505);
or U7724 (N_7724,N_5634,N_3884);
nand U7725 (N_7725,N_3762,N_5685);
nor U7726 (N_7726,N_5537,N_4902);
and U7727 (N_7727,N_5182,N_4628);
nand U7728 (N_7728,N_4690,N_4660);
nand U7729 (N_7729,N_4744,N_4468);
nand U7730 (N_7730,N_5908,N_4495);
nand U7731 (N_7731,N_3752,N_5930);
and U7732 (N_7732,N_5125,N_5017);
or U7733 (N_7733,N_3604,N_3783);
nor U7734 (N_7734,N_3756,N_5034);
and U7735 (N_7735,N_4916,N_4709);
nand U7736 (N_7736,N_3226,N_5740);
nand U7737 (N_7737,N_4678,N_4323);
nor U7738 (N_7738,N_5164,N_3033);
nor U7739 (N_7739,N_4687,N_4149);
nor U7740 (N_7740,N_4847,N_3973);
and U7741 (N_7741,N_5775,N_4022);
or U7742 (N_7742,N_5509,N_5422);
xor U7743 (N_7743,N_4821,N_4827);
or U7744 (N_7744,N_3667,N_5008);
and U7745 (N_7745,N_3524,N_5090);
or U7746 (N_7746,N_4728,N_5201);
nand U7747 (N_7747,N_4324,N_4373);
and U7748 (N_7748,N_4814,N_3074);
nand U7749 (N_7749,N_3052,N_3479);
and U7750 (N_7750,N_5244,N_3732);
or U7751 (N_7751,N_3853,N_5091);
xnor U7752 (N_7752,N_5536,N_5743);
xnor U7753 (N_7753,N_4601,N_5973);
nor U7754 (N_7754,N_4172,N_5037);
and U7755 (N_7755,N_5153,N_5301);
nor U7756 (N_7756,N_3702,N_5112);
nor U7757 (N_7757,N_5487,N_5717);
and U7758 (N_7758,N_5191,N_5768);
or U7759 (N_7759,N_5141,N_5138);
or U7760 (N_7760,N_3441,N_4442);
nor U7761 (N_7761,N_5440,N_3936);
and U7762 (N_7762,N_3967,N_3199);
nand U7763 (N_7763,N_5756,N_5005);
nand U7764 (N_7764,N_3496,N_4389);
or U7765 (N_7765,N_4745,N_4530);
or U7766 (N_7766,N_4616,N_4343);
or U7767 (N_7767,N_4149,N_3412);
or U7768 (N_7768,N_4821,N_4241);
or U7769 (N_7769,N_4040,N_5453);
nor U7770 (N_7770,N_5752,N_4646);
nor U7771 (N_7771,N_3030,N_4763);
nand U7772 (N_7772,N_3209,N_3119);
nand U7773 (N_7773,N_3715,N_3457);
and U7774 (N_7774,N_3022,N_5322);
nor U7775 (N_7775,N_5406,N_3028);
nor U7776 (N_7776,N_4922,N_3124);
or U7777 (N_7777,N_5809,N_4377);
nor U7778 (N_7778,N_5491,N_4211);
nor U7779 (N_7779,N_4187,N_4119);
nor U7780 (N_7780,N_4608,N_5767);
nor U7781 (N_7781,N_3796,N_4253);
or U7782 (N_7782,N_5920,N_5760);
or U7783 (N_7783,N_5814,N_4041);
nand U7784 (N_7784,N_3239,N_3822);
or U7785 (N_7785,N_5167,N_3290);
nor U7786 (N_7786,N_5455,N_4332);
nor U7787 (N_7787,N_5543,N_4953);
nor U7788 (N_7788,N_4938,N_5616);
xnor U7789 (N_7789,N_3333,N_5535);
or U7790 (N_7790,N_4620,N_4305);
or U7791 (N_7791,N_3511,N_5741);
and U7792 (N_7792,N_3985,N_5533);
and U7793 (N_7793,N_4968,N_3276);
or U7794 (N_7794,N_5042,N_3768);
and U7795 (N_7795,N_3429,N_4860);
xnor U7796 (N_7796,N_5301,N_3387);
or U7797 (N_7797,N_4111,N_4404);
nand U7798 (N_7798,N_3543,N_5462);
nand U7799 (N_7799,N_4792,N_4094);
and U7800 (N_7800,N_4928,N_3683);
and U7801 (N_7801,N_3852,N_4496);
nand U7802 (N_7802,N_4089,N_3086);
or U7803 (N_7803,N_5725,N_4575);
and U7804 (N_7804,N_4487,N_5968);
nand U7805 (N_7805,N_4733,N_4233);
or U7806 (N_7806,N_4857,N_4020);
nor U7807 (N_7807,N_4200,N_4633);
nand U7808 (N_7808,N_4450,N_5040);
nor U7809 (N_7809,N_3008,N_5624);
nand U7810 (N_7810,N_5305,N_4055);
nor U7811 (N_7811,N_5052,N_5400);
nand U7812 (N_7812,N_5930,N_3378);
and U7813 (N_7813,N_3056,N_5290);
or U7814 (N_7814,N_3635,N_4941);
nor U7815 (N_7815,N_3302,N_4333);
nand U7816 (N_7816,N_4174,N_5694);
nand U7817 (N_7817,N_4060,N_3453);
nand U7818 (N_7818,N_4434,N_4015);
xnor U7819 (N_7819,N_5748,N_3827);
or U7820 (N_7820,N_5832,N_3613);
nor U7821 (N_7821,N_5342,N_3103);
nor U7822 (N_7822,N_3679,N_5073);
nand U7823 (N_7823,N_3303,N_5783);
nor U7824 (N_7824,N_5046,N_5849);
nand U7825 (N_7825,N_5903,N_3699);
nand U7826 (N_7826,N_5205,N_4548);
xnor U7827 (N_7827,N_5131,N_4179);
and U7828 (N_7828,N_3422,N_3899);
and U7829 (N_7829,N_4864,N_3265);
nor U7830 (N_7830,N_4797,N_3583);
nand U7831 (N_7831,N_4147,N_5458);
nand U7832 (N_7832,N_4828,N_3729);
xor U7833 (N_7833,N_3142,N_5385);
and U7834 (N_7834,N_3647,N_5811);
nand U7835 (N_7835,N_5604,N_4022);
nand U7836 (N_7836,N_5669,N_4610);
nor U7837 (N_7837,N_4500,N_3115);
or U7838 (N_7838,N_5798,N_5880);
and U7839 (N_7839,N_3269,N_3797);
or U7840 (N_7840,N_5400,N_4641);
and U7841 (N_7841,N_4668,N_3366);
or U7842 (N_7842,N_4999,N_5822);
nor U7843 (N_7843,N_5813,N_5769);
nand U7844 (N_7844,N_4451,N_5183);
xnor U7845 (N_7845,N_4710,N_5322);
or U7846 (N_7846,N_4266,N_3377);
nand U7847 (N_7847,N_4170,N_5389);
or U7848 (N_7848,N_4234,N_3365);
or U7849 (N_7849,N_4181,N_4453);
nand U7850 (N_7850,N_4817,N_5565);
nor U7851 (N_7851,N_3720,N_4241);
nand U7852 (N_7852,N_4997,N_4974);
nand U7853 (N_7853,N_5796,N_4089);
or U7854 (N_7854,N_5181,N_5700);
nor U7855 (N_7855,N_4577,N_5105);
or U7856 (N_7856,N_4367,N_5126);
nand U7857 (N_7857,N_5662,N_3457);
nand U7858 (N_7858,N_5040,N_4941);
or U7859 (N_7859,N_4323,N_4018);
or U7860 (N_7860,N_3017,N_4100);
and U7861 (N_7861,N_4439,N_4957);
and U7862 (N_7862,N_3856,N_4684);
nor U7863 (N_7863,N_4146,N_3685);
nand U7864 (N_7864,N_3140,N_3124);
nor U7865 (N_7865,N_4754,N_3398);
nor U7866 (N_7866,N_4891,N_3441);
nor U7867 (N_7867,N_4721,N_3702);
nor U7868 (N_7868,N_5183,N_4018);
nand U7869 (N_7869,N_4048,N_5548);
nor U7870 (N_7870,N_3461,N_5724);
nor U7871 (N_7871,N_4886,N_4573);
or U7872 (N_7872,N_4929,N_4047);
nand U7873 (N_7873,N_5087,N_4904);
and U7874 (N_7874,N_5223,N_3255);
and U7875 (N_7875,N_5970,N_5511);
or U7876 (N_7876,N_5499,N_5477);
or U7877 (N_7877,N_5058,N_3235);
or U7878 (N_7878,N_4088,N_4442);
nor U7879 (N_7879,N_5614,N_5172);
and U7880 (N_7880,N_5044,N_5792);
or U7881 (N_7881,N_3504,N_3057);
nand U7882 (N_7882,N_4120,N_3824);
nor U7883 (N_7883,N_3890,N_4133);
or U7884 (N_7884,N_3857,N_4206);
and U7885 (N_7885,N_3765,N_3539);
nand U7886 (N_7886,N_4066,N_3387);
nor U7887 (N_7887,N_5318,N_3071);
nor U7888 (N_7888,N_3733,N_5105);
and U7889 (N_7889,N_4415,N_3534);
or U7890 (N_7890,N_3780,N_5655);
and U7891 (N_7891,N_5479,N_3009);
and U7892 (N_7892,N_4123,N_4091);
nor U7893 (N_7893,N_4822,N_4814);
nand U7894 (N_7894,N_5576,N_4297);
or U7895 (N_7895,N_4356,N_3369);
nor U7896 (N_7896,N_5548,N_4629);
nand U7897 (N_7897,N_4080,N_5693);
nand U7898 (N_7898,N_5508,N_3696);
nand U7899 (N_7899,N_5896,N_3227);
nand U7900 (N_7900,N_4924,N_5634);
or U7901 (N_7901,N_4649,N_4402);
nor U7902 (N_7902,N_4569,N_4183);
or U7903 (N_7903,N_4611,N_3564);
nand U7904 (N_7904,N_5685,N_5130);
nor U7905 (N_7905,N_4967,N_4957);
nor U7906 (N_7906,N_4193,N_4798);
nor U7907 (N_7907,N_5974,N_5983);
nand U7908 (N_7908,N_4912,N_5752);
or U7909 (N_7909,N_3345,N_3360);
and U7910 (N_7910,N_5625,N_3865);
or U7911 (N_7911,N_3460,N_4803);
and U7912 (N_7912,N_5252,N_5136);
and U7913 (N_7913,N_3894,N_3120);
and U7914 (N_7914,N_4399,N_3772);
or U7915 (N_7915,N_4244,N_3539);
nor U7916 (N_7916,N_4590,N_4407);
nor U7917 (N_7917,N_4369,N_5114);
or U7918 (N_7918,N_4997,N_4597);
or U7919 (N_7919,N_5756,N_5452);
nand U7920 (N_7920,N_5682,N_3877);
and U7921 (N_7921,N_4542,N_3294);
and U7922 (N_7922,N_4495,N_4777);
or U7923 (N_7923,N_3078,N_3579);
and U7924 (N_7924,N_3442,N_4915);
and U7925 (N_7925,N_3860,N_5525);
nand U7926 (N_7926,N_4729,N_3172);
nor U7927 (N_7927,N_5272,N_4971);
or U7928 (N_7928,N_5985,N_3750);
nand U7929 (N_7929,N_5302,N_5616);
or U7930 (N_7930,N_5805,N_3259);
or U7931 (N_7931,N_5112,N_5782);
and U7932 (N_7932,N_5893,N_3310);
and U7933 (N_7933,N_3551,N_4339);
nor U7934 (N_7934,N_5195,N_4594);
nand U7935 (N_7935,N_3975,N_3304);
nand U7936 (N_7936,N_3078,N_5256);
nand U7937 (N_7937,N_3736,N_3872);
nor U7938 (N_7938,N_4828,N_4218);
nor U7939 (N_7939,N_3730,N_3959);
nand U7940 (N_7940,N_5684,N_4954);
and U7941 (N_7941,N_3766,N_4610);
nand U7942 (N_7942,N_4082,N_4351);
nor U7943 (N_7943,N_4639,N_5976);
nand U7944 (N_7944,N_4355,N_4323);
or U7945 (N_7945,N_4514,N_4106);
and U7946 (N_7946,N_4520,N_4686);
nor U7947 (N_7947,N_3313,N_5243);
nor U7948 (N_7948,N_4641,N_5036);
or U7949 (N_7949,N_3738,N_4538);
nand U7950 (N_7950,N_3524,N_3800);
or U7951 (N_7951,N_3101,N_3890);
nand U7952 (N_7952,N_5548,N_4539);
nor U7953 (N_7953,N_5894,N_3929);
or U7954 (N_7954,N_3084,N_3907);
nor U7955 (N_7955,N_4918,N_4886);
nor U7956 (N_7956,N_5731,N_5154);
nand U7957 (N_7957,N_4355,N_4170);
and U7958 (N_7958,N_3897,N_4596);
nor U7959 (N_7959,N_3970,N_5321);
and U7960 (N_7960,N_4701,N_4842);
nor U7961 (N_7961,N_3737,N_5441);
nor U7962 (N_7962,N_5181,N_5370);
and U7963 (N_7963,N_3590,N_3565);
nor U7964 (N_7964,N_5734,N_5043);
nor U7965 (N_7965,N_4832,N_3206);
nand U7966 (N_7966,N_3212,N_3528);
and U7967 (N_7967,N_5435,N_4135);
nor U7968 (N_7968,N_3975,N_5296);
nand U7969 (N_7969,N_4992,N_4280);
and U7970 (N_7970,N_5168,N_4713);
nand U7971 (N_7971,N_3077,N_4379);
nor U7972 (N_7972,N_5603,N_4284);
or U7973 (N_7973,N_4702,N_4272);
nor U7974 (N_7974,N_5626,N_4024);
nor U7975 (N_7975,N_4455,N_3492);
nor U7976 (N_7976,N_3856,N_5604);
nor U7977 (N_7977,N_3425,N_5497);
nor U7978 (N_7978,N_4808,N_4846);
xor U7979 (N_7979,N_5148,N_5405);
or U7980 (N_7980,N_4768,N_3986);
nand U7981 (N_7981,N_5207,N_3785);
and U7982 (N_7982,N_5385,N_5423);
or U7983 (N_7983,N_5646,N_3724);
nor U7984 (N_7984,N_5392,N_3551);
nor U7985 (N_7985,N_5324,N_4922);
and U7986 (N_7986,N_5205,N_5665);
or U7987 (N_7987,N_5352,N_4846);
xnor U7988 (N_7988,N_3710,N_4289);
or U7989 (N_7989,N_3295,N_4046);
nand U7990 (N_7990,N_3783,N_3973);
or U7991 (N_7991,N_4644,N_4325);
or U7992 (N_7992,N_4339,N_5413);
or U7993 (N_7993,N_4997,N_4922);
or U7994 (N_7994,N_5808,N_5745);
or U7995 (N_7995,N_3954,N_4835);
nand U7996 (N_7996,N_4439,N_3741);
or U7997 (N_7997,N_3498,N_4740);
or U7998 (N_7998,N_3292,N_4592);
and U7999 (N_7999,N_5615,N_5569);
or U8000 (N_8000,N_5285,N_5432);
nand U8001 (N_8001,N_4511,N_4989);
or U8002 (N_8002,N_4771,N_4089);
nand U8003 (N_8003,N_5788,N_5638);
nor U8004 (N_8004,N_4090,N_3943);
and U8005 (N_8005,N_5415,N_3977);
or U8006 (N_8006,N_4455,N_5426);
nor U8007 (N_8007,N_4245,N_3503);
or U8008 (N_8008,N_3680,N_5901);
or U8009 (N_8009,N_4797,N_5080);
nand U8010 (N_8010,N_3273,N_5680);
nor U8011 (N_8011,N_4492,N_3307);
nand U8012 (N_8012,N_3376,N_4158);
or U8013 (N_8013,N_5029,N_3840);
or U8014 (N_8014,N_5890,N_3458);
nand U8015 (N_8015,N_5228,N_5953);
xnor U8016 (N_8016,N_3005,N_3423);
nand U8017 (N_8017,N_4105,N_3117);
nor U8018 (N_8018,N_4502,N_4324);
nor U8019 (N_8019,N_5890,N_3089);
or U8020 (N_8020,N_4941,N_3108);
or U8021 (N_8021,N_5777,N_3235);
and U8022 (N_8022,N_5126,N_4940);
nand U8023 (N_8023,N_3390,N_5670);
and U8024 (N_8024,N_3926,N_3101);
nand U8025 (N_8025,N_5298,N_3008);
or U8026 (N_8026,N_4285,N_4854);
or U8027 (N_8027,N_5197,N_5433);
nor U8028 (N_8028,N_4836,N_5191);
nand U8029 (N_8029,N_3984,N_5679);
nand U8030 (N_8030,N_4163,N_3277);
and U8031 (N_8031,N_5304,N_3320);
nor U8032 (N_8032,N_3819,N_5621);
nor U8033 (N_8033,N_4549,N_3466);
and U8034 (N_8034,N_4267,N_5548);
nand U8035 (N_8035,N_4194,N_4436);
nand U8036 (N_8036,N_5675,N_4742);
nor U8037 (N_8037,N_3776,N_3853);
nor U8038 (N_8038,N_3393,N_3025);
and U8039 (N_8039,N_5731,N_4050);
nand U8040 (N_8040,N_4359,N_4210);
or U8041 (N_8041,N_3664,N_3265);
nand U8042 (N_8042,N_3218,N_3035);
and U8043 (N_8043,N_4769,N_5292);
and U8044 (N_8044,N_4948,N_5749);
nor U8045 (N_8045,N_3258,N_5269);
or U8046 (N_8046,N_4315,N_3580);
nor U8047 (N_8047,N_5882,N_3218);
nand U8048 (N_8048,N_5919,N_5063);
and U8049 (N_8049,N_3745,N_3343);
nor U8050 (N_8050,N_3756,N_4882);
or U8051 (N_8051,N_3843,N_3658);
nand U8052 (N_8052,N_3709,N_3433);
or U8053 (N_8053,N_4740,N_4952);
or U8054 (N_8054,N_5635,N_3657);
nand U8055 (N_8055,N_4412,N_3163);
nand U8056 (N_8056,N_4462,N_4949);
xnor U8057 (N_8057,N_5364,N_4313);
nor U8058 (N_8058,N_5746,N_3548);
and U8059 (N_8059,N_4043,N_4845);
or U8060 (N_8060,N_5635,N_5838);
or U8061 (N_8061,N_4964,N_3438);
nor U8062 (N_8062,N_4787,N_5277);
nor U8063 (N_8063,N_3450,N_5970);
nand U8064 (N_8064,N_4452,N_4667);
and U8065 (N_8065,N_3763,N_5869);
xor U8066 (N_8066,N_4172,N_5390);
and U8067 (N_8067,N_3927,N_3039);
nor U8068 (N_8068,N_5547,N_5593);
nand U8069 (N_8069,N_3258,N_4671);
nor U8070 (N_8070,N_5967,N_5806);
nor U8071 (N_8071,N_5462,N_4561);
nand U8072 (N_8072,N_3079,N_5119);
and U8073 (N_8073,N_4217,N_5043);
nor U8074 (N_8074,N_3199,N_5102);
or U8075 (N_8075,N_3961,N_4718);
nor U8076 (N_8076,N_3748,N_3609);
nor U8077 (N_8077,N_3690,N_5515);
and U8078 (N_8078,N_3980,N_5664);
nor U8079 (N_8079,N_3223,N_3404);
and U8080 (N_8080,N_4604,N_4961);
nand U8081 (N_8081,N_3172,N_5050);
nor U8082 (N_8082,N_3165,N_5794);
nand U8083 (N_8083,N_3458,N_3329);
nand U8084 (N_8084,N_5089,N_4890);
or U8085 (N_8085,N_5525,N_5951);
or U8086 (N_8086,N_4681,N_5588);
nand U8087 (N_8087,N_4498,N_4871);
nor U8088 (N_8088,N_4266,N_3707);
and U8089 (N_8089,N_3408,N_4118);
nor U8090 (N_8090,N_4077,N_3475);
nor U8091 (N_8091,N_3922,N_4053);
nand U8092 (N_8092,N_4367,N_5894);
and U8093 (N_8093,N_5734,N_5649);
or U8094 (N_8094,N_4009,N_3265);
nor U8095 (N_8095,N_5737,N_4079);
or U8096 (N_8096,N_5713,N_5045);
nand U8097 (N_8097,N_3176,N_4056);
nor U8098 (N_8098,N_3823,N_4011);
nand U8099 (N_8099,N_5363,N_3054);
and U8100 (N_8100,N_5988,N_5954);
nand U8101 (N_8101,N_5592,N_5362);
nor U8102 (N_8102,N_5903,N_5263);
and U8103 (N_8103,N_4166,N_4482);
nand U8104 (N_8104,N_5131,N_3525);
and U8105 (N_8105,N_4505,N_5335);
or U8106 (N_8106,N_3265,N_4675);
and U8107 (N_8107,N_3935,N_4819);
xor U8108 (N_8108,N_4480,N_3297);
or U8109 (N_8109,N_5220,N_3561);
or U8110 (N_8110,N_4123,N_3742);
and U8111 (N_8111,N_5628,N_4707);
or U8112 (N_8112,N_4662,N_4500);
or U8113 (N_8113,N_5604,N_3097);
and U8114 (N_8114,N_5647,N_3547);
and U8115 (N_8115,N_4413,N_3586);
nor U8116 (N_8116,N_4538,N_3513);
or U8117 (N_8117,N_4608,N_5213);
and U8118 (N_8118,N_3428,N_5791);
nand U8119 (N_8119,N_5947,N_4251);
or U8120 (N_8120,N_3458,N_5920);
and U8121 (N_8121,N_3843,N_4038);
nor U8122 (N_8122,N_3254,N_5617);
nand U8123 (N_8123,N_4935,N_3740);
nand U8124 (N_8124,N_3393,N_4695);
or U8125 (N_8125,N_4510,N_4289);
or U8126 (N_8126,N_5945,N_5782);
or U8127 (N_8127,N_4550,N_5005);
nand U8128 (N_8128,N_3795,N_3541);
or U8129 (N_8129,N_5505,N_4813);
or U8130 (N_8130,N_3427,N_5956);
and U8131 (N_8131,N_3912,N_3642);
nand U8132 (N_8132,N_5732,N_3019);
and U8133 (N_8133,N_3011,N_4940);
and U8134 (N_8134,N_3367,N_5680);
or U8135 (N_8135,N_4863,N_3113);
nand U8136 (N_8136,N_4493,N_4272);
or U8137 (N_8137,N_5268,N_5900);
nor U8138 (N_8138,N_3142,N_3167);
and U8139 (N_8139,N_3199,N_5172);
or U8140 (N_8140,N_5093,N_4460);
and U8141 (N_8141,N_5620,N_4394);
and U8142 (N_8142,N_3151,N_3251);
or U8143 (N_8143,N_5999,N_5396);
nor U8144 (N_8144,N_5503,N_3104);
nand U8145 (N_8145,N_5960,N_5151);
or U8146 (N_8146,N_3088,N_5244);
or U8147 (N_8147,N_5043,N_3270);
or U8148 (N_8148,N_3003,N_3962);
or U8149 (N_8149,N_4088,N_4794);
nand U8150 (N_8150,N_5616,N_5444);
nand U8151 (N_8151,N_4858,N_3987);
nor U8152 (N_8152,N_5567,N_3843);
and U8153 (N_8153,N_4976,N_5459);
nand U8154 (N_8154,N_3852,N_4325);
or U8155 (N_8155,N_3677,N_5182);
xnor U8156 (N_8156,N_4185,N_5885);
nor U8157 (N_8157,N_3298,N_3017);
xnor U8158 (N_8158,N_4622,N_5955);
and U8159 (N_8159,N_3332,N_4087);
nand U8160 (N_8160,N_5607,N_3799);
nand U8161 (N_8161,N_4112,N_4192);
or U8162 (N_8162,N_5068,N_4760);
and U8163 (N_8163,N_4145,N_5041);
and U8164 (N_8164,N_3215,N_5214);
or U8165 (N_8165,N_5582,N_3292);
or U8166 (N_8166,N_4303,N_3287);
nand U8167 (N_8167,N_3658,N_4186);
nand U8168 (N_8168,N_5167,N_5218);
nor U8169 (N_8169,N_3004,N_5615);
and U8170 (N_8170,N_3142,N_3089);
nor U8171 (N_8171,N_5340,N_5829);
or U8172 (N_8172,N_5906,N_3437);
and U8173 (N_8173,N_5738,N_5252);
or U8174 (N_8174,N_3670,N_3951);
nor U8175 (N_8175,N_5035,N_3208);
nor U8176 (N_8176,N_3971,N_5732);
nor U8177 (N_8177,N_3782,N_5990);
and U8178 (N_8178,N_3796,N_4134);
nor U8179 (N_8179,N_5572,N_4628);
nor U8180 (N_8180,N_5064,N_3345);
or U8181 (N_8181,N_5563,N_4089);
nor U8182 (N_8182,N_4264,N_5710);
nor U8183 (N_8183,N_3069,N_4309);
nand U8184 (N_8184,N_4882,N_5666);
and U8185 (N_8185,N_5510,N_5496);
nand U8186 (N_8186,N_4363,N_3708);
and U8187 (N_8187,N_4954,N_3589);
nand U8188 (N_8188,N_5837,N_4822);
nor U8189 (N_8189,N_5262,N_5120);
and U8190 (N_8190,N_5091,N_3287);
or U8191 (N_8191,N_5813,N_3247);
nand U8192 (N_8192,N_5128,N_4705);
xor U8193 (N_8193,N_4911,N_3962);
and U8194 (N_8194,N_4733,N_3818);
nand U8195 (N_8195,N_4723,N_3766);
nand U8196 (N_8196,N_5475,N_3335);
nand U8197 (N_8197,N_4930,N_5921);
nand U8198 (N_8198,N_4862,N_3651);
or U8199 (N_8199,N_3061,N_4382);
and U8200 (N_8200,N_5710,N_4278);
nand U8201 (N_8201,N_4802,N_5820);
nor U8202 (N_8202,N_4433,N_5357);
nor U8203 (N_8203,N_5434,N_3484);
or U8204 (N_8204,N_5637,N_5017);
or U8205 (N_8205,N_5010,N_4319);
or U8206 (N_8206,N_5612,N_4979);
or U8207 (N_8207,N_4417,N_5462);
nor U8208 (N_8208,N_4494,N_3206);
nor U8209 (N_8209,N_3824,N_3051);
or U8210 (N_8210,N_3450,N_3996);
nor U8211 (N_8211,N_4313,N_5720);
nor U8212 (N_8212,N_5065,N_5537);
and U8213 (N_8213,N_4267,N_5071);
nand U8214 (N_8214,N_3822,N_4472);
or U8215 (N_8215,N_3830,N_4278);
nand U8216 (N_8216,N_3390,N_3236);
nor U8217 (N_8217,N_5219,N_3391);
nor U8218 (N_8218,N_4631,N_5889);
nand U8219 (N_8219,N_5134,N_4914);
and U8220 (N_8220,N_4485,N_3616);
xnor U8221 (N_8221,N_5390,N_5993);
and U8222 (N_8222,N_4051,N_3207);
nand U8223 (N_8223,N_4473,N_3577);
and U8224 (N_8224,N_4444,N_5329);
nor U8225 (N_8225,N_4919,N_3295);
or U8226 (N_8226,N_5390,N_5497);
nor U8227 (N_8227,N_4095,N_4189);
or U8228 (N_8228,N_4930,N_3648);
and U8229 (N_8229,N_3138,N_3344);
nor U8230 (N_8230,N_3318,N_4124);
and U8231 (N_8231,N_4530,N_4251);
or U8232 (N_8232,N_4345,N_3836);
and U8233 (N_8233,N_4831,N_3002);
xor U8234 (N_8234,N_5165,N_3253);
and U8235 (N_8235,N_3313,N_5909);
nor U8236 (N_8236,N_5679,N_4043);
and U8237 (N_8237,N_5636,N_3041);
or U8238 (N_8238,N_5329,N_3049);
and U8239 (N_8239,N_5668,N_5430);
and U8240 (N_8240,N_3136,N_3678);
nor U8241 (N_8241,N_3932,N_3557);
xnor U8242 (N_8242,N_5100,N_3398);
nand U8243 (N_8243,N_3377,N_4312);
nor U8244 (N_8244,N_4651,N_5894);
or U8245 (N_8245,N_5441,N_4439);
or U8246 (N_8246,N_3409,N_5591);
and U8247 (N_8247,N_3133,N_5881);
and U8248 (N_8248,N_3145,N_5869);
nand U8249 (N_8249,N_4533,N_4553);
or U8250 (N_8250,N_5052,N_5272);
nand U8251 (N_8251,N_5548,N_3172);
nor U8252 (N_8252,N_4099,N_4420);
and U8253 (N_8253,N_3084,N_5166);
nand U8254 (N_8254,N_3128,N_4657);
xor U8255 (N_8255,N_4330,N_5746);
nor U8256 (N_8256,N_3926,N_5756);
or U8257 (N_8257,N_5169,N_3275);
nor U8258 (N_8258,N_4157,N_3585);
nand U8259 (N_8259,N_5510,N_4455);
nand U8260 (N_8260,N_3847,N_4560);
or U8261 (N_8261,N_4167,N_3067);
or U8262 (N_8262,N_3723,N_5297);
and U8263 (N_8263,N_5479,N_4486);
and U8264 (N_8264,N_3545,N_3275);
and U8265 (N_8265,N_3556,N_4692);
nand U8266 (N_8266,N_4261,N_5347);
nor U8267 (N_8267,N_4264,N_5239);
or U8268 (N_8268,N_4302,N_5024);
or U8269 (N_8269,N_5711,N_4380);
nor U8270 (N_8270,N_5410,N_3464);
and U8271 (N_8271,N_5087,N_4718);
nand U8272 (N_8272,N_4684,N_4245);
nand U8273 (N_8273,N_5874,N_3568);
nand U8274 (N_8274,N_3255,N_3053);
or U8275 (N_8275,N_4293,N_3256);
xor U8276 (N_8276,N_3690,N_4782);
or U8277 (N_8277,N_4160,N_5621);
nand U8278 (N_8278,N_4709,N_3048);
or U8279 (N_8279,N_3529,N_4218);
and U8280 (N_8280,N_3035,N_4509);
nor U8281 (N_8281,N_5546,N_4105);
nand U8282 (N_8282,N_3947,N_4286);
or U8283 (N_8283,N_4342,N_5193);
and U8284 (N_8284,N_5421,N_3521);
nor U8285 (N_8285,N_3712,N_5883);
xnor U8286 (N_8286,N_5564,N_5467);
nand U8287 (N_8287,N_4014,N_4425);
nor U8288 (N_8288,N_4026,N_3264);
nor U8289 (N_8289,N_5324,N_5712);
or U8290 (N_8290,N_3496,N_5263);
or U8291 (N_8291,N_3900,N_4100);
and U8292 (N_8292,N_5445,N_3408);
nor U8293 (N_8293,N_4391,N_3059);
xor U8294 (N_8294,N_4635,N_5377);
or U8295 (N_8295,N_5686,N_4919);
xnor U8296 (N_8296,N_3207,N_4977);
nor U8297 (N_8297,N_3766,N_4681);
or U8298 (N_8298,N_3245,N_4036);
nor U8299 (N_8299,N_5938,N_5780);
nand U8300 (N_8300,N_5050,N_4380);
or U8301 (N_8301,N_5562,N_5028);
nor U8302 (N_8302,N_3764,N_4702);
or U8303 (N_8303,N_3750,N_5933);
nand U8304 (N_8304,N_3724,N_5413);
nor U8305 (N_8305,N_4473,N_5710);
nand U8306 (N_8306,N_3325,N_4618);
or U8307 (N_8307,N_5166,N_3489);
nor U8308 (N_8308,N_5606,N_5544);
and U8309 (N_8309,N_4561,N_5854);
nor U8310 (N_8310,N_5439,N_3078);
and U8311 (N_8311,N_4702,N_4057);
nor U8312 (N_8312,N_5227,N_4069);
and U8313 (N_8313,N_3281,N_4583);
nand U8314 (N_8314,N_4249,N_4462);
nand U8315 (N_8315,N_4202,N_3876);
nor U8316 (N_8316,N_3124,N_4730);
or U8317 (N_8317,N_4606,N_5329);
nand U8318 (N_8318,N_4324,N_3577);
and U8319 (N_8319,N_5518,N_5766);
nor U8320 (N_8320,N_4512,N_3624);
nor U8321 (N_8321,N_5430,N_4907);
nand U8322 (N_8322,N_4627,N_5719);
or U8323 (N_8323,N_4742,N_4611);
nand U8324 (N_8324,N_4423,N_5142);
and U8325 (N_8325,N_3796,N_4916);
nand U8326 (N_8326,N_5632,N_3100);
nand U8327 (N_8327,N_3936,N_4274);
nand U8328 (N_8328,N_4382,N_3383);
and U8329 (N_8329,N_3723,N_3058);
nor U8330 (N_8330,N_4470,N_5358);
and U8331 (N_8331,N_5682,N_5427);
or U8332 (N_8332,N_3659,N_5534);
nand U8333 (N_8333,N_3492,N_5194);
or U8334 (N_8334,N_5149,N_4915);
and U8335 (N_8335,N_3091,N_4614);
or U8336 (N_8336,N_5389,N_3809);
and U8337 (N_8337,N_4202,N_4281);
nand U8338 (N_8338,N_4961,N_5914);
nand U8339 (N_8339,N_3514,N_5668);
or U8340 (N_8340,N_4400,N_4926);
and U8341 (N_8341,N_5983,N_4731);
or U8342 (N_8342,N_4496,N_4191);
nand U8343 (N_8343,N_4956,N_5372);
nor U8344 (N_8344,N_4526,N_5044);
or U8345 (N_8345,N_4289,N_3730);
or U8346 (N_8346,N_3619,N_3224);
or U8347 (N_8347,N_3955,N_3798);
and U8348 (N_8348,N_3663,N_3394);
or U8349 (N_8349,N_3051,N_3495);
or U8350 (N_8350,N_5518,N_4844);
or U8351 (N_8351,N_5758,N_4827);
nor U8352 (N_8352,N_4617,N_5895);
nand U8353 (N_8353,N_4153,N_5777);
xnor U8354 (N_8354,N_5304,N_3756);
or U8355 (N_8355,N_4881,N_3446);
or U8356 (N_8356,N_5248,N_3801);
nand U8357 (N_8357,N_5596,N_4245);
nor U8358 (N_8358,N_4458,N_3402);
and U8359 (N_8359,N_4179,N_4281);
nand U8360 (N_8360,N_3802,N_4229);
nand U8361 (N_8361,N_3170,N_3729);
and U8362 (N_8362,N_4203,N_5517);
and U8363 (N_8363,N_3655,N_3830);
nor U8364 (N_8364,N_3268,N_3809);
or U8365 (N_8365,N_3091,N_5502);
and U8366 (N_8366,N_4650,N_4662);
nor U8367 (N_8367,N_4168,N_3226);
nand U8368 (N_8368,N_3527,N_5477);
nand U8369 (N_8369,N_5893,N_4216);
nor U8370 (N_8370,N_5392,N_3425);
and U8371 (N_8371,N_3704,N_3863);
and U8372 (N_8372,N_5355,N_3099);
and U8373 (N_8373,N_4841,N_5347);
and U8374 (N_8374,N_4289,N_4888);
and U8375 (N_8375,N_5966,N_4650);
or U8376 (N_8376,N_3342,N_5818);
or U8377 (N_8377,N_5988,N_4184);
or U8378 (N_8378,N_4037,N_4443);
or U8379 (N_8379,N_5832,N_3086);
and U8380 (N_8380,N_3055,N_5520);
nor U8381 (N_8381,N_5936,N_5752);
and U8382 (N_8382,N_3002,N_4941);
nor U8383 (N_8383,N_5551,N_5236);
nand U8384 (N_8384,N_3753,N_3408);
and U8385 (N_8385,N_4997,N_3925);
or U8386 (N_8386,N_3961,N_4506);
nor U8387 (N_8387,N_3148,N_3338);
or U8388 (N_8388,N_4243,N_5127);
nor U8389 (N_8389,N_4675,N_4232);
and U8390 (N_8390,N_3045,N_3604);
and U8391 (N_8391,N_4822,N_3715);
or U8392 (N_8392,N_5417,N_5095);
nand U8393 (N_8393,N_4326,N_3968);
nor U8394 (N_8394,N_5298,N_3980);
or U8395 (N_8395,N_3603,N_4838);
nand U8396 (N_8396,N_3172,N_4211);
nor U8397 (N_8397,N_3788,N_3392);
or U8398 (N_8398,N_5813,N_4060);
or U8399 (N_8399,N_4879,N_5139);
nand U8400 (N_8400,N_4803,N_4926);
or U8401 (N_8401,N_3899,N_3415);
or U8402 (N_8402,N_4290,N_4102);
or U8403 (N_8403,N_4528,N_5501);
nor U8404 (N_8404,N_5054,N_4209);
and U8405 (N_8405,N_5372,N_3501);
nor U8406 (N_8406,N_3651,N_4011);
or U8407 (N_8407,N_4087,N_4413);
xor U8408 (N_8408,N_5990,N_5176);
nand U8409 (N_8409,N_5882,N_4596);
nor U8410 (N_8410,N_3422,N_5498);
nor U8411 (N_8411,N_3061,N_5422);
or U8412 (N_8412,N_3184,N_4130);
nor U8413 (N_8413,N_5323,N_4525);
nand U8414 (N_8414,N_3139,N_4579);
or U8415 (N_8415,N_5885,N_3705);
or U8416 (N_8416,N_5200,N_3328);
and U8417 (N_8417,N_5745,N_4163);
nand U8418 (N_8418,N_4996,N_4114);
and U8419 (N_8419,N_3412,N_4156);
nor U8420 (N_8420,N_3458,N_3672);
nor U8421 (N_8421,N_3957,N_3708);
or U8422 (N_8422,N_5261,N_5802);
xnor U8423 (N_8423,N_4770,N_3652);
or U8424 (N_8424,N_5302,N_5876);
nand U8425 (N_8425,N_3349,N_4459);
and U8426 (N_8426,N_4020,N_4936);
nor U8427 (N_8427,N_3346,N_4718);
and U8428 (N_8428,N_5417,N_3742);
nand U8429 (N_8429,N_3714,N_5062);
or U8430 (N_8430,N_3187,N_3341);
or U8431 (N_8431,N_3368,N_5605);
nand U8432 (N_8432,N_5467,N_5343);
or U8433 (N_8433,N_4273,N_3978);
or U8434 (N_8434,N_3861,N_5239);
nor U8435 (N_8435,N_4845,N_5400);
nor U8436 (N_8436,N_3314,N_4616);
nor U8437 (N_8437,N_3826,N_5667);
or U8438 (N_8438,N_3777,N_4647);
nor U8439 (N_8439,N_5249,N_4464);
nor U8440 (N_8440,N_4585,N_5491);
nor U8441 (N_8441,N_5976,N_4275);
nor U8442 (N_8442,N_3171,N_3732);
nand U8443 (N_8443,N_3311,N_4666);
or U8444 (N_8444,N_5239,N_5816);
and U8445 (N_8445,N_5039,N_5340);
nor U8446 (N_8446,N_4245,N_4979);
or U8447 (N_8447,N_5378,N_4792);
and U8448 (N_8448,N_5088,N_5873);
nor U8449 (N_8449,N_3726,N_5036);
and U8450 (N_8450,N_4750,N_3864);
nand U8451 (N_8451,N_3960,N_5590);
nand U8452 (N_8452,N_5578,N_4621);
nor U8453 (N_8453,N_3388,N_4663);
and U8454 (N_8454,N_3108,N_3706);
nor U8455 (N_8455,N_5177,N_3689);
nor U8456 (N_8456,N_3492,N_4312);
nor U8457 (N_8457,N_4604,N_5443);
or U8458 (N_8458,N_5222,N_4211);
nor U8459 (N_8459,N_5068,N_5223);
xor U8460 (N_8460,N_3050,N_3327);
or U8461 (N_8461,N_5490,N_4818);
nand U8462 (N_8462,N_5674,N_3253);
nand U8463 (N_8463,N_4230,N_5592);
and U8464 (N_8464,N_3678,N_3279);
nor U8465 (N_8465,N_4846,N_5975);
nor U8466 (N_8466,N_5468,N_5940);
nor U8467 (N_8467,N_5354,N_3179);
or U8468 (N_8468,N_3609,N_5873);
or U8469 (N_8469,N_5819,N_3194);
or U8470 (N_8470,N_3393,N_5547);
or U8471 (N_8471,N_4452,N_5685);
nand U8472 (N_8472,N_5738,N_3457);
and U8473 (N_8473,N_4435,N_5741);
or U8474 (N_8474,N_4247,N_4763);
and U8475 (N_8475,N_4429,N_5907);
nor U8476 (N_8476,N_5838,N_5109);
nor U8477 (N_8477,N_3221,N_3541);
nor U8478 (N_8478,N_3646,N_5827);
nand U8479 (N_8479,N_4346,N_5495);
nor U8480 (N_8480,N_5312,N_3762);
xor U8481 (N_8481,N_4523,N_3205);
or U8482 (N_8482,N_4102,N_4042);
nand U8483 (N_8483,N_4016,N_3170);
nor U8484 (N_8484,N_5290,N_5308);
nor U8485 (N_8485,N_4885,N_3006);
nor U8486 (N_8486,N_3693,N_5478);
and U8487 (N_8487,N_5863,N_5269);
nand U8488 (N_8488,N_4530,N_3161);
or U8489 (N_8489,N_5485,N_3988);
nor U8490 (N_8490,N_3319,N_3785);
and U8491 (N_8491,N_4271,N_3038);
xnor U8492 (N_8492,N_4716,N_3941);
nor U8493 (N_8493,N_4862,N_3494);
nand U8494 (N_8494,N_5048,N_5584);
nor U8495 (N_8495,N_3465,N_5516);
or U8496 (N_8496,N_4488,N_4358);
nand U8497 (N_8497,N_3019,N_3725);
or U8498 (N_8498,N_5826,N_4223);
nand U8499 (N_8499,N_4360,N_3702);
nor U8500 (N_8500,N_4246,N_5415);
or U8501 (N_8501,N_4574,N_4717);
nor U8502 (N_8502,N_4216,N_5120);
nand U8503 (N_8503,N_4632,N_4501);
and U8504 (N_8504,N_5665,N_5562);
or U8505 (N_8505,N_3321,N_4407);
xor U8506 (N_8506,N_3175,N_3272);
or U8507 (N_8507,N_3345,N_4781);
and U8508 (N_8508,N_3174,N_4395);
nor U8509 (N_8509,N_4736,N_4898);
or U8510 (N_8510,N_4314,N_5431);
xnor U8511 (N_8511,N_4605,N_5890);
nand U8512 (N_8512,N_3445,N_5228);
nor U8513 (N_8513,N_5656,N_3389);
nand U8514 (N_8514,N_5636,N_3389);
or U8515 (N_8515,N_3294,N_3153);
and U8516 (N_8516,N_3308,N_3825);
nand U8517 (N_8517,N_5480,N_4469);
and U8518 (N_8518,N_4334,N_4237);
and U8519 (N_8519,N_3801,N_3252);
nor U8520 (N_8520,N_3990,N_5176);
nor U8521 (N_8521,N_4558,N_3936);
xor U8522 (N_8522,N_3004,N_4650);
nor U8523 (N_8523,N_5333,N_3200);
and U8524 (N_8524,N_3476,N_5585);
or U8525 (N_8525,N_5280,N_5563);
nand U8526 (N_8526,N_5384,N_4973);
nor U8527 (N_8527,N_5189,N_3589);
and U8528 (N_8528,N_4938,N_3099);
and U8529 (N_8529,N_4168,N_3908);
and U8530 (N_8530,N_4080,N_3923);
and U8531 (N_8531,N_4713,N_3298);
nor U8532 (N_8532,N_5655,N_3587);
or U8533 (N_8533,N_4879,N_5241);
nor U8534 (N_8534,N_4923,N_4398);
nor U8535 (N_8535,N_5673,N_5614);
nor U8536 (N_8536,N_3822,N_3437);
and U8537 (N_8537,N_4767,N_3816);
nor U8538 (N_8538,N_3379,N_3276);
nand U8539 (N_8539,N_3369,N_3600);
or U8540 (N_8540,N_4013,N_3321);
nor U8541 (N_8541,N_5207,N_3136);
or U8542 (N_8542,N_4120,N_3032);
nand U8543 (N_8543,N_5153,N_3361);
or U8544 (N_8544,N_3007,N_5172);
or U8545 (N_8545,N_4959,N_5917);
or U8546 (N_8546,N_4126,N_5272);
and U8547 (N_8547,N_5675,N_3409);
or U8548 (N_8548,N_3452,N_5220);
and U8549 (N_8549,N_5174,N_5006);
and U8550 (N_8550,N_3408,N_5427);
nor U8551 (N_8551,N_5719,N_3659);
nor U8552 (N_8552,N_4543,N_4627);
nand U8553 (N_8553,N_5269,N_3801);
nand U8554 (N_8554,N_4316,N_4456);
nand U8555 (N_8555,N_3959,N_5802);
or U8556 (N_8556,N_5406,N_4709);
nor U8557 (N_8557,N_3278,N_5497);
nand U8558 (N_8558,N_5319,N_4867);
nand U8559 (N_8559,N_5106,N_5248);
nand U8560 (N_8560,N_5087,N_3390);
and U8561 (N_8561,N_3933,N_5247);
nor U8562 (N_8562,N_5766,N_3536);
and U8563 (N_8563,N_4503,N_3037);
nor U8564 (N_8564,N_4498,N_5429);
nand U8565 (N_8565,N_4177,N_4954);
and U8566 (N_8566,N_3536,N_5789);
and U8567 (N_8567,N_3215,N_4957);
nand U8568 (N_8568,N_3020,N_3424);
nand U8569 (N_8569,N_3075,N_5501);
and U8570 (N_8570,N_5274,N_5863);
nand U8571 (N_8571,N_5487,N_3190);
nor U8572 (N_8572,N_4387,N_5718);
nand U8573 (N_8573,N_3619,N_4568);
nand U8574 (N_8574,N_5796,N_3240);
nor U8575 (N_8575,N_5498,N_3324);
or U8576 (N_8576,N_3962,N_3580);
and U8577 (N_8577,N_3168,N_4379);
or U8578 (N_8578,N_4684,N_3908);
nand U8579 (N_8579,N_3227,N_5681);
and U8580 (N_8580,N_4555,N_3653);
nand U8581 (N_8581,N_3860,N_5164);
or U8582 (N_8582,N_4387,N_4106);
or U8583 (N_8583,N_4472,N_5899);
nand U8584 (N_8584,N_3001,N_4592);
nor U8585 (N_8585,N_3677,N_5399);
or U8586 (N_8586,N_5648,N_4835);
nand U8587 (N_8587,N_4417,N_3135);
nand U8588 (N_8588,N_5742,N_4785);
nor U8589 (N_8589,N_5394,N_4814);
nand U8590 (N_8590,N_4183,N_3487);
nand U8591 (N_8591,N_3748,N_5016);
and U8592 (N_8592,N_3939,N_3857);
and U8593 (N_8593,N_3175,N_5227);
or U8594 (N_8594,N_4112,N_4425);
xor U8595 (N_8595,N_5481,N_4690);
nor U8596 (N_8596,N_3734,N_3567);
and U8597 (N_8597,N_4209,N_4466);
nor U8598 (N_8598,N_5201,N_3301);
or U8599 (N_8599,N_4993,N_5631);
nor U8600 (N_8600,N_3959,N_3823);
nand U8601 (N_8601,N_3328,N_3957);
or U8602 (N_8602,N_3785,N_4056);
and U8603 (N_8603,N_4993,N_3105);
and U8604 (N_8604,N_3755,N_4603);
or U8605 (N_8605,N_5010,N_3745);
nand U8606 (N_8606,N_3255,N_5844);
nand U8607 (N_8607,N_4405,N_5444);
and U8608 (N_8608,N_5819,N_4199);
and U8609 (N_8609,N_5958,N_5631);
nor U8610 (N_8610,N_4043,N_5841);
and U8611 (N_8611,N_5208,N_4100);
and U8612 (N_8612,N_5867,N_3562);
nand U8613 (N_8613,N_3651,N_4836);
nor U8614 (N_8614,N_3746,N_5274);
or U8615 (N_8615,N_5431,N_5868);
or U8616 (N_8616,N_3441,N_4371);
nand U8617 (N_8617,N_3118,N_4453);
nand U8618 (N_8618,N_3486,N_5787);
or U8619 (N_8619,N_3422,N_5796);
nand U8620 (N_8620,N_4691,N_4310);
and U8621 (N_8621,N_5888,N_5229);
xnor U8622 (N_8622,N_5500,N_3831);
and U8623 (N_8623,N_4867,N_5543);
and U8624 (N_8624,N_4542,N_3895);
or U8625 (N_8625,N_4912,N_5616);
or U8626 (N_8626,N_5142,N_4269);
and U8627 (N_8627,N_4958,N_3353);
or U8628 (N_8628,N_4842,N_5091);
or U8629 (N_8629,N_3256,N_4935);
and U8630 (N_8630,N_4259,N_3509);
nand U8631 (N_8631,N_5450,N_5709);
or U8632 (N_8632,N_5408,N_5788);
nor U8633 (N_8633,N_3173,N_4396);
and U8634 (N_8634,N_4551,N_3608);
and U8635 (N_8635,N_5012,N_4599);
nor U8636 (N_8636,N_3057,N_5287);
or U8637 (N_8637,N_3827,N_4704);
nor U8638 (N_8638,N_5792,N_4586);
and U8639 (N_8639,N_3708,N_3907);
nor U8640 (N_8640,N_4447,N_4517);
nor U8641 (N_8641,N_3528,N_3951);
and U8642 (N_8642,N_3088,N_4022);
nand U8643 (N_8643,N_3436,N_3387);
nor U8644 (N_8644,N_4120,N_3779);
xor U8645 (N_8645,N_4270,N_3336);
nand U8646 (N_8646,N_5619,N_5705);
or U8647 (N_8647,N_3668,N_4834);
nand U8648 (N_8648,N_3769,N_4747);
nor U8649 (N_8649,N_5523,N_4647);
nand U8650 (N_8650,N_5601,N_4587);
nor U8651 (N_8651,N_3098,N_4653);
and U8652 (N_8652,N_3578,N_4624);
nand U8653 (N_8653,N_4726,N_4573);
and U8654 (N_8654,N_5074,N_5076);
nor U8655 (N_8655,N_3878,N_5102);
nor U8656 (N_8656,N_3129,N_5021);
nand U8657 (N_8657,N_5542,N_4059);
nor U8658 (N_8658,N_5742,N_4471);
xnor U8659 (N_8659,N_4285,N_5439);
and U8660 (N_8660,N_5704,N_4730);
or U8661 (N_8661,N_4589,N_5605);
and U8662 (N_8662,N_4042,N_3544);
nor U8663 (N_8663,N_3671,N_3295);
nor U8664 (N_8664,N_4903,N_5541);
nand U8665 (N_8665,N_3258,N_4424);
or U8666 (N_8666,N_3495,N_5869);
or U8667 (N_8667,N_4092,N_5024);
nand U8668 (N_8668,N_5438,N_5078);
and U8669 (N_8669,N_5582,N_5787);
or U8670 (N_8670,N_4099,N_4637);
or U8671 (N_8671,N_5788,N_5837);
nand U8672 (N_8672,N_5074,N_4147);
or U8673 (N_8673,N_5674,N_4560);
or U8674 (N_8674,N_4968,N_5987);
nor U8675 (N_8675,N_4836,N_4391);
nand U8676 (N_8676,N_5802,N_5630);
or U8677 (N_8677,N_4347,N_3790);
xnor U8678 (N_8678,N_4418,N_3131);
nand U8679 (N_8679,N_3581,N_3615);
or U8680 (N_8680,N_3849,N_3797);
nand U8681 (N_8681,N_5172,N_3136);
or U8682 (N_8682,N_4548,N_4082);
nor U8683 (N_8683,N_3386,N_4502);
or U8684 (N_8684,N_5969,N_5879);
nor U8685 (N_8685,N_5040,N_3358);
nor U8686 (N_8686,N_4043,N_3671);
and U8687 (N_8687,N_5410,N_4204);
nor U8688 (N_8688,N_5767,N_4939);
and U8689 (N_8689,N_4174,N_4059);
nand U8690 (N_8690,N_3091,N_4651);
xor U8691 (N_8691,N_4467,N_5420);
xnor U8692 (N_8692,N_4476,N_5427);
nor U8693 (N_8693,N_3044,N_5095);
nor U8694 (N_8694,N_4783,N_5466);
and U8695 (N_8695,N_4719,N_5965);
and U8696 (N_8696,N_5958,N_5515);
or U8697 (N_8697,N_3424,N_5536);
and U8698 (N_8698,N_5888,N_5105);
nand U8699 (N_8699,N_3284,N_5628);
nor U8700 (N_8700,N_3346,N_5498);
or U8701 (N_8701,N_5817,N_4754);
nor U8702 (N_8702,N_5541,N_4516);
and U8703 (N_8703,N_3283,N_3181);
nor U8704 (N_8704,N_5688,N_3041);
or U8705 (N_8705,N_3789,N_3712);
and U8706 (N_8706,N_3801,N_4788);
nor U8707 (N_8707,N_4512,N_4866);
nor U8708 (N_8708,N_4139,N_4801);
and U8709 (N_8709,N_4089,N_3859);
and U8710 (N_8710,N_3615,N_4540);
nand U8711 (N_8711,N_4997,N_5404);
nand U8712 (N_8712,N_3886,N_3897);
nand U8713 (N_8713,N_4712,N_3011);
or U8714 (N_8714,N_5520,N_5983);
and U8715 (N_8715,N_5891,N_5924);
or U8716 (N_8716,N_4554,N_3067);
nand U8717 (N_8717,N_4546,N_4024);
nand U8718 (N_8718,N_5375,N_4341);
xor U8719 (N_8719,N_4328,N_4842);
and U8720 (N_8720,N_4431,N_3921);
and U8721 (N_8721,N_4822,N_4747);
or U8722 (N_8722,N_5879,N_5685);
and U8723 (N_8723,N_4570,N_4239);
nor U8724 (N_8724,N_3376,N_5858);
nor U8725 (N_8725,N_5724,N_5492);
and U8726 (N_8726,N_3047,N_5381);
nor U8727 (N_8727,N_3220,N_4362);
or U8728 (N_8728,N_4524,N_3608);
and U8729 (N_8729,N_5331,N_5774);
or U8730 (N_8730,N_4573,N_3710);
nand U8731 (N_8731,N_3383,N_3324);
nand U8732 (N_8732,N_5686,N_3699);
or U8733 (N_8733,N_4893,N_5389);
and U8734 (N_8734,N_5090,N_5526);
nor U8735 (N_8735,N_4747,N_3119);
or U8736 (N_8736,N_4262,N_5882);
and U8737 (N_8737,N_4491,N_5795);
nor U8738 (N_8738,N_4095,N_4741);
or U8739 (N_8739,N_3326,N_5999);
xor U8740 (N_8740,N_3459,N_4702);
or U8741 (N_8741,N_5519,N_3382);
or U8742 (N_8742,N_3513,N_5597);
nor U8743 (N_8743,N_3221,N_5419);
or U8744 (N_8744,N_3388,N_5451);
or U8745 (N_8745,N_3067,N_5141);
or U8746 (N_8746,N_4710,N_5974);
and U8747 (N_8747,N_3618,N_3667);
nand U8748 (N_8748,N_3524,N_4768);
nor U8749 (N_8749,N_5166,N_4531);
or U8750 (N_8750,N_3018,N_5967);
nor U8751 (N_8751,N_3830,N_3338);
and U8752 (N_8752,N_3326,N_5960);
nand U8753 (N_8753,N_4423,N_5818);
nor U8754 (N_8754,N_4532,N_5335);
or U8755 (N_8755,N_5263,N_3358);
nand U8756 (N_8756,N_4547,N_4132);
or U8757 (N_8757,N_5033,N_4810);
and U8758 (N_8758,N_3315,N_4587);
and U8759 (N_8759,N_3855,N_3002);
nand U8760 (N_8760,N_5293,N_3469);
and U8761 (N_8761,N_3481,N_3483);
and U8762 (N_8762,N_5512,N_5944);
nor U8763 (N_8763,N_5264,N_4168);
and U8764 (N_8764,N_5340,N_3254);
nor U8765 (N_8765,N_4265,N_5968);
and U8766 (N_8766,N_5891,N_5309);
nand U8767 (N_8767,N_5694,N_4865);
or U8768 (N_8768,N_3637,N_4321);
nor U8769 (N_8769,N_3855,N_5881);
or U8770 (N_8770,N_3548,N_4647);
nor U8771 (N_8771,N_4074,N_4323);
nand U8772 (N_8772,N_5178,N_3677);
nand U8773 (N_8773,N_5460,N_4297);
and U8774 (N_8774,N_5359,N_5593);
or U8775 (N_8775,N_3862,N_4373);
xnor U8776 (N_8776,N_4168,N_4412);
and U8777 (N_8777,N_4791,N_4419);
and U8778 (N_8778,N_4389,N_5660);
or U8779 (N_8779,N_5144,N_5203);
and U8780 (N_8780,N_4923,N_4020);
xor U8781 (N_8781,N_4148,N_4678);
nor U8782 (N_8782,N_5608,N_5508);
nor U8783 (N_8783,N_3680,N_4494);
nand U8784 (N_8784,N_5356,N_5881);
and U8785 (N_8785,N_5376,N_5027);
nor U8786 (N_8786,N_4335,N_3257);
and U8787 (N_8787,N_5981,N_4600);
nand U8788 (N_8788,N_5147,N_3105);
nor U8789 (N_8789,N_5918,N_4888);
nand U8790 (N_8790,N_5426,N_4775);
nor U8791 (N_8791,N_4856,N_4822);
nand U8792 (N_8792,N_4398,N_4465);
nand U8793 (N_8793,N_5631,N_4257);
or U8794 (N_8794,N_5220,N_5580);
nor U8795 (N_8795,N_5232,N_4616);
or U8796 (N_8796,N_4439,N_5716);
nor U8797 (N_8797,N_4989,N_5003);
or U8798 (N_8798,N_3988,N_5826);
or U8799 (N_8799,N_5353,N_3144);
nand U8800 (N_8800,N_4056,N_5163);
or U8801 (N_8801,N_4470,N_5029);
and U8802 (N_8802,N_4935,N_3592);
nor U8803 (N_8803,N_4056,N_3880);
nor U8804 (N_8804,N_3678,N_5179);
nand U8805 (N_8805,N_5540,N_3769);
or U8806 (N_8806,N_3358,N_5927);
and U8807 (N_8807,N_3209,N_5151);
or U8808 (N_8808,N_3289,N_5941);
nand U8809 (N_8809,N_4355,N_5137);
xor U8810 (N_8810,N_5283,N_3783);
and U8811 (N_8811,N_3552,N_3073);
and U8812 (N_8812,N_5096,N_4050);
or U8813 (N_8813,N_3874,N_4730);
nor U8814 (N_8814,N_5354,N_3080);
nand U8815 (N_8815,N_5658,N_5814);
nand U8816 (N_8816,N_4848,N_5677);
nor U8817 (N_8817,N_5498,N_4373);
nor U8818 (N_8818,N_5667,N_5964);
nor U8819 (N_8819,N_3783,N_5653);
or U8820 (N_8820,N_4497,N_4667);
nor U8821 (N_8821,N_5802,N_4880);
nor U8822 (N_8822,N_5277,N_4300);
and U8823 (N_8823,N_4853,N_4822);
and U8824 (N_8824,N_4106,N_3232);
and U8825 (N_8825,N_5520,N_5172);
or U8826 (N_8826,N_5117,N_5574);
and U8827 (N_8827,N_5199,N_4612);
nand U8828 (N_8828,N_3782,N_3991);
or U8829 (N_8829,N_5592,N_3641);
nand U8830 (N_8830,N_3786,N_5538);
nor U8831 (N_8831,N_5457,N_3175);
nor U8832 (N_8832,N_4571,N_3116);
nor U8833 (N_8833,N_3779,N_3354);
or U8834 (N_8834,N_4612,N_3052);
and U8835 (N_8835,N_4133,N_3527);
nand U8836 (N_8836,N_4554,N_5114);
nand U8837 (N_8837,N_4915,N_4599);
nor U8838 (N_8838,N_3405,N_3440);
nor U8839 (N_8839,N_5684,N_4641);
or U8840 (N_8840,N_3083,N_3730);
and U8841 (N_8841,N_3523,N_4409);
or U8842 (N_8842,N_5358,N_5933);
nor U8843 (N_8843,N_5195,N_5529);
and U8844 (N_8844,N_3504,N_4350);
or U8845 (N_8845,N_5375,N_4833);
and U8846 (N_8846,N_4163,N_4138);
and U8847 (N_8847,N_4755,N_4635);
and U8848 (N_8848,N_4080,N_5452);
or U8849 (N_8849,N_4670,N_3053);
and U8850 (N_8850,N_3042,N_5133);
or U8851 (N_8851,N_4232,N_5175);
or U8852 (N_8852,N_3840,N_3126);
nand U8853 (N_8853,N_4807,N_4340);
xnor U8854 (N_8854,N_4670,N_4039);
or U8855 (N_8855,N_3048,N_4577);
or U8856 (N_8856,N_5608,N_5210);
or U8857 (N_8857,N_5474,N_4668);
or U8858 (N_8858,N_3769,N_3286);
nor U8859 (N_8859,N_3512,N_4632);
nor U8860 (N_8860,N_3026,N_4834);
xnor U8861 (N_8861,N_4683,N_5498);
and U8862 (N_8862,N_4426,N_5983);
nor U8863 (N_8863,N_4186,N_3627);
nor U8864 (N_8864,N_3080,N_5315);
nand U8865 (N_8865,N_3341,N_4774);
xnor U8866 (N_8866,N_5497,N_3233);
or U8867 (N_8867,N_5040,N_5524);
nor U8868 (N_8868,N_4627,N_5628);
nor U8869 (N_8869,N_4847,N_5646);
and U8870 (N_8870,N_3112,N_4420);
and U8871 (N_8871,N_5564,N_5499);
nand U8872 (N_8872,N_3971,N_4550);
and U8873 (N_8873,N_3243,N_5870);
and U8874 (N_8874,N_5024,N_5282);
nand U8875 (N_8875,N_4295,N_3082);
xnor U8876 (N_8876,N_4542,N_4448);
nand U8877 (N_8877,N_3835,N_4550);
nor U8878 (N_8878,N_5394,N_4328);
or U8879 (N_8879,N_3291,N_3054);
and U8880 (N_8880,N_4146,N_5760);
nand U8881 (N_8881,N_3236,N_5864);
and U8882 (N_8882,N_4680,N_4638);
nand U8883 (N_8883,N_5382,N_3920);
or U8884 (N_8884,N_4500,N_5252);
nor U8885 (N_8885,N_3575,N_5484);
nand U8886 (N_8886,N_4180,N_4008);
and U8887 (N_8887,N_3490,N_4438);
and U8888 (N_8888,N_5028,N_4865);
or U8889 (N_8889,N_5896,N_3063);
nand U8890 (N_8890,N_3304,N_5514);
nand U8891 (N_8891,N_3148,N_3369);
or U8892 (N_8892,N_3595,N_3931);
nand U8893 (N_8893,N_5873,N_4163);
and U8894 (N_8894,N_4798,N_5890);
or U8895 (N_8895,N_4341,N_3083);
and U8896 (N_8896,N_5811,N_5749);
nand U8897 (N_8897,N_4542,N_4900);
xor U8898 (N_8898,N_3211,N_3314);
nor U8899 (N_8899,N_5825,N_3712);
or U8900 (N_8900,N_5974,N_4701);
and U8901 (N_8901,N_4947,N_4853);
nand U8902 (N_8902,N_4101,N_3686);
nand U8903 (N_8903,N_5200,N_5359);
nand U8904 (N_8904,N_5474,N_5152);
and U8905 (N_8905,N_4201,N_3051);
nand U8906 (N_8906,N_5115,N_3751);
nor U8907 (N_8907,N_3480,N_4660);
and U8908 (N_8908,N_5600,N_4787);
nand U8909 (N_8909,N_5616,N_3484);
nor U8910 (N_8910,N_5367,N_3547);
or U8911 (N_8911,N_5582,N_5542);
nor U8912 (N_8912,N_4168,N_4977);
nand U8913 (N_8913,N_5091,N_3573);
nor U8914 (N_8914,N_4701,N_3569);
or U8915 (N_8915,N_5930,N_4387);
nor U8916 (N_8916,N_5638,N_3390);
nand U8917 (N_8917,N_3494,N_5079);
nor U8918 (N_8918,N_3949,N_4748);
nand U8919 (N_8919,N_4361,N_5051);
and U8920 (N_8920,N_3647,N_5789);
nor U8921 (N_8921,N_4289,N_4780);
and U8922 (N_8922,N_3304,N_5143);
or U8923 (N_8923,N_3451,N_3286);
or U8924 (N_8924,N_3809,N_4452);
or U8925 (N_8925,N_3122,N_3422);
nor U8926 (N_8926,N_4490,N_3872);
and U8927 (N_8927,N_5258,N_3983);
or U8928 (N_8928,N_4904,N_4413);
nor U8929 (N_8929,N_5189,N_5247);
nor U8930 (N_8930,N_4741,N_4164);
nor U8931 (N_8931,N_4948,N_5240);
nor U8932 (N_8932,N_4147,N_3144);
nand U8933 (N_8933,N_4052,N_5516);
nand U8934 (N_8934,N_5629,N_5977);
nor U8935 (N_8935,N_5585,N_4264);
xor U8936 (N_8936,N_3138,N_5872);
nor U8937 (N_8937,N_3834,N_3917);
and U8938 (N_8938,N_5439,N_5517);
and U8939 (N_8939,N_5822,N_3456);
or U8940 (N_8940,N_5175,N_5767);
nand U8941 (N_8941,N_5482,N_5891);
nand U8942 (N_8942,N_3181,N_4913);
nand U8943 (N_8943,N_5781,N_4825);
nor U8944 (N_8944,N_5533,N_3056);
nor U8945 (N_8945,N_5617,N_5210);
and U8946 (N_8946,N_4130,N_5536);
or U8947 (N_8947,N_4063,N_3779);
and U8948 (N_8948,N_5870,N_5468);
nor U8949 (N_8949,N_5761,N_3213);
and U8950 (N_8950,N_5650,N_3647);
nor U8951 (N_8951,N_4895,N_4325);
nor U8952 (N_8952,N_4778,N_5264);
xor U8953 (N_8953,N_3556,N_3685);
or U8954 (N_8954,N_3143,N_4105);
nand U8955 (N_8955,N_4035,N_3735);
nor U8956 (N_8956,N_3623,N_4393);
and U8957 (N_8957,N_5300,N_4552);
nor U8958 (N_8958,N_3611,N_5442);
and U8959 (N_8959,N_4439,N_3002);
nor U8960 (N_8960,N_3820,N_4103);
xor U8961 (N_8961,N_4168,N_5322);
or U8962 (N_8962,N_3808,N_5443);
nand U8963 (N_8963,N_3792,N_5517);
nand U8964 (N_8964,N_5267,N_4624);
or U8965 (N_8965,N_5284,N_4370);
nand U8966 (N_8966,N_4351,N_4939);
nor U8967 (N_8967,N_5186,N_5528);
xor U8968 (N_8968,N_4881,N_5628);
and U8969 (N_8969,N_5093,N_3270);
nand U8970 (N_8970,N_3727,N_5626);
xnor U8971 (N_8971,N_4880,N_5403);
and U8972 (N_8972,N_5059,N_5868);
or U8973 (N_8973,N_4026,N_5046);
and U8974 (N_8974,N_5677,N_5651);
and U8975 (N_8975,N_3870,N_4437);
and U8976 (N_8976,N_5927,N_5644);
nand U8977 (N_8977,N_5630,N_4212);
or U8978 (N_8978,N_3492,N_3134);
nand U8979 (N_8979,N_4425,N_3189);
nor U8980 (N_8980,N_4648,N_3244);
nor U8981 (N_8981,N_3557,N_4237);
nor U8982 (N_8982,N_3750,N_5930);
or U8983 (N_8983,N_4455,N_5421);
nor U8984 (N_8984,N_4596,N_5379);
and U8985 (N_8985,N_3115,N_5867);
or U8986 (N_8986,N_5021,N_4599);
nand U8987 (N_8987,N_5366,N_3227);
and U8988 (N_8988,N_3848,N_5391);
or U8989 (N_8989,N_4917,N_3287);
nor U8990 (N_8990,N_5283,N_5316);
nand U8991 (N_8991,N_5331,N_3015);
or U8992 (N_8992,N_3392,N_5274);
or U8993 (N_8993,N_5395,N_5141);
nor U8994 (N_8994,N_5854,N_3784);
nand U8995 (N_8995,N_5633,N_5329);
and U8996 (N_8996,N_5481,N_3774);
nand U8997 (N_8997,N_5733,N_3241);
or U8998 (N_8998,N_5241,N_5069);
or U8999 (N_8999,N_3049,N_4563);
nand U9000 (N_9000,N_7761,N_8672);
or U9001 (N_9001,N_8349,N_6217);
nand U9002 (N_9002,N_6844,N_7991);
or U9003 (N_9003,N_8350,N_8867);
and U9004 (N_9004,N_6654,N_6470);
nand U9005 (N_9005,N_7777,N_6629);
nand U9006 (N_9006,N_7268,N_7569);
and U9007 (N_9007,N_6040,N_8066);
and U9008 (N_9008,N_6863,N_8243);
and U9009 (N_9009,N_8206,N_7898);
and U9010 (N_9010,N_7771,N_7190);
and U9011 (N_9011,N_8965,N_7403);
nor U9012 (N_9012,N_7257,N_8214);
nand U9013 (N_9013,N_8938,N_6353);
nand U9014 (N_9014,N_6072,N_6609);
and U9015 (N_9015,N_8664,N_6797);
or U9016 (N_9016,N_6801,N_6739);
and U9017 (N_9017,N_6909,N_6548);
xnor U9018 (N_9018,N_7920,N_6652);
nand U9019 (N_9019,N_6299,N_8132);
nand U9020 (N_9020,N_6558,N_6443);
nor U9021 (N_9021,N_8401,N_7361);
nand U9022 (N_9022,N_7576,N_6897);
nor U9023 (N_9023,N_7938,N_7187);
or U9024 (N_9024,N_8986,N_6850);
nor U9025 (N_9025,N_7559,N_6700);
nor U9026 (N_9026,N_7947,N_7234);
nand U9027 (N_9027,N_8949,N_7389);
or U9028 (N_9028,N_6529,N_8930);
nand U9029 (N_9029,N_7445,N_8038);
and U9030 (N_9030,N_7285,N_7504);
or U9031 (N_9031,N_7850,N_7732);
nand U9032 (N_9032,N_6900,N_8115);
and U9033 (N_9033,N_7435,N_8203);
and U9034 (N_9034,N_8872,N_7049);
and U9035 (N_9035,N_6263,N_8688);
or U9036 (N_9036,N_6424,N_8495);
and U9037 (N_9037,N_7451,N_7260);
and U9038 (N_9038,N_8530,N_7349);
nand U9039 (N_9039,N_8735,N_8476);
nand U9040 (N_9040,N_8659,N_6525);
nand U9041 (N_9041,N_8977,N_8674);
or U9042 (N_9042,N_8760,N_7527);
and U9043 (N_9043,N_8900,N_7604);
nor U9044 (N_9044,N_7314,N_6378);
and U9045 (N_9045,N_7873,N_6054);
nand U9046 (N_9046,N_6685,N_6199);
nand U9047 (N_9047,N_7002,N_6163);
nor U9048 (N_9048,N_7201,N_8817);
nor U9049 (N_9049,N_7994,N_8703);
nor U9050 (N_9050,N_7607,N_7958);
nor U9051 (N_9051,N_8962,N_8791);
nor U9052 (N_9052,N_6522,N_8311);
and U9053 (N_9053,N_6971,N_8542);
or U9054 (N_9054,N_7829,N_8671);
and U9055 (N_9055,N_7337,N_8597);
or U9056 (N_9056,N_6584,N_6273);
or U9057 (N_9057,N_6912,N_7172);
nand U9058 (N_9058,N_7238,N_8314);
and U9059 (N_9059,N_8711,N_8380);
or U9060 (N_9060,N_7969,N_7227);
or U9061 (N_9061,N_8549,N_8513);
and U9062 (N_9062,N_6058,N_7459);
nor U9063 (N_9063,N_7714,N_6240);
and U9064 (N_9064,N_7057,N_7622);
and U9065 (N_9065,N_6032,N_8886);
xor U9066 (N_9066,N_6095,N_6143);
or U9067 (N_9067,N_7155,N_7617);
nor U9068 (N_9068,N_8830,N_6567);
nor U9069 (N_9069,N_6330,N_6042);
nand U9070 (N_9070,N_7375,N_6021);
nand U9071 (N_9071,N_6406,N_7768);
xor U9072 (N_9072,N_8546,N_7409);
or U9073 (N_9073,N_6446,N_8563);
and U9074 (N_9074,N_8719,N_6591);
nand U9075 (N_9075,N_6890,N_8718);
nor U9076 (N_9076,N_6827,N_8839);
nor U9077 (N_9077,N_8357,N_8754);
or U9078 (N_9078,N_7779,N_6628);
or U9079 (N_9079,N_6917,N_8544);
nor U9080 (N_9080,N_7264,N_6796);
xnor U9081 (N_9081,N_8560,N_6921);
nor U9082 (N_9082,N_6483,N_6869);
nand U9083 (N_9083,N_7140,N_8063);
nor U9084 (N_9084,N_6288,N_6445);
or U9085 (N_9085,N_7654,N_8741);
nand U9086 (N_9086,N_7970,N_7022);
and U9087 (N_9087,N_8358,N_7119);
nor U9088 (N_9088,N_8072,N_7081);
nand U9089 (N_9089,N_7594,N_7426);
or U9090 (N_9090,N_8590,N_6212);
nand U9091 (N_9091,N_6216,N_8832);
nand U9092 (N_9092,N_8390,N_7490);
nor U9093 (N_9093,N_7399,N_6825);
and U9094 (N_9094,N_8406,N_7668);
and U9095 (N_9095,N_7987,N_7997);
nor U9096 (N_9096,N_7376,N_7046);
nor U9097 (N_9097,N_6762,N_8606);
and U9098 (N_9098,N_6998,N_7808);
or U9099 (N_9099,N_8870,N_6510);
and U9100 (N_9100,N_8047,N_7858);
xor U9101 (N_9101,N_8103,N_6784);
nand U9102 (N_9102,N_7674,N_8764);
or U9103 (N_9103,N_7304,N_8275);
and U9104 (N_9104,N_7014,N_7996);
nand U9105 (N_9105,N_8890,N_8693);
nand U9106 (N_9106,N_7791,N_8681);
nor U9107 (N_9107,N_8141,N_8086);
and U9108 (N_9108,N_8224,N_8685);
nand U9109 (N_9109,N_8241,N_8716);
xor U9110 (N_9110,N_7918,N_8228);
nand U9111 (N_9111,N_7064,N_6806);
and U9112 (N_9112,N_8407,N_6368);
nand U9113 (N_9113,N_6104,N_8852);
nor U9114 (N_9114,N_8222,N_7070);
or U9115 (N_9115,N_7683,N_8581);
or U9116 (N_9116,N_6868,N_8185);
nor U9117 (N_9117,N_6956,N_8759);
and U9118 (N_9118,N_6624,N_7783);
nor U9119 (N_9119,N_6943,N_7378);
nor U9120 (N_9120,N_7432,N_8985);
and U9121 (N_9121,N_6933,N_8457);
nand U9122 (N_9122,N_6901,N_8950);
nor U9123 (N_9123,N_7041,N_8437);
or U9124 (N_9124,N_6246,N_8005);
or U9125 (N_9125,N_7466,N_6154);
nand U9126 (N_9126,N_8580,N_6575);
or U9127 (N_9127,N_8013,N_7967);
and U9128 (N_9128,N_6644,N_8212);
or U9129 (N_9129,N_6012,N_6655);
and U9130 (N_9130,N_6767,N_8289);
or U9131 (N_9131,N_7083,N_7018);
nor U9132 (N_9132,N_8814,N_6551);
nand U9133 (N_9133,N_8745,N_8248);
and U9134 (N_9134,N_7862,N_6907);
nand U9135 (N_9135,N_8118,N_6803);
nand U9136 (N_9136,N_6795,N_6794);
nor U9137 (N_9137,N_7501,N_7878);
nand U9138 (N_9138,N_6047,N_8253);
nand U9139 (N_9139,N_6476,N_7185);
nor U9140 (N_9140,N_8533,N_8129);
and U9141 (N_9141,N_6602,N_8936);
nand U9142 (N_9142,N_7618,N_6536);
or U9143 (N_9143,N_7439,N_8720);
nor U9144 (N_9144,N_8677,N_7724);
and U9145 (N_9145,N_8998,N_7306);
and U9146 (N_9146,N_6607,N_6265);
nand U9147 (N_9147,N_8687,N_6307);
and U9148 (N_9148,N_7675,N_7123);
nand U9149 (N_9149,N_7692,N_6277);
xnor U9150 (N_9150,N_6127,N_8299);
nand U9151 (N_9151,N_8270,N_7927);
and U9152 (N_9152,N_6218,N_8502);
or U9153 (N_9153,N_8413,N_8761);
and U9154 (N_9154,N_6948,N_6405);
and U9155 (N_9155,N_8307,N_8082);
or U9156 (N_9156,N_8097,N_8249);
or U9157 (N_9157,N_7799,N_7186);
nand U9158 (N_9158,N_6695,N_7735);
or U9159 (N_9159,N_8566,N_7658);
nor U9160 (N_9160,N_7343,N_8440);
or U9161 (N_9161,N_8381,N_6589);
and U9162 (N_9162,N_6489,N_6701);
xnor U9163 (N_9163,N_8925,N_7999);
and U9164 (N_9164,N_6671,N_8956);
and U9165 (N_9165,N_6229,N_7300);
and U9166 (N_9166,N_7952,N_8062);
or U9167 (N_9167,N_6696,N_6592);
or U9168 (N_9168,N_7525,N_8026);
or U9169 (N_9169,N_6281,N_6922);
nor U9170 (N_9170,N_7224,N_7008);
nor U9171 (N_9171,N_7897,N_7117);
or U9172 (N_9172,N_8445,N_6219);
nor U9173 (N_9173,N_8922,N_8098);
and U9174 (N_9174,N_7101,N_6531);
nor U9175 (N_9175,N_8901,N_8859);
or U9176 (N_9176,N_8699,N_7762);
nand U9177 (N_9177,N_7701,N_6732);
and U9178 (N_9178,N_8827,N_8242);
or U9179 (N_9179,N_6730,N_7077);
nor U9180 (N_9180,N_7621,N_6515);
xor U9181 (N_9181,N_7367,N_8015);
and U9182 (N_9182,N_8067,N_6464);
and U9183 (N_9183,N_6289,N_7354);
nand U9184 (N_9184,N_6455,N_8747);
nor U9185 (N_9185,N_8993,N_8004);
nor U9186 (N_9186,N_6244,N_6395);
or U9187 (N_9187,N_6512,N_8539);
nand U9188 (N_9188,N_6003,N_7784);
and U9189 (N_9189,N_6761,N_7360);
or U9190 (N_9190,N_7637,N_7239);
and U9191 (N_9191,N_8154,N_6503);
nor U9192 (N_9192,N_6735,N_7757);
nand U9193 (N_9193,N_6559,N_8351);
nor U9194 (N_9194,N_6731,N_7442);
nor U9195 (N_9195,N_7011,N_8421);
and U9196 (N_9196,N_8712,N_8377);
and U9197 (N_9197,N_8807,N_6486);
or U9198 (N_9198,N_7158,N_8702);
or U9199 (N_9199,N_8447,N_6996);
nor U9200 (N_9200,N_7189,N_7464);
nor U9201 (N_9201,N_6383,N_8497);
and U9202 (N_9202,N_6411,N_7096);
or U9203 (N_9203,N_7339,N_7847);
nor U9204 (N_9204,N_7831,N_6133);
nor U9205 (N_9205,N_8419,N_7549);
or U9206 (N_9206,N_7250,N_7720);
nand U9207 (N_9207,N_8803,N_7192);
nand U9208 (N_9208,N_6360,N_7157);
and U9209 (N_9209,N_8891,N_7145);
nand U9210 (N_9210,N_7323,N_7864);
or U9211 (N_9211,N_7523,N_6672);
nand U9212 (N_9212,N_7254,N_7796);
nor U9213 (N_9213,N_6285,N_7785);
nand U9214 (N_9214,N_8967,N_8060);
or U9215 (N_9215,N_8435,N_6543);
nor U9216 (N_9216,N_6019,N_7148);
nand U9217 (N_9217,N_7910,N_8861);
or U9218 (N_9218,N_6995,N_7372);
or U9219 (N_9219,N_8823,N_8519);
nor U9220 (N_9220,N_7136,N_6679);
xor U9221 (N_9221,N_6164,N_7362);
and U9222 (N_9222,N_8194,N_6849);
nor U9223 (N_9223,N_6439,N_8011);
xor U9224 (N_9224,N_7826,N_7957);
nand U9225 (N_9225,N_6247,N_7792);
nand U9226 (N_9226,N_8575,N_6600);
nand U9227 (N_9227,N_6842,N_7919);
or U9228 (N_9228,N_8752,N_6699);
or U9229 (N_9229,N_8984,N_6684);
or U9230 (N_9230,N_8928,N_7861);
or U9231 (N_9231,N_7695,N_8648);
nand U9232 (N_9232,N_8298,N_8442);
or U9233 (N_9233,N_6898,N_7028);
nor U9234 (N_9234,N_7039,N_6793);
and U9235 (N_9235,N_7905,N_7547);
nand U9236 (N_9236,N_8053,N_8085);
or U9237 (N_9237,N_8518,N_8087);
nor U9238 (N_9238,N_7258,N_6804);
and U9239 (N_9239,N_7382,N_7840);
nand U9240 (N_9240,N_6179,N_7038);
or U9241 (N_9241,N_6328,N_7043);
and U9242 (N_9242,N_8520,N_6677);
and U9243 (N_9243,N_6430,N_6810);
or U9244 (N_9244,N_8918,N_8835);
and U9245 (N_9245,N_7823,N_6755);
nand U9246 (N_9246,N_7122,N_6829);
and U9247 (N_9247,N_8731,N_8904);
nor U9248 (N_9248,N_8051,N_6860);
nand U9249 (N_9249,N_6335,N_6769);
nor U9250 (N_9250,N_6322,N_7556);
nor U9251 (N_9251,N_8090,N_7244);
nor U9252 (N_9252,N_8216,N_6450);
and U9253 (N_9253,N_6749,N_7428);
and U9254 (N_9254,N_6135,N_6286);
or U9255 (N_9255,N_8866,N_7803);
or U9256 (N_9256,N_8199,N_6595);
nor U9257 (N_9257,N_6474,N_8468);
nand U9258 (N_9258,N_7537,N_8170);
nor U9259 (N_9259,N_8075,N_6471);
nand U9260 (N_9260,N_6283,N_6858);
nand U9261 (N_9261,N_6945,N_7310);
and U9262 (N_9262,N_6018,N_8286);
xnor U9263 (N_9263,N_7591,N_8198);
and U9264 (N_9264,N_6968,N_6932);
and U9265 (N_9265,N_7587,N_6924);
nor U9266 (N_9266,N_7972,N_7265);
and U9267 (N_9267,N_6751,N_7699);
xor U9268 (N_9268,N_8217,N_6087);
nand U9269 (N_9269,N_6076,N_6402);
nor U9270 (N_9270,N_8151,N_7742);
and U9271 (N_9271,N_8422,N_6970);
nor U9272 (N_9272,N_6560,N_8610);
and U9273 (N_9273,N_7857,N_8283);
nand U9274 (N_9274,N_6305,N_6715);
and U9275 (N_9275,N_8055,N_7709);
nand U9276 (N_9276,N_6946,N_6852);
nand U9277 (N_9277,N_6243,N_8376);
and U9278 (N_9278,N_8880,N_6190);
nand U9279 (N_9279,N_6657,N_6991);
or U9280 (N_9280,N_7819,N_8816);
or U9281 (N_9281,N_6332,N_7769);
or U9282 (N_9282,N_6582,N_8043);
nor U9283 (N_9283,N_7468,N_8439);
nor U9284 (N_9284,N_6656,N_7739);
nand U9285 (N_9285,N_8698,N_8319);
nand U9286 (N_9286,N_8410,N_8924);
or U9287 (N_9287,N_8364,N_6653);
or U9288 (N_9288,N_6459,N_6209);
or U9289 (N_9289,N_7383,N_8997);
nor U9290 (N_9290,N_8465,N_8080);
nor U9291 (N_9291,N_6027,N_7210);
nor U9292 (N_9292,N_7960,N_6440);
nand U9293 (N_9293,N_7109,N_6638);
and U9294 (N_9294,N_6557,N_7945);
and U9295 (N_9295,N_7753,N_6588);
nor U9296 (N_9296,N_7072,N_8460);
nand U9297 (N_9297,N_7270,N_7390);
nand U9298 (N_9298,N_6119,N_6640);
nor U9299 (N_9299,N_7429,N_7998);
and U9300 (N_9300,N_8981,N_8430);
and U9301 (N_9301,N_6905,N_7191);
or U9302 (N_9302,N_7213,N_6276);
or U9303 (N_9303,N_8205,N_8767);
nand U9304 (N_9304,N_7004,N_7906);
and U9305 (N_9305,N_7029,N_7651);
nand U9306 (N_9306,N_6051,N_8142);
or U9307 (N_9307,N_6437,N_8802);
nor U9308 (N_9308,N_7682,N_6091);
and U9309 (N_9309,N_8751,N_7402);
or U9310 (N_9310,N_6747,N_8521);
and U9311 (N_9311,N_7763,N_7040);
nor U9312 (N_9312,N_8774,N_8140);
or U9313 (N_9313,N_7939,N_6848);
nor U9314 (N_9314,N_7685,N_6130);
or U9315 (N_9315,N_8078,N_8436);
or U9316 (N_9316,N_8596,N_6181);
and U9317 (N_9317,N_7843,N_8303);
xnor U9318 (N_9318,N_7180,N_7794);
nand U9319 (N_9319,N_6815,N_7838);
and U9320 (N_9320,N_8424,N_6310);
or U9321 (N_9321,N_6166,N_7240);
xnor U9322 (N_9322,N_6903,N_8130);
nor U9323 (N_9323,N_7131,N_7931);
nand U9324 (N_9324,N_7641,N_7955);
and U9325 (N_9325,N_7759,N_6052);
or U9326 (N_9326,N_6986,N_7216);
or U9327 (N_9327,N_7017,N_7849);
nor U9328 (N_9328,N_8039,N_8854);
and U9329 (N_9329,N_6385,N_6239);
and U9330 (N_9330,N_8598,N_8279);
and U9331 (N_9331,N_6542,N_8257);
or U9332 (N_9332,N_7333,N_7448);
or U9333 (N_9333,N_6785,N_6547);
and U9334 (N_9334,N_7722,N_8446);
and U9335 (N_9335,N_7068,N_8244);
nor U9336 (N_9336,N_8683,N_8679);
nand U9337 (N_9337,N_6999,N_6641);
and U9338 (N_9338,N_8510,N_7539);
nand U9339 (N_9339,N_7859,N_6663);
or U9340 (N_9340,N_8669,N_7635);
or U9341 (N_9341,N_8869,N_7916);
xnor U9342 (N_9342,N_7454,N_6646);
xor U9343 (N_9343,N_7434,N_7252);
and U9344 (N_9344,N_8775,N_7624);
nand U9345 (N_9345,N_8344,N_8846);
and U9346 (N_9346,N_8779,N_6981);
or U9347 (N_9347,N_7817,N_8336);
nor U9348 (N_9348,N_8148,N_7295);
nor U9349 (N_9349,N_6833,N_7359);
nor U9350 (N_9350,N_8695,N_6121);
nor U9351 (N_9351,N_8232,N_8980);
and U9352 (N_9352,N_6538,N_8696);
nand U9353 (N_9353,N_6528,N_8149);
nand U9354 (N_9354,N_6098,N_8161);
and U9355 (N_9355,N_8739,N_7369);
nand U9356 (N_9356,N_8027,N_7659);
and U9357 (N_9357,N_7384,N_6422);
or U9358 (N_9358,N_7166,N_6908);
nand U9359 (N_9359,N_6182,N_6223);
or U9360 (N_9360,N_7542,N_8639);
and U9361 (N_9361,N_6851,N_8461);
nor U9362 (N_9362,N_7262,N_8804);
and U9363 (N_9363,N_6053,N_8907);
nor U9364 (N_9364,N_7853,N_8902);
nand U9365 (N_9365,N_8105,N_8632);
nor U9366 (N_9366,N_8534,N_7413);
and U9367 (N_9367,N_8507,N_6992);
and U9368 (N_9368,N_8793,N_7697);
or U9369 (N_9369,N_6936,N_7942);
or U9370 (N_9370,N_7610,N_6585);
or U9371 (N_9371,N_6065,N_7748);
nand U9372 (N_9372,N_7577,N_7645);
nor U9373 (N_9373,N_8272,N_8577);
and U9374 (N_9374,N_8554,N_6469);
nand U9375 (N_9375,N_6669,N_8167);
and U9376 (N_9376,N_8262,N_8813);
or U9377 (N_9377,N_8361,N_7342);
and U9378 (N_9378,N_6963,N_7476);
and U9379 (N_9379,N_7112,N_8858);
or U9380 (N_9380,N_7872,N_7626);
or U9381 (N_9381,N_8061,N_6911);
nand U9382 (N_9382,N_7400,N_7740);
and U9383 (N_9383,N_7221,N_7058);
or U9384 (N_9384,N_8010,N_6726);
or U9385 (N_9385,N_6085,N_8841);
nand U9386 (N_9386,N_6195,N_7608);
xor U9387 (N_9387,N_7143,N_8694);
nor U9388 (N_9388,N_8372,N_6934);
nor U9389 (N_9389,N_7822,N_8007);
and U9390 (N_9390,N_8076,N_7346);
or U9391 (N_9391,N_8193,N_7968);
nand U9392 (N_9392,N_7506,N_8294);
and U9393 (N_9393,N_6612,N_7477);
or U9394 (N_9394,N_8266,N_7115);
or U9395 (N_9395,N_7900,N_7449);
or U9396 (N_9396,N_7755,N_7782);
and U9397 (N_9397,N_6895,N_8240);
nor U9398 (N_9398,N_7188,N_7470);
and U9399 (N_9399,N_7089,N_8605);
and U9400 (N_9400,N_8874,N_8729);
nor U9401 (N_9401,N_8983,N_8146);
and U9402 (N_9402,N_6084,N_6577);
or U9403 (N_9403,N_8124,N_7632);
and U9404 (N_9404,N_6752,N_8293);
or U9405 (N_9405,N_6140,N_7907);
nand U9406 (N_9406,N_8789,N_8164);
nand U9407 (N_9407,N_6350,N_6165);
and U9408 (N_9408,N_6633,N_6108);
nor U9409 (N_9409,N_7025,N_8282);
nand U9410 (N_9410,N_6847,N_7596);
nor U9411 (N_9411,N_7666,N_7456);
or U9412 (N_9412,N_8996,N_7548);
nor U9413 (N_9413,N_6409,N_7135);
nor U9414 (N_9414,N_8658,N_7937);
xnor U9415 (N_9415,N_8656,N_6938);
xor U9416 (N_9416,N_7377,N_8678);
nor U9417 (N_9417,N_7540,N_6498);
nor U9418 (N_9418,N_6703,N_6710);
and U9419 (N_9419,N_7237,N_8200);
nor U9420 (N_9420,N_7243,N_8035);
nor U9421 (N_9421,N_8602,N_7107);
and U9422 (N_9422,N_6102,N_7461);
nand U9423 (N_9423,N_6782,N_8278);
nand U9424 (N_9424,N_6826,N_8946);
nand U9425 (N_9425,N_6566,N_6011);
and U9426 (N_9426,N_6708,N_7223);
nor U9427 (N_9427,N_7855,N_6959);
and U9428 (N_9428,N_7743,N_8989);
and U9429 (N_9429,N_6495,N_8943);
and U9430 (N_9430,N_6315,N_7567);
and U9431 (N_9431,N_6365,N_6606);
and U9432 (N_9432,N_7198,N_6442);
and U9433 (N_9433,N_6507,N_7214);
and U9434 (N_9434,N_6253,N_6105);
or U9435 (N_9435,N_6855,N_7248);
nand U9436 (N_9436,N_8139,N_7092);
and U9437 (N_9437,N_6064,N_8790);
and U9438 (N_9438,N_6312,N_8618);
nor U9439 (N_9439,N_6337,N_7446);
nor U9440 (N_9440,N_7793,N_7706);
nor U9441 (N_9441,N_8389,N_8144);
and U9442 (N_9442,N_8002,N_6928);
or U9443 (N_9443,N_7328,N_6024);
nand U9444 (N_9444,N_7356,N_6993);
and U9445 (N_9445,N_7329,N_8068);
nand U9446 (N_9446,N_6122,N_7655);
or U9447 (N_9447,N_7447,N_7228);
nor U9448 (N_9448,N_7042,N_7138);
nor U9449 (N_9449,N_6777,N_8366);
nand U9450 (N_9450,N_6293,N_6291);
and U9451 (N_9451,N_7475,N_7259);
and U9452 (N_9452,N_6242,N_7698);
and U9453 (N_9453,N_8196,N_7749);
or U9454 (N_9454,N_7868,N_8260);
or U9455 (N_9455,N_8528,N_7357);
and U9456 (N_9456,N_8123,N_6431);
or U9457 (N_9457,N_8210,N_7964);
xnor U9458 (N_9458,N_6729,N_8318);
nand U9459 (N_9459,N_6436,N_7275);
nor U9460 (N_9460,N_6448,N_7639);
or U9461 (N_9461,N_7084,N_7584);
and U9462 (N_9462,N_8589,N_7756);
and U9463 (N_9463,N_6960,N_6658);
xnor U9464 (N_9464,N_7544,N_7113);
or U9465 (N_9465,N_6904,N_8420);
nand U9466 (N_9466,N_6651,N_8786);
nand U9467 (N_9467,N_6568,N_6840);
and U9468 (N_9468,N_6327,N_8663);
or U9469 (N_9469,N_6834,N_7097);
nand U9470 (N_9470,N_8969,N_7892);
and U9471 (N_9471,N_8909,N_6808);
or U9472 (N_9472,N_8730,N_6925);
and U9473 (N_9473,N_8572,N_8360);
nand U9474 (N_9474,N_8339,N_8576);
nor U9475 (N_9475,N_8312,N_6838);
and U9476 (N_9476,N_6723,N_8523);
and U9477 (N_9477,N_6982,N_6613);
and U9478 (N_9478,N_8820,N_8255);
nor U9479 (N_9479,N_6026,N_7633);
and U9480 (N_9480,N_7325,N_6103);
nor U9481 (N_9481,N_8689,N_8021);
nand U9482 (N_9482,N_8717,N_6879);
xnor U9483 (N_9483,N_6241,N_7586);
nor U9484 (N_9484,N_6947,N_6579);
nor U9485 (N_9485,N_8583,N_6357);
and U9486 (N_9486,N_8635,N_6812);
and U9487 (N_9487,N_6728,N_6670);
nor U9488 (N_9488,N_7124,N_7851);
nand U9489 (N_9489,N_6514,N_7775);
and U9490 (N_9490,N_7269,N_6680);
or U9491 (N_9491,N_6033,N_7299);
and U9492 (N_9492,N_7572,N_7394);
xor U9493 (N_9493,N_8432,N_7168);
and U9494 (N_9494,N_6394,N_8882);
and U9495 (N_9495,N_7846,N_8819);
or U9496 (N_9496,N_6349,N_8675);
and U9497 (N_9497,N_7568,N_6080);
nor U9498 (N_9498,N_8825,N_8230);
and U9499 (N_9499,N_7047,N_6627);
and U9500 (N_9500,N_7730,N_7789);
nor U9501 (N_9501,N_7904,N_6683);
nand U9502 (N_9502,N_8746,N_8322);
nand U9503 (N_9503,N_7079,N_8443);
or U9504 (N_9504,N_7209,N_8231);
nor U9505 (N_9505,N_6974,N_7962);
nor U9506 (N_9506,N_6413,N_6472);
nor U9507 (N_9507,N_8175,N_7174);
nor U9508 (N_9508,N_7713,N_8961);
and U9509 (N_9509,N_8184,N_6191);
and U9510 (N_9510,N_6381,N_8955);
and U9511 (N_9511,N_8875,N_6799);
nor U9512 (N_9512,N_8765,N_6271);
nand U9513 (N_9513,N_7163,N_8171);
and U9514 (N_9514,N_8885,N_7781);
nand U9515 (N_9515,N_7911,N_8463);
or U9516 (N_9516,N_6180,N_8207);
xor U9517 (N_9517,N_8611,N_7580);
or U9518 (N_9518,N_8088,N_7592);
or U9519 (N_9519,N_7094,N_7035);
nor U9520 (N_9520,N_6261,N_7978);
and U9521 (N_9521,N_7984,N_8582);
nand U9522 (N_9522,N_7917,N_6206);
nand U9523 (N_9523,N_7553,N_8951);
or U9524 (N_9524,N_7886,N_8444);
and U9525 (N_9525,N_7233,N_6225);
nand U9526 (N_9526,N_7280,N_6137);
nand U9527 (N_9527,N_8926,N_7552);
nand U9528 (N_9528,N_7206,N_6738);
nand U9529 (N_9529,N_8849,N_6144);
and U9530 (N_9530,N_7737,N_8108);
nand U9531 (N_9531,N_7116,N_8792);
nand U9532 (N_9532,N_6372,N_6871);
nand U9533 (N_9533,N_7073,N_8603);
or U9534 (N_9534,N_7647,N_6099);
nor U9535 (N_9535,N_6036,N_7319);
nor U9536 (N_9536,N_6979,N_7102);
nand U9537 (N_9537,N_6964,N_7764);
nor U9538 (N_9538,N_7979,N_8706);
nand U9539 (N_9539,N_6720,N_7696);
xor U9540 (N_9540,N_8873,N_7474);
or U9541 (N_9541,N_7033,N_8726);
nand U9542 (N_9542,N_7640,N_8722);
or U9543 (N_9543,N_6113,N_8012);
nand U9544 (N_9544,N_6918,N_8238);
and U9545 (N_9545,N_8479,N_6043);
or U9546 (N_9546,N_8960,N_7989);
or U9547 (N_9547,N_6718,N_8050);
nand U9548 (N_9548,N_8391,N_7992);
nor U9549 (N_9549,N_7286,N_6620);
or U9550 (N_9550,N_6831,N_7393);
or U9551 (N_9551,N_8268,N_8769);
or U9552 (N_9552,N_6967,N_8968);
or U9553 (N_9553,N_8935,N_8482);
nand U9554 (N_9554,N_8809,N_8083);
and U9555 (N_9555,N_8405,N_6269);
nand U9556 (N_9556,N_6552,N_6038);
nand U9557 (N_9557,N_7121,N_8512);
nand U9558 (N_9558,N_7725,N_8315);
nand U9559 (N_9559,N_8174,N_7561);
nand U9560 (N_9560,N_6294,N_6088);
nor U9561 (N_9561,N_8190,N_7059);
xor U9562 (N_9562,N_6523,N_7313);
nand U9563 (N_9563,N_6200,N_8697);
nor U9564 (N_9564,N_6147,N_8821);
nor U9565 (N_9565,N_7691,N_7001);
and U9566 (N_9566,N_7496,N_8310);
nor U9567 (N_9567,N_7412,N_7932);
or U9568 (N_9568,N_6083,N_7149);
and U9569 (N_9569,N_7060,N_8213);
nor U9570 (N_9570,N_8971,N_6404);
and U9571 (N_9571,N_6006,N_8548);
or U9572 (N_9572,N_8888,N_8824);
nand U9573 (N_9573,N_8234,N_6989);
or U9574 (N_9574,N_6230,N_6321);
or U9575 (N_9575,N_7520,N_7289);
and U9576 (N_9576,N_6454,N_6174);
nor U9577 (N_9577,N_6766,N_7162);
nor U9578 (N_9578,N_6484,N_6603);
nand U9579 (N_9579,N_7982,N_7293);
and U9580 (N_9580,N_7871,N_7512);
nand U9581 (N_9581,N_6382,N_6231);
and U9582 (N_9582,N_6460,N_8288);
nor U9583 (N_9583,N_7603,N_8383);
nand U9584 (N_9584,N_7869,N_6391);
and U9585 (N_9585,N_6134,N_7205);
or U9586 (N_9586,N_8836,N_7667);
and U9587 (N_9587,N_6177,N_7108);
nor U9588 (N_9588,N_8628,N_6778);
nor U9589 (N_9589,N_8462,N_8114);
or U9590 (N_9590,N_7814,N_7277);
and U9591 (N_9591,N_8034,N_7754);
or U9592 (N_9592,N_8899,N_6030);
or U9593 (N_9593,N_7810,N_7194);
or U9594 (N_9594,N_8020,N_7051);
and U9595 (N_9595,N_8469,N_6705);
and U9596 (N_9596,N_7616,N_7723);
or U9597 (N_9597,N_7184,N_6876);
nand U9598 (N_9598,N_6973,N_8617);
or U9599 (N_9599,N_7845,N_8487);
nand U9600 (N_9600,N_7780,N_7220);
nand U9601 (N_9601,N_7401,N_8158);
and U9602 (N_9602,N_6881,N_7307);
nand U9603 (N_9603,N_8223,N_6082);
nor U9604 (N_9604,N_8177,N_7318);
or U9605 (N_9605,N_6714,N_6961);
nand U9606 (N_9606,N_7211,N_8599);
or U9607 (N_9607,N_6407,N_6549);
nand U9608 (N_9608,N_7075,N_8458);
or U9609 (N_9609,N_6513,N_8452);
nand U9610 (N_9610,N_6681,N_6724);
and U9611 (N_9611,N_7335,N_8600);
or U9612 (N_9612,N_8584,N_8428);
and U9613 (N_9613,N_6574,N_8195);
or U9614 (N_9614,N_8186,N_6820);
and U9615 (N_9615,N_8459,N_8058);
or U9616 (N_9616,N_6988,N_8626);
nand U9617 (N_9617,N_8089,N_6611);
or U9618 (N_9618,N_8737,N_7195);
or U9619 (N_9619,N_7054,N_7598);
or U9620 (N_9620,N_8555,N_8649);
and U9621 (N_9621,N_6167,N_7882);
nand U9622 (N_9622,N_6625,N_6110);
nor U9623 (N_9623,N_6880,N_7518);
or U9624 (N_9624,N_7712,N_6814);
nor U9625 (N_9625,N_8895,N_8192);
nor U9626 (N_9626,N_6790,N_6865);
nor U9627 (N_9627,N_8048,N_7327);
or U9628 (N_9628,N_7179,N_7574);
or U9629 (N_9629,N_6074,N_7835);
or U9630 (N_9630,N_6220,N_8493);
or U9631 (N_9631,N_6342,N_6532);
nand U9632 (N_9632,N_8914,N_6415);
nand U9633 (N_9633,N_8454,N_6224);
nand U9634 (N_9634,N_8806,N_6069);
or U9635 (N_9635,N_6867,N_6887);
or U9636 (N_9636,N_6758,N_7545);
or U9637 (N_9637,N_7636,N_7261);
or U9638 (N_9638,N_6425,N_7127);
nor U9639 (N_9639,N_6304,N_7818);
nand U9640 (N_9640,N_8107,N_7371);
and U9641 (N_9641,N_6770,N_7802);
nor U9642 (N_9642,N_6071,N_6910);
nand U9643 (N_9643,N_6746,N_8838);
nor U9644 (N_9644,N_8277,N_6093);
or U9645 (N_9645,N_8488,N_8837);
nand U9646 (N_9646,N_8101,N_6913);
or U9647 (N_9647,N_7881,N_6530);
nand U9648 (N_9648,N_6990,N_7164);
nand U9649 (N_9649,N_8438,N_7801);
or U9650 (N_9650,N_6444,N_6668);
nand U9651 (N_9651,N_7010,N_6045);
nor U9652 (N_9652,N_7330,N_8994);
nor U9653 (N_9653,N_7809,N_6951);
and U9654 (N_9654,N_6857,N_6853);
nand U9655 (N_9655,N_7657,N_8733);
or U9656 (N_9656,N_6587,N_6870);
nor U9657 (N_9657,N_6475,N_6189);
or U9658 (N_9658,N_7452,N_7813);
or U9659 (N_9659,N_8680,N_7833);
and U9660 (N_9660,N_8545,N_8906);
or U9661 (N_9661,N_8046,N_6623);
nand U9662 (N_9662,N_8889,N_6524);
nor U9663 (N_9663,N_7276,N_7225);
nand U9664 (N_9664,N_7745,N_8787);
or U9665 (N_9665,N_7585,N_8017);
nand U9666 (N_9666,N_6650,N_7896);
and U9667 (N_9667,N_6753,N_6396);
or U9668 (N_9668,N_7628,N_8978);
nand U9669 (N_9669,N_6356,N_8134);
and U9670 (N_9670,N_8074,N_8798);
nor U9671 (N_9671,N_6028,N_7161);
and U9672 (N_9672,N_8096,N_6287);
or U9673 (N_9673,N_6354,N_8707);
or U9674 (N_9674,N_6173,N_8550);
nand U9675 (N_9675,N_7729,N_6387);
nor U9676 (N_9676,N_6158,N_7993);
and U9677 (N_9677,N_8220,N_7538);
or U9678 (N_9678,N_6941,N_6118);
or U9679 (N_9679,N_6478,N_6333);
and U9680 (N_9680,N_8300,N_7746);
xor U9681 (N_9681,N_6075,N_7566);
and U9682 (N_9682,N_8415,N_8947);
or U9683 (N_9683,N_8547,N_6204);
nor U9684 (N_9684,N_7665,N_7006);
nand U9685 (N_9685,N_7928,N_7492);
nand U9686 (N_9686,N_8354,N_8368);
or U9687 (N_9687,N_8917,N_6211);
nor U9688 (N_9688,N_6233,N_8095);
or U9689 (N_9689,N_7772,N_8477);
nand U9690 (N_9690,N_7863,N_7629);
nor U9691 (N_9691,N_6346,N_7983);
and U9692 (N_9692,N_6434,N_7332);
or U9693 (N_9693,N_7133,N_8271);
nand U9694 (N_9694,N_8676,N_7926);
nor U9695 (N_9695,N_8499,N_7643);
nor U9696 (N_9696,N_6994,N_8749);
nand U9697 (N_9697,N_8109,N_6846);
or U9698 (N_9698,N_6234,N_6598);
nor U9699 (N_9699,N_6859,N_7877);
and U9700 (N_9700,N_8250,N_6236);
and U9701 (N_9701,N_8974,N_8333);
nand U9702 (N_9702,N_7336,N_8615);
nand U9703 (N_9703,N_8069,N_7142);
or U9704 (N_9704,N_7884,N_7550);
and U9705 (N_9705,N_7642,N_6416);
nor U9706 (N_9706,N_7705,N_6397);
nand U9707 (N_9707,N_8652,N_6061);
nand U9708 (N_9708,N_7595,N_6323);
nor U9709 (N_9709,N_8723,N_7024);
and U9710 (N_9710,N_6013,N_6920);
nand U9711 (N_9711,N_7848,N_7555);
nand U9712 (N_9712,N_8408,N_8896);
nor U9713 (N_9713,N_6719,N_8532);
and U9714 (N_9714,N_6935,N_8152);
nand U9715 (N_9715,N_6420,N_6073);
and U9716 (N_9716,N_6124,N_7508);
and U9717 (N_9717,N_8504,N_8348);
nand U9718 (N_9718,N_8157,N_6183);
nand U9719 (N_9719,N_7106,N_6813);
nor U9720 (N_9720,N_8166,N_6150);
or U9721 (N_9721,N_6886,N_6237);
nor U9722 (N_9722,N_8373,N_7126);
and U9723 (N_9723,N_7350,N_6884);
nand U9724 (N_9724,N_6340,N_6520);
or U9725 (N_9725,N_8147,N_8126);
and U9726 (N_9726,N_7291,N_6953);
or U9727 (N_9727,N_6516,N_7128);
nand U9728 (N_9728,N_6055,N_8274);
nor U9729 (N_9729,N_8168,N_7934);
or U9730 (N_9730,N_8397,N_6314);
nand U9731 (N_9731,N_8091,N_6818);
or U9732 (N_9732,N_6329,N_7348);
or U9733 (N_9733,N_7312,N_8850);
nand U9734 (N_9734,N_8952,N_8056);
nor U9735 (N_9735,N_7694,N_8860);
nor U9736 (N_9736,N_6160,N_6873);
and U9737 (N_9737,N_6453,N_8133);
nand U9738 (N_9738,N_6194,N_6573);
or U9739 (N_9739,N_8023,N_7410);
or U9740 (N_9740,N_8219,N_8338);
and U9741 (N_9741,N_6580,N_8226);
nor U9742 (N_9742,N_8715,N_8018);
nand U9743 (N_9743,N_8258,N_8834);
nor U9744 (N_9744,N_7480,N_8948);
and U9745 (N_9745,N_6107,N_7602);
and U9746 (N_9746,N_7153,N_7533);
or U9747 (N_9747,N_6016,N_6817);
and U9748 (N_9748,N_6148,N_7795);
nand U9749 (N_9749,N_6343,N_7478);
nor U9750 (N_9750,N_6494,N_6977);
or U9751 (N_9751,N_8799,N_6320);
and U9752 (N_9752,N_8742,N_7433);
and U9753 (N_9753,N_8579,N_8755);
nand U9754 (N_9754,N_8201,N_6352);
and U9755 (N_9755,N_7620,N_6334);
and U9756 (N_9756,N_7943,N_6081);
nor U9757 (N_9757,N_8225,N_7020);
or U9758 (N_9758,N_6358,N_6618);
and U9759 (N_9759,N_6090,N_6249);
nand U9760 (N_9760,N_7973,N_8708);
nor U9761 (N_9761,N_7457,N_6112);
nand U9762 (N_9762,N_8106,N_6937);
nand U9763 (N_9763,N_7774,N_7093);
nor U9764 (N_9764,N_8831,N_8173);
and U9765 (N_9765,N_6734,N_7649);
or U9766 (N_9766,N_8862,N_8910);
and U9767 (N_9767,N_6185,N_6149);
nor U9768 (N_9768,N_7811,N_7551);
nand U9769 (N_9769,N_6771,N_6264);
nor U9770 (N_9770,N_8857,N_8863);
or U9771 (N_9771,N_6954,N_7830);
nand U9772 (N_9772,N_8399,N_6787);
nand U9773 (N_9773,N_6046,N_6141);
nand U9774 (N_9774,N_8040,N_7631);
or U9775 (N_9775,N_7605,N_6693);
nand U9776 (N_9776,N_8209,N_6742);
or U9777 (N_9777,N_6980,N_6316);
or U9778 (N_9778,N_6213,N_8337);
and U9779 (N_9779,N_7103,N_6563);
and U9780 (N_9780,N_6421,N_7913);
nand U9781 (N_9781,N_8941,N_8921);
nand U9782 (N_9782,N_7027,N_7425);
nand U9783 (N_9783,N_7381,N_8578);
nor U9784 (N_9784,N_8165,N_7253);
or U9785 (N_9785,N_7950,N_8393);
xnor U9786 (N_9786,N_6126,N_7193);
nand U9787 (N_9787,N_7690,N_6914);
nor U9788 (N_9788,N_7946,N_8475);
nand U9789 (N_9789,N_6152,N_6717);
nand U9790 (N_9790,N_6756,N_7485);
nand U9791 (N_9791,N_6227,N_6070);
or U9792 (N_9792,N_8662,N_6649);
and U9793 (N_9793,N_8001,N_6596);
nand U9794 (N_9794,N_8117,N_6891);
nor U9795 (N_9795,N_8916,N_8254);
and U9796 (N_9796,N_7680,N_7170);
nand U9797 (N_9797,N_7090,N_7975);
nor U9798 (N_9798,N_8973,N_7440);
or U9799 (N_9799,N_6041,N_7521);
nand U9800 (N_9800,N_6639,N_7676);
or U9801 (N_9801,N_6517,N_6153);
or U9802 (N_9802,N_6260,N_8884);
and U9803 (N_9803,N_7719,N_8059);
or U9804 (N_9804,N_8394,N_6637);
or U9805 (N_9805,N_7509,N_6682);
nand U9806 (N_9806,N_6845,N_8567);
nand U9807 (N_9807,N_8571,N_7673);
nor U9808 (N_9808,N_8734,N_6768);
nor U9809 (N_9809,N_6800,N_8093);
and U9810 (N_9810,N_6196,N_6392);
nand U9811 (N_9811,N_6972,N_8363);
nor U9812 (N_9812,N_8267,N_8763);
and U9813 (N_9813,N_7100,N_7171);
or U9814 (N_9814,N_8116,N_8848);
nor U9815 (N_9815,N_8302,N_8022);
or U9816 (N_9816,N_8102,N_8370);
nor U9817 (N_9817,N_7944,N_7634);
nor U9818 (N_9818,N_6697,N_8833);
or U9819 (N_9819,N_6645,N_8434);
and U9820 (N_9820,N_8016,N_8306);
and U9821 (N_9821,N_6059,N_7052);
nor U9822 (N_9822,N_6306,N_6727);
and U9823 (N_9823,N_8490,N_6186);
or U9824 (N_9824,N_7797,N_7301);
nand U9825 (N_9825,N_6744,N_7340);
nand U9826 (N_9826,N_8145,N_6632);
xor U9827 (N_9827,N_6050,N_8281);
xor U9828 (N_9828,N_6039,N_7095);
nor U9829 (N_9829,N_7546,N_7575);
or U9830 (N_9830,N_8506,N_7294);
nor U9831 (N_9831,N_6789,N_6203);
or U9832 (N_9832,N_7895,N_7317);
and U9833 (N_9833,N_7511,N_6037);
nor U9834 (N_9834,N_8402,N_7397);
nor U9835 (N_9835,N_8263,N_7578);
or U9836 (N_9836,N_6590,N_8912);
and U9837 (N_9837,N_8897,N_6419);
and U9838 (N_9838,N_8531,N_8690);
and U9839 (N_9839,N_6282,N_6721);
xor U9840 (N_9840,N_7758,N_7866);
nand U9841 (N_9841,N_7747,N_8954);
nand U9842 (N_9842,N_6691,N_8481);
nor U9843 (N_9843,N_8384,N_6702);
or U9844 (N_9844,N_8218,N_7980);
nor U9845 (N_9845,N_6014,N_8137);
nand U9846 (N_9846,N_7693,N_7226);
nor U9847 (N_9847,N_7351,N_6210);
and U9848 (N_9848,N_7247,N_8753);
nand U9849 (N_9849,N_8673,N_7279);
and U9850 (N_9850,N_7599,N_6284);
and U9851 (N_9851,N_8525,N_6711);
or U9852 (N_9852,N_6930,N_7130);
or U9853 (N_9853,N_7807,N_7644);
and U9854 (N_9854,N_8188,N_8684);
or U9855 (N_9855,N_7703,N_8645);
or U9856 (N_9856,N_7582,N_6519);
and U9857 (N_9857,N_6272,N_7110);
nor U9858 (N_9858,N_8153,N_6296);
nor U9859 (N_9859,N_7085,N_7914);
and U9860 (N_9860,N_8776,N_6479);
nor U9861 (N_9861,N_8670,N_8379);
or U9862 (N_9862,N_8296,N_7650);
nor U9863 (N_9863,N_6508,N_8471);
and U9864 (N_9864,N_6092,N_6020);
or U9865 (N_9865,N_6426,N_7053);
or U9866 (N_9866,N_8908,N_6518);
nand U9867 (N_9867,N_6765,N_7613);
nand U9868 (N_9868,N_8728,N_8797);
or U9869 (N_9869,N_7689,N_7326);
or U9870 (N_9870,N_8536,N_6534);
or U9871 (N_9871,N_6722,N_7912);
nand U9872 (N_9872,N_7953,N_6151);
or U9873 (N_9873,N_6202,N_7623);
and U9874 (N_9874,N_7949,N_7165);
nor U9875 (N_9875,N_6408,N_8607);
and U9876 (N_9876,N_7066,N_6599);
nor U9877 (N_9877,N_6535,N_6608);
and U9878 (N_9878,N_7507,N_7612);
and U9879 (N_9879,N_6198,N_8202);
and U9880 (N_9880,N_8359,N_7062);
or U9881 (N_9881,N_6712,N_8427);
nand U9882 (N_9882,N_8565,N_8113);
nor U9883 (N_9883,N_8433,N_7954);
nand U9884 (N_9884,N_7660,N_6379);
nand U9885 (N_9885,N_8744,N_7707);
or U9886 (N_9886,N_8812,N_7661);
nor U9887 (N_9887,N_7874,N_8472);
and U9888 (N_9888,N_7935,N_7483);
nand U9889 (N_9889,N_6667,N_6376);
and U9890 (N_9890,N_8593,N_7593);
or U9891 (N_9891,N_6889,N_7263);
or U9892 (N_9892,N_8423,N_6029);
nor U9893 (N_9893,N_8633,N_7717);
nor U9894 (N_9894,N_6809,N_8127);
nand U9895 (N_9895,N_8033,N_7773);
or U9896 (N_9896,N_8375,N_8425);
and U9897 (N_9897,N_7738,N_7274);
or U9898 (N_9898,N_7614,N_7815);
and U9899 (N_9899,N_8541,N_7986);
and U9900 (N_9900,N_8757,N_6005);
nor U9901 (N_9901,N_8538,N_6488);
nand U9902 (N_9902,N_8176,N_6958);
nand U9903 (N_9903,N_7700,N_6745);
or U9904 (N_9904,N_6878,N_8614);
or U9905 (N_9905,N_8019,N_6393);
nor U9906 (N_9906,N_6115,N_7776);
nand U9907 (N_9907,N_7030,N_7411);
nand U9908 (N_9908,N_8100,N_8556);
and U9909 (N_9909,N_7308,N_8784);
and U9910 (N_9910,N_8251,N_7903);
and U9911 (N_9911,N_8937,N_6159);
nand U9912 (N_9912,N_6969,N_8505);
nor U9913 (N_9913,N_7366,N_7365);
nand U9914 (N_9914,N_8570,N_8622);
and U9915 (N_9915,N_8261,N_7806);
or U9916 (N_9916,N_7355,N_8842);
or U9917 (N_9917,N_6215,N_6791);
and U9918 (N_9918,N_6388,N_8162);
or U9919 (N_9919,N_7726,N_7812);
or U9920 (N_9920,N_7924,N_7888);
and U9921 (N_9921,N_6274,N_6676);
or U9922 (N_9922,N_8829,N_7368);
and U9923 (N_9923,N_6540,N_8092);
nand U9924 (N_9924,N_6001,N_6615);
nor U9925 (N_9925,N_7876,N_8844);
nor U9926 (N_9926,N_6781,N_8594);
or U9927 (N_9927,N_8416,N_7421);
nor U9928 (N_9928,N_6576,N_7995);
or U9929 (N_9929,N_8623,N_6364);
nand U9930 (N_9930,N_6931,N_6841);
nand U9931 (N_9931,N_8725,N_8041);
nor U9932 (N_9932,N_7290,N_6280);
nor U9933 (N_9933,N_8568,N_8933);
or U9934 (N_9934,N_8543,N_6664);
nand U9935 (N_9935,N_8478,N_8156);
nand U9936 (N_9936,N_6116,N_7150);
nand U9937 (N_9937,N_7686,N_8295);
nor U9938 (N_9938,N_8325,N_8448);
nand U9939 (N_9939,N_8285,N_7894);
or U9940 (N_9940,N_7579,N_8982);
nor U9941 (N_9941,N_7486,N_6690);
nand U9942 (N_9942,N_8898,N_6326);
or U9943 (N_9943,N_6302,N_6377);
or U9944 (N_9944,N_7437,N_7679);
and U9945 (N_9945,N_6317,N_7481);
and U9946 (N_9946,N_8738,N_8591);
nor U9947 (N_9947,N_6390,N_8028);
or U9948 (N_9948,N_8772,N_8245);
nor U9949 (N_9949,N_7284,N_8637);
nor U9950 (N_9950,N_8768,N_8343);
and U9951 (N_9951,N_7406,N_7590);
nor U9952 (N_9952,N_6266,N_8342);
nand U9953 (N_9953,N_7891,N_7414);
nor U9954 (N_9954,N_7203,N_6067);
nor U9955 (N_9955,N_8794,N_6049);
nor U9956 (N_9956,N_7303,N_8647);
and U9957 (N_9957,N_7646,N_8128);
nand U9958 (N_9958,N_7255,N_6197);
nor U9959 (N_9959,N_7990,N_7484);
or U9960 (N_9960,N_6386,N_8111);
nor U9961 (N_9961,N_8800,N_8485);
or U9962 (N_9962,N_8071,N_7741);
nor U9963 (N_9963,N_7118,N_6571);
nor U9964 (N_9964,N_6111,N_7517);
and U9965 (N_9965,N_7199,N_8612);
or U9966 (N_9966,N_7272,N_8211);
and U9967 (N_9967,N_6172,N_7472);
nor U9968 (N_9968,N_7798,N_8169);
nor U9969 (N_9969,N_8783,N_6944);
nand U9970 (N_9970,N_7526,N_8187);
nand U9971 (N_9971,N_7322,N_7821);
nand U9972 (N_9972,N_6581,N_6068);
nand U9973 (N_9973,N_8650,N_8378);
nand U9974 (N_9974,N_8624,N_6978);
or U9975 (N_9975,N_7499,N_8815);
or U9976 (N_9976,N_6145,N_8341);
and U9977 (N_9977,N_7334,N_8621);
nor U9978 (N_9978,N_7498,N_8332);
or U9979 (N_9979,N_6309,N_6497);
nand U9980 (N_9980,N_7767,N_7044);
and U9981 (N_9981,N_7208,N_8516);
nor U9982 (N_9982,N_6779,N_7839);
or U9983 (N_9983,N_7222,N_8498);
or U9984 (N_9984,N_7921,N_7296);
or U9985 (N_9985,N_8345,N_8273);
and U9986 (N_9986,N_6874,N_8327);
and U9987 (N_9987,N_6268,N_6120);
or U9988 (N_9988,N_6222,N_6255);
xnor U9989 (N_9989,N_7364,N_6187);
or U9990 (N_9990,N_6987,N_7557);
nand U9991 (N_9991,N_6836,N_6648);
nand U9992 (N_9992,N_7930,N_8411);
and U9993 (N_9993,N_7708,N_7977);
nor U9994 (N_9994,N_6616,N_8409);
or U9995 (N_9995,N_7687,N_8592);
and U9996 (N_9996,N_7497,N_8159);
nor U9997 (N_9997,N_7056,N_8451);
nor U9998 (N_9998,N_7321,N_8927);
or U9999 (N_9999,N_6776,N_6673);
or U10000 (N_10000,N_7899,N_7246);
nand U10001 (N_10001,N_6002,N_8045);
nand U10002 (N_10002,N_6458,N_7436);
and U10003 (N_10003,N_6146,N_8893);
nand U10004 (N_10004,N_6432,N_7974);
and U10005 (N_10005,N_8084,N_6926);
or U10006 (N_10006,N_8771,N_7023);
or U10007 (N_10007,N_8979,N_6984);
nor U10008 (N_10008,N_7305,N_7519);
nand U10009 (N_10009,N_8065,N_8509);
and U10010 (N_10010,N_6949,N_7005);
nor U10011 (N_10011,N_7236,N_8181);
and U10012 (N_10012,N_6290,N_6292);
nor U10013 (N_10013,N_6750,N_8191);
or U10014 (N_10014,N_6642,N_7182);
or U10015 (N_10015,N_7563,N_6355);
or U10016 (N_10016,N_7215,N_6438);
or U10017 (N_10017,N_7804,N_8456);
and U10018 (N_10018,N_8208,N_8121);
nand U10019 (N_10019,N_8651,N_8155);
or U10020 (N_10020,N_7408,N_6610);
nor U10021 (N_10021,N_8355,N_7879);
nand U10022 (N_10022,N_7071,N_8535);
nand U10023 (N_10023,N_8009,N_6089);
nor U10024 (N_10024,N_6894,N_6939);
or U10025 (N_10025,N_7731,N_8099);
or U10026 (N_10026,N_7852,N_8524);
and U10027 (N_10027,N_6123,N_8330);
and U10028 (N_10028,N_6345,N_6614);
or U10029 (N_10029,N_6830,N_6389);
and U10030 (N_10030,N_7832,N_8467);
nor U10031 (N_10031,N_8508,N_6660);
nor U10032 (N_10032,N_6902,N_6816);
and U10033 (N_10033,N_6544,N_8845);
or U10034 (N_10034,N_7144,N_7744);
or U10035 (N_10035,N_7453,N_8879);
and U10036 (N_10036,N_8903,N_7045);
nor U10037 (N_10037,N_7710,N_6007);
nor U10038 (N_10038,N_7528,N_8501);
xor U10039 (N_10039,N_8049,N_7570);
nor U10040 (N_10040,N_6862,N_8331);
nor U10041 (N_10041,N_8588,N_8247);
nand U10042 (N_10042,N_8486,N_6313);
and U10043 (N_10043,N_7000,N_6193);
nor U10044 (N_10044,N_8864,N_7026);
and U10045 (N_10045,N_8704,N_8031);
and U10046 (N_10046,N_8496,N_6000);
nor U10047 (N_10047,N_6593,N_8335);
and U10048 (N_10048,N_7581,N_6733);
and U10049 (N_10049,N_7311,N_8006);
nor U10050 (N_10050,N_8634,N_7370);
and U10051 (N_10051,N_6433,N_6570);
nand U10052 (N_10052,N_6057,N_8290);
or U10053 (N_10053,N_6096,N_6184);
nand U10054 (N_10054,N_6201,N_7141);
or U10055 (N_10055,N_7324,N_7320);
or U10056 (N_10056,N_6208,N_8229);
nor U10057 (N_10057,N_8178,N_7503);
and U10058 (N_10058,N_7147,N_6341);
nor U10059 (N_10059,N_6687,N_7420);
nand U10060 (N_10060,N_8362,N_7048);
or U10061 (N_10061,N_7893,N_7407);
nand U10062 (N_10062,N_6864,N_6207);
nor U10063 (N_10063,N_8808,N_6493);
nor U10064 (N_10064,N_7207,N_8052);
and U10065 (N_10065,N_7245,N_7494);
nor U10066 (N_10066,N_8644,N_8911);
nand U10067 (N_10067,N_6452,N_6539);
and U10068 (N_10068,N_8773,N_7902);
nand U10069 (N_10069,N_7653,N_6228);
or U10070 (N_10070,N_7063,N_8641);
and U10071 (N_10071,N_6463,N_7465);
and U10072 (N_10072,N_7656,N_8395);
and U10073 (N_10073,N_6399,N_6139);
and U10074 (N_10074,N_8110,N_6578);
nand U10075 (N_10075,N_8037,N_7790);
nand U10076 (N_10076,N_8094,N_7923);
or U10077 (N_10077,N_6117,N_6636);
and U10078 (N_10078,N_6952,N_6142);
and U10079 (N_10079,N_7455,N_8398);
and U10080 (N_10080,N_6843,N_7460);
or U10081 (N_10081,N_6772,N_6835);
nor U10082 (N_10082,N_6966,N_7589);
nor U10083 (N_10083,N_8944,N_7836);
or U10084 (N_10084,N_7601,N_8667);
nand U10085 (N_10085,N_7232,N_8483);
or U10086 (N_10086,N_8431,N_6605);
nor U10087 (N_10087,N_7513,N_8371);
xnor U10088 (N_10088,N_6561,N_8822);
nand U10089 (N_10089,N_6056,N_6348);
and U10090 (N_10090,N_7534,N_8595);
and U10091 (N_10091,N_6662,N_6919);
nand U10092 (N_10092,N_7287,N_8291);
nor U10093 (N_10093,N_6811,N_7890);
and U10094 (N_10094,N_8480,N_8387);
and U10095 (N_10095,N_7385,N_6214);
nand U10096 (N_10096,N_7627,N_8929);
and U10097 (N_10097,N_6361,N_8305);
or U10098 (N_10098,N_6366,N_8736);
and U10099 (N_10099,N_6832,N_6764);
nand U10100 (N_10100,N_6347,N_6526);
and U10101 (N_10101,N_6788,N_8077);
or U10102 (N_10102,N_6429,N_7860);
nand U10103 (N_10103,N_8700,N_6015);
and U10104 (N_10104,N_6965,N_7625);
nor U10105 (N_10105,N_7315,N_8915);
or U10106 (N_10106,N_8135,N_7736);
xor U10107 (N_10107,N_6866,N_7181);
nand U10108 (N_10108,N_8643,N_6686);
and U10109 (N_10109,N_8215,N_7345);
nor U10110 (N_10110,N_8365,N_7114);
nand U10111 (N_10111,N_8940,N_7202);
or U10112 (N_10112,N_8608,N_6940);
and U10113 (N_10113,N_7541,N_7176);
nor U10114 (N_10114,N_7443,N_8221);
nand U10115 (N_10115,N_6048,N_8732);
nand U10116 (N_10116,N_6725,N_6480);
and U10117 (N_10117,N_7529,N_6491);
or U10118 (N_10118,N_8713,N_8801);
nand U10119 (N_10119,N_8313,N_7733);
nand U10120 (N_10120,N_6748,N_8517);
or U10121 (N_10121,N_7536,N_7760);
nor U10122 (N_10122,N_7915,N_6802);
xnor U10123 (N_10123,N_6492,N_6128);
nand U10124 (N_10124,N_8855,N_6311);
or U10125 (N_10125,N_7431,N_7702);
or U10126 (N_10126,N_8453,N_6044);
or U10127 (N_10127,N_6359,N_7816);
xor U10128 (N_10128,N_8256,N_6773);
nand U10129 (N_10129,N_7505,N_6462);
and U10130 (N_10130,N_8905,N_7292);
and U10131 (N_10131,N_8682,N_7441);
or U10132 (N_10132,N_7134,N_6010);
nand U10133 (N_10133,N_8727,N_6872);
or U10134 (N_10134,N_6754,N_8418);
and U10135 (N_10135,N_8527,N_6643);
or U10136 (N_10136,N_7159,N_6461);
nor U10137 (N_10137,N_7600,N_8450);
nor U10138 (N_10138,N_7516,N_6506);
nor U10139 (N_10139,N_6819,N_6896);
nand U10140 (N_10140,N_6303,N_8710);
and U10141 (N_10141,N_7111,N_6270);
nand U10142 (N_10142,N_8064,N_8782);
nand U10143 (N_10143,N_6235,N_8721);
and U10144 (N_10144,N_7219,N_6401);
and U10145 (N_10145,N_6251,N_8104);
nor U10146 (N_10146,N_6647,N_6295);
and U10147 (N_10147,N_8160,N_8292);
or U10148 (N_10148,N_8122,N_7273);
xor U10149 (N_10149,N_6318,N_8492);
or U10150 (N_10150,N_8795,N_7391);
and U10151 (N_10151,N_7309,N_8923);
and U10152 (N_10152,N_7688,N_6985);
nand U10153 (N_10153,N_8382,N_8367);
and U10154 (N_10154,N_6906,N_6565);
nand U10155 (N_10155,N_8871,N_8204);
xnor U10156 (N_10156,N_8227,N_6562);
and U10157 (N_10157,N_8008,N_6275);
or U10158 (N_10158,N_7438,N_8029);
nor U10159 (N_10159,N_6155,N_6500);
or U10160 (N_10160,N_7217,N_6400);
nand U10161 (N_10161,N_6553,N_8449);
nor U10162 (N_10162,N_7825,N_8613);
nand U10163 (N_10163,N_8780,N_8881);
nand U10164 (N_10164,N_6774,N_8470);
or U10165 (N_10165,N_8609,N_8934);
xnor U10166 (N_10166,N_7105,N_6527);
nand U10167 (N_10167,N_8932,N_8329);
nor U10168 (N_10168,N_8970,N_6485);
and U10169 (N_10169,N_7200,N_7031);
or U10170 (N_10170,N_6798,N_6521);
nor U10171 (N_10171,N_7251,N_6583);
nand U10172 (N_10172,N_7936,N_7948);
nand U10173 (N_10173,N_8352,N_7985);
and U10174 (N_10174,N_8564,N_7597);
and U10175 (N_10175,N_6861,N_8604);
nor U10176 (N_10176,N_8259,N_8740);
nand U10177 (N_10177,N_6757,N_6248);
nor U10178 (N_10178,N_6892,N_7734);
nor U10179 (N_10179,N_8403,N_7088);
nand U10180 (N_10180,N_7450,N_8280);
nand U10181 (N_10181,N_7976,N_6367);
or U10182 (N_10182,N_6384,N_7611);
and U10183 (N_10183,N_7241,N_7565);
xnor U10184 (N_10184,N_7865,N_8586);
nand U10185 (N_10185,N_7271,N_7463);
or U10186 (N_10186,N_7638,N_6783);
and U10187 (N_10187,N_7415,N_6418);
nor U10188 (N_10188,N_7788,N_8638);
and U10189 (N_10189,N_7125,N_6077);
nor U10190 (N_10190,N_8308,N_7341);
nand U10191 (N_10191,N_7778,N_8748);
nand U10192 (N_10192,N_7671,N_6875);
or U10193 (N_10193,N_7524,N_7373);
nor U10194 (N_10194,N_7422,N_6854);
nor U10195 (N_10195,N_6792,N_8138);
nand U10196 (N_10196,N_8972,N_6621);
nor U10197 (N_10197,N_6630,N_7489);
or U10198 (N_10198,N_8356,N_6466);
or U10199 (N_10199,N_7560,N_7353);
xor U10200 (N_10200,N_7606,N_8426);
nand U10201 (N_10201,N_6035,N_8003);
nand U10202 (N_10202,N_8939,N_6821);
and U10203 (N_10203,N_6245,N_8958);
and U10204 (N_10204,N_6617,N_7473);
nor U10205 (N_10205,N_6572,N_7458);
nand U10206 (N_10206,N_7842,N_7530);
nor U10207 (N_10207,N_6499,N_7386);
nor U10208 (N_10208,N_8265,N_8179);
nand U10209 (N_10209,N_6063,N_8054);
nand U10210 (N_10210,N_6449,N_6062);
and U10211 (N_10211,N_8287,N_8236);
nand U10212 (N_10212,N_6665,N_6279);
nor U10213 (N_10213,N_6267,N_7281);
and U10214 (N_10214,N_7901,N_8320);
and U10215 (N_10215,N_6564,N_7834);
nor U10216 (N_10216,N_7854,N_7965);
xor U10217 (N_10217,N_7765,N_8276);
nor U10218 (N_10218,N_6300,N_6161);
nand U10219 (N_10219,N_8826,N_7078);
nand U10220 (N_10220,N_7302,N_6232);
nor U10221 (N_10221,N_8347,N_8112);
or U10222 (N_10222,N_7242,N_6957);
or U10223 (N_10223,N_8553,N_7146);
nand U10224 (N_10224,N_6477,N_6171);
nand U10225 (N_10225,N_7098,N_6175);
and U10226 (N_10226,N_7178,N_6427);
nor U10227 (N_10227,N_7019,N_7880);
and U10228 (N_10228,N_7358,N_8762);
nand U10229 (N_10229,N_6371,N_7664);
and U10230 (N_10230,N_6256,N_6129);
nor U10231 (N_10231,N_6008,N_8558);
and U10232 (N_10232,N_8374,N_7820);
nand U10233 (N_10233,N_6336,N_6856);
or U10234 (N_10234,N_7167,N_6916);
nor U10235 (N_10235,N_7069,N_8964);
nor U10236 (N_10236,N_8913,N_7331);
nor U10237 (N_10237,N_8627,N_6132);
xnor U10238 (N_10238,N_8284,N_7531);
or U10239 (N_10239,N_8919,N_7177);
nand U10240 (N_10240,N_7966,N_6688);
nand U10241 (N_10241,N_6162,N_7256);
nand U10242 (N_10242,N_6569,N_7824);
or U10243 (N_10243,N_6157,N_8587);
nor U10244 (N_10244,N_7500,N_6259);
and U10245 (N_10245,N_8992,N_6374);
nand U10246 (N_10246,N_6017,N_6325);
nor U10247 (N_10247,N_7396,N_6447);
nor U10248 (N_10248,N_6131,N_6807);
nand U10249 (N_10249,N_8429,N_6743);
or U10250 (N_10250,N_8619,N_7424);
or U10251 (N_10251,N_6976,N_6060);
and U10252 (N_10252,N_8392,N_6034);
nand U10253 (N_10253,N_7721,N_6136);
nor U10254 (N_10254,N_8750,N_7493);
xor U10255 (N_10255,N_8766,N_8321);
and U10256 (N_10256,N_8653,N_6205);
nor U10257 (N_10257,N_8851,N_7514);
and U10258 (N_10258,N_7352,N_6674);
nand U10259 (N_10259,N_8894,N_8892);
or U10260 (N_10260,N_6373,N_8143);
nand U10261 (N_10261,N_6505,N_7129);
and U10262 (N_10262,N_8876,N_7338);
xnor U10263 (N_10263,N_8636,N_7387);
nand U10264 (N_10264,N_7067,N_6250);
or U10265 (N_10265,N_7885,N_6252);
nand U10266 (N_10266,N_6004,N_7137);
and U10267 (N_10267,N_7388,N_6997);
and U10268 (N_10268,N_6839,N_6496);
nor U10269 (N_10269,N_7562,N_7663);
and U10270 (N_10270,N_7419,N_6828);
nor U10271 (N_10271,N_6533,N_8484);
or U10272 (N_10272,N_6983,N_8235);
nand U10273 (N_10273,N_8079,N_8865);
or U10274 (N_10274,N_7212,N_6176);
nand U10275 (N_10275,N_7065,N_6501);
nand U10276 (N_10276,N_8297,N_8995);
nor U10277 (N_10277,N_8665,N_7728);
or U10278 (N_10278,N_8070,N_8323);
or U10279 (N_10279,N_6414,N_8514);
nor U10280 (N_10280,N_8686,N_6504);
and U10281 (N_10281,N_6666,N_6339);
or U10282 (N_10282,N_6556,N_8000);
nand U10283 (N_10283,N_6915,N_7487);
and U10284 (N_10284,N_7961,N_8887);
nor U10285 (N_10285,N_8999,N_8559);
or U10286 (N_10286,N_8396,N_7909);
nand U10287 (N_10287,N_8692,N_8805);
or U10288 (N_10288,N_8966,N_7395);
and U10289 (N_10289,N_6022,N_7282);
or U10290 (N_10290,N_8625,N_8551);
and U10291 (N_10291,N_7956,N_7502);
and U10292 (N_10292,N_7183,N_8569);
and U10293 (N_10293,N_6950,N_6740);
and U10294 (N_10294,N_6226,N_6106);
or U10295 (N_10295,N_8705,N_6675);
and U10296 (N_10296,N_6899,N_7805);
nor U10297 (N_10297,N_8988,N_7230);
or U10298 (N_10298,N_7681,N_8136);
xnor U10299 (N_10299,N_6009,N_8620);
or U10300 (N_10300,N_6114,N_8334);
or U10301 (N_10301,N_6101,N_8957);
nand U10302 (N_10302,N_7471,N_7055);
xor U10303 (N_10303,N_8856,N_6482);
nor U10304 (N_10304,N_8466,N_8264);
nand U10305 (N_10305,N_7021,N_6713);
and U10306 (N_10306,N_7380,N_6546);
nor U10307 (N_10307,N_6369,N_8326);
nand U10308 (N_10308,N_6824,N_7564);
nor U10309 (N_10309,N_6955,N_8758);
and U10310 (N_10310,N_7941,N_8464);
nand U10311 (N_10311,N_8237,N_6601);
and U10312 (N_10312,N_8975,N_8585);
nand U10313 (N_10313,N_7196,N_6716);
and U10314 (N_10314,N_6188,N_6545);
nand U10315 (N_10315,N_8868,N_7648);
nor U10316 (N_10316,N_7482,N_7278);
and U10317 (N_10317,N_8853,N_7652);
nand U10318 (N_10318,N_8172,N_8150);
nand U10319 (N_10319,N_6597,N_7491);
nor U10320 (N_10320,N_8441,N_7875);
nor U10321 (N_10321,N_8630,N_8473);
or U10322 (N_10322,N_6403,N_6837);
nand U10323 (N_10323,N_6490,N_7086);
nand U10324 (N_10324,N_7266,N_7662);
nor U10325 (N_10325,N_6412,N_7363);
or U10326 (N_10326,N_7786,N_8877);
and U10327 (N_10327,N_7495,N_8511);
and U10328 (N_10328,N_7704,N_8119);
and U10329 (N_10329,N_6094,N_8976);
nand U10330 (N_10330,N_7173,N_6156);
or U10331 (N_10331,N_6278,N_8788);
nor U10332 (N_10332,N_6375,N_6079);
nand U10333 (N_10333,N_7933,N_7751);
and U10334 (N_10334,N_8120,N_7398);
or U10335 (N_10335,N_6221,N_8404);
nand U10336 (N_10336,N_7175,N_6502);
nand U10337 (N_10337,N_6923,N_8840);
nand U10338 (N_10338,N_6706,N_7669);
nor U10339 (N_10339,N_8529,N_8963);
nor U10340 (N_10340,N_8796,N_7615);
nor U10341 (N_10341,N_6659,N_8540);
and U10342 (N_10342,N_8417,N_6257);
and U10343 (N_10343,N_8990,N_7036);
or U10344 (N_10344,N_8131,N_6877);
xor U10345 (N_10345,N_6554,N_8655);
or U10346 (N_10346,N_7374,N_6736);
and U10347 (N_10347,N_7297,N_8269);
and U10348 (N_10348,N_6410,N_7867);
or U10349 (N_10349,N_8024,N_8959);
nor U10350 (N_10350,N_7750,N_6622);
xor U10351 (N_10351,N_6380,N_7711);
and U10352 (N_10352,N_6631,N_7479);
nor U10353 (N_10353,N_6759,N_6823);
or U10354 (N_10354,N_8810,N_8503);
nor U10355 (N_10355,N_8660,N_7104);
nand U10356 (N_10356,N_7837,N_6541);
and U10357 (N_10357,N_7283,N_8920);
or U10358 (N_10358,N_8987,N_8573);
or U10359 (N_10359,N_7050,N_7344);
or U10360 (N_10360,N_7929,N_8770);
nor U10361 (N_10361,N_7416,N_7515);
and U10362 (N_10362,N_8057,N_6786);
nand U10363 (N_10363,N_8304,N_8701);
nand U10364 (N_10364,N_8183,N_8042);
nand U10365 (N_10365,N_8030,N_6344);
nor U10366 (N_10366,N_6362,N_8557);
and U10367 (N_10367,N_7316,N_7922);
and U10368 (N_10368,N_8724,N_7951);
or U10369 (N_10369,N_7418,N_7554);
nor U10370 (N_10370,N_7430,N_7154);
xnor U10371 (N_10371,N_6078,N_6885);
or U10372 (N_10372,N_8654,N_7156);
nor U10373 (N_10373,N_7298,N_7870);
and U10374 (N_10374,N_7132,N_8455);
or U10375 (N_10375,N_6883,N_6398);
nand U10376 (N_10376,N_7015,N_7677);
and U10377 (N_10377,N_7012,N_7981);
and U10378 (N_10378,N_7488,N_6692);
or U10379 (N_10379,N_8601,N_8991);
or U10380 (N_10380,N_8163,N_8781);
nor U10381 (N_10381,N_6661,N_7034);
nor U10382 (N_10382,N_6707,N_8353);
nor U10383 (N_10383,N_6023,N_7003);
nor U10384 (N_10384,N_7160,N_8883);
or U10385 (N_10385,N_8317,N_7959);
nand U10386 (N_10386,N_8489,N_6468);
nor U10387 (N_10387,N_7076,N_7267);
and U10388 (N_10388,N_7152,N_6694);
or U10389 (N_10389,N_6324,N_7032);
nand U10390 (N_10390,N_8642,N_7787);
and U10391 (N_10391,N_6805,N_8252);
and U10392 (N_10392,N_8515,N_6301);
nand U10393 (N_10393,N_7715,N_6481);
or U10394 (N_10394,N_7883,N_6741);
nor U10395 (N_10395,N_8328,N_7971);
or U10396 (N_10396,N_6888,N_7404);
nand U10397 (N_10397,N_6297,N_7925);
or U10398 (N_10398,N_8388,N_7249);
nand U10399 (N_10399,N_7080,N_6192);
nand U10400 (N_10400,N_7197,N_7583);
or U10401 (N_10401,N_6169,N_8073);
nor U10402 (N_10402,N_7571,N_7609);
and U10403 (N_10403,N_6929,N_8500);
nor U10404 (N_10404,N_7672,N_6097);
and U10405 (N_10405,N_6298,N_7684);
nand U10406 (N_10406,N_6086,N_6351);
or U10407 (N_10407,N_6457,N_7462);
or U10408 (N_10408,N_7908,N_6537);
or U10409 (N_10409,N_7061,N_8316);
nor U10410 (N_10410,N_7074,N_7392);
nor U10411 (N_10411,N_7007,N_8036);
or U10412 (N_10412,N_7379,N_8032);
or U10413 (N_10413,N_7828,N_7588);
nand U10414 (N_10414,N_8661,N_8847);
nand U10415 (N_10415,N_7469,N_8522);
nand U10416 (N_10416,N_6689,N_8743);
or U10417 (N_10417,N_8691,N_6775);
or U10418 (N_10418,N_8014,N_8931);
and U10419 (N_10419,N_7423,N_6262);
nor U10420 (N_10420,N_7573,N_8189);
nand U10421 (N_10421,N_7218,N_7099);
and U10422 (N_10422,N_6594,N_8197);
and U10423 (N_10423,N_6238,N_6822);
or U10424 (N_10424,N_8246,N_7151);
and U10425 (N_10425,N_8945,N_6586);
nor U10426 (N_10426,N_7727,N_8494);
nand U10427 (N_10427,N_8709,N_8346);
and U10428 (N_10428,N_6025,N_6109);
nor U10429 (N_10429,N_8309,N_8369);
nand U10430 (N_10430,N_7522,N_8777);
nor U10431 (N_10431,N_6760,N_6882);
nor U10432 (N_10432,N_8640,N_7009);
and U10433 (N_10433,N_6619,N_6942);
nand U10434 (N_10434,N_6555,N_8385);
and U10435 (N_10435,N_6780,N_7827);
or U10436 (N_10436,N_8646,N_8025);
nor U10437 (N_10437,N_7716,N_6465);
and U10438 (N_10438,N_8414,N_8301);
nor U10439 (N_10439,N_8953,N_7856);
or U10440 (N_10440,N_8239,N_8657);
and U10441 (N_10441,N_6441,N_6178);
nor U10442 (N_10442,N_6363,N_6417);
nand U10443 (N_10443,N_6473,N_8474);
or U10444 (N_10444,N_8818,N_7766);
or U10445 (N_10445,N_8125,N_6370);
nor U10446 (N_10446,N_6331,N_7082);
nand U10447 (N_10447,N_8400,N_8785);
nor U10448 (N_10448,N_7013,N_8491);
nand U10449 (N_10449,N_8714,N_6634);
nor U10450 (N_10450,N_6487,N_7444);
nand U10451 (N_10451,N_7139,N_6737);
nand U10452 (N_10452,N_8340,N_6927);
nor U10453 (N_10453,N_6456,N_8828);
nand U10454 (N_10454,N_7204,N_6626);
and U10455 (N_10455,N_7800,N_7630);
or U10456 (N_10456,N_7467,N_6975);
or U10457 (N_10457,N_6254,N_7841);
nor U10458 (N_10458,N_8616,N_8843);
nand U10459 (N_10459,N_7169,N_6451);
or U10460 (N_10460,N_8811,N_7091);
and U10461 (N_10461,N_7087,N_7678);
or U10462 (N_10462,N_6704,N_7417);
nand U10463 (N_10463,N_8629,N_6962);
and U10464 (N_10464,N_8552,N_8324);
nand U10465 (N_10465,N_8562,N_6893);
nand U10466 (N_10466,N_6511,N_7120);
and U10467 (N_10467,N_8878,N_7535);
nor U10468 (N_10468,N_8561,N_6168);
nor U10469 (N_10469,N_8386,N_6428);
or U10470 (N_10470,N_7558,N_6258);
nor U10471 (N_10471,N_6423,N_6467);
nand U10472 (N_10472,N_7940,N_7427);
nor U10473 (N_10473,N_8233,N_6338);
nor U10474 (N_10474,N_7844,N_7532);
nor U10475 (N_10475,N_7016,N_8537);
or U10476 (N_10476,N_7889,N_7670);
and U10477 (N_10477,N_7037,N_6604);
xnor U10478 (N_10478,N_8044,N_6635);
or U10479 (N_10479,N_7988,N_8526);
or U10480 (N_10480,N_7770,N_8668);
or U10481 (N_10481,N_6763,N_6435);
or U10482 (N_10482,N_7752,N_7229);
or U10483 (N_10483,N_6100,N_8574);
nor U10484 (N_10484,N_7887,N_8182);
nor U10485 (N_10485,N_7543,N_7347);
nand U10486 (N_10486,N_8180,N_8942);
and U10487 (N_10487,N_6698,N_8412);
and U10488 (N_10488,N_6031,N_6138);
nand U10489 (N_10489,N_8778,N_7510);
nand U10490 (N_10490,N_6709,N_6125);
nand U10491 (N_10491,N_6678,N_6319);
and U10492 (N_10492,N_6509,N_6550);
nand U10493 (N_10493,N_7619,N_7235);
nand U10494 (N_10494,N_7231,N_7963);
nor U10495 (N_10495,N_6066,N_8081);
nor U10496 (N_10496,N_6170,N_6308);
nand U10497 (N_10497,N_7405,N_8756);
or U10498 (N_10498,N_7718,N_8631);
nor U10499 (N_10499,N_8666,N_7288);
and U10500 (N_10500,N_6815,N_8720);
and U10501 (N_10501,N_8485,N_6204);
nand U10502 (N_10502,N_6561,N_6408);
or U10503 (N_10503,N_6709,N_8027);
xnor U10504 (N_10504,N_6664,N_6037);
or U10505 (N_10505,N_6791,N_8181);
or U10506 (N_10506,N_7741,N_7528);
nand U10507 (N_10507,N_6410,N_7934);
or U10508 (N_10508,N_7830,N_8795);
or U10509 (N_10509,N_6190,N_6536);
nor U10510 (N_10510,N_7921,N_7153);
or U10511 (N_10511,N_7462,N_8065);
nand U10512 (N_10512,N_8896,N_8196);
and U10513 (N_10513,N_6310,N_7345);
xnor U10514 (N_10514,N_6656,N_7882);
or U10515 (N_10515,N_7019,N_7734);
nand U10516 (N_10516,N_6643,N_7100);
nand U10517 (N_10517,N_6680,N_6767);
nor U10518 (N_10518,N_7847,N_7622);
and U10519 (N_10519,N_6459,N_8512);
and U10520 (N_10520,N_6792,N_6778);
nand U10521 (N_10521,N_8188,N_8218);
and U10522 (N_10522,N_7859,N_6519);
xnor U10523 (N_10523,N_6408,N_7843);
nor U10524 (N_10524,N_8904,N_6470);
and U10525 (N_10525,N_8211,N_6470);
nand U10526 (N_10526,N_6107,N_7349);
or U10527 (N_10527,N_6054,N_8265);
nand U10528 (N_10528,N_8639,N_8150);
or U10529 (N_10529,N_6537,N_8580);
nand U10530 (N_10530,N_8005,N_8164);
nor U10531 (N_10531,N_8552,N_7154);
nand U10532 (N_10532,N_6929,N_8954);
or U10533 (N_10533,N_8075,N_7890);
xnor U10534 (N_10534,N_6415,N_7359);
xor U10535 (N_10535,N_8358,N_6744);
nor U10536 (N_10536,N_7273,N_6626);
and U10537 (N_10537,N_6478,N_7115);
nand U10538 (N_10538,N_8239,N_8207);
or U10539 (N_10539,N_6815,N_6590);
nand U10540 (N_10540,N_7443,N_7608);
nand U10541 (N_10541,N_6983,N_7385);
nor U10542 (N_10542,N_7892,N_7989);
or U10543 (N_10543,N_7688,N_6231);
or U10544 (N_10544,N_7087,N_6486);
nor U10545 (N_10545,N_8339,N_8287);
nor U10546 (N_10546,N_8209,N_6486);
nand U10547 (N_10547,N_8852,N_7990);
nand U10548 (N_10548,N_6496,N_8827);
nand U10549 (N_10549,N_8664,N_8205);
xnor U10550 (N_10550,N_8748,N_6261);
or U10551 (N_10551,N_7947,N_8520);
and U10552 (N_10552,N_7096,N_6164);
nor U10553 (N_10553,N_7742,N_6445);
nand U10554 (N_10554,N_8831,N_6004);
and U10555 (N_10555,N_6303,N_7920);
nand U10556 (N_10556,N_8342,N_7480);
nand U10557 (N_10557,N_7919,N_8184);
nor U10558 (N_10558,N_7492,N_7475);
nand U10559 (N_10559,N_8103,N_6058);
nand U10560 (N_10560,N_6004,N_8110);
nand U10561 (N_10561,N_6686,N_7869);
or U10562 (N_10562,N_7434,N_6252);
or U10563 (N_10563,N_8438,N_6815);
nand U10564 (N_10564,N_7530,N_7762);
or U10565 (N_10565,N_7710,N_6082);
and U10566 (N_10566,N_8352,N_6318);
or U10567 (N_10567,N_8044,N_8573);
or U10568 (N_10568,N_6564,N_8791);
nor U10569 (N_10569,N_7687,N_8303);
or U10570 (N_10570,N_7445,N_8766);
and U10571 (N_10571,N_6913,N_8614);
nor U10572 (N_10572,N_6749,N_7061);
or U10573 (N_10573,N_6141,N_7159);
nand U10574 (N_10574,N_6594,N_8658);
or U10575 (N_10575,N_8296,N_6192);
nor U10576 (N_10576,N_7960,N_6740);
nor U10577 (N_10577,N_6384,N_6471);
nand U10578 (N_10578,N_6893,N_6041);
and U10579 (N_10579,N_8992,N_7748);
nand U10580 (N_10580,N_8268,N_7436);
and U10581 (N_10581,N_7078,N_8801);
nand U10582 (N_10582,N_8403,N_7991);
xor U10583 (N_10583,N_8345,N_6569);
or U10584 (N_10584,N_7579,N_8409);
or U10585 (N_10585,N_6730,N_6685);
nand U10586 (N_10586,N_8251,N_8125);
nor U10587 (N_10587,N_7881,N_7271);
or U10588 (N_10588,N_7380,N_6035);
nand U10589 (N_10589,N_8508,N_8291);
nand U10590 (N_10590,N_8164,N_8627);
nor U10591 (N_10591,N_8937,N_7108);
nand U10592 (N_10592,N_8974,N_6228);
and U10593 (N_10593,N_7066,N_7678);
nand U10594 (N_10594,N_6447,N_8056);
or U10595 (N_10595,N_6448,N_6943);
nand U10596 (N_10596,N_8517,N_8773);
or U10597 (N_10597,N_6807,N_6298);
nor U10598 (N_10598,N_7070,N_6344);
and U10599 (N_10599,N_7707,N_6125);
xnor U10600 (N_10600,N_6226,N_7304);
nor U10601 (N_10601,N_8057,N_7296);
or U10602 (N_10602,N_8731,N_8922);
and U10603 (N_10603,N_8736,N_8165);
or U10604 (N_10604,N_8357,N_6513);
nor U10605 (N_10605,N_6202,N_7151);
or U10606 (N_10606,N_8866,N_7000);
or U10607 (N_10607,N_6758,N_6259);
or U10608 (N_10608,N_8140,N_6050);
or U10609 (N_10609,N_7249,N_6588);
nand U10610 (N_10610,N_6354,N_8834);
or U10611 (N_10611,N_6656,N_7108);
and U10612 (N_10612,N_6843,N_7194);
or U10613 (N_10613,N_8149,N_7625);
xnor U10614 (N_10614,N_6771,N_8273);
nand U10615 (N_10615,N_8203,N_7437);
nor U10616 (N_10616,N_8471,N_8934);
and U10617 (N_10617,N_7641,N_7963);
nor U10618 (N_10618,N_7481,N_7021);
and U10619 (N_10619,N_7747,N_8179);
nand U10620 (N_10620,N_7042,N_8625);
nand U10621 (N_10621,N_7885,N_7454);
nor U10622 (N_10622,N_7480,N_7838);
or U10623 (N_10623,N_6974,N_6336);
and U10624 (N_10624,N_7130,N_6053);
and U10625 (N_10625,N_7164,N_7313);
or U10626 (N_10626,N_7751,N_7778);
and U10627 (N_10627,N_6482,N_6069);
or U10628 (N_10628,N_6929,N_8278);
or U10629 (N_10629,N_6976,N_8829);
nand U10630 (N_10630,N_7529,N_6907);
nor U10631 (N_10631,N_8594,N_7337);
and U10632 (N_10632,N_7178,N_8519);
nor U10633 (N_10633,N_7439,N_6621);
xnor U10634 (N_10634,N_7820,N_7142);
and U10635 (N_10635,N_8047,N_8508);
nor U10636 (N_10636,N_8694,N_8791);
nand U10637 (N_10637,N_7320,N_7672);
nand U10638 (N_10638,N_8189,N_6828);
xor U10639 (N_10639,N_6869,N_8657);
nor U10640 (N_10640,N_6769,N_8806);
and U10641 (N_10641,N_7658,N_7345);
nor U10642 (N_10642,N_7860,N_6319);
or U10643 (N_10643,N_7292,N_7547);
nor U10644 (N_10644,N_7942,N_8592);
nor U10645 (N_10645,N_7266,N_6859);
xor U10646 (N_10646,N_8044,N_6227);
nand U10647 (N_10647,N_8560,N_6888);
nor U10648 (N_10648,N_7324,N_7592);
nor U10649 (N_10649,N_8408,N_6313);
and U10650 (N_10650,N_8483,N_7164);
nand U10651 (N_10651,N_7093,N_7762);
and U10652 (N_10652,N_7407,N_8825);
xnor U10653 (N_10653,N_6575,N_7925);
nor U10654 (N_10654,N_8458,N_8758);
nor U10655 (N_10655,N_8305,N_7219);
nor U10656 (N_10656,N_8548,N_6877);
nor U10657 (N_10657,N_6168,N_8101);
nor U10658 (N_10658,N_8033,N_7086);
or U10659 (N_10659,N_8216,N_7355);
and U10660 (N_10660,N_7919,N_8579);
and U10661 (N_10661,N_8486,N_8535);
nand U10662 (N_10662,N_7553,N_6808);
nor U10663 (N_10663,N_6403,N_8710);
nand U10664 (N_10664,N_7754,N_7506);
or U10665 (N_10665,N_7707,N_7548);
or U10666 (N_10666,N_8737,N_8490);
or U10667 (N_10667,N_6821,N_6026);
nor U10668 (N_10668,N_7064,N_8832);
and U10669 (N_10669,N_6712,N_8910);
nand U10670 (N_10670,N_8341,N_8258);
nand U10671 (N_10671,N_8693,N_8597);
or U10672 (N_10672,N_6809,N_8743);
and U10673 (N_10673,N_6250,N_7368);
and U10674 (N_10674,N_6527,N_7328);
nor U10675 (N_10675,N_8687,N_8338);
nand U10676 (N_10676,N_6500,N_8291);
nand U10677 (N_10677,N_6575,N_6752);
or U10678 (N_10678,N_8708,N_8514);
and U10679 (N_10679,N_7452,N_8420);
and U10680 (N_10680,N_7129,N_6200);
or U10681 (N_10681,N_6692,N_6450);
or U10682 (N_10682,N_7254,N_6061);
nor U10683 (N_10683,N_7736,N_7045);
nor U10684 (N_10684,N_6754,N_8715);
nand U10685 (N_10685,N_7417,N_8397);
xor U10686 (N_10686,N_8165,N_6290);
nand U10687 (N_10687,N_7010,N_8057);
nand U10688 (N_10688,N_6359,N_6913);
nand U10689 (N_10689,N_6091,N_6512);
nand U10690 (N_10690,N_6985,N_8724);
and U10691 (N_10691,N_7237,N_8259);
nand U10692 (N_10692,N_8857,N_8747);
and U10693 (N_10693,N_7588,N_8298);
or U10694 (N_10694,N_7644,N_7504);
or U10695 (N_10695,N_6325,N_8005);
xnor U10696 (N_10696,N_8724,N_8935);
and U10697 (N_10697,N_7151,N_8088);
nand U10698 (N_10698,N_6510,N_6608);
or U10699 (N_10699,N_8378,N_6923);
and U10700 (N_10700,N_6585,N_8838);
and U10701 (N_10701,N_6535,N_8534);
nor U10702 (N_10702,N_7155,N_6575);
and U10703 (N_10703,N_6975,N_7507);
nor U10704 (N_10704,N_7542,N_6989);
nand U10705 (N_10705,N_8173,N_6350);
and U10706 (N_10706,N_7089,N_6159);
or U10707 (N_10707,N_7343,N_7976);
nor U10708 (N_10708,N_7716,N_6996);
and U10709 (N_10709,N_6407,N_7494);
or U10710 (N_10710,N_6818,N_7694);
nand U10711 (N_10711,N_6067,N_7797);
nor U10712 (N_10712,N_8443,N_7792);
nor U10713 (N_10713,N_7133,N_8974);
and U10714 (N_10714,N_7157,N_8653);
nor U10715 (N_10715,N_8577,N_7840);
or U10716 (N_10716,N_8336,N_8037);
and U10717 (N_10717,N_6018,N_6758);
xor U10718 (N_10718,N_8524,N_6509);
and U10719 (N_10719,N_8669,N_6689);
nand U10720 (N_10720,N_8812,N_6847);
or U10721 (N_10721,N_8070,N_6753);
or U10722 (N_10722,N_8208,N_7410);
nor U10723 (N_10723,N_8778,N_7741);
nor U10724 (N_10724,N_6486,N_7384);
or U10725 (N_10725,N_7805,N_6066);
nand U10726 (N_10726,N_8443,N_7313);
nand U10727 (N_10727,N_8822,N_7848);
nand U10728 (N_10728,N_7846,N_8267);
or U10729 (N_10729,N_7857,N_8665);
nor U10730 (N_10730,N_8542,N_6243);
nor U10731 (N_10731,N_6039,N_8416);
or U10732 (N_10732,N_8393,N_7135);
and U10733 (N_10733,N_6136,N_7482);
nand U10734 (N_10734,N_7456,N_7102);
nor U10735 (N_10735,N_6434,N_7845);
or U10736 (N_10736,N_7896,N_8477);
or U10737 (N_10737,N_8920,N_7379);
and U10738 (N_10738,N_8271,N_7785);
and U10739 (N_10739,N_7518,N_6766);
or U10740 (N_10740,N_6954,N_6300);
nor U10741 (N_10741,N_6484,N_6644);
nor U10742 (N_10742,N_8056,N_7664);
xor U10743 (N_10743,N_8457,N_6267);
and U10744 (N_10744,N_8543,N_7225);
nand U10745 (N_10745,N_6515,N_7414);
or U10746 (N_10746,N_8216,N_7905);
xnor U10747 (N_10747,N_7104,N_6501);
or U10748 (N_10748,N_7183,N_6494);
nand U10749 (N_10749,N_6619,N_8214);
and U10750 (N_10750,N_8415,N_6327);
nor U10751 (N_10751,N_8194,N_8827);
nand U10752 (N_10752,N_8216,N_6217);
nor U10753 (N_10753,N_8836,N_8129);
nor U10754 (N_10754,N_6600,N_7128);
xnor U10755 (N_10755,N_6635,N_7320);
nand U10756 (N_10756,N_8029,N_7880);
nor U10757 (N_10757,N_7650,N_6920);
or U10758 (N_10758,N_6458,N_6755);
and U10759 (N_10759,N_6885,N_6175);
and U10760 (N_10760,N_7086,N_8990);
nand U10761 (N_10761,N_6919,N_7257);
and U10762 (N_10762,N_8764,N_8293);
or U10763 (N_10763,N_6725,N_6952);
or U10764 (N_10764,N_6408,N_7755);
nand U10765 (N_10765,N_6374,N_6599);
or U10766 (N_10766,N_6988,N_6248);
nor U10767 (N_10767,N_8597,N_6715);
and U10768 (N_10768,N_8514,N_7147);
nand U10769 (N_10769,N_6106,N_6797);
nand U10770 (N_10770,N_7901,N_7394);
nand U10771 (N_10771,N_7304,N_7213);
and U10772 (N_10772,N_7897,N_8324);
and U10773 (N_10773,N_8756,N_6571);
or U10774 (N_10774,N_6477,N_8004);
nor U10775 (N_10775,N_6542,N_8864);
nand U10776 (N_10776,N_7646,N_8450);
or U10777 (N_10777,N_8444,N_6625);
xnor U10778 (N_10778,N_8692,N_6826);
nand U10779 (N_10779,N_7369,N_8582);
nand U10780 (N_10780,N_6986,N_7202);
nand U10781 (N_10781,N_7485,N_7129);
nor U10782 (N_10782,N_7962,N_6549);
nand U10783 (N_10783,N_8516,N_8179);
or U10784 (N_10784,N_7307,N_8249);
nand U10785 (N_10785,N_8590,N_7554);
nor U10786 (N_10786,N_8844,N_6682);
or U10787 (N_10787,N_8263,N_6796);
and U10788 (N_10788,N_7844,N_8704);
nor U10789 (N_10789,N_6961,N_7896);
or U10790 (N_10790,N_8106,N_8035);
nor U10791 (N_10791,N_6663,N_6836);
nor U10792 (N_10792,N_6135,N_6352);
nor U10793 (N_10793,N_7155,N_7164);
or U10794 (N_10794,N_8116,N_7764);
nand U10795 (N_10795,N_8071,N_6077);
and U10796 (N_10796,N_8044,N_6263);
nor U10797 (N_10797,N_7296,N_6809);
nand U10798 (N_10798,N_8203,N_8603);
nor U10799 (N_10799,N_8681,N_6734);
and U10800 (N_10800,N_8119,N_6737);
nand U10801 (N_10801,N_8344,N_8245);
and U10802 (N_10802,N_8797,N_7968);
and U10803 (N_10803,N_6041,N_7619);
nor U10804 (N_10804,N_7030,N_8196);
xnor U10805 (N_10805,N_7484,N_8022);
or U10806 (N_10806,N_6305,N_7642);
and U10807 (N_10807,N_8731,N_8026);
nor U10808 (N_10808,N_6694,N_6742);
or U10809 (N_10809,N_6853,N_6384);
and U10810 (N_10810,N_7258,N_8599);
or U10811 (N_10811,N_8993,N_8999);
or U10812 (N_10812,N_8918,N_8210);
nor U10813 (N_10813,N_8167,N_6013);
nor U10814 (N_10814,N_7598,N_8434);
or U10815 (N_10815,N_6931,N_7032);
nand U10816 (N_10816,N_7799,N_6209);
nand U10817 (N_10817,N_8513,N_7462);
nor U10818 (N_10818,N_7668,N_8218);
and U10819 (N_10819,N_6712,N_7554);
or U10820 (N_10820,N_8390,N_7776);
nor U10821 (N_10821,N_6671,N_7895);
nand U10822 (N_10822,N_8408,N_7796);
nor U10823 (N_10823,N_8177,N_8016);
xor U10824 (N_10824,N_8269,N_8362);
nor U10825 (N_10825,N_8279,N_6639);
nand U10826 (N_10826,N_6603,N_8905);
nor U10827 (N_10827,N_8959,N_8482);
or U10828 (N_10828,N_8782,N_7391);
or U10829 (N_10829,N_7621,N_7381);
or U10830 (N_10830,N_8274,N_6400);
nor U10831 (N_10831,N_8934,N_7403);
xor U10832 (N_10832,N_8217,N_6774);
or U10833 (N_10833,N_8657,N_7994);
and U10834 (N_10834,N_8730,N_6848);
and U10835 (N_10835,N_8422,N_6742);
and U10836 (N_10836,N_6388,N_8347);
and U10837 (N_10837,N_8147,N_7777);
nand U10838 (N_10838,N_7765,N_6445);
nand U10839 (N_10839,N_8289,N_8823);
nand U10840 (N_10840,N_8925,N_6630);
nand U10841 (N_10841,N_6705,N_7701);
or U10842 (N_10842,N_7660,N_6693);
nor U10843 (N_10843,N_7534,N_7104);
or U10844 (N_10844,N_6504,N_7532);
nor U10845 (N_10845,N_8576,N_6337);
or U10846 (N_10846,N_7073,N_7754);
or U10847 (N_10847,N_8437,N_6835);
and U10848 (N_10848,N_6070,N_6359);
nand U10849 (N_10849,N_8219,N_7647);
nor U10850 (N_10850,N_7872,N_8215);
or U10851 (N_10851,N_7779,N_7206);
nand U10852 (N_10852,N_6360,N_6062);
nand U10853 (N_10853,N_8006,N_8882);
and U10854 (N_10854,N_6295,N_7340);
nor U10855 (N_10855,N_8759,N_7882);
nor U10856 (N_10856,N_8118,N_7067);
nand U10857 (N_10857,N_7123,N_8977);
or U10858 (N_10858,N_8693,N_7322);
nor U10859 (N_10859,N_8056,N_6575);
or U10860 (N_10860,N_6613,N_6305);
and U10861 (N_10861,N_6870,N_6090);
and U10862 (N_10862,N_6678,N_7629);
nor U10863 (N_10863,N_8463,N_8967);
nand U10864 (N_10864,N_8451,N_6571);
and U10865 (N_10865,N_8588,N_7794);
or U10866 (N_10866,N_6446,N_6664);
xnor U10867 (N_10867,N_6787,N_6223);
nor U10868 (N_10868,N_7973,N_6673);
xnor U10869 (N_10869,N_6704,N_8255);
nand U10870 (N_10870,N_7518,N_7843);
nand U10871 (N_10871,N_8475,N_6348);
nand U10872 (N_10872,N_7325,N_8051);
nor U10873 (N_10873,N_8095,N_6176);
or U10874 (N_10874,N_8687,N_7599);
or U10875 (N_10875,N_6980,N_8649);
or U10876 (N_10876,N_8367,N_8045);
nor U10877 (N_10877,N_8579,N_6196);
or U10878 (N_10878,N_7183,N_8205);
or U10879 (N_10879,N_6772,N_6998);
and U10880 (N_10880,N_7171,N_8930);
nand U10881 (N_10881,N_8665,N_6155);
or U10882 (N_10882,N_6270,N_8921);
and U10883 (N_10883,N_7522,N_6615);
nor U10884 (N_10884,N_7970,N_6041);
or U10885 (N_10885,N_6949,N_7640);
nand U10886 (N_10886,N_7325,N_6690);
nor U10887 (N_10887,N_7615,N_6075);
or U10888 (N_10888,N_6052,N_6255);
nor U10889 (N_10889,N_7989,N_6080);
nand U10890 (N_10890,N_7220,N_6445);
nand U10891 (N_10891,N_6917,N_8058);
and U10892 (N_10892,N_8484,N_7026);
and U10893 (N_10893,N_6618,N_8001);
nand U10894 (N_10894,N_8861,N_7498);
and U10895 (N_10895,N_7274,N_6049);
and U10896 (N_10896,N_6992,N_7317);
nor U10897 (N_10897,N_7715,N_6681);
or U10898 (N_10898,N_8533,N_7226);
nor U10899 (N_10899,N_6612,N_6985);
or U10900 (N_10900,N_6190,N_7811);
or U10901 (N_10901,N_7606,N_7638);
or U10902 (N_10902,N_8709,N_8836);
and U10903 (N_10903,N_6018,N_6239);
xor U10904 (N_10904,N_7293,N_8863);
nand U10905 (N_10905,N_6458,N_7068);
or U10906 (N_10906,N_6947,N_6534);
or U10907 (N_10907,N_8446,N_8897);
or U10908 (N_10908,N_6343,N_6174);
or U10909 (N_10909,N_8755,N_6959);
and U10910 (N_10910,N_8172,N_6716);
nand U10911 (N_10911,N_8092,N_7573);
nor U10912 (N_10912,N_8506,N_6402);
or U10913 (N_10913,N_7821,N_6105);
and U10914 (N_10914,N_6679,N_6303);
xor U10915 (N_10915,N_8113,N_7497);
and U10916 (N_10916,N_6327,N_7357);
and U10917 (N_10917,N_7997,N_6565);
and U10918 (N_10918,N_6169,N_7117);
nor U10919 (N_10919,N_8363,N_8837);
or U10920 (N_10920,N_6538,N_6267);
or U10921 (N_10921,N_8747,N_8108);
and U10922 (N_10922,N_6287,N_8950);
nor U10923 (N_10923,N_6011,N_6357);
or U10924 (N_10924,N_8546,N_6420);
or U10925 (N_10925,N_7685,N_6981);
nor U10926 (N_10926,N_8136,N_8783);
nand U10927 (N_10927,N_7837,N_8340);
nor U10928 (N_10928,N_7415,N_6776);
nor U10929 (N_10929,N_8339,N_6248);
or U10930 (N_10930,N_7210,N_6494);
nand U10931 (N_10931,N_6464,N_7382);
nand U10932 (N_10932,N_7231,N_6359);
or U10933 (N_10933,N_8670,N_6485);
nand U10934 (N_10934,N_7821,N_7046);
nand U10935 (N_10935,N_6458,N_8269);
nand U10936 (N_10936,N_6429,N_8830);
or U10937 (N_10937,N_8790,N_8410);
nand U10938 (N_10938,N_8082,N_8107);
or U10939 (N_10939,N_8748,N_8860);
or U10940 (N_10940,N_7302,N_8758);
and U10941 (N_10941,N_8147,N_7871);
nor U10942 (N_10942,N_7845,N_8022);
or U10943 (N_10943,N_6165,N_7263);
nand U10944 (N_10944,N_6383,N_8117);
or U10945 (N_10945,N_6302,N_7459);
and U10946 (N_10946,N_6683,N_8624);
nor U10947 (N_10947,N_8926,N_8252);
nand U10948 (N_10948,N_8168,N_6403);
and U10949 (N_10949,N_8191,N_6203);
or U10950 (N_10950,N_6221,N_7620);
and U10951 (N_10951,N_7140,N_8674);
and U10952 (N_10952,N_6226,N_6246);
nand U10953 (N_10953,N_8377,N_6593);
and U10954 (N_10954,N_6063,N_8821);
nor U10955 (N_10955,N_7401,N_6588);
nor U10956 (N_10956,N_6823,N_8178);
nor U10957 (N_10957,N_6008,N_6370);
nor U10958 (N_10958,N_6643,N_7340);
nand U10959 (N_10959,N_8362,N_7398);
and U10960 (N_10960,N_8155,N_6196);
nand U10961 (N_10961,N_8648,N_6510);
nor U10962 (N_10962,N_8741,N_6194);
nor U10963 (N_10963,N_6361,N_8727);
nand U10964 (N_10964,N_6318,N_6920);
or U10965 (N_10965,N_6115,N_7871);
or U10966 (N_10966,N_6792,N_6571);
xor U10967 (N_10967,N_8397,N_6113);
nor U10968 (N_10968,N_7429,N_7049);
nor U10969 (N_10969,N_7688,N_8005);
xnor U10970 (N_10970,N_8601,N_8956);
nor U10971 (N_10971,N_7703,N_8359);
nor U10972 (N_10972,N_7065,N_8294);
nand U10973 (N_10973,N_8454,N_6691);
or U10974 (N_10974,N_8295,N_6077);
nor U10975 (N_10975,N_6210,N_7055);
nor U10976 (N_10976,N_6867,N_7717);
or U10977 (N_10977,N_8714,N_8270);
xnor U10978 (N_10978,N_7156,N_7711);
or U10979 (N_10979,N_8365,N_6461);
nor U10980 (N_10980,N_6569,N_8970);
nand U10981 (N_10981,N_7214,N_7367);
and U10982 (N_10982,N_7060,N_6390);
or U10983 (N_10983,N_8303,N_7705);
nor U10984 (N_10984,N_6421,N_7659);
xnor U10985 (N_10985,N_6784,N_6264);
and U10986 (N_10986,N_6647,N_8857);
nand U10987 (N_10987,N_8377,N_8341);
nand U10988 (N_10988,N_8726,N_8538);
nor U10989 (N_10989,N_8116,N_8350);
nand U10990 (N_10990,N_7635,N_7469);
nand U10991 (N_10991,N_8008,N_7313);
nor U10992 (N_10992,N_8595,N_6298);
nand U10993 (N_10993,N_6937,N_6267);
nor U10994 (N_10994,N_6858,N_8741);
xor U10995 (N_10995,N_6713,N_7509);
xnor U10996 (N_10996,N_6258,N_7276);
nor U10997 (N_10997,N_6304,N_7823);
and U10998 (N_10998,N_6053,N_7537);
nor U10999 (N_10999,N_8250,N_7824);
or U11000 (N_11000,N_7207,N_7334);
and U11001 (N_11001,N_6466,N_6151);
nand U11002 (N_11002,N_7023,N_6512);
nor U11003 (N_11003,N_8051,N_8714);
nand U11004 (N_11004,N_8348,N_7441);
or U11005 (N_11005,N_6145,N_7515);
nor U11006 (N_11006,N_6306,N_7717);
nand U11007 (N_11007,N_8062,N_7232);
nor U11008 (N_11008,N_8518,N_7909);
and U11009 (N_11009,N_8158,N_7885);
nor U11010 (N_11010,N_8699,N_6465);
nand U11011 (N_11011,N_8405,N_6947);
nand U11012 (N_11012,N_8019,N_7531);
nor U11013 (N_11013,N_6002,N_8031);
nand U11014 (N_11014,N_6541,N_7171);
nor U11015 (N_11015,N_8623,N_7636);
and U11016 (N_11016,N_8303,N_8006);
and U11017 (N_11017,N_8411,N_7883);
or U11018 (N_11018,N_8873,N_8370);
nor U11019 (N_11019,N_7347,N_6141);
and U11020 (N_11020,N_6962,N_7202);
nor U11021 (N_11021,N_6046,N_6652);
nor U11022 (N_11022,N_7130,N_8878);
nor U11023 (N_11023,N_7055,N_8445);
or U11024 (N_11024,N_7611,N_6448);
or U11025 (N_11025,N_7706,N_8526);
and U11026 (N_11026,N_8299,N_6681);
nand U11027 (N_11027,N_7087,N_7860);
nor U11028 (N_11028,N_7116,N_6396);
nand U11029 (N_11029,N_6648,N_8339);
nand U11030 (N_11030,N_6068,N_6346);
and U11031 (N_11031,N_7776,N_8959);
nor U11032 (N_11032,N_8032,N_7703);
nand U11033 (N_11033,N_6960,N_8282);
nor U11034 (N_11034,N_6718,N_6338);
or U11035 (N_11035,N_6068,N_8385);
nand U11036 (N_11036,N_7747,N_8834);
nand U11037 (N_11037,N_7096,N_8587);
or U11038 (N_11038,N_7780,N_6437);
or U11039 (N_11039,N_8643,N_6827);
and U11040 (N_11040,N_6633,N_8821);
nor U11041 (N_11041,N_7944,N_6693);
nand U11042 (N_11042,N_6785,N_6985);
nor U11043 (N_11043,N_6563,N_6608);
nor U11044 (N_11044,N_6803,N_6894);
or U11045 (N_11045,N_8422,N_8125);
nor U11046 (N_11046,N_6511,N_6255);
or U11047 (N_11047,N_8201,N_7786);
and U11048 (N_11048,N_7074,N_6608);
nand U11049 (N_11049,N_8035,N_7759);
nand U11050 (N_11050,N_7925,N_8999);
nand U11051 (N_11051,N_8401,N_6807);
and U11052 (N_11052,N_7062,N_8448);
nand U11053 (N_11053,N_7929,N_6045);
nor U11054 (N_11054,N_8199,N_8993);
nor U11055 (N_11055,N_7083,N_8384);
and U11056 (N_11056,N_6772,N_8912);
and U11057 (N_11057,N_6887,N_6817);
and U11058 (N_11058,N_6526,N_8488);
and U11059 (N_11059,N_6746,N_6427);
nor U11060 (N_11060,N_6209,N_8112);
nand U11061 (N_11061,N_6740,N_7430);
or U11062 (N_11062,N_6397,N_7645);
and U11063 (N_11063,N_7380,N_8756);
nand U11064 (N_11064,N_8373,N_7153);
nor U11065 (N_11065,N_8951,N_6285);
or U11066 (N_11066,N_6234,N_7816);
nand U11067 (N_11067,N_7962,N_6976);
and U11068 (N_11068,N_6711,N_7829);
or U11069 (N_11069,N_6446,N_6682);
nor U11070 (N_11070,N_7534,N_8534);
and U11071 (N_11071,N_8254,N_8957);
or U11072 (N_11072,N_7584,N_7426);
or U11073 (N_11073,N_6480,N_6491);
or U11074 (N_11074,N_7228,N_6307);
nand U11075 (N_11075,N_8051,N_8707);
nor U11076 (N_11076,N_6522,N_7763);
nand U11077 (N_11077,N_8895,N_6189);
nand U11078 (N_11078,N_7352,N_8347);
and U11079 (N_11079,N_7214,N_8919);
and U11080 (N_11080,N_7473,N_6466);
xnor U11081 (N_11081,N_8075,N_6833);
nor U11082 (N_11082,N_8923,N_7135);
nor U11083 (N_11083,N_7519,N_8034);
nand U11084 (N_11084,N_6136,N_6882);
nor U11085 (N_11085,N_6842,N_7858);
or U11086 (N_11086,N_8162,N_6019);
nor U11087 (N_11087,N_7421,N_8307);
or U11088 (N_11088,N_8322,N_7260);
nand U11089 (N_11089,N_8629,N_6272);
and U11090 (N_11090,N_8577,N_7338);
nand U11091 (N_11091,N_8312,N_6223);
or U11092 (N_11092,N_8711,N_8392);
xor U11093 (N_11093,N_8183,N_6951);
or U11094 (N_11094,N_8668,N_6806);
nand U11095 (N_11095,N_7887,N_6403);
nor U11096 (N_11096,N_7116,N_7860);
nor U11097 (N_11097,N_6621,N_8660);
or U11098 (N_11098,N_8043,N_6047);
nand U11099 (N_11099,N_6740,N_7105);
and U11100 (N_11100,N_6700,N_8219);
nand U11101 (N_11101,N_8082,N_8267);
nor U11102 (N_11102,N_6273,N_8396);
or U11103 (N_11103,N_8461,N_6354);
and U11104 (N_11104,N_7076,N_8335);
or U11105 (N_11105,N_8760,N_8158);
nand U11106 (N_11106,N_7838,N_7959);
or U11107 (N_11107,N_8731,N_8073);
nand U11108 (N_11108,N_7761,N_6469);
nand U11109 (N_11109,N_7001,N_7356);
and U11110 (N_11110,N_6731,N_8382);
or U11111 (N_11111,N_6431,N_6758);
nand U11112 (N_11112,N_7899,N_7600);
and U11113 (N_11113,N_7187,N_8605);
or U11114 (N_11114,N_6627,N_7594);
nor U11115 (N_11115,N_7101,N_7615);
or U11116 (N_11116,N_6153,N_6004);
and U11117 (N_11117,N_6680,N_8020);
and U11118 (N_11118,N_6572,N_8653);
nor U11119 (N_11119,N_7348,N_7651);
and U11120 (N_11120,N_8825,N_8277);
nor U11121 (N_11121,N_7386,N_6594);
and U11122 (N_11122,N_8362,N_8523);
nand U11123 (N_11123,N_6296,N_7788);
or U11124 (N_11124,N_8776,N_7417);
nand U11125 (N_11125,N_7949,N_8618);
and U11126 (N_11126,N_8825,N_6238);
and U11127 (N_11127,N_6181,N_7425);
and U11128 (N_11128,N_6022,N_8288);
and U11129 (N_11129,N_8351,N_7433);
xnor U11130 (N_11130,N_6335,N_6823);
nor U11131 (N_11131,N_6044,N_8866);
and U11132 (N_11132,N_6706,N_8288);
nor U11133 (N_11133,N_6111,N_6263);
or U11134 (N_11134,N_7050,N_8356);
or U11135 (N_11135,N_7136,N_7135);
nand U11136 (N_11136,N_6472,N_8746);
nand U11137 (N_11137,N_7766,N_8999);
and U11138 (N_11138,N_6785,N_7109);
and U11139 (N_11139,N_7407,N_7644);
and U11140 (N_11140,N_6313,N_7235);
or U11141 (N_11141,N_7835,N_6833);
nand U11142 (N_11142,N_6715,N_7945);
nor U11143 (N_11143,N_6281,N_7891);
nand U11144 (N_11144,N_7186,N_6578);
and U11145 (N_11145,N_8152,N_6904);
nor U11146 (N_11146,N_7966,N_6383);
and U11147 (N_11147,N_7833,N_8790);
nand U11148 (N_11148,N_6170,N_6788);
or U11149 (N_11149,N_8608,N_6089);
or U11150 (N_11150,N_6847,N_6317);
or U11151 (N_11151,N_8874,N_8474);
nor U11152 (N_11152,N_7898,N_6379);
or U11153 (N_11153,N_6688,N_7104);
xor U11154 (N_11154,N_7442,N_6371);
and U11155 (N_11155,N_6792,N_6258);
nand U11156 (N_11156,N_6905,N_8956);
or U11157 (N_11157,N_7865,N_8529);
or U11158 (N_11158,N_6828,N_8198);
or U11159 (N_11159,N_6966,N_8566);
or U11160 (N_11160,N_8948,N_8541);
or U11161 (N_11161,N_6083,N_6344);
and U11162 (N_11162,N_7952,N_6644);
and U11163 (N_11163,N_7668,N_6678);
and U11164 (N_11164,N_7512,N_7337);
or U11165 (N_11165,N_6126,N_7415);
nand U11166 (N_11166,N_8988,N_8749);
nor U11167 (N_11167,N_7661,N_6473);
and U11168 (N_11168,N_8444,N_8921);
and U11169 (N_11169,N_7435,N_7351);
and U11170 (N_11170,N_6728,N_7787);
and U11171 (N_11171,N_8941,N_8082);
or U11172 (N_11172,N_8212,N_8754);
nand U11173 (N_11173,N_6936,N_6151);
nand U11174 (N_11174,N_7093,N_6873);
xnor U11175 (N_11175,N_6866,N_6101);
and U11176 (N_11176,N_8208,N_6360);
or U11177 (N_11177,N_8581,N_7695);
nor U11178 (N_11178,N_6966,N_7365);
or U11179 (N_11179,N_7453,N_7845);
nand U11180 (N_11180,N_7950,N_8503);
or U11181 (N_11181,N_6511,N_6236);
or U11182 (N_11182,N_7137,N_6595);
and U11183 (N_11183,N_8997,N_6259);
and U11184 (N_11184,N_7452,N_7124);
and U11185 (N_11185,N_8624,N_6987);
or U11186 (N_11186,N_8508,N_7842);
or U11187 (N_11187,N_6306,N_7983);
and U11188 (N_11188,N_6500,N_8123);
and U11189 (N_11189,N_7481,N_7787);
and U11190 (N_11190,N_6711,N_6772);
nor U11191 (N_11191,N_8486,N_6696);
nand U11192 (N_11192,N_7508,N_7085);
nand U11193 (N_11193,N_8931,N_8436);
nand U11194 (N_11194,N_7744,N_8083);
and U11195 (N_11195,N_6352,N_8475);
nor U11196 (N_11196,N_7426,N_8688);
nand U11197 (N_11197,N_6574,N_7381);
nor U11198 (N_11198,N_8220,N_7716);
or U11199 (N_11199,N_6950,N_7011);
nand U11200 (N_11200,N_6541,N_7949);
nor U11201 (N_11201,N_8580,N_6605);
nand U11202 (N_11202,N_8249,N_7352);
nor U11203 (N_11203,N_6473,N_8405);
nor U11204 (N_11204,N_8736,N_8030);
nand U11205 (N_11205,N_8264,N_6158);
or U11206 (N_11206,N_8197,N_7662);
nand U11207 (N_11207,N_7153,N_6110);
and U11208 (N_11208,N_6641,N_6474);
nand U11209 (N_11209,N_6998,N_7283);
nand U11210 (N_11210,N_6115,N_6140);
and U11211 (N_11211,N_7114,N_8668);
nand U11212 (N_11212,N_8026,N_6221);
or U11213 (N_11213,N_7182,N_7268);
and U11214 (N_11214,N_7926,N_6333);
and U11215 (N_11215,N_7120,N_8784);
or U11216 (N_11216,N_7861,N_8495);
nor U11217 (N_11217,N_6381,N_6807);
nor U11218 (N_11218,N_6271,N_8266);
and U11219 (N_11219,N_6427,N_6632);
xnor U11220 (N_11220,N_6885,N_8392);
nor U11221 (N_11221,N_6466,N_7274);
nor U11222 (N_11222,N_8423,N_6072);
nor U11223 (N_11223,N_8553,N_6052);
nand U11224 (N_11224,N_6731,N_8472);
or U11225 (N_11225,N_8191,N_6835);
nor U11226 (N_11226,N_6682,N_6235);
and U11227 (N_11227,N_7116,N_6257);
nand U11228 (N_11228,N_6126,N_7446);
and U11229 (N_11229,N_7331,N_7862);
or U11230 (N_11230,N_7352,N_8923);
nor U11231 (N_11231,N_8782,N_6432);
nand U11232 (N_11232,N_6770,N_7177);
nand U11233 (N_11233,N_8541,N_8608);
and U11234 (N_11234,N_6976,N_7620);
or U11235 (N_11235,N_6746,N_6793);
and U11236 (N_11236,N_7095,N_6950);
and U11237 (N_11237,N_7687,N_7053);
and U11238 (N_11238,N_6988,N_7837);
and U11239 (N_11239,N_8133,N_8277);
and U11240 (N_11240,N_8303,N_8850);
xor U11241 (N_11241,N_6065,N_6573);
or U11242 (N_11242,N_6328,N_6436);
and U11243 (N_11243,N_6260,N_7775);
nand U11244 (N_11244,N_8680,N_6746);
or U11245 (N_11245,N_8604,N_8885);
or U11246 (N_11246,N_7903,N_6244);
or U11247 (N_11247,N_6925,N_8195);
or U11248 (N_11248,N_6968,N_7548);
and U11249 (N_11249,N_6876,N_6692);
or U11250 (N_11250,N_6042,N_8447);
or U11251 (N_11251,N_8057,N_7722);
nor U11252 (N_11252,N_7854,N_6598);
and U11253 (N_11253,N_7998,N_6952);
nand U11254 (N_11254,N_8145,N_7095);
and U11255 (N_11255,N_7916,N_8489);
nand U11256 (N_11256,N_7722,N_6642);
and U11257 (N_11257,N_6697,N_7522);
nand U11258 (N_11258,N_6703,N_7716);
nor U11259 (N_11259,N_7607,N_7667);
xnor U11260 (N_11260,N_8500,N_8591);
and U11261 (N_11261,N_8875,N_8947);
nor U11262 (N_11262,N_6042,N_8944);
nand U11263 (N_11263,N_8476,N_8496);
and U11264 (N_11264,N_7347,N_7699);
nand U11265 (N_11265,N_7456,N_6007);
or U11266 (N_11266,N_7625,N_6648);
and U11267 (N_11267,N_6016,N_7039);
nand U11268 (N_11268,N_7059,N_8580);
nand U11269 (N_11269,N_6969,N_8276);
nand U11270 (N_11270,N_6888,N_6368);
or U11271 (N_11271,N_8258,N_6120);
and U11272 (N_11272,N_7799,N_6695);
nor U11273 (N_11273,N_8153,N_6728);
and U11274 (N_11274,N_8613,N_8920);
nand U11275 (N_11275,N_6277,N_6999);
nand U11276 (N_11276,N_6037,N_6996);
nor U11277 (N_11277,N_7337,N_6266);
or U11278 (N_11278,N_7048,N_8890);
and U11279 (N_11279,N_8808,N_7082);
nand U11280 (N_11280,N_6616,N_7566);
nand U11281 (N_11281,N_7335,N_8059);
nor U11282 (N_11282,N_7819,N_6588);
and U11283 (N_11283,N_6978,N_6316);
or U11284 (N_11284,N_7068,N_6806);
nand U11285 (N_11285,N_8423,N_6522);
and U11286 (N_11286,N_7748,N_7708);
nor U11287 (N_11287,N_7756,N_7387);
nand U11288 (N_11288,N_7420,N_6384);
nor U11289 (N_11289,N_7765,N_6594);
nand U11290 (N_11290,N_7200,N_8415);
or U11291 (N_11291,N_6557,N_6778);
nor U11292 (N_11292,N_7591,N_6725);
nor U11293 (N_11293,N_6356,N_6404);
nand U11294 (N_11294,N_7944,N_8898);
nor U11295 (N_11295,N_7847,N_6285);
xor U11296 (N_11296,N_7524,N_6344);
nand U11297 (N_11297,N_6314,N_6500);
and U11298 (N_11298,N_8188,N_8704);
nand U11299 (N_11299,N_8477,N_7853);
nand U11300 (N_11300,N_6500,N_8668);
nor U11301 (N_11301,N_6375,N_7002);
nor U11302 (N_11302,N_6310,N_6915);
and U11303 (N_11303,N_8746,N_7592);
nor U11304 (N_11304,N_6030,N_6420);
or U11305 (N_11305,N_7911,N_6713);
and U11306 (N_11306,N_6078,N_7242);
and U11307 (N_11307,N_6973,N_6968);
or U11308 (N_11308,N_8649,N_6541);
nand U11309 (N_11309,N_7253,N_8598);
or U11310 (N_11310,N_7808,N_7736);
nand U11311 (N_11311,N_8877,N_7045);
and U11312 (N_11312,N_6421,N_8938);
nand U11313 (N_11313,N_8181,N_8359);
nor U11314 (N_11314,N_6283,N_8785);
nor U11315 (N_11315,N_6904,N_8833);
and U11316 (N_11316,N_8578,N_6392);
nor U11317 (N_11317,N_7766,N_6387);
or U11318 (N_11318,N_8658,N_6704);
nand U11319 (N_11319,N_8625,N_8560);
and U11320 (N_11320,N_8846,N_6607);
nand U11321 (N_11321,N_6939,N_7424);
nor U11322 (N_11322,N_8170,N_8565);
nand U11323 (N_11323,N_8995,N_7354);
nand U11324 (N_11324,N_8940,N_6952);
or U11325 (N_11325,N_7487,N_7963);
nor U11326 (N_11326,N_6882,N_7040);
nand U11327 (N_11327,N_7945,N_7804);
and U11328 (N_11328,N_7196,N_8995);
nor U11329 (N_11329,N_8183,N_7489);
or U11330 (N_11330,N_6062,N_8970);
or U11331 (N_11331,N_8716,N_6572);
or U11332 (N_11332,N_7313,N_8770);
nor U11333 (N_11333,N_6804,N_6083);
or U11334 (N_11334,N_7188,N_7987);
or U11335 (N_11335,N_7340,N_7938);
or U11336 (N_11336,N_8344,N_7779);
and U11337 (N_11337,N_7190,N_6989);
nand U11338 (N_11338,N_7965,N_7376);
nand U11339 (N_11339,N_7990,N_6892);
nor U11340 (N_11340,N_7201,N_6250);
nor U11341 (N_11341,N_6919,N_7554);
nand U11342 (N_11342,N_6282,N_8234);
and U11343 (N_11343,N_8885,N_8706);
or U11344 (N_11344,N_8882,N_7138);
or U11345 (N_11345,N_7148,N_7217);
nand U11346 (N_11346,N_7463,N_7164);
nor U11347 (N_11347,N_7577,N_7968);
nor U11348 (N_11348,N_6709,N_6916);
and U11349 (N_11349,N_8394,N_8353);
nor U11350 (N_11350,N_8446,N_6417);
or U11351 (N_11351,N_7274,N_7728);
xnor U11352 (N_11352,N_6092,N_8742);
nand U11353 (N_11353,N_8259,N_8703);
and U11354 (N_11354,N_7952,N_7287);
or U11355 (N_11355,N_8572,N_7800);
nor U11356 (N_11356,N_7751,N_7620);
xnor U11357 (N_11357,N_8904,N_7737);
nand U11358 (N_11358,N_7867,N_7933);
nand U11359 (N_11359,N_6499,N_6936);
nand U11360 (N_11360,N_7764,N_6604);
or U11361 (N_11361,N_7484,N_8063);
nor U11362 (N_11362,N_8657,N_7831);
and U11363 (N_11363,N_8919,N_8383);
nand U11364 (N_11364,N_7593,N_7976);
nor U11365 (N_11365,N_6694,N_7494);
or U11366 (N_11366,N_7065,N_8760);
nor U11367 (N_11367,N_6173,N_6920);
nor U11368 (N_11368,N_8727,N_6614);
xor U11369 (N_11369,N_6843,N_8269);
or U11370 (N_11370,N_8873,N_8827);
or U11371 (N_11371,N_8110,N_6277);
nand U11372 (N_11372,N_7673,N_8466);
nor U11373 (N_11373,N_7407,N_6536);
nor U11374 (N_11374,N_6482,N_7894);
nand U11375 (N_11375,N_6707,N_7907);
nand U11376 (N_11376,N_6882,N_6891);
nand U11377 (N_11377,N_8230,N_6997);
nand U11378 (N_11378,N_8093,N_6163);
and U11379 (N_11379,N_6445,N_7149);
and U11380 (N_11380,N_6052,N_6963);
nor U11381 (N_11381,N_7789,N_6511);
nor U11382 (N_11382,N_6403,N_6982);
nor U11383 (N_11383,N_7791,N_8532);
or U11384 (N_11384,N_7663,N_6016);
xor U11385 (N_11385,N_8372,N_8815);
and U11386 (N_11386,N_6723,N_8588);
nor U11387 (N_11387,N_6092,N_7723);
nand U11388 (N_11388,N_8324,N_6302);
and U11389 (N_11389,N_8365,N_7259);
nand U11390 (N_11390,N_8898,N_8596);
or U11391 (N_11391,N_6500,N_6965);
and U11392 (N_11392,N_6798,N_6590);
and U11393 (N_11393,N_7597,N_6227);
nand U11394 (N_11394,N_7967,N_8963);
or U11395 (N_11395,N_8700,N_8745);
nor U11396 (N_11396,N_7769,N_6006);
nand U11397 (N_11397,N_6339,N_6247);
and U11398 (N_11398,N_8593,N_8179);
or U11399 (N_11399,N_7344,N_6976);
or U11400 (N_11400,N_8435,N_8255);
nand U11401 (N_11401,N_6135,N_7392);
and U11402 (N_11402,N_6155,N_6790);
nand U11403 (N_11403,N_7184,N_7467);
nand U11404 (N_11404,N_6484,N_8993);
and U11405 (N_11405,N_6590,N_7243);
nand U11406 (N_11406,N_6456,N_6449);
and U11407 (N_11407,N_7941,N_7178);
nand U11408 (N_11408,N_6308,N_7024);
nand U11409 (N_11409,N_7070,N_6053);
nor U11410 (N_11410,N_8081,N_6730);
and U11411 (N_11411,N_8646,N_7787);
or U11412 (N_11412,N_7953,N_8242);
and U11413 (N_11413,N_8688,N_7236);
or U11414 (N_11414,N_6913,N_6012);
nor U11415 (N_11415,N_8273,N_7207);
and U11416 (N_11416,N_7789,N_7366);
nor U11417 (N_11417,N_8593,N_8076);
nor U11418 (N_11418,N_6627,N_7007);
nor U11419 (N_11419,N_8253,N_6810);
nor U11420 (N_11420,N_7795,N_7907);
and U11421 (N_11421,N_8120,N_7097);
and U11422 (N_11422,N_6872,N_8550);
nand U11423 (N_11423,N_8078,N_8294);
nor U11424 (N_11424,N_7616,N_7211);
and U11425 (N_11425,N_7167,N_7620);
xnor U11426 (N_11426,N_7113,N_8491);
and U11427 (N_11427,N_8542,N_7637);
or U11428 (N_11428,N_7921,N_7355);
nor U11429 (N_11429,N_7985,N_8400);
and U11430 (N_11430,N_7615,N_6907);
nand U11431 (N_11431,N_8249,N_8662);
and U11432 (N_11432,N_8426,N_7630);
and U11433 (N_11433,N_7599,N_6224);
nand U11434 (N_11434,N_8455,N_6181);
or U11435 (N_11435,N_8180,N_7714);
and U11436 (N_11436,N_7233,N_8615);
or U11437 (N_11437,N_8107,N_7257);
nand U11438 (N_11438,N_8865,N_8177);
or U11439 (N_11439,N_6987,N_7746);
nand U11440 (N_11440,N_8285,N_6686);
and U11441 (N_11441,N_7520,N_8325);
or U11442 (N_11442,N_7164,N_8092);
or U11443 (N_11443,N_7659,N_7758);
nor U11444 (N_11444,N_6881,N_7343);
nor U11445 (N_11445,N_6798,N_8433);
and U11446 (N_11446,N_7472,N_6832);
or U11447 (N_11447,N_8253,N_8622);
nand U11448 (N_11448,N_6503,N_6046);
or U11449 (N_11449,N_6059,N_6687);
nor U11450 (N_11450,N_8393,N_8196);
and U11451 (N_11451,N_6922,N_6350);
nand U11452 (N_11452,N_7801,N_7041);
xor U11453 (N_11453,N_8293,N_8738);
and U11454 (N_11454,N_7347,N_6966);
nor U11455 (N_11455,N_7946,N_7082);
nor U11456 (N_11456,N_8198,N_6082);
or U11457 (N_11457,N_8986,N_6584);
nand U11458 (N_11458,N_7321,N_6919);
nand U11459 (N_11459,N_8303,N_7484);
nor U11460 (N_11460,N_6855,N_6131);
or U11461 (N_11461,N_8783,N_6893);
and U11462 (N_11462,N_7978,N_7870);
nor U11463 (N_11463,N_7015,N_8345);
nand U11464 (N_11464,N_8230,N_6376);
xor U11465 (N_11465,N_6578,N_6750);
and U11466 (N_11466,N_8931,N_6175);
nor U11467 (N_11467,N_8777,N_8783);
and U11468 (N_11468,N_7192,N_6203);
and U11469 (N_11469,N_7839,N_7982);
nor U11470 (N_11470,N_7769,N_6521);
and U11471 (N_11471,N_8541,N_6487);
and U11472 (N_11472,N_7903,N_6876);
and U11473 (N_11473,N_7996,N_7981);
nor U11474 (N_11474,N_8634,N_8607);
nand U11475 (N_11475,N_8903,N_8223);
or U11476 (N_11476,N_8844,N_8324);
nor U11477 (N_11477,N_6627,N_7252);
and U11478 (N_11478,N_8981,N_8296);
nand U11479 (N_11479,N_8772,N_7641);
nand U11480 (N_11480,N_7167,N_8522);
or U11481 (N_11481,N_7408,N_7019);
nor U11482 (N_11482,N_7919,N_7867);
nand U11483 (N_11483,N_7366,N_7589);
and U11484 (N_11484,N_6617,N_6210);
nand U11485 (N_11485,N_8550,N_7398);
and U11486 (N_11486,N_7483,N_7053);
or U11487 (N_11487,N_6488,N_8505);
nand U11488 (N_11488,N_6237,N_6686);
and U11489 (N_11489,N_7153,N_6111);
nor U11490 (N_11490,N_7732,N_7764);
nand U11491 (N_11491,N_8009,N_7936);
or U11492 (N_11492,N_6092,N_6558);
or U11493 (N_11493,N_7025,N_6568);
or U11494 (N_11494,N_7346,N_6250);
xor U11495 (N_11495,N_6418,N_7376);
nor U11496 (N_11496,N_8754,N_8545);
nand U11497 (N_11497,N_6879,N_6601);
or U11498 (N_11498,N_8602,N_8910);
and U11499 (N_11499,N_6522,N_6180);
nand U11500 (N_11500,N_7552,N_8476);
nand U11501 (N_11501,N_7421,N_7732);
nor U11502 (N_11502,N_6149,N_6760);
or U11503 (N_11503,N_7064,N_7910);
and U11504 (N_11504,N_8704,N_8510);
nand U11505 (N_11505,N_7719,N_7563);
and U11506 (N_11506,N_8694,N_8065);
xor U11507 (N_11507,N_8812,N_8421);
xor U11508 (N_11508,N_8796,N_8865);
xor U11509 (N_11509,N_6689,N_6037);
nand U11510 (N_11510,N_8694,N_8850);
or U11511 (N_11511,N_7244,N_6892);
and U11512 (N_11512,N_8552,N_8198);
nor U11513 (N_11513,N_7063,N_6764);
or U11514 (N_11514,N_7417,N_7432);
or U11515 (N_11515,N_6159,N_7466);
or U11516 (N_11516,N_6073,N_6411);
and U11517 (N_11517,N_7238,N_8827);
and U11518 (N_11518,N_8632,N_6332);
nand U11519 (N_11519,N_6838,N_6048);
and U11520 (N_11520,N_8594,N_8985);
and U11521 (N_11521,N_7176,N_6384);
nor U11522 (N_11522,N_6924,N_7052);
or U11523 (N_11523,N_7437,N_8141);
or U11524 (N_11524,N_8960,N_7953);
nor U11525 (N_11525,N_6154,N_6782);
nor U11526 (N_11526,N_7961,N_6805);
and U11527 (N_11527,N_7226,N_6327);
and U11528 (N_11528,N_6184,N_6498);
nand U11529 (N_11529,N_7583,N_6742);
and U11530 (N_11530,N_8466,N_7033);
nor U11531 (N_11531,N_7198,N_7378);
and U11532 (N_11532,N_6125,N_7979);
xnor U11533 (N_11533,N_6786,N_6469);
and U11534 (N_11534,N_6281,N_8622);
or U11535 (N_11535,N_7499,N_8665);
and U11536 (N_11536,N_8228,N_8630);
and U11537 (N_11537,N_6950,N_8647);
or U11538 (N_11538,N_7059,N_6339);
nand U11539 (N_11539,N_8739,N_7587);
or U11540 (N_11540,N_8114,N_7636);
nor U11541 (N_11541,N_8066,N_8450);
and U11542 (N_11542,N_7089,N_8961);
nor U11543 (N_11543,N_6473,N_7515);
and U11544 (N_11544,N_6530,N_7571);
nand U11545 (N_11545,N_6344,N_7176);
xor U11546 (N_11546,N_8743,N_8630);
and U11547 (N_11547,N_8590,N_6849);
nor U11548 (N_11548,N_8601,N_6676);
nor U11549 (N_11549,N_6121,N_8066);
and U11550 (N_11550,N_7664,N_8250);
or U11551 (N_11551,N_7563,N_7677);
and U11552 (N_11552,N_7926,N_7613);
nand U11553 (N_11553,N_6245,N_8917);
nor U11554 (N_11554,N_8777,N_6033);
or U11555 (N_11555,N_6952,N_6507);
nor U11556 (N_11556,N_7682,N_7104);
and U11557 (N_11557,N_6340,N_7268);
and U11558 (N_11558,N_8511,N_6135);
or U11559 (N_11559,N_8596,N_6930);
nand U11560 (N_11560,N_6659,N_8289);
and U11561 (N_11561,N_7409,N_6693);
nand U11562 (N_11562,N_6998,N_8907);
nand U11563 (N_11563,N_6331,N_7060);
or U11564 (N_11564,N_7402,N_7230);
and U11565 (N_11565,N_8046,N_8842);
nor U11566 (N_11566,N_6603,N_7283);
nand U11567 (N_11567,N_8186,N_6430);
nand U11568 (N_11568,N_7927,N_7309);
and U11569 (N_11569,N_8703,N_8552);
and U11570 (N_11570,N_6875,N_6751);
nor U11571 (N_11571,N_7644,N_6449);
nor U11572 (N_11572,N_6375,N_8721);
nand U11573 (N_11573,N_8024,N_6722);
nand U11574 (N_11574,N_6702,N_7714);
nand U11575 (N_11575,N_6678,N_8356);
nand U11576 (N_11576,N_7565,N_6896);
or U11577 (N_11577,N_8607,N_8291);
nor U11578 (N_11578,N_6468,N_6624);
nand U11579 (N_11579,N_6131,N_8351);
nand U11580 (N_11580,N_8086,N_6550);
or U11581 (N_11581,N_6976,N_6040);
nor U11582 (N_11582,N_7327,N_6395);
and U11583 (N_11583,N_8741,N_8325);
or U11584 (N_11584,N_8341,N_6620);
or U11585 (N_11585,N_6274,N_6204);
or U11586 (N_11586,N_6949,N_8602);
nand U11587 (N_11587,N_8933,N_7002);
and U11588 (N_11588,N_6599,N_7959);
nor U11589 (N_11589,N_7478,N_8440);
or U11590 (N_11590,N_7499,N_6270);
or U11591 (N_11591,N_6935,N_7755);
xor U11592 (N_11592,N_8519,N_7097);
nand U11593 (N_11593,N_7195,N_7650);
nand U11594 (N_11594,N_7261,N_6841);
nor U11595 (N_11595,N_7198,N_7237);
or U11596 (N_11596,N_8369,N_7994);
or U11597 (N_11597,N_8551,N_7662);
nor U11598 (N_11598,N_8379,N_7549);
or U11599 (N_11599,N_8636,N_6468);
or U11600 (N_11600,N_8819,N_7803);
and U11601 (N_11601,N_6157,N_8904);
nor U11602 (N_11602,N_7022,N_6898);
and U11603 (N_11603,N_8593,N_6989);
nand U11604 (N_11604,N_6320,N_7009);
nand U11605 (N_11605,N_6313,N_8024);
nand U11606 (N_11606,N_8353,N_6376);
nand U11607 (N_11607,N_8551,N_7407);
nand U11608 (N_11608,N_8631,N_8305);
or U11609 (N_11609,N_6073,N_8645);
and U11610 (N_11610,N_8863,N_8205);
nand U11611 (N_11611,N_6487,N_6285);
or U11612 (N_11612,N_8661,N_7759);
and U11613 (N_11613,N_6218,N_8779);
or U11614 (N_11614,N_6207,N_8461);
and U11615 (N_11615,N_7427,N_7395);
nor U11616 (N_11616,N_6494,N_6186);
nand U11617 (N_11617,N_7343,N_7932);
nand U11618 (N_11618,N_6349,N_7415);
and U11619 (N_11619,N_8497,N_7489);
nand U11620 (N_11620,N_7901,N_7933);
and U11621 (N_11621,N_6886,N_8688);
nand U11622 (N_11622,N_6236,N_6594);
nor U11623 (N_11623,N_8172,N_7875);
and U11624 (N_11624,N_7161,N_8680);
or U11625 (N_11625,N_7540,N_8132);
nand U11626 (N_11626,N_7421,N_7832);
nor U11627 (N_11627,N_7579,N_8162);
nor U11628 (N_11628,N_6655,N_6899);
nor U11629 (N_11629,N_8274,N_8169);
and U11630 (N_11630,N_6737,N_6972);
nand U11631 (N_11631,N_8975,N_7542);
and U11632 (N_11632,N_7442,N_6978);
or U11633 (N_11633,N_7232,N_7721);
and U11634 (N_11634,N_6391,N_7911);
nand U11635 (N_11635,N_8760,N_7054);
nand U11636 (N_11636,N_8195,N_7452);
nand U11637 (N_11637,N_6281,N_8105);
nand U11638 (N_11638,N_8331,N_7632);
or U11639 (N_11639,N_8143,N_8923);
nand U11640 (N_11640,N_8052,N_6680);
and U11641 (N_11641,N_7085,N_6348);
nand U11642 (N_11642,N_6791,N_6792);
and U11643 (N_11643,N_7113,N_7061);
nor U11644 (N_11644,N_8858,N_7832);
and U11645 (N_11645,N_8037,N_7244);
or U11646 (N_11646,N_8387,N_6428);
nor U11647 (N_11647,N_7165,N_6504);
xnor U11648 (N_11648,N_6044,N_7446);
and U11649 (N_11649,N_6539,N_7346);
and U11650 (N_11650,N_7144,N_8703);
nor U11651 (N_11651,N_6074,N_6996);
or U11652 (N_11652,N_8633,N_7171);
and U11653 (N_11653,N_6030,N_8549);
nor U11654 (N_11654,N_6014,N_7911);
or U11655 (N_11655,N_8784,N_6518);
nor U11656 (N_11656,N_6151,N_8515);
or U11657 (N_11657,N_6290,N_7495);
or U11658 (N_11658,N_7281,N_8431);
nor U11659 (N_11659,N_6857,N_8272);
nor U11660 (N_11660,N_8742,N_8117);
nor U11661 (N_11661,N_6955,N_8255);
xor U11662 (N_11662,N_6597,N_6236);
and U11663 (N_11663,N_6075,N_7232);
nor U11664 (N_11664,N_7276,N_6288);
nor U11665 (N_11665,N_8732,N_7091);
and U11666 (N_11666,N_6030,N_8015);
xnor U11667 (N_11667,N_7383,N_8238);
or U11668 (N_11668,N_8482,N_6718);
nor U11669 (N_11669,N_7895,N_8936);
nor U11670 (N_11670,N_7907,N_6568);
and U11671 (N_11671,N_7667,N_8030);
nand U11672 (N_11672,N_8852,N_6373);
or U11673 (N_11673,N_6324,N_6820);
and U11674 (N_11674,N_6452,N_6808);
nand U11675 (N_11675,N_7547,N_6842);
nand U11676 (N_11676,N_8330,N_7115);
and U11677 (N_11677,N_6881,N_6197);
and U11678 (N_11678,N_7914,N_7991);
and U11679 (N_11679,N_8024,N_7774);
and U11680 (N_11680,N_7311,N_6922);
nor U11681 (N_11681,N_8337,N_7224);
or U11682 (N_11682,N_6392,N_7005);
or U11683 (N_11683,N_6415,N_7246);
xor U11684 (N_11684,N_6368,N_7260);
nor U11685 (N_11685,N_8270,N_7600);
nor U11686 (N_11686,N_8439,N_7955);
or U11687 (N_11687,N_7771,N_6725);
nor U11688 (N_11688,N_6696,N_8854);
nor U11689 (N_11689,N_6838,N_7915);
or U11690 (N_11690,N_7013,N_6929);
nand U11691 (N_11691,N_6268,N_8498);
or U11692 (N_11692,N_6438,N_6977);
and U11693 (N_11693,N_8608,N_8451);
nor U11694 (N_11694,N_7498,N_8659);
or U11695 (N_11695,N_8466,N_8183);
and U11696 (N_11696,N_6716,N_6047);
or U11697 (N_11697,N_8334,N_7677);
nand U11698 (N_11698,N_6349,N_8199);
nor U11699 (N_11699,N_7163,N_8153);
or U11700 (N_11700,N_8972,N_6484);
and U11701 (N_11701,N_7178,N_7973);
and U11702 (N_11702,N_7612,N_6243);
nand U11703 (N_11703,N_6639,N_6484);
nand U11704 (N_11704,N_6475,N_6351);
nor U11705 (N_11705,N_6639,N_8371);
nor U11706 (N_11706,N_7761,N_8584);
nand U11707 (N_11707,N_6391,N_6971);
nand U11708 (N_11708,N_8700,N_7047);
or U11709 (N_11709,N_6169,N_7166);
and U11710 (N_11710,N_8140,N_8100);
nor U11711 (N_11711,N_6344,N_8816);
or U11712 (N_11712,N_6621,N_8943);
and U11713 (N_11713,N_7662,N_6351);
nand U11714 (N_11714,N_7935,N_6778);
nor U11715 (N_11715,N_8723,N_6319);
and U11716 (N_11716,N_7904,N_6411);
nand U11717 (N_11717,N_8422,N_8639);
or U11718 (N_11718,N_7016,N_8726);
nor U11719 (N_11719,N_7024,N_7474);
nand U11720 (N_11720,N_6828,N_8998);
nand U11721 (N_11721,N_8974,N_8601);
and U11722 (N_11722,N_6296,N_8531);
or U11723 (N_11723,N_6591,N_6919);
nand U11724 (N_11724,N_7347,N_7630);
nand U11725 (N_11725,N_6557,N_6495);
or U11726 (N_11726,N_8748,N_6075);
nand U11727 (N_11727,N_7948,N_7394);
and U11728 (N_11728,N_8587,N_7976);
or U11729 (N_11729,N_6339,N_8403);
nand U11730 (N_11730,N_6024,N_8217);
nor U11731 (N_11731,N_8439,N_6785);
xor U11732 (N_11732,N_8670,N_6392);
nor U11733 (N_11733,N_7845,N_7432);
or U11734 (N_11734,N_6499,N_8669);
or U11735 (N_11735,N_6404,N_6593);
or U11736 (N_11736,N_8467,N_7595);
or U11737 (N_11737,N_7199,N_8261);
or U11738 (N_11738,N_6886,N_6558);
or U11739 (N_11739,N_7832,N_6321);
nand U11740 (N_11740,N_6500,N_6353);
nor U11741 (N_11741,N_8561,N_6530);
or U11742 (N_11742,N_7192,N_6377);
nand U11743 (N_11743,N_7926,N_6510);
nand U11744 (N_11744,N_6626,N_6997);
or U11745 (N_11745,N_8802,N_7268);
nand U11746 (N_11746,N_8522,N_6619);
or U11747 (N_11747,N_7225,N_7064);
and U11748 (N_11748,N_6035,N_8271);
nand U11749 (N_11749,N_7668,N_8902);
and U11750 (N_11750,N_8986,N_6951);
or U11751 (N_11751,N_8042,N_8277);
and U11752 (N_11752,N_6679,N_7231);
nor U11753 (N_11753,N_8125,N_6020);
and U11754 (N_11754,N_8650,N_6491);
nand U11755 (N_11755,N_8944,N_6491);
nand U11756 (N_11756,N_7542,N_8934);
nor U11757 (N_11757,N_7578,N_7503);
nand U11758 (N_11758,N_7787,N_7504);
or U11759 (N_11759,N_7851,N_8265);
xor U11760 (N_11760,N_7163,N_6315);
nand U11761 (N_11761,N_7144,N_6730);
and U11762 (N_11762,N_6778,N_8465);
nor U11763 (N_11763,N_8980,N_8705);
and U11764 (N_11764,N_6457,N_6475);
nand U11765 (N_11765,N_7576,N_8010);
or U11766 (N_11766,N_7446,N_7545);
nand U11767 (N_11767,N_8108,N_7751);
and U11768 (N_11768,N_6369,N_8297);
nor U11769 (N_11769,N_8764,N_6560);
nand U11770 (N_11770,N_6365,N_6526);
nor U11771 (N_11771,N_7352,N_6083);
or U11772 (N_11772,N_7504,N_8122);
nand U11773 (N_11773,N_8177,N_7850);
nand U11774 (N_11774,N_8285,N_7463);
nand U11775 (N_11775,N_7947,N_7366);
or U11776 (N_11776,N_7001,N_8864);
nand U11777 (N_11777,N_8924,N_6813);
or U11778 (N_11778,N_6345,N_7516);
nand U11779 (N_11779,N_8674,N_8693);
or U11780 (N_11780,N_6111,N_8588);
or U11781 (N_11781,N_7638,N_7928);
or U11782 (N_11782,N_8494,N_8408);
or U11783 (N_11783,N_8150,N_6536);
nor U11784 (N_11784,N_8380,N_6243);
nand U11785 (N_11785,N_6435,N_8875);
nand U11786 (N_11786,N_7481,N_7577);
and U11787 (N_11787,N_8850,N_6166);
or U11788 (N_11788,N_7263,N_7173);
nor U11789 (N_11789,N_8029,N_7167);
or U11790 (N_11790,N_7935,N_6668);
or U11791 (N_11791,N_8168,N_6866);
nor U11792 (N_11792,N_7106,N_6557);
nand U11793 (N_11793,N_8764,N_7501);
or U11794 (N_11794,N_7833,N_7594);
nor U11795 (N_11795,N_8953,N_8001);
or U11796 (N_11796,N_6397,N_6714);
nand U11797 (N_11797,N_8305,N_6553);
nor U11798 (N_11798,N_6774,N_8507);
or U11799 (N_11799,N_8662,N_8372);
or U11800 (N_11800,N_7527,N_6418);
and U11801 (N_11801,N_6987,N_7568);
and U11802 (N_11802,N_6176,N_6216);
or U11803 (N_11803,N_7746,N_7576);
nor U11804 (N_11804,N_8810,N_8206);
nor U11805 (N_11805,N_6094,N_8596);
or U11806 (N_11806,N_8575,N_6575);
and U11807 (N_11807,N_8739,N_7294);
nand U11808 (N_11808,N_7646,N_7605);
or U11809 (N_11809,N_7643,N_8199);
nand U11810 (N_11810,N_8800,N_8414);
nor U11811 (N_11811,N_8584,N_6816);
or U11812 (N_11812,N_8530,N_8187);
nor U11813 (N_11813,N_7005,N_6647);
nor U11814 (N_11814,N_6236,N_7165);
xor U11815 (N_11815,N_7330,N_8971);
nand U11816 (N_11816,N_7221,N_8172);
and U11817 (N_11817,N_7445,N_7838);
nor U11818 (N_11818,N_7511,N_7746);
or U11819 (N_11819,N_7240,N_7998);
xnor U11820 (N_11820,N_6169,N_7855);
and U11821 (N_11821,N_8011,N_8677);
nor U11822 (N_11822,N_6474,N_6936);
and U11823 (N_11823,N_8645,N_8231);
nand U11824 (N_11824,N_6755,N_6935);
and U11825 (N_11825,N_8751,N_8486);
or U11826 (N_11826,N_8352,N_6504);
nor U11827 (N_11827,N_7413,N_8281);
nand U11828 (N_11828,N_7813,N_7256);
or U11829 (N_11829,N_7749,N_7664);
and U11830 (N_11830,N_8503,N_8329);
nor U11831 (N_11831,N_7261,N_8873);
or U11832 (N_11832,N_6189,N_6164);
and U11833 (N_11833,N_8317,N_8362);
nor U11834 (N_11834,N_8741,N_7674);
nor U11835 (N_11835,N_8674,N_7827);
and U11836 (N_11836,N_6461,N_7063);
nand U11837 (N_11837,N_7890,N_8044);
or U11838 (N_11838,N_6349,N_6465);
and U11839 (N_11839,N_8101,N_8782);
or U11840 (N_11840,N_6644,N_8045);
nor U11841 (N_11841,N_7364,N_7776);
or U11842 (N_11842,N_6643,N_8343);
nand U11843 (N_11843,N_6646,N_6398);
or U11844 (N_11844,N_8966,N_7682);
nand U11845 (N_11845,N_8769,N_7959);
and U11846 (N_11846,N_7122,N_7218);
and U11847 (N_11847,N_6153,N_7260);
and U11848 (N_11848,N_7974,N_6737);
or U11849 (N_11849,N_6191,N_6359);
nor U11850 (N_11850,N_8646,N_8764);
nand U11851 (N_11851,N_7656,N_6852);
xnor U11852 (N_11852,N_6805,N_7351);
nor U11853 (N_11853,N_6604,N_6197);
nand U11854 (N_11854,N_7601,N_8321);
and U11855 (N_11855,N_8500,N_8224);
and U11856 (N_11856,N_8554,N_7795);
or U11857 (N_11857,N_7463,N_8989);
or U11858 (N_11858,N_6377,N_8399);
nor U11859 (N_11859,N_7353,N_6508);
xor U11860 (N_11860,N_8018,N_8250);
and U11861 (N_11861,N_6337,N_7177);
and U11862 (N_11862,N_8991,N_7584);
or U11863 (N_11863,N_8649,N_7364);
nor U11864 (N_11864,N_6193,N_6085);
nor U11865 (N_11865,N_7399,N_7044);
nand U11866 (N_11866,N_8410,N_8967);
nand U11867 (N_11867,N_7833,N_8736);
nor U11868 (N_11868,N_7970,N_8147);
or U11869 (N_11869,N_8218,N_6648);
and U11870 (N_11870,N_8478,N_7616);
or U11871 (N_11871,N_7058,N_8333);
nand U11872 (N_11872,N_6822,N_7524);
and U11873 (N_11873,N_7471,N_6134);
or U11874 (N_11874,N_6275,N_7281);
and U11875 (N_11875,N_7154,N_6524);
nand U11876 (N_11876,N_7058,N_7690);
nor U11877 (N_11877,N_6093,N_7247);
or U11878 (N_11878,N_7808,N_7008);
nand U11879 (N_11879,N_8029,N_7301);
and U11880 (N_11880,N_7358,N_6828);
nand U11881 (N_11881,N_6648,N_6639);
or U11882 (N_11882,N_8989,N_7976);
nand U11883 (N_11883,N_6430,N_6415);
xor U11884 (N_11884,N_7507,N_6750);
xnor U11885 (N_11885,N_7026,N_8238);
or U11886 (N_11886,N_8202,N_7755);
or U11887 (N_11887,N_8944,N_6822);
nand U11888 (N_11888,N_7487,N_7945);
nand U11889 (N_11889,N_7926,N_7883);
nor U11890 (N_11890,N_7910,N_6784);
nor U11891 (N_11891,N_7346,N_7434);
nand U11892 (N_11892,N_7360,N_6838);
or U11893 (N_11893,N_7291,N_7480);
nor U11894 (N_11894,N_8734,N_7719);
nand U11895 (N_11895,N_8661,N_6553);
and U11896 (N_11896,N_6426,N_6040);
nor U11897 (N_11897,N_6963,N_6773);
nor U11898 (N_11898,N_6937,N_7281);
or U11899 (N_11899,N_7930,N_8669);
or U11900 (N_11900,N_6416,N_7012);
or U11901 (N_11901,N_8167,N_6039);
nand U11902 (N_11902,N_7225,N_7767);
or U11903 (N_11903,N_8935,N_8270);
nor U11904 (N_11904,N_8576,N_8120);
nand U11905 (N_11905,N_7803,N_6194);
nor U11906 (N_11906,N_8558,N_6351);
nand U11907 (N_11907,N_7039,N_6047);
nand U11908 (N_11908,N_8456,N_8303);
nor U11909 (N_11909,N_8754,N_8830);
and U11910 (N_11910,N_8284,N_6866);
and U11911 (N_11911,N_8089,N_7659);
nor U11912 (N_11912,N_7824,N_6684);
nor U11913 (N_11913,N_6264,N_8580);
nand U11914 (N_11914,N_6957,N_6798);
and U11915 (N_11915,N_6275,N_6460);
nand U11916 (N_11916,N_6478,N_6005);
and U11917 (N_11917,N_8759,N_7838);
or U11918 (N_11918,N_8883,N_8263);
nand U11919 (N_11919,N_8544,N_7617);
or U11920 (N_11920,N_8389,N_8295);
nor U11921 (N_11921,N_6974,N_7128);
or U11922 (N_11922,N_8471,N_8309);
nand U11923 (N_11923,N_7174,N_6860);
or U11924 (N_11924,N_6881,N_7339);
nor U11925 (N_11925,N_6315,N_6650);
nor U11926 (N_11926,N_7125,N_8795);
and U11927 (N_11927,N_7526,N_6142);
and U11928 (N_11928,N_8033,N_6123);
and U11929 (N_11929,N_7036,N_7157);
or U11930 (N_11930,N_6684,N_8087);
nand U11931 (N_11931,N_6577,N_6622);
and U11932 (N_11932,N_8989,N_8009);
nor U11933 (N_11933,N_7839,N_6823);
or U11934 (N_11934,N_6637,N_7434);
and U11935 (N_11935,N_6317,N_7109);
nand U11936 (N_11936,N_8164,N_6472);
or U11937 (N_11937,N_8138,N_8536);
or U11938 (N_11938,N_8808,N_8866);
or U11939 (N_11939,N_7194,N_8048);
and U11940 (N_11940,N_6045,N_8330);
or U11941 (N_11941,N_8250,N_7761);
and U11942 (N_11942,N_6947,N_8128);
nor U11943 (N_11943,N_8967,N_8136);
and U11944 (N_11944,N_7493,N_7925);
and U11945 (N_11945,N_6765,N_7418);
nand U11946 (N_11946,N_8812,N_8431);
or U11947 (N_11947,N_8039,N_6850);
and U11948 (N_11948,N_7012,N_8802);
nand U11949 (N_11949,N_7609,N_7666);
nor U11950 (N_11950,N_7592,N_6063);
and U11951 (N_11951,N_8845,N_7817);
and U11952 (N_11952,N_8032,N_8976);
and U11953 (N_11953,N_6021,N_6714);
nor U11954 (N_11954,N_7965,N_6420);
or U11955 (N_11955,N_7007,N_6695);
or U11956 (N_11956,N_7184,N_6345);
nor U11957 (N_11957,N_6387,N_7226);
or U11958 (N_11958,N_7379,N_8471);
or U11959 (N_11959,N_8958,N_6012);
nor U11960 (N_11960,N_8055,N_8879);
or U11961 (N_11961,N_8539,N_6928);
xnor U11962 (N_11962,N_7756,N_8691);
xnor U11963 (N_11963,N_6968,N_8227);
nand U11964 (N_11964,N_7201,N_6868);
or U11965 (N_11965,N_6739,N_8155);
nor U11966 (N_11966,N_6302,N_6368);
nand U11967 (N_11967,N_6819,N_7860);
or U11968 (N_11968,N_8674,N_6812);
or U11969 (N_11969,N_6076,N_7309);
nor U11970 (N_11970,N_8161,N_7164);
nor U11971 (N_11971,N_7159,N_8925);
nand U11972 (N_11972,N_6231,N_7502);
nand U11973 (N_11973,N_7368,N_6686);
nand U11974 (N_11974,N_6314,N_7293);
and U11975 (N_11975,N_8685,N_7304);
xor U11976 (N_11976,N_7754,N_6766);
and U11977 (N_11977,N_8800,N_8490);
nand U11978 (N_11978,N_8210,N_6231);
nand U11979 (N_11979,N_6032,N_7683);
and U11980 (N_11980,N_7517,N_8669);
nand U11981 (N_11981,N_7749,N_8502);
nand U11982 (N_11982,N_7191,N_7834);
or U11983 (N_11983,N_8135,N_8016);
or U11984 (N_11984,N_7647,N_6515);
or U11985 (N_11985,N_6183,N_7792);
and U11986 (N_11986,N_7103,N_7099);
or U11987 (N_11987,N_6292,N_6605);
nor U11988 (N_11988,N_8416,N_6320);
nand U11989 (N_11989,N_7238,N_8823);
or U11990 (N_11990,N_7334,N_7283);
nor U11991 (N_11991,N_6204,N_7562);
nand U11992 (N_11992,N_8149,N_6648);
or U11993 (N_11993,N_6692,N_6827);
or U11994 (N_11994,N_8882,N_7470);
or U11995 (N_11995,N_8487,N_8933);
nor U11996 (N_11996,N_7868,N_6321);
or U11997 (N_11997,N_8718,N_8028);
or U11998 (N_11998,N_6741,N_6780);
or U11999 (N_11999,N_8043,N_6391);
nor U12000 (N_12000,N_11302,N_10887);
or U12001 (N_12001,N_10476,N_10403);
or U12002 (N_12002,N_11985,N_10024);
nor U12003 (N_12003,N_11466,N_9881);
nor U12004 (N_12004,N_10845,N_9554);
nand U12005 (N_12005,N_10123,N_11654);
nor U12006 (N_12006,N_11024,N_10780);
nor U12007 (N_12007,N_10092,N_11841);
nand U12008 (N_12008,N_10440,N_10379);
nor U12009 (N_12009,N_9491,N_11130);
or U12010 (N_12010,N_11432,N_11366);
or U12011 (N_12011,N_11154,N_11825);
nand U12012 (N_12012,N_10049,N_9242);
and U12013 (N_12013,N_10304,N_11604);
nand U12014 (N_12014,N_9176,N_10270);
nand U12015 (N_12015,N_10474,N_9490);
and U12016 (N_12016,N_10982,N_11289);
or U12017 (N_12017,N_10583,N_9227);
nor U12018 (N_12018,N_9671,N_11078);
or U12019 (N_12019,N_10328,N_10171);
and U12020 (N_12020,N_10636,N_10807);
and U12021 (N_12021,N_9178,N_9469);
and U12022 (N_12022,N_10165,N_11542);
and U12023 (N_12023,N_9087,N_11279);
nand U12024 (N_12024,N_11545,N_10541);
nor U12025 (N_12025,N_11874,N_9878);
and U12026 (N_12026,N_11226,N_10813);
nand U12027 (N_12027,N_11193,N_10779);
or U12028 (N_12028,N_9263,N_10785);
xor U12029 (N_12029,N_9349,N_11535);
nand U12030 (N_12030,N_9136,N_10215);
and U12031 (N_12031,N_11408,N_10009);
nor U12032 (N_12032,N_10930,N_11810);
and U12033 (N_12033,N_10968,N_10265);
xor U12034 (N_12034,N_11107,N_10053);
and U12035 (N_12035,N_9326,N_10726);
and U12036 (N_12036,N_11555,N_9317);
and U12037 (N_12037,N_11666,N_11603);
nor U12038 (N_12038,N_11591,N_11904);
nand U12039 (N_12039,N_10701,N_10922);
nor U12040 (N_12040,N_9782,N_11830);
or U12041 (N_12041,N_9185,N_11506);
or U12042 (N_12042,N_11702,N_11381);
nand U12043 (N_12043,N_10828,N_9094);
and U12044 (N_12044,N_11971,N_11230);
nor U12045 (N_12045,N_10467,N_11079);
or U12046 (N_12046,N_9809,N_11897);
nor U12047 (N_12047,N_11657,N_10788);
nand U12048 (N_12048,N_10586,N_9007);
and U12049 (N_12049,N_10759,N_9436);
nor U12050 (N_12050,N_10926,N_9851);
or U12051 (N_12051,N_10499,N_10030);
and U12052 (N_12052,N_9420,N_10959);
and U12053 (N_12053,N_10515,N_11636);
and U12054 (N_12054,N_11334,N_9464);
or U12055 (N_12055,N_9064,N_11724);
nor U12056 (N_12056,N_9157,N_10255);
and U12057 (N_12057,N_10717,N_9238);
and U12058 (N_12058,N_9223,N_9067);
nand U12059 (N_12059,N_9365,N_10498);
and U12060 (N_12060,N_9456,N_10649);
nand U12061 (N_12061,N_9999,N_9408);
and U12062 (N_12062,N_10212,N_9510);
nand U12063 (N_12063,N_9724,N_11561);
and U12064 (N_12064,N_11885,N_10682);
nor U12065 (N_12065,N_9002,N_10455);
or U12066 (N_12066,N_9149,N_9864);
nand U12067 (N_12067,N_10249,N_10589);
nand U12068 (N_12068,N_9247,N_10272);
and U12069 (N_12069,N_10851,N_10456);
nand U12070 (N_12070,N_9976,N_9827);
nand U12071 (N_12071,N_9333,N_11426);
nand U12072 (N_12072,N_10156,N_9519);
and U12073 (N_12073,N_11609,N_11246);
and U12074 (N_12074,N_10316,N_11779);
and U12075 (N_12075,N_9353,N_11800);
nor U12076 (N_12076,N_9310,N_10015);
nor U12077 (N_12077,N_9741,N_11084);
nor U12078 (N_12078,N_10007,N_11301);
and U12079 (N_12079,N_10524,N_10776);
or U12080 (N_12080,N_11490,N_11801);
nand U12081 (N_12081,N_10039,N_9980);
and U12082 (N_12082,N_11339,N_11350);
nor U12083 (N_12083,N_11071,N_9346);
or U12084 (N_12084,N_9729,N_10923);
nand U12085 (N_12085,N_11846,N_9857);
and U12086 (N_12086,N_9587,N_10219);
xnor U12087 (N_12087,N_11626,N_11397);
or U12088 (N_12088,N_11546,N_9425);
nor U12089 (N_12089,N_11291,N_9563);
nor U12090 (N_12090,N_10734,N_9774);
and U12091 (N_12091,N_11069,N_9192);
nand U12092 (N_12092,N_9177,N_9240);
nor U12093 (N_12093,N_11455,N_9319);
nor U12094 (N_12094,N_11930,N_11832);
nor U12095 (N_12095,N_11136,N_9793);
nor U12096 (N_12096,N_9288,N_10060);
nand U12097 (N_12097,N_9191,N_11621);
and U12098 (N_12098,N_11762,N_10050);
and U12099 (N_12099,N_11596,N_9700);
or U12100 (N_12100,N_9831,N_10837);
nand U12101 (N_12101,N_10337,N_11096);
nand U12102 (N_12102,N_11676,N_9059);
nor U12103 (N_12103,N_10364,N_11976);
or U12104 (N_12104,N_9115,N_10979);
nand U12105 (N_12105,N_9367,N_11638);
or U12106 (N_12106,N_11593,N_9642);
nand U12107 (N_12107,N_11489,N_9706);
and U12108 (N_12108,N_9139,N_9093);
xnor U12109 (N_12109,N_10825,N_10234);
and U12110 (N_12110,N_9614,N_11693);
xor U12111 (N_12111,N_11217,N_10948);
or U12112 (N_12112,N_11739,N_11091);
or U12113 (N_12113,N_10262,N_9400);
and U12114 (N_12114,N_10975,N_10812);
and U12115 (N_12115,N_10471,N_11652);
or U12116 (N_12116,N_9988,N_11590);
or U12117 (N_12117,N_10327,N_10067);
nand U12118 (N_12118,N_9052,N_11367);
and U12119 (N_12119,N_9434,N_9968);
or U12120 (N_12120,N_10016,N_9508);
or U12121 (N_12121,N_10590,N_10210);
nand U12122 (N_12122,N_11095,N_11415);
nand U12123 (N_12123,N_11627,N_9388);
nor U12124 (N_12124,N_9625,N_10973);
nand U12125 (N_12125,N_9032,N_9561);
or U12126 (N_12126,N_11139,N_11320);
or U12127 (N_12127,N_9668,N_11077);
and U12128 (N_12128,N_11290,N_9651);
or U12129 (N_12129,N_11059,N_11420);
nand U12130 (N_12130,N_9682,N_10027);
or U12131 (N_12131,N_10076,N_11674);
or U12132 (N_12132,N_10281,N_10634);
xor U12133 (N_12133,N_11733,N_10872);
nand U12134 (N_12134,N_9171,N_10928);
or U12135 (N_12135,N_10205,N_10106);
or U12136 (N_12136,N_11135,N_11966);
nor U12137 (N_12137,N_11922,N_11991);
nor U12138 (N_12138,N_11713,N_11766);
nor U12139 (N_12139,N_9600,N_10939);
and U12140 (N_12140,N_9132,N_9633);
nand U12141 (N_12141,N_10412,N_10965);
or U12142 (N_12142,N_10461,N_9475);
and U12143 (N_12143,N_9483,N_11808);
nand U12144 (N_12144,N_11053,N_9452);
nand U12145 (N_12145,N_9041,N_9663);
or U12146 (N_12146,N_11871,N_10633);
and U12147 (N_12147,N_9040,N_10670);
or U12148 (N_12148,N_9787,N_10905);
nor U12149 (N_12149,N_10302,N_11065);
nand U12150 (N_12150,N_10142,N_9536);
nor U12151 (N_12151,N_10104,N_11896);
and U12152 (N_12152,N_10534,N_10560);
nand U12153 (N_12153,N_10850,N_11026);
nor U12154 (N_12154,N_11647,N_9296);
or U12155 (N_12155,N_9858,N_9039);
and U12156 (N_12156,N_10018,N_11806);
nor U12157 (N_12157,N_11181,N_9842);
nand U12158 (N_12158,N_10147,N_11559);
and U12159 (N_12159,N_10111,N_11039);
nand U12160 (N_12160,N_9197,N_9818);
or U12161 (N_12161,N_11696,N_11496);
or U12162 (N_12162,N_11834,N_10258);
nand U12163 (N_12163,N_9450,N_9797);
nor U12164 (N_12164,N_10619,N_9429);
nor U12165 (N_12165,N_10115,N_10324);
nand U12166 (N_12166,N_9082,N_11949);
and U12167 (N_12167,N_11278,N_10429);
and U12168 (N_12168,N_9538,N_10859);
or U12169 (N_12169,N_10036,N_9414);
nand U12170 (N_12170,N_11359,N_9233);
and U12171 (N_12171,N_11034,N_10709);
xor U12172 (N_12172,N_11964,N_11893);
and U12173 (N_12173,N_11736,N_11630);
nand U12174 (N_12174,N_10688,N_9591);
or U12175 (N_12175,N_11168,N_10692);
and U12176 (N_12176,N_10635,N_10750);
and U12177 (N_12177,N_11171,N_11681);
nor U12178 (N_12178,N_9424,N_11369);
nand U12179 (N_12179,N_9664,N_11788);
or U12180 (N_12180,N_11441,N_10382);
or U12181 (N_12181,N_11510,N_9439);
and U12182 (N_12182,N_9199,N_11500);
or U12183 (N_12183,N_9919,N_9397);
nor U12184 (N_12184,N_10436,N_11057);
nor U12185 (N_12185,N_10735,N_10108);
or U12186 (N_12186,N_10164,N_11140);
nor U12187 (N_12187,N_9658,N_9730);
or U12188 (N_12188,N_11121,N_9876);
nor U12189 (N_12189,N_11649,N_10553);
and U12190 (N_12190,N_9243,N_9846);
and U12191 (N_12191,N_10808,N_10190);
and U12192 (N_12192,N_9896,N_10862);
and U12193 (N_12193,N_10416,N_9764);
and U12194 (N_12194,N_11514,N_9042);
and U12195 (N_12195,N_9552,N_11507);
and U12196 (N_12196,N_9843,N_11850);
nand U12197 (N_12197,N_11575,N_10090);
and U12198 (N_12198,N_10962,N_9448);
nor U12199 (N_12199,N_11642,N_10334);
or U12200 (N_12200,N_9293,N_9043);
and U12201 (N_12201,N_10604,N_9295);
or U12202 (N_12202,N_11137,N_11195);
or U12203 (N_12203,N_11730,N_11128);
nand U12204 (N_12204,N_10293,N_9503);
nand U12205 (N_12205,N_11973,N_11436);
xor U12206 (N_12206,N_9862,N_11665);
or U12207 (N_12207,N_11016,N_10453);
nand U12208 (N_12208,N_9799,N_11267);
or U12209 (N_12209,N_9286,N_10149);
nor U12210 (N_12210,N_9328,N_11111);
nand U12211 (N_12211,N_10847,N_10620);
nand U12212 (N_12212,N_10626,N_10796);
and U12213 (N_12213,N_9211,N_9337);
nor U12214 (N_12214,N_9596,N_9673);
and U12215 (N_12215,N_10197,N_9410);
nand U12216 (N_12216,N_10241,N_10805);
and U12217 (N_12217,N_10662,N_11775);
xnor U12218 (N_12218,N_9249,N_9909);
nand U12219 (N_12219,N_10511,N_10013);
or U12220 (N_12220,N_11858,N_11308);
and U12221 (N_12221,N_10001,N_9321);
and U12222 (N_12222,N_10211,N_9075);
nand U12223 (N_12223,N_10180,N_10724);
nand U12224 (N_12224,N_10623,N_9099);
nor U12225 (N_12225,N_9119,N_11684);
and U12226 (N_12226,N_9237,N_10786);
nand U12227 (N_12227,N_11223,N_9543);
and U12228 (N_12228,N_9704,N_11635);
or U12229 (N_12229,N_11158,N_10587);
nor U12230 (N_12230,N_11812,N_9735);
or U12231 (N_12231,N_10607,N_10512);
nand U12232 (N_12232,N_10591,N_9792);
nor U12233 (N_12233,N_9060,N_9234);
and U12234 (N_12234,N_10366,N_10519);
or U12235 (N_12235,N_11761,N_9783);
and U12236 (N_12236,N_10562,N_10774);
nand U12237 (N_12237,N_10213,N_9879);
nor U12238 (N_12238,N_10625,N_10117);
or U12239 (N_12239,N_10244,N_11502);
nor U12240 (N_12240,N_9021,N_10310);
and U12241 (N_12241,N_10765,N_9357);
nor U12242 (N_12242,N_9144,N_11229);
nor U12243 (N_12243,N_10680,N_10003);
nor U12244 (N_12244,N_11325,N_11117);
xnor U12245 (N_12245,N_11047,N_9212);
nand U12246 (N_12246,N_10487,N_11050);
and U12247 (N_12247,N_9161,N_10656);
and U12248 (N_12248,N_10072,N_10818);
nor U12249 (N_12249,N_9235,N_11857);
or U12250 (N_12250,N_9551,N_9101);
or U12251 (N_12251,N_9079,N_9727);
and U12252 (N_12252,N_10609,N_9455);
and U12253 (N_12253,N_9355,N_11934);
and U12254 (N_12254,N_9811,N_11605);
and U12255 (N_12255,N_10983,N_11040);
nand U12256 (N_12256,N_11074,N_11873);
nor U12257 (N_12257,N_9418,N_10853);
and U12258 (N_12258,N_10086,N_9051);
or U12259 (N_12259,N_10323,N_11892);
nand U12260 (N_12260,N_10497,N_11745);
or U12261 (N_12261,N_11321,N_10863);
and U12262 (N_12262,N_9252,N_11254);
or U12263 (N_12263,N_11183,N_11062);
or U12264 (N_12264,N_10354,N_9720);
nand U12265 (N_12265,N_10658,N_9123);
xor U12266 (N_12266,N_11145,N_11357);
or U12267 (N_12267,N_9748,N_10953);
nand U12268 (N_12268,N_9710,N_10313);
and U12269 (N_12269,N_9125,N_10010);
and U12270 (N_12270,N_10058,N_10134);
or U12271 (N_12271,N_10345,N_10322);
or U12272 (N_12272,N_9517,N_9865);
or U12273 (N_12273,N_11423,N_10955);
and U12274 (N_12274,N_11282,N_9269);
and U12275 (N_12275,N_9494,N_10362);
and U12276 (N_12276,N_9686,N_11109);
nor U12277 (N_12277,N_11103,N_10761);
and U12278 (N_12278,N_11394,N_9555);
or U12279 (N_12279,N_9189,N_9696);
xnor U12280 (N_12280,N_10643,N_9849);
nand U12281 (N_12281,N_10209,N_10787);
and U12282 (N_12282,N_11299,N_10909);
and U12283 (N_12283,N_9761,N_11917);
nor U12284 (N_12284,N_11554,N_11743);
or U12285 (N_12285,N_9246,N_10326);
and U12286 (N_12286,N_10738,N_9081);
nor U12287 (N_12287,N_10889,N_9913);
or U12288 (N_12288,N_11807,N_9360);
or U12289 (N_12289,N_11097,N_10120);
or U12290 (N_12290,N_11169,N_9732);
nor U12291 (N_12291,N_9670,N_10972);
nand U12292 (N_12292,N_10064,N_10729);
or U12293 (N_12293,N_9932,N_11669);
nand U12294 (N_12294,N_10296,N_10093);
nor U12295 (N_12295,N_11756,N_11188);
and U12296 (N_12296,N_10603,N_10199);
nand U12297 (N_12297,N_10198,N_9050);
or U12298 (N_12298,N_11721,N_9880);
nand U12299 (N_12299,N_11710,N_10061);
nor U12300 (N_12300,N_11623,N_9151);
nor U12301 (N_12301,N_10230,N_9411);
nor U12302 (N_12302,N_9169,N_9325);
and U12303 (N_12303,N_9259,N_10528);
nand U12304 (N_12304,N_11755,N_9655);
nor U12305 (N_12305,N_10996,N_9105);
and U12306 (N_12306,N_11965,N_11588);
or U12307 (N_12307,N_10668,N_10087);
or U12308 (N_12308,N_9541,N_11319);
nand U12309 (N_12309,N_9894,N_9055);
or U12310 (N_12310,N_9726,N_11821);
and U12311 (N_12311,N_11232,N_10391);
nand U12312 (N_12312,N_9091,N_9767);
and U12313 (N_12313,N_10394,N_10756);
or U12314 (N_12314,N_10183,N_11335);
nand U12315 (N_12315,N_10742,N_9405);
or U12316 (N_12316,N_9701,N_11550);
and U12317 (N_12317,N_11951,N_11203);
nand U12318 (N_12318,N_9672,N_9564);
nand U12319 (N_12319,N_11045,N_9037);
and U12320 (N_12320,N_11618,N_9559);
and U12321 (N_12321,N_11388,N_10950);
nor U12322 (N_12322,N_9111,N_9058);
nor U12323 (N_12323,N_10914,N_10752);
and U12324 (N_12324,N_9389,N_10593);
nand U12325 (N_12325,N_9725,N_11296);
nand U12326 (N_12326,N_11351,N_9683);
nor U12327 (N_12327,N_9332,N_9933);
nor U12328 (N_12328,N_9721,N_11374);
or U12329 (N_12329,N_9952,N_10458);
nand U12330 (N_12330,N_10426,N_9497);
or U12331 (N_12331,N_10159,N_11478);
nor U12332 (N_12332,N_11481,N_9970);
and U12333 (N_12333,N_11586,N_11304);
nand U12334 (N_12334,N_10358,N_10194);
xor U12335 (N_12335,N_11539,N_9861);
nand U12336 (N_12336,N_9165,N_10409);
nand U12337 (N_12337,N_11895,N_10538);
nor U12338 (N_12338,N_11716,N_11119);
nand U12339 (N_12339,N_11541,N_11480);
nand U12340 (N_12340,N_10848,N_10493);
or U12341 (N_12341,N_11014,N_9048);
nand U12342 (N_12342,N_9283,N_9402);
nand U12343 (N_12343,N_10208,N_9219);
nor U12344 (N_12344,N_10946,N_9751);
or U12345 (N_12345,N_9206,N_10744);
nor U12346 (N_12346,N_10686,N_9649);
or U12347 (N_12347,N_9231,N_9184);
nor U12348 (N_12348,N_10886,N_11134);
nand U12349 (N_12349,N_11337,N_10338);
or U12350 (N_12350,N_9030,N_9141);
and U12351 (N_12351,N_10827,N_11698);
nor U12352 (N_12352,N_11753,N_9344);
nor U12353 (N_12353,N_11386,N_10174);
nand U12354 (N_12354,N_9172,N_11405);
or U12355 (N_12355,N_9431,N_11600);
nor U12356 (N_12356,N_10306,N_11701);
or U12357 (N_12357,N_11943,N_9553);
nand U12358 (N_12358,N_9709,N_9468);
and U12359 (N_12359,N_10011,N_10000);
nand U12360 (N_12360,N_11720,N_9722);
and U12361 (N_12361,N_9816,N_10931);
nand U12362 (N_12362,N_9585,N_9903);
and U12363 (N_12363,N_10916,N_9602);
and U12364 (N_12364,N_11164,N_9540);
or U12365 (N_12365,N_9681,N_10713);
or U12366 (N_12366,N_10703,N_10871);
and U12367 (N_12367,N_9945,N_10333);
or U12368 (N_12368,N_10842,N_9122);
and U12369 (N_12369,N_10114,N_9794);
nor U12370 (N_12370,N_10413,N_11905);
and U12371 (N_12371,N_9631,N_11439);
and U12372 (N_12372,N_9925,N_9356);
nor U12373 (N_12373,N_11607,N_9624);
nand U12374 (N_12374,N_10999,N_9447);
and U12375 (N_12375,N_9035,N_9549);
or U12376 (N_12376,N_9100,N_10986);
and U12377 (N_12377,N_9329,N_9940);
or U12378 (N_12378,N_9640,N_10112);
nor U12379 (N_12379,N_10820,N_11629);
nor U12380 (N_12380,N_10763,N_9962);
nand U12381 (N_12381,N_9392,N_11574);
nand U12382 (N_12382,N_10268,N_9373);
nor U12383 (N_12383,N_10582,N_11678);
or U12384 (N_12384,N_11473,N_11360);
nand U12385 (N_12385,N_10672,N_11688);
or U12386 (N_12386,N_10980,N_11066);
nand U12387 (N_12387,N_11963,N_9084);
nand U12388 (N_12388,N_11073,N_10263);
nand U12389 (N_12389,N_10824,N_10732);
and U12390 (N_12390,N_10094,N_9590);
nor U12391 (N_12391,N_9530,N_9106);
nor U12392 (N_12392,N_10925,N_10532);
or U12393 (N_12393,N_11692,N_11151);
or U12394 (N_12394,N_10279,N_9085);
nand U12395 (N_12395,N_9487,N_11872);
or U12396 (N_12396,N_9505,N_9959);
nor U12397 (N_12397,N_9440,N_9979);
xor U12398 (N_12398,N_9711,N_10089);
nand U12399 (N_12399,N_9377,N_9776);
nor U12400 (N_12400,N_9824,N_10745);
or U12401 (N_12401,N_10631,N_10563);
or U12402 (N_12402,N_11003,N_11576);
or U12403 (N_12403,N_11814,N_10554);
and U12404 (N_12404,N_11737,N_11634);
nor U12405 (N_12405,N_11968,N_11332);
nor U12406 (N_12406,N_11712,N_9376);
nand U12407 (N_12407,N_10764,N_9905);
nand U12408 (N_12408,N_11553,N_9921);
or U12409 (N_12409,N_9303,N_11780);
or U12410 (N_12410,N_11578,N_9391);
or U12411 (N_12411,N_11012,N_9331);
or U12412 (N_12412,N_9918,N_11854);
nand U12413 (N_12413,N_9719,N_9595);
nand U12414 (N_12414,N_10690,N_9302);
nand U12415 (N_12415,N_11373,N_11061);
xor U12416 (N_12416,N_9364,N_10835);
nand U12417 (N_12417,N_11551,N_9599);
or U12418 (N_12418,N_9795,N_9513);
and U12419 (N_12419,N_9800,N_11025);
and U12420 (N_12420,N_11659,N_9415);
nor U12421 (N_12421,N_10287,N_9347);
nor U12422 (N_12422,N_10126,N_10144);
nand U12423 (N_12423,N_10119,N_9545);
or U12424 (N_12424,N_11064,N_9790);
and U12425 (N_12425,N_11051,N_9944);
nand U12426 (N_12426,N_10103,N_11768);
or U12427 (N_12427,N_9802,N_9619);
and U12428 (N_12428,N_9598,N_10526);
and U12429 (N_12429,N_11148,N_11903);
or U12430 (N_12430,N_11384,N_10008);
nand U12431 (N_12431,N_10261,N_9078);
or U12432 (N_12432,N_9788,N_10970);
nor U12433 (N_12433,N_10856,N_9594);
nand U12434 (N_12434,N_10739,N_10439);
nor U12435 (N_12435,N_9244,N_10466);
nor U12436 (N_12436,N_9068,N_11820);
or U12437 (N_12437,N_10880,N_11058);
or U12438 (N_12438,N_11132,N_11915);
or U12439 (N_12439,N_9969,N_11249);
nor U12440 (N_12440,N_10430,N_10961);
or U12441 (N_12441,N_9926,N_10196);
nand U12442 (N_12442,N_11942,N_9224);
nor U12443 (N_12443,N_9386,N_9928);
nand U12444 (N_12444,N_10908,N_10195);
nand U12445 (N_12445,N_11880,N_9550);
and U12446 (N_12446,N_11902,N_11243);
nor U12447 (N_12447,N_11453,N_9383);
and U12448 (N_12448,N_9027,N_10794);
nor U12449 (N_12449,N_11992,N_10665);
and U12450 (N_12450,N_10711,N_10852);
nand U12451 (N_12451,N_10290,N_9837);
and U12452 (N_12452,N_11310,N_9167);
nor U12453 (N_12453,N_10666,N_9703);
nor U12454 (N_12454,N_9758,N_9897);
or U12455 (N_12455,N_10629,N_9983);
nand U12456 (N_12456,N_9380,N_11271);
or U12457 (N_12457,N_11222,N_9305);
or U12458 (N_12458,N_11115,N_10383);
and U12459 (N_12459,N_9187,N_9635);
nand U12460 (N_12460,N_9180,N_11567);
and U12461 (N_12461,N_9736,N_10879);
nand U12462 (N_12462,N_11485,N_10184);
and U12463 (N_12463,N_11189,N_9278);
and U12464 (N_12464,N_9766,N_10570);
nor U12465 (N_12465,N_11498,N_10846);
or U12466 (N_12466,N_11201,N_11185);
or U12467 (N_12467,N_9656,N_11843);
or U12468 (N_12468,N_10700,N_9971);
nand U12469 (N_12469,N_9422,N_10091);
nor U12470 (N_12470,N_9716,N_9112);
and U12471 (N_12471,N_11338,N_9140);
nand U12472 (N_12472,N_10271,N_11105);
nand U12473 (N_12473,N_9524,N_9715);
or U12474 (N_12474,N_11430,N_11999);
nor U12475 (N_12475,N_9128,N_11606);
and U12476 (N_12476,N_11512,N_10288);
and U12477 (N_12477,N_9110,N_11356);
or U12478 (N_12478,N_10661,N_9648);
nor U12479 (N_12479,N_10292,N_11361);
nor U12480 (N_12480,N_10695,N_9282);
nor U12481 (N_12481,N_9798,N_11826);
and U12482 (N_12482,N_10274,N_10598);
nand U12483 (N_12483,N_10378,N_9941);
nor U12484 (N_12484,N_11706,N_9019);
or U12485 (N_12485,N_11831,N_9998);
nand U12486 (N_12486,N_11216,N_10055);
nand U12487 (N_12487,N_11163,N_10841);
or U12488 (N_12488,N_10934,N_10051);
nor U12489 (N_12489,N_9982,N_10130);
nand U12490 (N_12490,N_9092,N_11364);
and U12491 (N_12491,N_10694,N_11285);
xor U12492 (N_12492,N_9583,N_11354);
or U12493 (N_12493,N_11110,N_9385);
and U12494 (N_12494,N_11752,N_11632);
nand U12495 (N_12495,N_10992,N_9834);
xnor U12496 (N_12496,N_11876,N_9867);
or U12497 (N_12497,N_11689,N_11429);
nand U12498 (N_12498,N_9182,N_9805);
nor U12499 (N_12499,N_11910,N_9276);
nor U12500 (N_12500,N_11068,N_11286);
and U12501 (N_12501,N_9129,N_10136);
and U12502 (N_12502,N_11474,N_9923);
xor U12503 (N_12503,N_11732,N_11637);
or U12504 (N_12504,N_9753,N_9613);
and U12505 (N_12505,N_9571,N_9739);
nor U12506 (N_12506,N_10350,N_11495);
nor U12507 (N_12507,N_11521,N_9166);
and U12508 (N_12508,N_9154,N_11728);
and U12509 (N_12509,N_11523,N_11002);
or U12510 (N_12510,N_9647,N_11522);
nand U12511 (N_12511,N_9204,N_11044);
nand U12512 (N_12512,N_11075,N_11443);
nand U12513 (N_12513,N_11100,N_11708);
nand U12514 (N_12514,N_10760,N_11925);
or U12515 (N_12515,N_9046,N_9742);
and U12516 (N_12516,N_11067,N_9713);
nor U12517 (N_12517,N_11771,N_10936);
or U12518 (N_12518,N_9898,N_11936);
or U12519 (N_12519,N_11888,N_11571);
nor U12520 (N_12520,N_10247,N_11021);
nor U12521 (N_12521,N_11776,N_10746);
nand U12522 (N_12522,N_9348,N_11234);
nand U12523 (N_12523,N_10691,N_11153);
or U12524 (N_12524,N_11220,N_11414);
or U12525 (N_12525,N_9338,N_10465);
nand U12526 (N_12526,N_9936,N_11152);
and U12527 (N_12527,N_9131,N_11362);
nand U12528 (N_12528,N_11957,N_11298);
or U12529 (N_12529,N_9279,N_9714);
or U12530 (N_12530,N_10510,N_11327);
nand U12531 (N_12531,N_9230,N_9636);
nor U12532 (N_12532,N_11984,N_9038);
nor U12533 (N_12533,N_10958,N_10683);
or U12534 (N_12534,N_11157,N_9899);
or U12535 (N_12535,N_9004,N_11518);
nor U12536 (N_12536,N_9768,N_11644);
nand U12537 (N_12537,N_11572,N_9572);
nor U12538 (N_12538,N_9835,N_9931);
nor U12539 (N_12539,N_11425,N_11528);
or U12540 (N_12540,N_10138,N_10239);
or U12541 (N_12541,N_11317,N_10594);
and U12542 (N_12542,N_10141,N_9107);
nor U12543 (N_12543,N_9089,N_9016);
nor U12544 (N_12544,N_11931,N_10755);
nand U12545 (N_12545,N_11479,N_11734);
nor U12546 (N_12546,N_9698,N_11087);
and U12547 (N_12547,N_9752,N_9891);
nor U12548 (N_12548,N_9914,N_9993);
and U12549 (N_12549,N_11941,N_11564);
and U12550 (N_12550,N_11239,N_10877);
and U12551 (N_12551,N_10462,N_10243);
xor U12552 (N_12552,N_10778,N_11190);
or U12553 (N_12553,N_9076,N_10564);
nor U12554 (N_12554,N_9274,N_10971);
and U12555 (N_12555,N_9675,N_11513);
and U12556 (N_12556,N_9229,N_10821);
and U12557 (N_12557,N_9744,N_9074);
nor U12558 (N_12558,N_10900,N_11424);
nor U12559 (N_12559,N_11348,N_9884);
nand U12560 (N_12560,N_11511,N_11900);
xnor U12561 (N_12561,N_11054,N_11923);
and U12562 (N_12562,N_10605,N_11783);
and U12563 (N_12563,N_10343,N_10608);
nor U12564 (N_12564,N_10838,N_9026);
nor U12565 (N_12565,N_9509,N_11856);
nand U12566 (N_12566,N_11594,N_11944);
nor U12567 (N_12567,N_9342,N_10963);
and U12568 (N_12568,N_9967,N_9202);
and U12569 (N_12569,N_10645,N_11093);
nor U12570 (N_12570,N_10494,N_9255);
and U12571 (N_12571,N_9641,N_9963);
or U12572 (N_12572,N_10784,N_9275);
nor U12573 (N_12573,N_9523,N_9868);
nand U12574 (N_12574,N_9841,N_10911);
and U12575 (N_12575,N_10771,N_9576);
and U12576 (N_12576,N_9785,N_11663);
xor U12577 (N_12577,N_11655,N_10482);
nand U12578 (N_12578,N_10109,N_11417);
nand U12579 (N_12579,N_9372,N_9063);
or U12580 (N_12580,N_10082,N_11009);
nand U12581 (N_12581,N_9208,N_9950);
and U12582 (N_12582,N_9615,N_9034);
nor U12583 (N_12583,N_11838,N_9750);
or U12584 (N_12584,N_10351,N_11661);
or U12585 (N_12585,N_10715,N_11845);
and U12586 (N_12586,N_10079,N_11465);
and U12587 (N_12587,N_10017,N_11123);
nor U12588 (N_12588,N_10721,N_9070);
and U12589 (N_12589,N_10177,N_9446);
and U12590 (N_12590,N_10956,N_10810);
or U12591 (N_12591,N_10101,N_10179);
or U12592 (N_12592,N_9791,N_9628);
or U12593 (N_12593,N_10985,N_9022);
or U12594 (N_12594,N_10521,N_11182);
nand U12595 (N_12595,N_10995,N_10415);
nand U12596 (N_12596,N_10699,N_9465);
nor U12597 (N_12597,N_9173,N_9872);
nor U12598 (N_12598,N_11894,N_11407);
nor U12599 (N_12599,N_10684,N_9956);
or U12600 (N_12600,N_11258,N_9678);
nor U12601 (N_12601,N_11272,N_11172);
nand U12602 (N_12602,N_10988,N_10723);
nand U12603 (N_12603,N_11884,N_10193);
nand U12604 (N_12604,N_9906,N_11878);
xnor U12605 (N_12605,N_9267,N_9975);
or U12606 (N_12606,N_9280,N_10990);
nor U12607 (N_12607,N_9512,N_9580);
nand U12608 (N_12608,N_11263,N_11198);
nand U12609 (N_12609,N_10469,N_10371);
and U12610 (N_12610,N_11456,N_9930);
or U12611 (N_12611,N_10253,N_11330);
nand U12612 (N_12612,N_11294,N_10537);
nor U12613 (N_12613,N_10031,N_10187);
or U12614 (N_12614,N_9147,N_9953);
and U12615 (N_12615,N_10168,N_11619);
nand U12616 (N_12616,N_11851,N_11251);
and U12617 (N_12617,N_11370,N_11328);
nand U12618 (N_12618,N_10506,N_9152);
or U12619 (N_12619,N_11410,N_10902);
nand U12620 (N_12620,N_9401,N_10496);
nor U12621 (N_12621,N_11210,N_11958);
and U12622 (N_12622,N_9755,N_9973);
nor U12623 (N_12623,N_10543,N_11581);
nand U12624 (N_12624,N_9239,N_10434);
or U12625 (N_12625,N_11517,N_10414);
nor U12626 (N_12626,N_10606,N_9480);
nor U12627 (N_12627,N_10137,N_11314);
and U12628 (N_12628,N_9216,N_11244);
nand U12629 (N_12629,N_11191,N_10459);
and U12630 (N_12630,N_10282,N_9622);
or U12631 (N_12631,N_10289,N_10552);
and U12632 (N_12632,N_10696,N_10269);
nor U12633 (N_12633,N_10984,N_11184);
and U12634 (N_12634,N_10200,N_10733);
nand U12635 (N_12635,N_11906,N_9061);
or U12636 (N_12636,N_11471,N_10275);
and U12637 (N_12637,N_11990,N_10819);
nor U12638 (N_12638,N_10783,N_11001);
nand U12639 (N_12639,N_10470,N_11980);
or U12640 (N_12640,N_9003,N_10023);
nor U12641 (N_12641,N_11494,N_11611);
or U12642 (N_12642,N_11703,N_9574);
or U12643 (N_12643,N_9784,N_10952);
or U12644 (N_12644,N_11916,N_10397);
nor U12645 (N_12645,N_9499,N_10580);
nor U12646 (N_12646,N_10478,N_10876);
nand U12647 (N_12647,N_11387,N_10758);
and U12648 (N_12648,N_10616,N_10475);
nand U12649 (N_12649,N_11613,N_11960);
nand U12650 (N_12650,N_10107,N_9674);
nand U12651 (N_12651,N_10319,N_9604);
and U12652 (N_12652,N_11744,N_9297);
nor U12653 (N_12653,N_10918,N_11565);
and U12654 (N_12654,N_9057,N_10381);
or U12655 (N_12655,N_10720,N_9853);
nand U12656 (N_12656,N_9882,N_9010);
xor U12657 (N_12657,N_11238,N_11919);
nand U12658 (N_12658,N_11467,N_9379);
nand U12659 (N_12659,N_10642,N_10280);
nand U12660 (N_12660,N_9033,N_9334);
nor U12661 (N_12661,N_11794,N_9660);
nor U12662 (N_12662,N_11178,N_11225);
nand U12663 (N_12663,N_10675,N_11179);
nand U12664 (N_12664,N_11406,N_9972);
nand U12665 (N_12665,N_11597,N_9426);
nor U12666 (N_12666,N_9320,N_9265);
or U12667 (N_12667,N_10559,N_11809);
nor U12668 (N_12668,N_11462,N_9775);
and U12669 (N_12669,N_10618,N_11847);
or U12670 (N_12670,N_10155,N_11566);
and U12671 (N_12671,N_10443,N_10062);
nor U12672 (N_12672,N_9939,N_11815);
nand U12673 (N_12673,N_9665,N_9220);
and U12674 (N_12674,N_10096,N_9168);
nor U12675 (N_12675,N_9533,N_9522);
or U12676 (N_12676,N_11470,N_11767);
nand U12677 (N_12677,N_10539,N_10227);
nand U12678 (N_12678,N_10647,N_9174);
nand U12679 (N_12679,N_10312,N_9213);
or U12680 (N_12680,N_9053,N_11667);
xor U12681 (N_12681,N_10592,N_11608);
and U12682 (N_12682,N_10654,N_11264);
or U12683 (N_12683,N_9667,N_10201);
and U12684 (N_12684,N_10793,N_11060);
nor U12685 (N_12685,N_9838,N_10595);
and U12686 (N_12686,N_10172,N_9096);
or U12687 (N_12687,N_9121,N_10585);
or U12688 (N_12688,N_9746,N_11377);
and U12689 (N_12689,N_11840,N_9623);
nor U12690 (N_12690,N_11601,N_11037);
or U12691 (N_12691,N_11503,N_10192);
nor U12692 (N_12692,N_9877,N_10259);
nand U12693 (N_12693,N_10944,N_11970);
nand U12694 (N_12694,N_10341,N_11624);
and U12695 (N_12695,N_9828,N_9771);
nor U12696 (N_12696,N_11648,N_9814);
nor U12697 (N_12697,N_11088,N_10782);
or U12698 (N_12698,N_10097,N_10920);
xnor U12699 (N_12699,N_10899,N_11640);
or U12700 (N_12700,N_9659,N_11962);
nor U12701 (N_12701,N_10385,N_9284);
and U12702 (N_12702,N_10099,N_9527);
nand U12703 (N_12703,N_9343,N_10402);
nor U12704 (N_12704,N_10420,N_11993);
and U12705 (N_12705,N_11316,N_10428);
and U12706 (N_12706,N_11937,N_10078);
nand U12707 (N_12707,N_11221,N_11700);
and U12708 (N_12708,N_10573,N_10869);
or U12709 (N_12709,N_11560,N_10588);
and U12710 (N_12710,N_9852,N_9693);
and U12711 (N_12711,N_9608,N_10809);
nand U12712 (N_12712,N_11804,N_9694);
and U12713 (N_12713,N_9777,N_11340);
nor U12714 (N_12714,N_9277,N_9108);
nand U12715 (N_12715,N_9695,N_9335);
and U12716 (N_12716,N_10442,N_10545);
nor U12717 (N_12717,N_11256,N_11927);
xor U12718 (N_12718,N_10260,N_10311);
nand U12719 (N_12719,N_11785,N_10754);
and U12720 (N_12720,N_10359,N_10189);
or U12721 (N_12721,N_9458,N_9306);
nand U12722 (N_12722,N_11803,N_11438);
nor U12723 (N_12723,N_10480,N_9985);
and U12724 (N_12724,N_11538,N_11409);
nand U12725 (N_12725,N_11844,N_9646);
nor U12726 (N_12726,N_10372,N_9813);
and U12727 (N_12727,N_10457,N_10286);
or U12728 (N_12728,N_9848,N_9560);
nand U12729 (N_12729,N_10004,N_10678);
and U12730 (N_12730,N_9427,N_10309);
or U12731 (N_12731,N_10175,N_10714);
or U12732 (N_12732,N_9323,N_11089);
nor U12733 (N_12733,N_10207,N_9581);
nor U12734 (N_12734,N_11475,N_10389);
and U12735 (N_12735,N_11488,N_10568);
nor U12736 (N_12736,N_9226,N_10681);
nand U12737 (N_12737,N_10997,N_11177);
and U12738 (N_12738,N_11376,N_10535);
or U12739 (N_12739,N_11219,N_9996);
nor U12740 (N_12740,N_9575,N_9856);
nand U12741 (N_12741,N_9413,N_9194);
and U12742 (N_12742,N_9546,N_9496);
nand U12743 (N_12743,N_10329,N_11995);
or U12744 (N_12744,N_11757,N_11516);
or U12745 (N_12745,N_9833,N_10374);
nor U12746 (N_12746,N_10468,N_10811);
nand U12747 (N_12747,N_9218,N_9680);
and U12748 (N_12748,N_11940,N_10802);
and U12749 (N_12749,N_11928,N_11952);
and U12750 (N_12750,N_9817,N_11445);
nor U12751 (N_12751,N_11950,N_11092);
nand U12752 (N_12752,N_9479,N_11391);
xnor U12753 (N_12753,N_9609,N_9368);
nor U12754 (N_12754,N_10332,N_11750);
or U12755 (N_12755,N_11908,N_11162);
and U12756 (N_12756,N_9937,N_9991);
or U12757 (N_12757,N_9029,N_10574);
and U12758 (N_12758,N_9083,N_10597);
nand U12759 (N_12759,N_11281,N_10960);
nand U12760 (N_12760,N_10858,N_9699);
nand U12761 (N_12761,N_10894,N_9907);
and U12762 (N_12762,N_9478,N_9045);
or U12763 (N_12763,N_11176,N_9117);
nor U12764 (N_12764,N_9954,N_10669);
nand U12765 (N_12765,N_10883,N_9304);
or U12766 (N_12766,N_9984,N_10427);
or U12767 (N_12767,N_11419,N_10297);
or U12768 (N_12768,N_11180,N_11789);
or U12769 (N_12769,N_11907,N_11782);
nor U12770 (N_12770,N_10702,N_11380);
and U12771 (N_12771,N_9485,N_10225);
nor U12772 (N_12772,N_9734,N_10581);
nand U12773 (N_12773,N_10166,N_11690);
or U12774 (N_12774,N_10612,N_10867);
nor U12775 (N_12775,N_11175,N_10229);
nor U12776 (N_12776,N_10806,N_9620);
or U12777 (N_12777,N_10798,N_9459);
or U12778 (N_12778,N_9528,N_10705);
and U12779 (N_12779,N_11280,N_10488);
and U12780 (N_12780,N_10408,N_11786);
and U12781 (N_12781,N_11988,N_9214);
nor U12782 (N_12782,N_9592,N_10865);
and U12783 (N_12783,N_10181,N_11717);
nand U12784 (N_12784,N_10473,N_9637);
nor U12785 (N_12785,N_11707,N_9474);
nand U12786 (N_12786,N_9428,N_9175);
nor U12787 (N_12787,N_11454,N_10300);
or U12788 (N_12788,N_11749,N_11197);
and U12789 (N_12789,N_10638,N_11795);
and U12790 (N_12790,N_11277,N_11534);
nor U12791 (N_12791,N_9514,N_11746);
xnor U12792 (N_12792,N_11011,N_10977);
and U12793 (N_12793,N_11598,N_10548);
nor U12794 (N_12794,N_9924,N_11187);
nand U12795 (N_12795,N_9395,N_10508);
nand U12796 (N_12796,N_11450,N_10348);
nor U12797 (N_12797,N_10770,N_9066);
and U12798 (N_12798,N_9516,N_10648);
and U12799 (N_12799,N_11760,N_11483);
and U12800 (N_12800,N_9020,N_10447);
and U12801 (N_12801,N_11979,N_10509);
nand U12802 (N_12802,N_9363,N_10489);
nor U12803 (N_12803,N_10864,N_9915);
nand U12804 (N_12804,N_11482,N_11956);
and U12805 (N_12805,N_11633,N_10291);
or U12806 (N_12806,N_11469,N_11961);
nand U12807 (N_12807,N_10317,N_9691);
nand U12808 (N_12808,N_11570,N_10674);
nand U12809 (N_12809,N_9137,N_9535);
nor U12810 (N_12810,N_11358,N_10932);
nand U12811 (N_12811,N_10516,N_10047);
or U12812 (N_12812,N_9869,N_11822);
or U12813 (N_12813,N_11199,N_11250);
or U12814 (N_12814,N_10401,N_10221);
nor U12815 (N_12815,N_9626,N_11240);
and U12816 (N_12816,N_11112,N_9215);
and U12817 (N_12817,N_9217,N_11104);
or U12818 (N_12818,N_10527,N_10712);
nor U12819 (N_12819,N_11435,N_9158);
and U12820 (N_12820,N_9438,N_11227);
or U12821 (N_12821,N_11612,N_10601);
nand U12822 (N_12822,N_9362,N_10320);
and U12823 (N_12823,N_10070,N_9525);
nand U12824 (N_12824,N_11126,N_11035);
or U12825 (N_12825,N_10223,N_9947);
nor U12826 (N_12826,N_10125,N_10831);
or U12827 (N_12827,N_9526,N_10020);
nor U12828 (N_12828,N_10002,N_9605);
or U12829 (N_12829,N_10940,N_11173);
nor U12830 (N_12830,N_9500,N_11063);
or U12831 (N_12831,N_9256,N_9629);
and U12832 (N_12832,N_9557,N_11270);
and U12833 (N_12833,N_11019,N_9717);
nand U12834 (N_12834,N_10520,N_10762);
xnor U12835 (N_12835,N_10085,N_10736);
or U12836 (N_12836,N_10578,N_9018);
nor U12837 (N_12837,N_10081,N_11543);
and U12838 (N_12838,N_9486,N_10657);
or U12839 (N_12839,N_10384,N_10561);
and U12840 (N_12840,N_10941,N_11138);
nor U12841 (N_12841,N_9883,N_9382);
nor U12842 (N_12842,N_9374,N_9120);
nand U12843 (N_12843,N_9179,N_11805);
nand U12844 (N_12844,N_11769,N_9989);
xnor U12845 (N_12845,N_11673,N_9203);
and U12846 (N_12846,N_10264,N_10373);
nand U12847 (N_12847,N_9113,N_11998);
nor U12848 (N_12848,N_9810,N_9300);
nand U12849 (N_12849,N_10365,N_11793);
nand U12850 (N_12850,N_10822,N_9781);
nor U12851 (N_12851,N_10555,N_11141);
nor U12852 (N_12852,N_9650,N_11579);
nand U12853 (N_12853,N_11042,N_10550);
nand U12854 (N_12854,N_11631,N_9393);
or U12855 (N_12855,N_11532,N_9762);
and U12856 (N_12856,N_9506,N_11877);
or U12857 (N_12857,N_10045,N_10006);
nor U12858 (N_12858,N_11368,N_11664);
nand U12859 (N_12859,N_11186,N_9484);
and U12860 (N_12860,N_11781,N_11932);
nand U12861 (N_12861,N_9690,N_9350);
nor U12862 (N_12862,N_9258,N_11276);
xor U12863 (N_12863,N_11056,N_9584);
or U12864 (N_12864,N_10222,N_10355);
or U12865 (N_12865,N_9025,N_10907);
nor U12866 (N_12866,N_11122,N_9718);
nor U12867 (N_12867,N_11926,N_11192);
or U12868 (N_12868,N_11646,N_11326);
nor U12869 (N_12869,N_10182,N_9416);
nand U12870 (N_12870,N_10048,N_10012);
nor U12871 (N_12871,N_11085,N_11323);
nand U12872 (N_12872,N_10989,N_10419);
and U12873 (N_12873,N_11048,N_10056);
nand U12874 (N_12874,N_11741,N_11444);
and U12875 (N_12875,N_10152,N_9481);
xnor U12876 (N_12876,N_10370,N_11914);
nand U12877 (N_12877,N_10284,N_9253);
nand U12878 (N_12878,N_10501,N_10530);
nor U12879 (N_12879,N_11383,N_9911);
and U12880 (N_12880,N_11848,N_9241);
and U12881 (N_12881,N_10285,N_11924);
and U12882 (N_12882,N_9627,N_11797);
or U12883 (N_12883,N_9073,N_11853);
nor U12884 (N_12884,N_10220,N_11525);
nand U12885 (N_12885,N_10611,N_10392);
xnor U12886 (N_12886,N_10237,N_11836);
nand U12887 (N_12887,N_9815,N_10360);
and U12888 (N_12888,N_10650,N_11165);
nand U12889 (N_12889,N_10445,N_9160);
nor U12890 (N_12890,N_9001,N_10518);
nor U12891 (N_12891,N_11155,N_9688);
nand U12892 (N_12892,N_11747,N_10652);
and U12893 (N_12893,N_9812,N_11569);
nor U12894 (N_12894,N_11010,N_10624);
xor U12895 (N_12895,N_11824,N_10202);
and U12896 (N_12896,N_9088,N_10919);
and U12897 (N_12897,N_11341,N_11889);
nand U12898 (N_12898,N_9754,N_11283);
nand U12899 (N_12899,N_9015,N_10162);
nor U12900 (N_12900,N_9193,N_9893);
or U12901 (N_12901,N_11860,N_10929);
and U12902 (N_12902,N_9747,N_9000);
nand U12903 (N_12903,N_11890,N_10356);
nor U12904 (N_12904,N_10565,N_11530);
nor U12905 (N_12905,N_11587,N_11891);
nand U12906 (N_12906,N_11651,N_9049);
nand U12907 (N_12907,N_9568,N_11656);
nand U12908 (N_12908,N_9130,N_9181);
and U12909 (N_12909,N_10128,N_11120);
and U12910 (N_12910,N_10873,N_9712);
or U12911 (N_12911,N_9423,N_9902);
nand U12912 (N_12912,N_11727,N_10844);
or U12913 (N_12913,N_9723,N_11113);
and U12914 (N_12914,N_10627,N_10301);
nand U12915 (N_12915,N_10866,N_10836);
or U12916 (N_12916,N_11463,N_10792);
nor U12917 (N_12917,N_9822,N_11997);
nor U12918 (N_12918,N_10186,N_10882);
or U12919 (N_12919,N_10113,N_11540);
or U12920 (N_12920,N_9270,N_10307);
nand U12921 (N_12921,N_10969,N_9210);
or U12922 (N_12922,N_9014,N_10231);
or U12923 (N_12923,N_9470,N_10749);
and U12924 (N_12924,N_11018,N_9011);
and U12925 (N_12925,N_10395,N_10933);
nand U12926 (N_12926,N_9531,N_10472);
and U12927 (N_12927,N_11491,N_9261);
nand U12928 (N_12928,N_10676,N_9955);
nand U12929 (N_12929,N_11504,N_9299);
xor U12930 (N_12930,N_10135,N_11437);
nand U12931 (N_12931,N_10122,N_10935);
or U12932 (N_12932,N_9489,N_11602);
nor U12933 (N_12933,N_10095,N_11156);
or U12934 (N_12934,N_11967,N_9582);
or U12935 (N_12935,N_10444,N_9432);
nand U12936 (N_12936,N_9786,N_10450);
and U12937 (N_12937,N_11643,N_11870);
nor U12938 (N_12938,N_9757,N_11265);
or U12939 (N_12939,N_10127,N_9807);
nor U12940 (N_12940,N_9669,N_10800);
nand U12941 (N_12941,N_10238,N_10340);
or U12942 (N_12942,N_11813,N_11449);
xnor U12943 (N_12943,N_9830,N_10423);
or U12944 (N_12944,N_9573,N_9821);
and U12945 (N_12945,N_9779,N_9430);
or U12946 (N_12946,N_10600,N_10737);
nand U12947 (N_12947,N_11452,N_11382);
and U12948 (N_12948,N_10170,N_9960);
or U12949 (N_12949,N_10875,N_11777);
nand U12950 (N_12950,N_9534,N_10025);
nor U12951 (N_12951,N_9188,N_9978);
nor U12952 (N_12952,N_10704,N_9632);
and U12953 (N_12953,N_10173,N_11729);
and U12954 (N_12954,N_11899,N_11763);
and U12955 (N_12955,N_9638,N_11072);
nor U12956 (N_12956,N_10267,N_11865);
or U12957 (N_12957,N_9272,N_10677);
or U12958 (N_12958,N_10449,N_9077);
or U12959 (N_12959,N_10719,N_11714);
or U12960 (N_12960,N_10240,N_11212);
and U12961 (N_12961,N_11983,N_11378);
or U12962 (N_12962,N_10651,N_11705);
or U12963 (N_12963,N_11792,N_9806);
xor U12964 (N_12964,N_9301,N_9345);
nand U12965 (N_12965,N_11231,N_11022);
and U12966 (N_12966,N_9065,N_10567);
nand U12967 (N_12967,N_10206,N_11043);
nand U12968 (N_12968,N_11167,N_11509);
nor U12969 (N_12969,N_9012,N_11670);
and U12970 (N_12970,N_9341,N_10751);
or U12971 (N_12971,N_9558,N_10363);
or U12972 (N_12972,N_11006,N_10769);
xor U12973 (N_12973,N_11174,N_11959);
nor U12974 (N_12974,N_11431,N_9209);
and U12975 (N_12975,N_10966,N_9886);
and U12976 (N_12976,N_10131,N_11675);
and U12977 (N_12977,N_11616,N_10906);
nand U12978 (N_12978,N_9248,N_9062);
nor U12979 (N_12979,N_11017,N_10660);
and U12980 (N_12980,N_10949,N_9162);
and U12981 (N_12981,N_10305,N_9044);
and U12982 (N_12982,N_11599,N_11790);
or U12983 (N_12983,N_10245,N_10927);
and U12984 (N_12984,N_10242,N_9387);
or U12985 (N_12985,N_11641,N_9645);
nor U12986 (N_12986,N_9607,N_11955);
and U12987 (N_12987,N_11515,N_10331);
nand U12988 (N_12988,N_9653,N_11082);
and U12989 (N_12989,N_9287,N_9887);
or U12990 (N_12990,N_11548,N_10422);
and U12991 (N_12991,N_9566,N_9443);
and U12992 (N_12992,N_10613,N_10276);
nor U12993 (N_12993,N_10707,N_11204);
or U12994 (N_12994,N_10250,N_10857);
or U12995 (N_12995,N_10357,N_9163);
and U12996 (N_12996,N_9705,N_11086);
nand U12997 (N_12997,N_11448,N_10140);
xor U12998 (N_12998,N_9763,N_10217);
and U12999 (N_12999,N_10728,N_11839);
or U13000 (N_13000,N_11206,N_9361);
or U13001 (N_13001,N_10448,N_9290);
nand U13002 (N_13002,N_10797,N_11013);
nor U13003 (N_13003,N_10052,N_11842);
nand U13004 (N_13004,N_10431,N_11774);
and U13005 (N_13005,N_9611,N_9330);
and U13006 (N_13006,N_9482,N_10855);
or U13007 (N_13007,N_10602,N_10361);
and U13008 (N_13008,N_9981,N_9770);
nor U13009 (N_13009,N_10901,N_9028);
and U13010 (N_13010,N_10967,N_9854);
or U13011 (N_13011,N_10663,N_10065);
nor U13012 (N_13012,N_10098,N_10502);
or U13013 (N_13013,N_10100,N_10224);
or U13014 (N_13014,N_10041,N_10435);
nor U13015 (N_13015,N_9997,N_11484);
or U13016 (N_13016,N_11295,N_10892);
nand U13017 (N_13017,N_9801,N_10158);
or U13018 (N_13018,N_10369,N_9309);
nor U13019 (N_13019,N_11875,N_9769);
nand U13020 (N_13020,N_10557,N_9222);
and U13021 (N_13021,N_9072,N_11911);
nand U13022 (N_13022,N_9850,N_11033);
and U13023 (N_13023,N_9127,N_9461);
nand U13024 (N_13024,N_9697,N_11080);
nand U13025 (N_13025,N_9866,N_11614);
nand U13026 (N_13026,N_9228,N_10766);
or U13027 (N_13027,N_10832,N_11722);
and U13028 (N_13028,N_10981,N_9987);
nor U13029 (N_13029,N_9460,N_9765);
or U13030 (N_13030,N_9495,N_10233);
or U13031 (N_13031,N_11459,N_11259);
or U13032 (N_13032,N_9148,N_9644);
or U13033 (N_13033,N_11422,N_11284);
and U13034 (N_13034,N_10904,N_10938);
and U13035 (N_13035,N_10697,N_10547);
nor U13036 (N_13036,N_9895,N_11379);
or U13037 (N_13037,N_11237,N_9069);
or U13038 (N_13038,N_11401,N_10947);
nor U13039 (N_13039,N_10777,N_9307);
nor U13040 (N_13040,N_10226,N_9031);
or U13041 (N_13041,N_10839,N_10640);
nand U13042 (N_13042,N_10367,N_9257);
or U13043 (N_13043,N_11837,N_10298);
or U13044 (N_13044,N_10740,N_9404);
and U13045 (N_13045,N_10163,N_10029);
xor U13046 (N_13046,N_11166,N_10028);
nand U13047 (N_13047,N_10005,N_9054);
or U13048 (N_13048,N_9603,N_9616);
or U13049 (N_13049,N_9929,N_11715);
or U13050 (N_13050,N_10503,N_10437);
and U13051 (N_13051,N_11413,N_9707);
nor U13052 (N_13052,N_10464,N_11557);
and U13053 (N_13053,N_10057,N_9371);
nor U13054 (N_13054,N_11389,N_9961);
nand U13055 (N_13055,N_11697,N_9863);
or U13056 (N_13056,N_11861,N_10485);
nor U13057 (N_13057,N_9621,N_10504);
nor U13058 (N_13058,N_11938,N_9466);
and U13059 (N_13059,N_10477,N_11544);
or U13060 (N_13060,N_9116,N_10804);
and U13061 (N_13061,N_10743,N_10256);
nor U13062 (N_13062,N_10671,N_10576);
nand U13063 (N_13063,N_10531,N_10884);
nand U13064 (N_13064,N_11653,N_10891);
or U13065 (N_13065,N_11660,N_9740);
nor U13066 (N_13066,N_10257,N_10251);
nor U13067 (N_13067,N_11773,N_9164);
xnor U13068 (N_13068,N_11823,N_9569);
and U13069 (N_13069,N_11709,N_10167);
xor U13070 (N_13070,N_11248,N_9832);
xnor U13071 (N_13071,N_9201,N_10716);
and U13072 (N_13072,N_11331,N_11798);
xnor U13073 (N_13073,N_9407,N_9351);
nand U13074 (N_13074,N_11260,N_11041);
nor U13075 (N_13075,N_11921,N_11954);
or U13076 (N_13076,N_9892,N_9366);
or U13077 (N_13077,N_11562,N_9654);
and U13078 (N_13078,N_10407,N_10577);
nand U13079 (N_13079,N_11020,N_10725);
and U13080 (N_13080,N_10718,N_9298);
and U13081 (N_13081,N_11537,N_9225);
nand U13082 (N_13082,N_11828,N_11996);
nand U13083 (N_13083,N_10110,N_11679);
xor U13084 (N_13084,N_11778,N_9266);
nor U13085 (N_13085,N_11353,N_11253);
or U13086 (N_13086,N_11255,N_10843);
and U13087 (N_13087,N_9804,N_11772);
nor U13088 (N_13088,N_9417,N_9118);
nand U13089 (N_13089,N_9917,N_9186);
or U13090 (N_13090,N_11305,N_11529);
nand U13091 (N_13091,N_9521,N_10342);
or U13092 (N_13092,N_10551,N_11242);
nand U13093 (N_13093,N_11143,N_11519);
nor U13094 (N_13094,N_10438,N_10888);
or U13095 (N_13095,N_9403,N_10621);
xor U13096 (N_13096,N_11247,N_10228);
and U13097 (N_13097,N_9803,N_9384);
and U13098 (N_13098,N_10393,N_10033);
and U13099 (N_13099,N_9657,N_11533);
and U13100 (N_13100,N_10942,N_9738);
nand U13101 (N_13101,N_10599,N_9630);
or U13102 (N_13102,N_11118,N_9143);
and U13103 (N_13103,N_10133,N_9823);
nor U13104 (N_13104,N_11833,N_9098);
nor U13105 (N_13105,N_9548,N_11421);
and U13106 (N_13106,N_9451,N_11497);
nor U13107 (N_13107,N_10706,N_10043);
and U13108 (N_13108,N_10895,N_10315);
nor U13109 (N_13109,N_11811,N_11129);
nand U13110 (N_13110,N_9339,N_9090);
and U13111 (N_13111,N_11392,N_11307);
nand U13112 (N_13112,N_11748,N_11508);
or U13113 (N_13113,N_10525,N_11269);
and U13114 (N_13114,N_11333,N_11194);
nor U13115 (N_13115,N_10945,N_9183);
or U13116 (N_13116,N_11881,N_9578);
nand U13117 (N_13117,N_9477,N_11036);
or U13118 (N_13118,N_9692,N_9685);
nand U13119 (N_13119,N_11855,N_9789);
and U13120 (N_13120,N_9437,N_9743);
nand U13121 (N_13121,N_11224,N_11883);
and U13122 (N_13122,N_9547,N_10622);
or U13123 (N_13123,N_10639,N_11385);
nor U13124 (N_13124,N_10318,N_9938);
or U13125 (N_13125,N_11200,N_11556);
or U13126 (N_13126,N_9570,N_10452);
or U13127 (N_13127,N_10790,N_9463);
nor U13128 (N_13128,N_11524,N_10486);
or U13129 (N_13129,N_9873,N_10817);
and U13130 (N_13130,N_10584,N_11127);
and U13131 (N_13131,N_10653,N_10885);
nor U13132 (N_13132,N_11948,N_9378);
and U13133 (N_13133,N_9922,N_10157);
and U13134 (N_13134,N_10390,N_10044);
and U13135 (N_13135,N_9327,N_10321);
or U13136 (N_13136,N_11683,N_9156);
and U13137 (N_13137,N_9589,N_9916);
nand U13138 (N_13138,N_9492,N_11252);
nor U13139 (N_13139,N_11886,N_10073);
and U13140 (N_13140,N_9358,N_10121);
or U13141 (N_13141,N_9159,N_10417);
nand U13142 (N_13142,N_9104,N_11329);
xnor U13143 (N_13143,N_10490,N_10731);
and U13144 (N_13144,N_11658,N_11526);
xnor U13145 (N_13145,N_10878,N_9760);
and U13146 (N_13146,N_9251,N_11447);
nand U13147 (N_13147,N_10151,N_9145);
or U13148 (N_13148,N_11233,N_10614);
and U13149 (N_13149,N_9150,N_11202);
and U13150 (N_13150,N_11215,N_9904);
nand U13151 (N_13151,N_9236,N_10533);
or U13152 (N_13152,N_10628,N_9036);
or U13153 (N_13153,N_11735,N_11622);
nor U13154 (N_13154,N_10277,N_10659);
or U13155 (N_13155,N_11929,N_11433);
and U13156 (N_13156,N_9273,N_10679);
or U13157 (N_13157,N_10748,N_11898);
or U13158 (N_13158,N_9908,N_10460);
or U13159 (N_13159,N_10795,N_11827);
nand U13160 (N_13160,N_9844,N_9593);
nand U13161 (N_13161,N_10463,N_10687);
and U13162 (N_13162,N_9520,N_11818);
and U13163 (N_13163,N_11355,N_11046);
and U13164 (N_13164,N_11411,N_11668);
or U13165 (N_13165,N_9859,N_10118);
nor U13166 (N_13166,N_11866,N_10046);
nand U13167 (N_13167,N_9467,N_9679);
nor U13168 (N_13168,N_11835,N_10921);
xor U13169 (N_13169,N_9994,N_9005);
nand U13170 (N_13170,N_11472,N_10664);
nor U13171 (N_13171,N_10747,N_9662);
and U13172 (N_13172,N_11796,N_9324);
and U13173 (N_13173,N_10148,N_10026);
or U13174 (N_13174,N_9756,N_9340);
and U13175 (N_13175,N_11863,N_10396);
and U13176 (N_13176,N_9995,N_11427);
or U13177 (N_13177,N_11558,N_11816);
or U13178 (N_13178,N_11589,N_11133);
nor U13179 (N_13179,N_11912,N_10915);
nand U13180 (N_13180,N_11819,N_10542);
nor U13181 (N_13181,N_9102,N_11343);
or U13182 (N_13182,N_10032,N_10254);
or U13183 (N_13183,N_11106,N_10132);
or U13184 (N_13184,N_10339,N_10150);
and U13185 (N_13185,N_11731,N_9454);
and U13186 (N_13186,N_10185,N_10823);
or U13187 (N_13187,N_9901,N_10937);
nor U13188 (N_13188,N_9095,N_11859);
or U13189 (N_13189,N_10801,N_9634);
or U13190 (N_13190,N_11493,N_9471);
nand U13191 (N_13191,N_11292,N_9759);
or U13192 (N_13192,N_9977,N_11365);
nand U13193 (N_13193,N_11342,N_10105);
and U13194 (N_13194,N_11862,N_11114);
or U13195 (N_13195,N_9056,N_10513);
nand U13196 (N_13196,N_10203,N_10421);
nor U13197 (N_13197,N_9221,N_10730);
nor U13198 (N_13198,N_9542,N_11867);
and U13199 (N_13199,N_10893,N_11235);
nor U13200 (N_13200,N_10630,N_11719);
nand U13201 (N_13201,N_10815,N_10481);
nand U13202 (N_13202,N_11218,N_11293);
nand U13203 (N_13203,N_10066,N_9820);
nand U13204 (N_13204,N_11262,N_9511);
nand U13205 (N_13205,N_9207,N_11303);
nand U13206 (N_13206,N_11196,N_10387);
or U13207 (N_13207,N_11953,N_11547);
nand U13208 (N_13208,N_9124,N_10998);
nand U13209 (N_13209,N_10994,N_9196);
or U13210 (N_13210,N_11399,N_10214);
nand U13211 (N_13211,N_10579,N_9170);
or U13212 (N_13212,N_10685,N_10833);
nand U13213 (N_13213,N_11029,N_11266);
nor U13214 (N_13214,N_10523,N_9268);
or U13215 (N_13215,N_10398,N_9153);
and U13216 (N_13216,N_11682,N_9504);
nor U13217 (N_13217,N_11150,N_11442);
and U13218 (N_13218,N_10432,N_9515);
nor U13219 (N_13219,N_9927,N_9133);
or U13220 (N_13220,N_10741,N_11864);
nor U13221 (N_13221,N_11205,N_11868);
nand U13222 (N_13222,N_10514,N_11592);
or U13223 (N_13223,N_9399,N_10246);
nand U13224 (N_13224,N_9449,N_10566);
nor U13225 (N_13225,N_11149,N_10336);
nor U13226 (N_13226,N_10154,N_11625);
nor U13227 (N_13227,N_10153,N_9610);
or U13228 (N_13228,N_9825,N_10295);
nor U13229 (N_13229,N_10722,N_9024);
nand U13230 (N_13230,N_11687,N_11536);
and U13231 (N_13231,N_11287,N_11375);
or U13232 (N_13232,N_9808,N_11935);
or U13233 (N_13233,N_9840,N_11849);
or U13234 (N_13234,N_9071,N_9772);
or U13235 (N_13235,N_11015,N_10912);
and U13236 (N_13236,N_10768,N_10829);
and U13237 (N_13237,N_9986,N_9006);
nand U13238 (N_13238,N_9874,N_10913);
and U13239 (N_13239,N_11672,N_9912);
nor U13240 (N_13240,N_9462,N_10897);
nor U13241 (N_13241,N_11977,N_10781);
nand U13242 (N_13242,N_9920,N_10491);
or U13243 (N_13243,N_11311,N_11989);
or U13244 (N_13244,N_11030,N_11000);
and U13245 (N_13245,N_9281,N_11125);
nor U13246 (N_13246,N_9544,N_10266);
nor U13247 (N_13247,N_10283,N_11974);
and U13248 (N_13248,N_11404,N_11770);
or U13249 (N_13249,N_9155,N_9198);
nor U13250 (N_13250,N_10637,N_11032);
nand U13251 (N_13251,N_10399,N_9677);
or U13252 (N_13252,N_9445,N_9109);
and U13253 (N_13253,N_11461,N_10976);
or U13254 (N_13254,N_10549,N_10380);
nand U13255 (N_13255,N_11933,N_11451);
and U13256 (N_13256,N_9990,N_11457);
or U13257 (N_13257,N_11352,N_11349);
or U13258 (N_13258,N_10974,N_11055);
or U13259 (N_13259,N_9476,N_10054);
nor U13260 (N_13260,N_10507,N_10278);
nand U13261 (N_13261,N_11147,N_10145);
and U13262 (N_13262,N_11131,N_11802);
nand U13263 (N_13263,N_9666,N_9126);
or U13264 (N_13264,N_11549,N_11336);
and U13265 (N_13265,N_9870,N_9336);
nor U13266 (N_13266,N_10479,N_9294);
and U13267 (N_13267,N_11344,N_10232);
nand U13268 (N_13268,N_10139,N_10019);
and U13269 (N_13269,N_11982,N_11492);
nor U13270 (N_13270,N_10075,N_11671);
and U13271 (N_13271,N_9639,N_10505);
nor U13272 (N_13272,N_11918,N_10991);
or U13273 (N_13273,N_10860,N_9579);
and U13274 (N_13274,N_11583,N_9567);
and U13275 (N_13275,N_10814,N_9565);
nand U13276 (N_13276,N_9114,N_11680);
or U13277 (N_13277,N_11939,N_9354);
or U13278 (N_13278,N_9562,N_9974);
and U13279 (N_13279,N_9396,N_11695);
nor U13280 (N_13280,N_9885,N_11458);
xnor U13281 (N_13281,N_11577,N_9359);
nor U13282 (N_13282,N_9369,N_10727);
and U13283 (N_13283,N_9142,N_10451);
or U13284 (N_13284,N_11585,N_11306);
nor U13285 (N_13285,N_10610,N_10353);
nor U13286 (N_13286,N_11160,N_11416);
and U13287 (N_13287,N_10646,N_10375);
nand U13288 (N_13288,N_10038,N_9684);
nor U13289 (N_13289,N_9289,N_11440);
nand U13290 (N_13290,N_11662,N_9617);
nor U13291 (N_13291,N_11920,N_11725);
nor U13292 (N_13292,N_10102,N_11257);
nor U13293 (N_13293,N_10484,N_9966);
and U13294 (N_13294,N_11685,N_10903);
or U13295 (N_13295,N_10870,N_9889);
nand U13296 (N_13296,N_11273,N_11309);
and U13297 (N_13297,N_11582,N_11946);
and U13298 (N_13298,N_10753,N_10816);
or U13299 (N_13299,N_10160,N_9232);
and U13300 (N_13300,N_11288,N_9606);
nor U13301 (N_13301,N_10987,N_9949);
or U13302 (N_13302,N_11008,N_11477);
nand U13303 (N_13303,N_11464,N_9855);
nor U13304 (N_13304,N_10325,N_11527);
xnor U13305 (N_13305,N_11213,N_11312);
xor U13306 (N_13306,N_11563,N_11817);
or U13307 (N_13307,N_11403,N_9406);
nand U13308 (N_13308,N_9195,N_11144);
or U13309 (N_13309,N_11617,N_11094);
or U13310 (N_13310,N_11116,N_11580);
nand U13311 (N_13311,N_9687,N_9412);
or U13312 (N_13312,N_9507,N_10377);
nand U13313 (N_13313,N_11142,N_10964);
and U13314 (N_13314,N_9586,N_11909);
or U13315 (N_13315,N_10068,N_10037);
or U13316 (N_13316,N_9318,N_10388);
or U13317 (N_13317,N_9398,N_10368);
nand U13318 (N_13318,N_9597,N_9433);
or U13319 (N_13319,N_10405,N_11418);
nor U13320 (N_13320,N_11520,N_10083);
nor U13321 (N_13321,N_9442,N_9737);
nor U13322 (N_13322,N_11108,N_9839);
nand U13323 (N_13323,N_11704,N_9829);
nor U13324 (N_13324,N_9888,N_10178);
or U13325 (N_13325,N_10881,N_11090);
and U13326 (N_13326,N_9501,N_10536);
nand U13327 (N_13327,N_10335,N_9708);
or U13328 (N_13328,N_10834,N_11620);
and U13329 (N_13329,N_9796,N_10803);
nor U13330 (N_13330,N_11363,N_10191);
nor U13331 (N_13331,N_11628,N_10517);
nor U13332 (N_13332,N_10088,N_10116);
or U13333 (N_13333,N_10188,N_11028);
nor U13334 (N_13334,N_10330,N_11098);
and U13335 (N_13335,N_10022,N_11791);
nand U13336 (N_13336,N_10708,N_9612);
and U13337 (N_13337,N_9942,N_11723);
or U13338 (N_13338,N_11879,N_11738);
nand U13339 (N_13339,N_10303,N_10957);
or U13340 (N_13340,N_9453,N_9910);
and U13341 (N_13341,N_11102,N_11552);
nand U13342 (N_13342,N_11208,N_11595);
nand U13343 (N_13343,N_11346,N_11070);
nand U13344 (N_13344,N_9871,N_11829);
nand U13345 (N_13345,N_9588,N_11297);
and U13346 (N_13346,N_11969,N_9264);
nand U13347 (N_13347,N_10632,N_10216);
and U13348 (N_13348,N_11268,N_10406);
and U13349 (N_13349,N_9731,N_11751);
nand U13350 (N_13350,N_9245,N_11531);
nor U13351 (N_13351,N_9370,N_11758);
and U13352 (N_13352,N_11468,N_9819);
and U13353 (N_13353,N_10791,N_11947);
xor U13354 (N_13354,N_11742,N_10404);
and U13355 (N_13355,N_9390,N_10252);
nor U13356 (N_13356,N_10993,N_9017);
nor U13357 (N_13357,N_10454,N_9518);
nand U13358 (N_13358,N_11398,N_10978);
nor U13359 (N_13359,N_9935,N_10558);
and U13360 (N_13360,N_10236,N_9409);
and U13361 (N_13361,N_9009,N_9146);
nand U13362 (N_13362,N_10689,N_11639);
and U13363 (N_13363,N_9965,N_9315);
and U13364 (N_13364,N_9008,N_11764);
xor U13365 (N_13365,N_10572,N_11573);
and U13366 (N_13366,N_10673,N_9134);
nor U13367 (N_13367,N_11371,N_11052);
or U13368 (N_13368,N_10775,N_10424);
nor U13369 (N_13369,N_9291,N_11005);
nor U13370 (N_13370,N_11322,N_11901);
nand U13371 (N_13371,N_9313,N_11083);
nand U13372 (N_13372,N_10400,N_9138);
nor U13373 (N_13373,N_10352,N_10176);
nor U13374 (N_13374,N_10034,N_11211);
nand U13375 (N_13375,N_11691,N_10410);
nor U13376 (N_13376,N_9577,N_11300);
nand U13377 (N_13377,N_9502,N_10299);
nand U13378 (N_13378,N_9943,N_11318);
nor U13379 (N_13379,N_9190,N_9539);
nor U13380 (N_13380,N_10042,N_11645);
nand U13381 (N_13381,N_9749,N_9733);
nor U13382 (N_13382,N_11887,N_9352);
nand U13383 (N_13383,N_10483,N_11584);
nor U13384 (N_13384,N_10218,N_11615);
nand U13385 (N_13385,N_11852,N_10500);
nor U13386 (N_13386,N_10767,N_10492);
and U13387 (N_13387,N_9322,N_10344);
nand U13388 (N_13388,N_11241,N_11315);
or U13389 (N_13389,N_11031,N_10308);
and U13390 (N_13390,N_10569,N_10868);
or U13391 (N_13391,N_10854,N_11913);
or U13392 (N_13392,N_11754,N_10861);
and U13393 (N_13393,N_9135,N_9900);
nand U13394 (N_13394,N_11787,N_9200);
nor U13395 (N_13395,N_9934,N_10710);
and U13396 (N_13396,N_9529,N_11677);
nor U13397 (N_13397,N_10346,N_10124);
and U13398 (N_13398,N_11313,N_11214);
or U13399 (N_13399,N_11986,N_10830);
and U13400 (N_13400,N_11726,N_9205);
nor U13401 (N_13401,N_11159,N_11686);
nand U13402 (N_13402,N_11393,N_9254);
or U13403 (N_13403,N_9103,N_9780);
nor U13404 (N_13404,N_11486,N_11987);
nor U13405 (N_13405,N_9394,N_10840);
nand U13406 (N_13406,N_11099,N_11972);
or U13407 (N_13407,N_9958,N_10433);
and U13408 (N_13408,N_11711,N_9381);
nor U13409 (N_13409,N_11460,N_10071);
and U13410 (N_13410,N_9086,N_9314);
nand U13411 (N_13411,N_10540,N_9778);
and U13412 (N_13412,N_10773,N_10698);
or U13413 (N_13413,N_10273,N_10084);
or U13414 (N_13414,N_10169,N_9957);
and U13415 (N_13415,N_10693,N_11446);
nor U13416 (N_13416,N_10021,N_9444);
nor U13417 (N_13417,N_9537,N_10617);
and U13418 (N_13418,N_9860,N_10441);
or U13419 (N_13419,N_11274,N_10951);
or U13420 (N_13420,N_11759,N_9890);
nand U13421 (N_13421,N_9773,N_11023);
nor U13422 (N_13422,N_9992,N_10667);
nor U13423 (N_13423,N_9946,N_11994);
nor U13424 (N_13424,N_11765,N_11345);
or U13425 (N_13425,N_9435,N_10129);
or U13426 (N_13426,N_10069,N_9285);
nand U13427 (N_13427,N_10204,N_9047);
nor U13428 (N_13428,N_11170,N_11007);
nor U13429 (N_13429,N_10074,N_9745);
and U13430 (N_13430,N_10954,N_11975);
nand U13431 (N_13431,N_11799,N_10063);
or U13432 (N_13432,N_10014,N_9311);
nand U13433 (N_13433,N_11869,N_9643);
and U13434 (N_13434,N_11390,N_10146);
and U13435 (N_13435,N_9441,N_11209);
nor U13436 (N_13436,N_11396,N_10040);
nor U13437 (N_13437,N_11699,N_9013);
or U13438 (N_13438,N_9421,N_9556);
nor U13439 (N_13439,N_10059,N_11650);
nand U13440 (N_13440,N_11324,N_11038);
or U13441 (N_13441,N_11076,N_11434);
nor U13442 (N_13442,N_11245,N_10910);
nor U13443 (N_13443,N_9826,N_9312);
nand U13444 (N_13444,N_11049,N_11476);
nand U13445 (N_13445,N_11945,N_9601);
nor U13446 (N_13446,N_9472,N_10446);
nand U13447 (N_13447,N_11146,N_10575);
nor U13448 (N_13448,N_10896,N_11610);
nor U13449 (N_13449,N_10376,N_9250);
nand U13450 (N_13450,N_9260,N_9316);
and U13451 (N_13451,N_10789,N_11161);
and U13452 (N_13452,N_10349,N_9618);
nor U13453 (N_13453,N_10544,N_11124);
or U13454 (N_13454,N_10294,N_10077);
and U13455 (N_13455,N_11347,N_9845);
nand U13456 (N_13456,N_10874,N_9676);
nor U13457 (N_13457,N_9532,N_11004);
nand U13458 (N_13458,N_10425,N_9080);
and U13459 (N_13459,N_10347,N_11978);
and U13460 (N_13460,N_9661,N_11487);
or U13461 (N_13461,N_11501,N_9262);
xnor U13462 (N_13462,N_9951,N_11372);
and U13463 (N_13463,N_11740,N_10314);
or U13464 (N_13464,N_11101,N_10161);
or U13465 (N_13465,N_11981,N_11568);
nand U13466 (N_13466,N_9473,N_10080);
or U13467 (N_13467,N_10757,N_9419);
nand U13468 (N_13468,N_11081,N_10826);
nand U13469 (N_13469,N_11428,N_10655);
nor U13470 (N_13470,N_9702,N_9836);
nand U13471 (N_13471,N_11395,N_11505);
nand U13472 (N_13472,N_10849,N_10035);
or U13473 (N_13473,N_10890,N_10386);
and U13474 (N_13474,N_10522,N_9375);
nand U13475 (N_13475,N_9875,N_9308);
or U13476 (N_13476,N_10772,N_10924);
nand U13477 (N_13477,N_10917,N_9292);
xnor U13478 (N_13478,N_10248,N_11207);
nand U13479 (N_13479,N_11027,N_10556);
and U13480 (N_13480,N_10943,N_11412);
nand U13481 (N_13481,N_11694,N_9847);
nand U13482 (N_13482,N_9498,N_11228);
xor U13483 (N_13483,N_9948,N_10411);
and U13484 (N_13484,N_11882,N_10143);
or U13485 (N_13485,N_10235,N_9097);
nand U13486 (N_13486,N_11400,N_11718);
and U13487 (N_13487,N_11275,N_10644);
and U13488 (N_13488,N_9488,N_10529);
nand U13489 (N_13489,N_9493,N_10596);
nand U13490 (N_13490,N_10898,N_10641);
nand U13491 (N_13491,N_11784,N_10546);
nor U13492 (N_13492,N_9023,N_9689);
or U13493 (N_13493,N_9457,N_10571);
nand U13494 (N_13494,N_9652,N_10418);
and U13495 (N_13495,N_9271,N_11499);
and U13496 (N_13496,N_10615,N_10799);
or U13497 (N_13497,N_11261,N_9728);
or U13498 (N_13498,N_10495,N_11236);
nor U13499 (N_13499,N_9964,N_11402);
nand U13500 (N_13500,N_9330,N_11367);
or U13501 (N_13501,N_11401,N_10129);
and U13502 (N_13502,N_11040,N_10251);
nor U13503 (N_13503,N_9962,N_11915);
and U13504 (N_13504,N_10553,N_10172);
nand U13505 (N_13505,N_10493,N_9110);
and U13506 (N_13506,N_10207,N_9530);
nor U13507 (N_13507,N_11578,N_10585);
nand U13508 (N_13508,N_9597,N_10273);
and U13509 (N_13509,N_11018,N_9988);
and U13510 (N_13510,N_11495,N_9676);
or U13511 (N_13511,N_10676,N_9228);
nor U13512 (N_13512,N_9284,N_10088);
or U13513 (N_13513,N_9836,N_9469);
nand U13514 (N_13514,N_9746,N_9585);
nand U13515 (N_13515,N_10060,N_11342);
nor U13516 (N_13516,N_11119,N_10805);
and U13517 (N_13517,N_10472,N_9077);
nand U13518 (N_13518,N_10843,N_11803);
or U13519 (N_13519,N_10218,N_10999);
nand U13520 (N_13520,N_9027,N_9457);
nand U13521 (N_13521,N_9252,N_10528);
nand U13522 (N_13522,N_9110,N_10992);
or U13523 (N_13523,N_10268,N_11821);
or U13524 (N_13524,N_9996,N_10383);
nor U13525 (N_13525,N_11699,N_9236);
nand U13526 (N_13526,N_11845,N_9576);
nor U13527 (N_13527,N_9357,N_11184);
and U13528 (N_13528,N_9051,N_9455);
and U13529 (N_13529,N_11385,N_10780);
nor U13530 (N_13530,N_11339,N_9953);
nor U13531 (N_13531,N_10702,N_9943);
nor U13532 (N_13532,N_11878,N_9079);
or U13533 (N_13533,N_10460,N_10421);
or U13534 (N_13534,N_9002,N_9394);
and U13535 (N_13535,N_11571,N_10646);
and U13536 (N_13536,N_11221,N_11347);
or U13537 (N_13537,N_9500,N_11940);
and U13538 (N_13538,N_10690,N_10905);
nand U13539 (N_13539,N_10435,N_9365);
nand U13540 (N_13540,N_11417,N_10572);
or U13541 (N_13541,N_10916,N_11871);
nor U13542 (N_13542,N_10600,N_9404);
or U13543 (N_13543,N_10450,N_9793);
and U13544 (N_13544,N_9490,N_10350);
and U13545 (N_13545,N_11941,N_9131);
and U13546 (N_13546,N_9111,N_11545);
and U13547 (N_13547,N_11502,N_10868);
nor U13548 (N_13548,N_9453,N_9783);
nand U13549 (N_13549,N_11960,N_9465);
or U13550 (N_13550,N_9401,N_11626);
nand U13551 (N_13551,N_10910,N_11139);
and U13552 (N_13552,N_9009,N_9299);
nor U13553 (N_13553,N_11812,N_11541);
nor U13554 (N_13554,N_11811,N_11785);
and U13555 (N_13555,N_10500,N_9382);
and U13556 (N_13556,N_9072,N_9315);
nand U13557 (N_13557,N_9758,N_9891);
and U13558 (N_13558,N_10646,N_10332);
and U13559 (N_13559,N_10294,N_9218);
and U13560 (N_13560,N_11191,N_11322);
or U13561 (N_13561,N_9551,N_9393);
nor U13562 (N_13562,N_10440,N_10735);
or U13563 (N_13563,N_9315,N_9963);
or U13564 (N_13564,N_10380,N_10586);
or U13565 (N_13565,N_11166,N_10586);
nand U13566 (N_13566,N_11137,N_9999);
or U13567 (N_13567,N_9374,N_10079);
and U13568 (N_13568,N_10855,N_10997);
and U13569 (N_13569,N_10405,N_10853);
or U13570 (N_13570,N_9813,N_10416);
nand U13571 (N_13571,N_10885,N_10707);
nand U13572 (N_13572,N_10572,N_11618);
or U13573 (N_13573,N_11230,N_11542);
xor U13574 (N_13574,N_9463,N_10807);
or U13575 (N_13575,N_9281,N_11982);
nand U13576 (N_13576,N_11218,N_11228);
and U13577 (N_13577,N_11551,N_11566);
and U13578 (N_13578,N_11901,N_9246);
nand U13579 (N_13579,N_9671,N_10912);
nand U13580 (N_13580,N_9767,N_11033);
nor U13581 (N_13581,N_11868,N_9483);
and U13582 (N_13582,N_9827,N_9160);
nor U13583 (N_13583,N_11445,N_9619);
nand U13584 (N_13584,N_9428,N_10441);
and U13585 (N_13585,N_10175,N_10987);
or U13586 (N_13586,N_10452,N_9810);
or U13587 (N_13587,N_9497,N_9009);
and U13588 (N_13588,N_11000,N_10535);
and U13589 (N_13589,N_10107,N_9320);
nand U13590 (N_13590,N_10757,N_10401);
or U13591 (N_13591,N_9220,N_11796);
and U13592 (N_13592,N_10045,N_10739);
nand U13593 (N_13593,N_11293,N_10694);
nand U13594 (N_13594,N_11159,N_10988);
nand U13595 (N_13595,N_10116,N_9693);
or U13596 (N_13596,N_9781,N_11484);
xnor U13597 (N_13597,N_11492,N_11099);
nor U13598 (N_13598,N_10241,N_10644);
xor U13599 (N_13599,N_10359,N_9708);
nand U13600 (N_13600,N_9526,N_9394);
nand U13601 (N_13601,N_11528,N_11140);
and U13602 (N_13602,N_9767,N_9949);
and U13603 (N_13603,N_9457,N_11680);
nand U13604 (N_13604,N_11714,N_11158);
and U13605 (N_13605,N_11200,N_11201);
nand U13606 (N_13606,N_9711,N_9514);
nor U13607 (N_13607,N_10106,N_9702);
nor U13608 (N_13608,N_10856,N_11092);
nand U13609 (N_13609,N_9462,N_11316);
nand U13610 (N_13610,N_10372,N_9325);
nor U13611 (N_13611,N_11727,N_9586);
and U13612 (N_13612,N_9899,N_9812);
and U13613 (N_13613,N_10220,N_10638);
or U13614 (N_13614,N_11289,N_10888);
nand U13615 (N_13615,N_11057,N_11011);
nor U13616 (N_13616,N_11680,N_10629);
xnor U13617 (N_13617,N_10245,N_11693);
and U13618 (N_13618,N_10687,N_9343);
or U13619 (N_13619,N_10698,N_11792);
nand U13620 (N_13620,N_10008,N_9672);
xor U13621 (N_13621,N_9990,N_10395);
and U13622 (N_13622,N_9414,N_11150);
or U13623 (N_13623,N_9249,N_11059);
nor U13624 (N_13624,N_11241,N_11174);
or U13625 (N_13625,N_10489,N_11251);
and U13626 (N_13626,N_11700,N_10495);
xor U13627 (N_13627,N_9208,N_11331);
or U13628 (N_13628,N_11681,N_9529);
nand U13629 (N_13629,N_10239,N_11428);
nand U13630 (N_13630,N_11653,N_9202);
or U13631 (N_13631,N_10174,N_9478);
nand U13632 (N_13632,N_9601,N_11410);
nor U13633 (N_13633,N_10278,N_11706);
or U13634 (N_13634,N_9033,N_9296);
or U13635 (N_13635,N_11048,N_11845);
nor U13636 (N_13636,N_9992,N_9466);
xnor U13637 (N_13637,N_10724,N_11983);
or U13638 (N_13638,N_10630,N_9438);
and U13639 (N_13639,N_10970,N_9796);
nor U13640 (N_13640,N_10052,N_10396);
nand U13641 (N_13641,N_10662,N_10394);
nor U13642 (N_13642,N_11272,N_9511);
nor U13643 (N_13643,N_11445,N_10991);
or U13644 (N_13644,N_9518,N_9564);
and U13645 (N_13645,N_9154,N_9818);
and U13646 (N_13646,N_9382,N_11924);
nor U13647 (N_13647,N_10920,N_11642);
and U13648 (N_13648,N_9000,N_11795);
or U13649 (N_13649,N_9758,N_11373);
and U13650 (N_13650,N_9379,N_10982);
and U13651 (N_13651,N_10094,N_10623);
nand U13652 (N_13652,N_10929,N_10919);
nand U13653 (N_13653,N_10342,N_11520);
and U13654 (N_13654,N_11359,N_10433);
or U13655 (N_13655,N_9569,N_10312);
and U13656 (N_13656,N_9869,N_9884);
nor U13657 (N_13657,N_11053,N_10931);
or U13658 (N_13658,N_11400,N_10909);
nor U13659 (N_13659,N_10538,N_9911);
or U13660 (N_13660,N_10740,N_9878);
and U13661 (N_13661,N_11019,N_9463);
and U13662 (N_13662,N_9469,N_10731);
nor U13663 (N_13663,N_11139,N_11369);
nand U13664 (N_13664,N_11921,N_9212);
nor U13665 (N_13665,N_9814,N_10972);
nand U13666 (N_13666,N_10940,N_11056);
nor U13667 (N_13667,N_11384,N_9355);
or U13668 (N_13668,N_11711,N_9488);
nor U13669 (N_13669,N_10307,N_11788);
and U13670 (N_13670,N_11735,N_10669);
nor U13671 (N_13671,N_9335,N_9164);
nand U13672 (N_13672,N_11692,N_11799);
and U13673 (N_13673,N_11507,N_10338);
or U13674 (N_13674,N_11112,N_10044);
or U13675 (N_13675,N_9466,N_10567);
nand U13676 (N_13676,N_9717,N_9028);
or U13677 (N_13677,N_11785,N_11246);
nand U13678 (N_13678,N_9102,N_11743);
nor U13679 (N_13679,N_9767,N_11692);
nand U13680 (N_13680,N_11704,N_9444);
and U13681 (N_13681,N_9642,N_10072);
or U13682 (N_13682,N_11367,N_11866);
nor U13683 (N_13683,N_11858,N_10601);
nand U13684 (N_13684,N_11630,N_11085);
or U13685 (N_13685,N_11405,N_10728);
nand U13686 (N_13686,N_10041,N_9041);
nor U13687 (N_13687,N_10659,N_10752);
nand U13688 (N_13688,N_10999,N_9916);
and U13689 (N_13689,N_11934,N_11843);
or U13690 (N_13690,N_9319,N_9469);
nand U13691 (N_13691,N_9403,N_11061);
nor U13692 (N_13692,N_9144,N_9132);
or U13693 (N_13693,N_10980,N_9609);
or U13694 (N_13694,N_9717,N_11405);
or U13695 (N_13695,N_11223,N_9898);
nand U13696 (N_13696,N_10705,N_9087);
and U13697 (N_13697,N_9453,N_9847);
nand U13698 (N_13698,N_10854,N_11069);
nand U13699 (N_13699,N_9127,N_11757);
or U13700 (N_13700,N_10491,N_9006);
nor U13701 (N_13701,N_11989,N_11055);
nor U13702 (N_13702,N_11021,N_9985);
and U13703 (N_13703,N_10310,N_10084);
nor U13704 (N_13704,N_9497,N_10570);
and U13705 (N_13705,N_10739,N_11312);
and U13706 (N_13706,N_11275,N_9810);
and U13707 (N_13707,N_10300,N_11750);
nor U13708 (N_13708,N_10613,N_11418);
nand U13709 (N_13709,N_9832,N_11345);
nand U13710 (N_13710,N_9097,N_10042);
xor U13711 (N_13711,N_11940,N_9048);
or U13712 (N_13712,N_10431,N_11533);
or U13713 (N_13713,N_11591,N_11624);
and U13714 (N_13714,N_9528,N_9160);
and U13715 (N_13715,N_10102,N_9920);
or U13716 (N_13716,N_11071,N_10187);
or U13717 (N_13717,N_9332,N_9129);
and U13718 (N_13718,N_10281,N_11739);
and U13719 (N_13719,N_11137,N_11380);
nand U13720 (N_13720,N_9316,N_11953);
nand U13721 (N_13721,N_10669,N_10609);
and U13722 (N_13722,N_11525,N_10819);
nand U13723 (N_13723,N_11616,N_9630);
nor U13724 (N_13724,N_11839,N_9158);
nand U13725 (N_13725,N_10902,N_11668);
nor U13726 (N_13726,N_11137,N_10422);
nand U13727 (N_13727,N_9277,N_10702);
nor U13728 (N_13728,N_9470,N_11531);
xnor U13729 (N_13729,N_9115,N_9122);
nor U13730 (N_13730,N_11697,N_9079);
nor U13731 (N_13731,N_9662,N_11672);
and U13732 (N_13732,N_11020,N_10201);
or U13733 (N_13733,N_11942,N_10411);
and U13734 (N_13734,N_11385,N_9325);
nor U13735 (N_13735,N_9545,N_11019);
and U13736 (N_13736,N_9012,N_10053);
or U13737 (N_13737,N_9427,N_10499);
or U13738 (N_13738,N_11359,N_10253);
nand U13739 (N_13739,N_10493,N_9548);
nand U13740 (N_13740,N_10780,N_10459);
nand U13741 (N_13741,N_9091,N_11691);
or U13742 (N_13742,N_11185,N_10025);
nand U13743 (N_13743,N_11966,N_10356);
and U13744 (N_13744,N_10369,N_11292);
nor U13745 (N_13745,N_10681,N_10999);
nor U13746 (N_13746,N_10018,N_9562);
nor U13747 (N_13747,N_10422,N_11288);
and U13748 (N_13748,N_10338,N_11919);
nand U13749 (N_13749,N_10751,N_9968);
nor U13750 (N_13750,N_10107,N_11432);
nand U13751 (N_13751,N_10765,N_11016);
nand U13752 (N_13752,N_9831,N_10263);
or U13753 (N_13753,N_9131,N_11297);
and U13754 (N_13754,N_9996,N_9373);
and U13755 (N_13755,N_9284,N_9838);
nand U13756 (N_13756,N_11616,N_10691);
nor U13757 (N_13757,N_9658,N_11715);
nand U13758 (N_13758,N_9565,N_9865);
nand U13759 (N_13759,N_11935,N_11083);
nand U13760 (N_13760,N_11027,N_10543);
nor U13761 (N_13761,N_11802,N_11839);
nor U13762 (N_13762,N_9585,N_11931);
or U13763 (N_13763,N_9818,N_11934);
nand U13764 (N_13764,N_10442,N_9343);
and U13765 (N_13765,N_9775,N_10074);
or U13766 (N_13766,N_10508,N_11091);
xnor U13767 (N_13767,N_10009,N_9507);
and U13768 (N_13768,N_9231,N_10403);
nand U13769 (N_13769,N_9257,N_10120);
nor U13770 (N_13770,N_10403,N_9675);
nor U13771 (N_13771,N_9835,N_10362);
nand U13772 (N_13772,N_11366,N_9564);
or U13773 (N_13773,N_11928,N_9632);
or U13774 (N_13774,N_9303,N_9152);
nor U13775 (N_13775,N_9366,N_9948);
nor U13776 (N_13776,N_9072,N_10468);
and U13777 (N_13777,N_9809,N_10966);
or U13778 (N_13778,N_9930,N_11946);
nor U13779 (N_13779,N_10247,N_9366);
nand U13780 (N_13780,N_9580,N_11710);
nand U13781 (N_13781,N_9963,N_9392);
nand U13782 (N_13782,N_11948,N_9753);
or U13783 (N_13783,N_11858,N_9726);
nand U13784 (N_13784,N_10430,N_10800);
and U13785 (N_13785,N_10819,N_9556);
and U13786 (N_13786,N_10468,N_10340);
nand U13787 (N_13787,N_9490,N_10526);
nand U13788 (N_13788,N_10588,N_11894);
and U13789 (N_13789,N_11121,N_9205);
and U13790 (N_13790,N_9088,N_9632);
nor U13791 (N_13791,N_11889,N_9353);
nor U13792 (N_13792,N_10958,N_11464);
or U13793 (N_13793,N_11870,N_9541);
nor U13794 (N_13794,N_9236,N_11195);
nor U13795 (N_13795,N_9531,N_9928);
nand U13796 (N_13796,N_11659,N_11034);
nand U13797 (N_13797,N_10227,N_11435);
or U13798 (N_13798,N_9126,N_11174);
nand U13799 (N_13799,N_9314,N_9715);
and U13800 (N_13800,N_11381,N_11635);
nor U13801 (N_13801,N_9613,N_10454);
nor U13802 (N_13802,N_11379,N_11773);
nor U13803 (N_13803,N_11010,N_11252);
and U13804 (N_13804,N_9126,N_11388);
or U13805 (N_13805,N_10083,N_11503);
or U13806 (N_13806,N_9212,N_9884);
nor U13807 (N_13807,N_9260,N_10993);
nand U13808 (N_13808,N_10956,N_10913);
nand U13809 (N_13809,N_11847,N_10655);
or U13810 (N_13810,N_9824,N_9208);
or U13811 (N_13811,N_10100,N_9056);
nand U13812 (N_13812,N_9640,N_9962);
and U13813 (N_13813,N_9887,N_10409);
and U13814 (N_13814,N_10052,N_10130);
nand U13815 (N_13815,N_9943,N_11566);
and U13816 (N_13816,N_11984,N_10020);
nand U13817 (N_13817,N_11878,N_9061);
nor U13818 (N_13818,N_11729,N_10516);
nor U13819 (N_13819,N_11029,N_11774);
nand U13820 (N_13820,N_10922,N_11060);
nand U13821 (N_13821,N_11384,N_10921);
nand U13822 (N_13822,N_9077,N_10410);
and U13823 (N_13823,N_9979,N_9976);
nand U13824 (N_13824,N_10797,N_9494);
nand U13825 (N_13825,N_9330,N_9500);
nor U13826 (N_13826,N_9302,N_10788);
nor U13827 (N_13827,N_10401,N_10962);
or U13828 (N_13828,N_9526,N_11697);
nand U13829 (N_13829,N_9090,N_11309);
or U13830 (N_13830,N_9316,N_11077);
or U13831 (N_13831,N_11262,N_9457);
xnor U13832 (N_13832,N_11487,N_9137);
and U13833 (N_13833,N_11234,N_11549);
or U13834 (N_13834,N_10745,N_10856);
nand U13835 (N_13835,N_10870,N_11299);
and U13836 (N_13836,N_11894,N_11920);
and U13837 (N_13837,N_9611,N_9543);
or U13838 (N_13838,N_10572,N_10867);
or U13839 (N_13839,N_10399,N_9828);
nand U13840 (N_13840,N_10684,N_9692);
or U13841 (N_13841,N_9938,N_9005);
nand U13842 (N_13842,N_10058,N_9560);
and U13843 (N_13843,N_9596,N_10430);
and U13844 (N_13844,N_9086,N_9682);
and U13845 (N_13845,N_9168,N_9682);
or U13846 (N_13846,N_11409,N_10650);
and U13847 (N_13847,N_10129,N_9047);
or U13848 (N_13848,N_10387,N_10995);
xor U13849 (N_13849,N_9645,N_9795);
or U13850 (N_13850,N_10742,N_10010);
or U13851 (N_13851,N_10624,N_10279);
and U13852 (N_13852,N_10743,N_11058);
nand U13853 (N_13853,N_11969,N_11200);
nor U13854 (N_13854,N_9396,N_11265);
nor U13855 (N_13855,N_10521,N_9215);
and U13856 (N_13856,N_10158,N_9746);
nand U13857 (N_13857,N_10776,N_9773);
nor U13858 (N_13858,N_11655,N_11498);
xor U13859 (N_13859,N_9323,N_9828);
nor U13860 (N_13860,N_10079,N_10830);
or U13861 (N_13861,N_9829,N_11902);
and U13862 (N_13862,N_11716,N_10696);
nor U13863 (N_13863,N_9477,N_9918);
and U13864 (N_13864,N_11539,N_9228);
or U13865 (N_13865,N_11979,N_11092);
and U13866 (N_13866,N_11517,N_10606);
nand U13867 (N_13867,N_9169,N_9918);
and U13868 (N_13868,N_10296,N_9883);
and U13869 (N_13869,N_10152,N_10626);
and U13870 (N_13870,N_9514,N_10953);
nor U13871 (N_13871,N_10817,N_9239);
or U13872 (N_13872,N_9900,N_11818);
or U13873 (N_13873,N_9061,N_11468);
nor U13874 (N_13874,N_11400,N_10878);
and U13875 (N_13875,N_11927,N_9439);
nand U13876 (N_13876,N_11017,N_10060);
nand U13877 (N_13877,N_10377,N_11500);
nand U13878 (N_13878,N_9534,N_9376);
nor U13879 (N_13879,N_9851,N_9288);
nand U13880 (N_13880,N_11293,N_9249);
nand U13881 (N_13881,N_11601,N_9520);
or U13882 (N_13882,N_9351,N_10996);
nand U13883 (N_13883,N_10253,N_10900);
xor U13884 (N_13884,N_11634,N_9909);
nand U13885 (N_13885,N_9581,N_9823);
or U13886 (N_13886,N_11872,N_11564);
nand U13887 (N_13887,N_9431,N_10927);
nor U13888 (N_13888,N_10446,N_9757);
nor U13889 (N_13889,N_10611,N_10412);
and U13890 (N_13890,N_11637,N_11916);
or U13891 (N_13891,N_10313,N_10333);
or U13892 (N_13892,N_10215,N_11641);
and U13893 (N_13893,N_10492,N_10261);
and U13894 (N_13894,N_11798,N_11026);
or U13895 (N_13895,N_11181,N_11443);
nor U13896 (N_13896,N_11679,N_10796);
and U13897 (N_13897,N_11347,N_11558);
and U13898 (N_13898,N_11841,N_10626);
and U13899 (N_13899,N_10134,N_11644);
nor U13900 (N_13900,N_9987,N_10892);
and U13901 (N_13901,N_9384,N_10027);
or U13902 (N_13902,N_11946,N_10524);
and U13903 (N_13903,N_9859,N_9430);
nor U13904 (N_13904,N_11763,N_11508);
nor U13905 (N_13905,N_11886,N_10316);
or U13906 (N_13906,N_9708,N_10990);
and U13907 (N_13907,N_10919,N_9092);
nand U13908 (N_13908,N_10006,N_11229);
or U13909 (N_13909,N_10121,N_11091);
and U13910 (N_13910,N_10571,N_10623);
or U13911 (N_13911,N_9076,N_11423);
nand U13912 (N_13912,N_10732,N_10598);
or U13913 (N_13913,N_11749,N_11944);
or U13914 (N_13914,N_9297,N_10502);
xnor U13915 (N_13915,N_9645,N_10951);
or U13916 (N_13916,N_9536,N_9229);
nand U13917 (N_13917,N_10356,N_10654);
nand U13918 (N_13918,N_11963,N_9861);
xnor U13919 (N_13919,N_10629,N_11125);
and U13920 (N_13920,N_10357,N_10538);
and U13921 (N_13921,N_9199,N_11877);
nand U13922 (N_13922,N_9314,N_10647);
and U13923 (N_13923,N_10858,N_9885);
or U13924 (N_13924,N_9859,N_10815);
nor U13925 (N_13925,N_9037,N_11842);
and U13926 (N_13926,N_11942,N_11812);
or U13927 (N_13927,N_11368,N_9191);
or U13928 (N_13928,N_9419,N_10788);
or U13929 (N_13929,N_10489,N_11200);
nor U13930 (N_13930,N_10584,N_9578);
nor U13931 (N_13931,N_9331,N_11865);
xnor U13932 (N_13932,N_10920,N_9412);
nand U13933 (N_13933,N_9814,N_11739);
nand U13934 (N_13934,N_9959,N_10081);
nand U13935 (N_13935,N_11786,N_9847);
nor U13936 (N_13936,N_9028,N_10806);
or U13937 (N_13937,N_11708,N_10546);
and U13938 (N_13938,N_11370,N_9536);
or U13939 (N_13939,N_10075,N_11737);
xor U13940 (N_13940,N_9691,N_11809);
or U13941 (N_13941,N_10214,N_10852);
and U13942 (N_13942,N_11976,N_10313);
nand U13943 (N_13943,N_10761,N_10748);
nor U13944 (N_13944,N_11258,N_10037);
nor U13945 (N_13945,N_11039,N_10127);
or U13946 (N_13946,N_10294,N_11644);
or U13947 (N_13947,N_11297,N_10299);
or U13948 (N_13948,N_10337,N_11781);
nor U13949 (N_13949,N_9974,N_9311);
and U13950 (N_13950,N_9976,N_10770);
or U13951 (N_13951,N_9827,N_11491);
and U13952 (N_13952,N_11657,N_10501);
nand U13953 (N_13953,N_9687,N_9339);
nand U13954 (N_13954,N_11402,N_10612);
nand U13955 (N_13955,N_11613,N_11096);
nor U13956 (N_13956,N_10162,N_11832);
or U13957 (N_13957,N_10462,N_11992);
and U13958 (N_13958,N_10724,N_11426);
and U13959 (N_13959,N_10063,N_10522);
nand U13960 (N_13960,N_11921,N_9801);
and U13961 (N_13961,N_9301,N_11811);
and U13962 (N_13962,N_11879,N_11036);
nand U13963 (N_13963,N_10388,N_11812);
and U13964 (N_13964,N_10359,N_11607);
nand U13965 (N_13965,N_11113,N_10743);
or U13966 (N_13966,N_10862,N_10483);
or U13967 (N_13967,N_10861,N_9745);
or U13968 (N_13968,N_9802,N_9157);
or U13969 (N_13969,N_10765,N_9862);
nor U13970 (N_13970,N_9170,N_10289);
nand U13971 (N_13971,N_11611,N_11521);
or U13972 (N_13972,N_11315,N_11689);
nor U13973 (N_13973,N_9615,N_9932);
or U13974 (N_13974,N_9212,N_10884);
and U13975 (N_13975,N_11316,N_9373);
or U13976 (N_13976,N_10386,N_10098);
nor U13977 (N_13977,N_9672,N_9627);
and U13978 (N_13978,N_10791,N_9546);
or U13979 (N_13979,N_10507,N_11015);
nand U13980 (N_13980,N_11216,N_9608);
xnor U13981 (N_13981,N_11136,N_9636);
or U13982 (N_13982,N_9901,N_9956);
and U13983 (N_13983,N_9437,N_11784);
or U13984 (N_13984,N_9345,N_9527);
or U13985 (N_13985,N_11170,N_11833);
and U13986 (N_13986,N_9710,N_11739);
nand U13987 (N_13987,N_9689,N_11786);
and U13988 (N_13988,N_11569,N_9653);
and U13989 (N_13989,N_10129,N_11732);
and U13990 (N_13990,N_10653,N_9326);
or U13991 (N_13991,N_10583,N_11466);
nand U13992 (N_13992,N_10317,N_9317);
or U13993 (N_13993,N_10894,N_9109);
and U13994 (N_13994,N_11981,N_9313);
nand U13995 (N_13995,N_9050,N_9007);
and U13996 (N_13996,N_11522,N_9220);
xnor U13997 (N_13997,N_9194,N_10685);
and U13998 (N_13998,N_9565,N_10389);
nor U13999 (N_13999,N_11763,N_11363);
and U14000 (N_14000,N_9642,N_11463);
or U14001 (N_14001,N_11035,N_10391);
and U14002 (N_14002,N_9057,N_10942);
nand U14003 (N_14003,N_9474,N_10774);
nor U14004 (N_14004,N_11475,N_11874);
nand U14005 (N_14005,N_10998,N_10070);
xnor U14006 (N_14006,N_10134,N_10091);
nand U14007 (N_14007,N_11477,N_9453);
nand U14008 (N_14008,N_9312,N_10426);
nor U14009 (N_14009,N_9557,N_9376);
nor U14010 (N_14010,N_11750,N_9684);
and U14011 (N_14011,N_11332,N_9085);
or U14012 (N_14012,N_9743,N_11428);
nand U14013 (N_14013,N_9846,N_10702);
nor U14014 (N_14014,N_11817,N_9976);
and U14015 (N_14015,N_10810,N_9434);
and U14016 (N_14016,N_11725,N_11635);
or U14017 (N_14017,N_10565,N_11996);
nand U14018 (N_14018,N_10471,N_10827);
or U14019 (N_14019,N_9140,N_10440);
or U14020 (N_14020,N_11678,N_10175);
xnor U14021 (N_14021,N_11403,N_11565);
or U14022 (N_14022,N_9248,N_10557);
xnor U14023 (N_14023,N_10669,N_10042);
and U14024 (N_14024,N_11773,N_10699);
or U14025 (N_14025,N_11888,N_11372);
and U14026 (N_14026,N_10541,N_9342);
nor U14027 (N_14027,N_9100,N_11504);
or U14028 (N_14028,N_11307,N_11094);
or U14029 (N_14029,N_9180,N_9248);
or U14030 (N_14030,N_10232,N_11316);
or U14031 (N_14031,N_11336,N_9101);
or U14032 (N_14032,N_11155,N_10244);
or U14033 (N_14033,N_10492,N_10828);
or U14034 (N_14034,N_10028,N_9099);
or U14035 (N_14035,N_9395,N_9125);
or U14036 (N_14036,N_9257,N_11841);
or U14037 (N_14037,N_11443,N_10876);
and U14038 (N_14038,N_9762,N_10893);
nand U14039 (N_14039,N_11999,N_11947);
nand U14040 (N_14040,N_9091,N_10502);
or U14041 (N_14041,N_10138,N_10175);
nand U14042 (N_14042,N_10395,N_9986);
and U14043 (N_14043,N_9945,N_9552);
or U14044 (N_14044,N_9901,N_11701);
or U14045 (N_14045,N_9179,N_9506);
xor U14046 (N_14046,N_11090,N_11975);
or U14047 (N_14047,N_11176,N_11738);
and U14048 (N_14048,N_10183,N_11910);
nor U14049 (N_14049,N_11495,N_10846);
and U14050 (N_14050,N_9563,N_11342);
nor U14051 (N_14051,N_9353,N_11380);
or U14052 (N_14052,N_11818,N_10640);
nor U14053 (N_14053,N_9990,N_9999);
nor U14054 (N_14054,N_10145,N_9467);
or U14055 (N_14055,N_9546,N_10422);
nand U14056 (N_14056,N_11937,N_9067);
or U14057 (N_14057,N_11320,N_9144);
and U14058 (N_14058,N_9651,N_10057);
or U14059 (N_14059,N_9260,N_9741);
or U14060 (N_14060,N_9019,N_9722);
nor U14061 (N_14061,N_10132,N_9133);
or U14062 (N_14062,N_11669,N_11830);
nand U14063 (N_14063,N_9982,N_11205);
or U14064 (N_14064,N_11051,N_10872);
xor U14065 (N_14065,N_11468,N_9963);
or U14066 (N_14066,N_10410,N_9836);
nor U14067 (N_14067,N_10734,N_9898);
or U14068 (N_14068,N_10076,N_10413);
xnor U14069 (N_14069,N_10985,N_10390);
and U14070 (N_14070,N_9326,N_11314);
nand U14071 (N_14071,N_10457,N_9355);
or U14072 (N_14072,N_10076,N_9992);
nor U14073 (N_14073,N_9459,N_9694);
nor U14074 (N_14074,N_10421,N_9158);
nand U14075 (N_14075,N_9620,N_10943);
nor U14076 (N_14076,N_9470,N_10407);
or U14077 (N_14077,N_11973,N_10766);
nor U14078 (N_14078,N_11968,N_9428);
and U14079 (N_14079,N_10154,N_11113);
and U14080 (N_14080,N_11384,N_10275);
and U14081 (N_14081,N_11866,N_11711);
nand U14082 (N_14082,N_9448,N_10562);
and U14083 (N_14083,N_9274,N_9358);
and U14084 (N_14084,N_9925,N_11384);
nor U14085 (N_14085,N_10095,N_10787);
nand U14086 (N_14086,N_9472,N_11223);
nor U14087 (N_14087,N_10448,N_9556);
and U14088 (N_14088,N_10770,N_11618);
nor U14089 (N_14089,N_10120,N_9035);
nor U14090 (N_14090,N_11235,N_10477);
or U14091 (N_14091,N_10925,N_10375);
nand U14092 (N_14092,N_11043,N_9077);
nor U14093 (N_14093,N_10955,N_10439);
or U14094 (N_14094,N_9167,N_9898);
nor U14095 (N_14095,N_9984,N_11849);
and U14096 (N_14096,N_10708,N_9479);
nand U14097 (N_14097,N_11757,N_11620);
nand U14098 (N_14098,N_9311,N_11374);
and U14099 (N_14099,N_11146,N_10010);
nor U14100 (N_14100,N_11001,N_10061);
or U14101 (N_14101,N_10078,N_9769);
nand U14102 (N_14102,N_10654,N_11090);
nor U14103 (N_14103,N_11600,N_9972);
and U14104 (N_14104,N_10713,N_9282);
or U14105 (N_14105,N_10588,N_9433);
nor U14106 (N_14106,N_9142,N_9445);
nor U14107 (N_14107,N_9066,N_11450);
nand U14108 (N_14108,N_10348,N_9707);
and U14109 (N_14109,N_10722,N_10451);
or U14110 (N_14110,N_9672,N_9575);
nand U14111 (N_14111,N_11108,N_10548);
nand U14112 (N_14112,N_9504,N_9793);
nor U14113 (N_14113,N_11275,N_9632);
nand U14114 (N_14114,N_9122,N_10363);
and U14115 (N_14115,N_10733,N_11799);
nor U14116 (N_14116,N_11917,N_9452);
nor U14117 (N_14117,N_11086,N_9605);
or U14118 (N_14118,N_11704,N_10137);
nand U14119 (N_14119,N_9170,N_9709);
and U14120 (N_14120,N_10219,N_10348);
nor U14121 (N_14121,N_10123,N_9674);
or U14122 (N_14122,N_9163,N_11722);
and U14123 (N_14123,N_9656,N_11799);
nand U14124 (N_14124,N_9987,N_11382);
nor U14125 (N_14125,N_11065,N_9970);
nand U14126 (N_14126,N_9168,N_11012);
nand U14127 (N_14127,N_9666,N_10701);
xnor U14128 (N_14128,N_10870,N_9503);
and U14129 (N_14129,N_10908,N_11919);
and U14130 (N_14130,N_10117,N_9252);
nand U14131 (N_14131,N_11298,N_10415);
nand U14132 (N_14132,N_10282,N_9014);
nor U14133 (N_14133,N_10019,N_10132);
and U14134 (N_14134,N_9691,N_10906);
nor U14135 (N_14135,N_11733,N_11957);
nand U14136 (N_14136,N_11179,N_11207);
nand U14137 (N_14137,N_10780,N_10728);
and U14138 (N_14138,N_10174,N_10547);
or U14139 (N_14139,N_10245,N_11675);
nand U14140 (N_14140,N_10294,N_11982);
nor U14141 (N_14141,N_9334,N_10639);
nor U14142 (N_14142,N_10892,N_10201);
or U14143 (N_14143,N_11083,N_11409);
or U14144 (N_14144,N_9254,N_10377);
nor U14145 (N_14145,N_11897,N_9979);
nand U14146 (N_14146,N_9960,N_11146);
nor U14147 (N_14147,N_10796,N_11463);
nand U14148 (N_14148,N_10069,N_10247);
nor U14149 (N_14149,N_9737,N_9100);
nand U14150 (N_14150,N_10121,N_9199);
or U14151 (N_14151,N_11573,N_9610);
nand U14152 (N_14152,N_10802,N_10160);
or U14153 (N_14153,N_10721,N_9540);
xor U14154 (N_14154,N_11607,N_10049);
and U14155 (N_14155,N_11270,N_11517);
and U14156 (N_14156,N_10252,N_10045);
nand U14157 (N_14157,N_9752,N_11991);
and U14158 (N_14158,N_10225,N_10204);
nand U14159 (N_14159,N_9189,N_10936);
or U14160 (N_14160,N_11040,N_11190);
and U14161 (N_14161,N_9176,N_10955);
nand U14162 (N_14162,N_11732,N_10339);
or U14163 (N_14163,N_9928,N_11210);
or U14164 (N_14164,N_9976,N_9454);
nor U14165 (N_14165,N_10622,N_9247);
nor U14166 (N_14166,N_10179,N_9937);
xor U14167 (N_14167,N_11512,N_9664);
and U14168 (N_14168,N_11486,N_9751);
nand U14169 (N_14169,N_9765,N_10398);
or U14170 (N_14170,N_10734,N_11430);
nor U14171 (N_14171,N_9411,N_10145);
nor U14172 (N_14172,N_11508,N_9778);
nand U14173 (N_14173,N_10093,N_9393);
nor U14174 (N_14174,N_11628,N_9870);
nor U14175 (N_14175,N_10649,N_11145);
or U14176 (N_14176,N_9871,N_9297);
and U14177 (N_14177,N_9084,N_9264);
nor U14178 (N_14178,N_10833,N_11467);
nand U14179 (N_14179,N_10585,N_11168);
and U14180 (N_14180,N_10133,N_11096);
nand U14181 (N_14181,N_11598,N_9118);
and U14182 (N_14182,N_9003,N_11960);
and U14183 (N_14183,N_10200,N_9220);
nand U14184 (N_14184,N_11932,N_10597);
or U14185 (N_14185,N_9385,N_9059);
nand U14186 (N_14186,N_9404,N_9524);
and U14187 (N_14187,N_9092,N_9965);
and U14188 (N_14188,N_11658,N_11361);
nor U14189 (N_14189,N_11642,N_10827);
nand U14190 (N_14190,N_11655,N_9313);
and U14191 (N_14191,N_11033,N_11787);
nand U14192 (N_14192,N_11760,N_9742);
and U14193 (N_14193,N_11998,N_10247);
nor U14194 (N_14194,N_10351,N_11062);
nor U14195 (N_14195,N_11975,N_11571);
nand U14196 (N_14196,N_11991,N_11985);
nor U14197 (N_14197,N_9051,N_10008);
and U14198 (N_14198,N_11567,N_11495);
and U14199 (N_14199,N_9619,N_10276);
and U14200 (N_14200,N_11523,N_11263);
or U14201 (N_14201,N_9831,N_9876);
or U14202 (N_14202,N_9691,N_11354);
nor U14203 (N_14203,N_10976,N_11481);
nand U14204 (N_14204,N_9185,N_11384);
nor U14205 (N_14205,N_10479,N_9618);
or U14206 (N_14206,N_9362,N_11572);
and U14207 (N_14207,N_11403,N_10520);
and U14208 (N_14208,N_9065,N_10762);
and U14209 (N_14209,N_10237,N_9532);
nor U14210 (N_14210,N_10694,N_10050);
nor U14211 (N_14211,N_9144,N_10851);
or U14212 (N_14212,N_9143,N_9607);
and U14213 (N_14213,N_9054,N_11994);
nand U14214 (N_14214,N_10168,N_10714);
or U14215 (N_14215,N_10428,N_11208);
and U14216 (N_14216,N_11200,N_11666);
nor U14217 (N_14217,N_11798,N_9265);
nand U14218 (N_14218,N_9390,N_10568);
or U14219 (N_14219,N_10765,N_9045);
or U14220 (N_14220,N_11993,N_10127);
and U14221 (N_14221,N_10180,N_9942);
nor U14222 (N_14222,N_11699,N_11601);
or U14223 (N_14223,N_10899,N_10849);
nor U14224 (N_14224,N_10745,N_10276);
nor U14225 (N_14225,N_10504,N_10617);
or U14226 (N_14226,N_11764,N_10024);
nand U14227 (N_14227,N_9863,N_9284);
and U14228 (N_14228,N_10309,N_9032);
and U14229 (N_14229,N_11069,N_10921);
and U14230 (N_14230,N_11322,N_11603);
nand U14231 (N_14231,N_10843,N_9854);
nand U14232 (N_14232,N_11913,N_9510);
nor U14233 (N_14233,N_11892,N_11379);
and U14234 (N_14234,N_10091,N_9970);
and U14235 (N_14235,N_11994,N_10319);
nand U14236 (N_14236,N_9328,N_9921);
and U14237 (N_14237,N_9122,N_11434);
and U14238 (N_14238,N_9414,N_10837);
nand U14239 (N_14239,N_10167,N_9893);
or U14240 (N_14240,N_10431,N_11622);
and U14241 (N_14241,N_10717,N_9059);
and U14242 (N_14242,N_9261,N_9683);
or U14243 (N_14243,N_10715,N_10652);
nand U14244 (N_14244,N_11467,N_9138);
nor U14245 (N_14245,N_9211,N_11827);
and U14246 (N_14246,N_10559,N_9323);
nor U14247 (N_14247,N_10241,N_9664);
and U14248 (N_14248,N_9130,N_10141);
nor U14249 (N_14249,N_10015,N_11481);
and U14250 (N_14250,N_9562,N_9320);
nor U14251 (N_14251,N_11835,N_11792);
and U14252 (N_14252,N_9153,N_11160);
and U14253 (N_14253,N_11526,N_10361);
or U14254 (N_14254,N_10557,N_10811);
or U14255 (N_14255,N_11521,N_10650);
and U14256 (N_14256,N_9814,N_9618);
nor U14257 (N_14257,N_10720,N_10853);
and U14258 (N_14258,N_10564,N_10700);
and U14259 (N_14259,N_10340,N_9427);
nor U14260 (N_14260,N_9093,N_10026);
nand U14261 (N_14261,N_10543,N_9822);
nand U14262 (N_14262,N_9657,N_9405);
nor U14263 (N_14263,N_11053,N_10856);
or U14264 (N_14264,N_9359,N_10538);
and U14265 (N_14265,N_10519,N_11182);
and U14266 (N_14266,N_11706,N_10117);
nand U14267 (N_14267,N_11248,N_10378);
nor U14268 (N_14268,N_10185,N_9068);
nor U14269 (N_14269,N_9671,N_9148);
or U14270 (N_14270,N_11240,N_10646);
nor U14271 (N_14271,N_11045,N_10612);
or U14272 (N_14272,N_9070,N_9703);
and U14273 (N_14273,N_9926,N_9147);
or U14274 (N_14274,N_10823,N_9859);
nor U14275 (N_14275,N_11121,N_11871);
xnor U14276 (N_14276,N_9207,N_9587);
and U14277 (N_14277,N_9523,N_10146);
and U14278 (N_14278,N_9527,N_11184);
nand U14279 (N_14279,N_10316,N_10736);
and U14280 (N_14280,N_9305,N_9654);
and U14281 (N_14281,N_9942,N_9191);
nand U14282 (N_14282,N_10697,N_10278);
nand U14283 (N_14283,N_11232,N_10353);
and U14284 (N_14284,N_9442,N_10729);
nand U14285 (N_14285,N_10869,N_9756);
nor U14286 (N_14286,N_11808,N_10517);
and U14287 (N_14287,N_10279,N_11955);
and U14288 (N_14288,N_11079,N_10193);
nor U14289 (N_14289,N_11327,N_9978);
xnor U14290 (N_14290,N_10494,N_10402);
nor U14291 (N_14291,N_11816,N_9647);
nor U14292 (N_14292,N_11781,N_9418);
or U14293 (N_14293,N_9868,N_11943);
or U14294 (N_14294,N_10981,N_10458);
or U14295 (N_14295,N_11755,N_9790);
nand U14296 (N_14296,N_10513,N_10691);
nand U14297 (N_14297,N_11155,N_10642);
or U14298 (N_14298,N_11119,N_9225);
nor U14299 (N_14299,N_11497,N_10858);
nand U14300 (N_14300,N_9395,N_11603);
or U14301 (N_14301,N_11225,N_9472);
and U14302 (N_14302,N_11535,N_11449);
nor U14303 (N_14303,N_11714,N_10759);
nor U14304 (N_14304,N_9015,N_9338);
or U14305 (N_14305,N_11147,N_9706);
and U14306 (N_14306,N_9852,N_10892);
and U14307 (N_14307,N_11074,N_9731);
nand U14308 (N_14308,N_11159,N_9601);
or U14309 (N_14309,N_10439,N_10495);
and U14310 (N_14310,N_9043,N_9809);
xor U14311 (N_14311,N_10260,N_10838);
and U14312 (N_14312,N_9600,N_10369);
and U14313 (N_14313,N_9762,N_11991);
and U14314 (N_14314,N_10800,N_10276);
or U14315 (N_14315,N_9928,N_9793);
nand U14316 (N_14316,N_9962,N_11145);
nand U14317 (N_14317,N_9118,N_11609);
and U14318 (N_14318,N_11918,N_11865);
nor U14319 (N_14319,N_10519,N_10181);
and U14320 (N_14320,N_9359,N_11222);
and U14321 (N_14321,N_11121,N_10429);
and U14322 (N_14322,N_11347,N_9460);
nor U14323 (N_14323,N_11208,N_11738);
or U14324 (N_14324,N_9766,N_11427);
and U14325 (N_14325,N_11810,N_9566);
nor U14326 (N_14326,N_11900,N_11969);
or U14327 (N_14327,N_9066,N_11196);
or U14328 (N_14328,N_10557,N_11230);
and U14329 (N_14329,N_10297,N_11536);
xor U14330 (N_14330,N_10718,N_11971);
or U14331 (N_14331,N_11910,N_9609);
or U14332 (N_14332,N_11930,N_10403);
or U14333 (N_14333,N_11865,N_9536);
nor U14334 (N_14334,N_11895,N_9126);
nor U14335 (N_14335,N_11802,N_9030);
and U14336 (N_14336,N_9662,N_9702);
nor U14337 (N_14337,N_9019,N_9274);
nor U14338 (N_14338,N_9184,N_9309);
nor U14339 (N_14339,N_9220,N_10659);
nand U14340 (N_14340,N_9953,N_11817);
nand U14341 (N_14341,N_10361,N_9269);
nor U14342 (N_14342,N_11587,N_9758);
and U14343 (N_14343,N_10284,N_10439);
nor U14344 (N_14344,N_11823,N_10633);
and U14345 (N_14345,N_9607,N_9638);
and U14346 (N_14346,N_11725,N_9187);
or U14347 (N_14347,N_11760,N_11947);
nor U14348 (N_14348,N_9519,N_10826);
or U14349 (N_14349,N_11830,N_10184);
or U14350 (N_14350,N_9192,N_10731);
and U14351 (N_14351,N_9833,N_10039);
nand U14352 (N_14352,N_11816,N_9534);
or U14353 (N_14353,N_10618,N_11753);
nor U14354 (N_14354,N_11409,N_11529);
nand U14355 (N_14355,N_11338,N_11576);
or U14356 (N_14356,N_10609,N_9839);
or U14357 (N_14357,N_11168,N_11239);
nor U14358 (N_14358,N_11452,N_11610);
or U14359 (N_14359,N_9747,N_11142);
and U14360 (N_14360,N_9831,N_9273);
xor U14361 (N_14361,N_11384,N_9139);
and U14362 (N_14362,N_11288,N_9720);
or U14363 (N_14363,N_9272,N_10413);
or U14364 (N_14364,N_11157,N_9047);
or U14365 (N_14365,N_10065,N_11563);
and U14366 (N_14366,N_9576,N_10574);
or U14367 (N_14367,N_11366,N_9111);
nor U14368 (N_14368,N_11126,N_9967);
nand U14369 (N_14369,N_10877,N_11957);
nand U14370 (N_14370,N_9059,N_11606);
or U14371 (N_14371,N_10163,N_10354);
and U14372 (N_14372,N_9175,N_10089);
xnor U14373 (N_14373,N_11705,N_11185);
nand U14374 (N_14374,N_11560,N_10813);
and U14375 (N_14375,N_9957,N_10970);
and U14376 (N_14376,N_11912,N_9468);
nand U14377 (N_14377,N_9927,N_9601);
and U14378 (N_14378,N_11608,N_11242);
or U14379 (N_14379,N_9388,N_10367);
nor U14380 (N_14380,N_11519,N_10516);
or U14381 (N_14381,N_10514,N_9040);
and U14382 (N_14382,N_10716,N_11626);
and U14383 (N_14383,N_10788,N_9683);
nand U14384 (N_14384,N_9406,N_9575);
nand U14385 (N_14385,N_11945,N_9296);
and U14386 (N_14386,N_11439,N_10066);
nand U14387 (N_14387,N_10773,N_9354);
nand U14388 (N_14388,N_9871,N_9735);
nand U14389 (N_14389,N_11310,N_11339);
and U14390 (N_14390,N_11710,N_11700);
or U14391 (N_14391,N_9231,N_10601);
nor U14392 (N_14392,N_10254,N_9871);
nor U14393 (N_14393,N_11751,N_11701);
and U14394 (N_14394,N_9566,N_9364);
nand U14395 (N_14395,N_11232,N_10677);
or U14396 (N_14396,N_11787,N_10375);
or U14397 (N_14397,N_9728,N_11188);
nor U14398 (N_14398,N_10542,N_9381);
or U14399 (N_14399,N_10890,N_9043);
or U14400 (N_14400,N_10589,N_11902);
or U14401 (N_14401,N_9270,N_11439);
and U14402 (N_14402,N_10292,N_10221);
or U14403 (N_14403,N_11018,N_10945);
nand U14404 (N_14404,N_9555,N_10569);
nand U14405 (N_14405,N_9145,N_11842);
nor U14406 (N_14406,N_9471,N_11326);
and U14407 (N_14407,N_9594,N_9886);
nand U14408 (N_14408,N_10401,N_9115);
nand U14409 (N_14409,N_9331,N_11785);
nand U14410 (N_14410,N_10846,N_9595);
or U14411 (N_14411,N_10510,N_9286);
or U14412 (N_14412,N_11641,N_9936);
or U14413 (N_14413,N_10267,N_11986);
or U14414 (N_14414,N_10780,N_11013);
nand U14415 (N_14415,N_10239,N_11048);
nand U14416 (N_14416,N_10527,N_11637);
nand U14417 (N_14417,N_9848,N_9857);
nand U14418 (N_14418,N_11160,N_9514);
and U14419 (N_14419,N_10185,N_11550);
nand U14420 (N_14420,N_10138,N_11336);
or U14421 (N_14421,N_10239,N_11569);
xor U14422 (N_14422,N_11633,N_9548);
or U14423 (N_14423,N_9164,N_10008);
and U14424 (N_14424,N_9329,N_10826);
or U14425 (N_14425,N_9354,N_9365);
nor U14426 (N_14426,N_9898,N_10552);
and U14427 (N_14427,N_10918,N_9487);
or U14428 (N_14428,N_11698,N_9554);
or U14429 (N_14429,N_10777,N_9236);
and U14430 (N_14430,N_9980,N_11219);
nor U14431 (N_14431,N_11441,N_10704);
and U14432 (N_14432,N_9683,N_11353);
nor U14433 (N_14433,N_10067,N_10875);
nor U14434 (N_14434,N_10087,N_10905);
nand U14435 (N_14435,N_9990,N_9012);
or U14436 (N_14436,N_9412,N_11784);
or U14437 (N_14437,N_9873,N_10308);
nand U14438 (N_14438,N_9503,N_10412);
or U14439 (N_14439,N_9247,N_9709);
or U14440 (N_14440,N_9311,N_11074);
nor U14441 (N_14441,N_10917,N_9975);
and U14442 (N_14442,N_10942,N_10062);
and U14443 (N_14443,N_11842,N_10155);
or U14444 (N_14444,N_9303,N_11221);
or U14445 (N_14445,N_11628,N_9637);
nand U14446 (N_14446,N_9103,N_11067);
nor U14447 (N_14447,N_9799,N_9746);
or U14448 (N_14448,N_9728,N_11621);
or U14449 (N_14449,N_10316,N_9583);
and U14450 (N_14450,N_10566,N_11471);
nand U14451 (N_14451,N_9449,N_9191);
nand U14452 (N_14452,N_10790,N_10113);
xor U14453 (N_14453,N_11301,N_10689);
nand U14454 (N_14454,N_11691,N_10471);
nand U14455 (N_14455,N_9535,N_11131);
nor U14456 (N_14456,N_9487,N_11590);
and U14457 (N_14457,N_11610,N_11456);
and U14458 (N_14458,N_9920,N_10215);
nor U14459 (N_14459,N_10089,N_11763);
and U14460 (N_14460,N_11497,N_9646);
or U14461 (N_14461,N_11193,N_9662);
and U14462 (N_14462,N_11509,N_9544);
and U14463 (N_14463,N_11183,N_10242);
and U14464 (N_14464,N_9693,N_11431);
nor U14465 (N_14465,N_10709,N_11640);
nand U14466 (N_14466,N_9819,N_11026);
nor U14467 (N_14467,N_9553,N_10203);
or U14468 (N_14468,N_10795,N_10283);
or U14469 (N_14469,N_10018,N_11972);
or U14470 (N_14470,N_11146,N_9169);
nor U14471 (N_14471,N_9984,N_9760);
nand U14472 (N_14472,N_9295,N_11685);
and U14473 (N_14473,N_9663,N_10967);
nand U14474 (N_14474,N_11713,N_11817);
nand U14475 (N_14475,N_11326,N_11364);
nand U14476 (N_14476,N_11623,N_11970);
nand U14477 (N_14477,N_9736,N_10297);
nor U14478 (N_14478,N_11088,N_11851);
nor U14479 (N_14479,N_10781,N_11811);
xor U14480 (N_14480,N_10234,N_9604);
and U14481 (N_14481,N_9046,N_11505);
nand U14482 (N_14482,N_11109,N_9111);
and U14483 (N_14483,N_9586,N_11643);
or U14484 (N_14484,N_9217,N_10498);
and U14485 (N_14485,N_9190,N_9186);
nor U14486 (N_14486,N_9276,N_11016);
and U14487 (N_14487,N_9116,N_10175);
nor U14488 (N_14488,N_11340,N_9800);
and U14489 (N_14489,N_10750,N_11101);
and U14490 (N_14490,N_10737,N_11041);
nand U14491 (N_14491,N_11746,N_9116);
nand U14492 (N_14492,N_9010,N_10036);
or U14493 (N_14493,N_11238,N_11414);
nor U14494 (N_14494,N_11140,N_10413);
nand U14495 (N_14495,N_9690,N_11825);
and U14496 (N_14496,N_9676,N_11839);
nand U14497 (N_14497,N_11066,N_9572);
or U14498 (N_14498,N_11019,N_9074);
and U14499 (N_14499,N_11223,N_10671);
xnor U14500 (N_14500,N_10701,N_10123);
nor U14501 (N_14501,N_9046,N_11673);
and U14502 (N_14502,N_10572,N_11229);
nor U14503 (N_14503,N_10773,N_9800);
nand U14504 (N_14504,N_11341,N_9446);
nor U14505 (N_14505,N_10796,N_10311);
and U14506 (N_14506,N_11448,N_9921);
or U14507 (N_14507,N_10560,N_9244);
nand U14508 (N_14508,N_11265,N_10831);
or U14509 (N_14509,N_11987,N_10090);
nor U14510 (N_14510,N_9053,N_9385);
nor U14511 (N_14511,N_9843,N_11420);
nor U14512 (N_14512,N_9816,N_11465);
or U14513 (N_14513,N_10823,N_9467);
or U14514 (N_14514,N_11657,N_10558);
nand U14515 (N_14515,N_10039,N_11505);
nand U14516 (N_14516,N_11552,N_10538);
nand U14517 (N_14517,N_10641,N_10807);
or U14518 (N_14518,N_11068,N_10473);
or U14519 (N_14519,N_10787,N_10078);
or U14520 (N_14520,N_9277,N_11090);
nor U14521 (N_14521,N_11963,N_10072);
nand U14522 (N_14522,N_10771,N_9827);
nor U14523 (N_14523,N_11768,N_9615);
and U14524 (N_14524,N_9594,N_10452);
nand U14525 (N_14525,N_11842,N_10597);
or U14526 (N_14526,N_11037,N_11167);
and U14527 (N_14527,N_11095,N_10733);
nand U14528 (N_14528,N_9414,N_9742);
or U14529 (N_14529,N_10021,N_10019);
nand U14530 (N_14530,N_9776,N_9756);
nor U14531 (N_14531,N_11736,N_9978);
nand U14532 (N_14532,N_9995,N_9374);
and U14533 (N_14533,N_11463,N_10933);
nand U14534 (N_14534,N_10718,N_10681);
and U14535 (N_14535,N_11253,N_10014);
nor U14536 (N_14536,N_9284,N_10660);
and U14537 (N_14537,N_11714,N_10576);
nor U14538 (N_14538,N_10094,N_11357);
or U14539 (N_14539,N_10619,N_11913);
xor U14540 (N_14540,N_11851,N_9215);
and U14541 (N_14541,N_9908,N_9240);
nor U14542 (N_14542,N_11387,N_10158);
or U14543 (N_14543,N_9994,N_9414);
xnor U14544 (N_14544,N_10167,N_9152);
and U14545 (N_14545,N_10665,N_10049);
and U14546 (N_14546,N_10959,N_10637);
nand U14547 (N_14547,N_11563,N_10583);
nor U14548 (N_14548,N_10219,N_11640);
nand U14549 (N_14549,N_9011,N_9954);
and U14550 (N_14550,N_9452,N_10509);
and U14551 (N_14551,N_9132,N_11668);
nand U14552 (N_14552,N_9376,N_9615);
or U14553 (N_14553,N_10816,N_9224);
or U14554 (N_14554,N_9705,N_11893);
nor U14555 (N_14555,N_11008,N_11954);
nor U14556 (N_14556,N_11330,N_9859);
nor U14557 (N_14557,N_10365,N_9745);
nor U14558 (N_14558,N_10667,N_11874);
nor U14559 (N_14559,N_11140,N_10184);
nand U14560 (N_14560,N_9922,N_9631);
nand U14561 (N_14561,N_9139,N_10526);
nand U14562 (N_14562,N_10945,N_10337);
or U14563 (N_14563,N_11212,N_9306);
and U14564 (N_14564,N_9569,N_10734);
nor U14565 (N_14565,N_10998,N_10378);
nand U14566 (N_14566,N_9729,N_10009);
and U14567 (N_14567,N_9454,N_10444);
xor U14568 (N_14568,N_9115,N_9505);
and U14569 (N_14569,N_11699,N_11060);
or U14570 (N_14570,N_10862,N_10070);
or U14571 (N_14571,N_10337,N_9916);
or U14572 (N_14572,N_9777,N_9899);
nand U14573 (N_14573,N_10177,N_9585);
nand U14574 (N_14574,N_10289,N_11441);
nand U14575 (N_14575,N_11285,N_10444);
or U14576 (N_14576,N_11934,N_10414);
nor U14577 (N_14577,N_9089,N_11330);
xor U14578 (N_14578,N_11145,N_11576);
nand U14579 (N_14579,N_11447,N_9578);
nand U14580 (N_14580,N_10103,N_9463);
and U14581 (N_14581,N_10763,N_9475);
xor U14582 (N_14582,N_11957,N_9838);
nor U14583 (N_14583,N_11659,N_11018);
or U14584 (N_14584,N_9684,N_11721);
or U14585 (N_14585,N_10234,N_11084);
nor U14586 (N_14586,N_10127,N_11418);
nor U14587 (N_14587,N_9364,N_10131);
and U14588 (N_14588,N_11376,N_10429);
or U14589 (N_14589,N_11033,N_11604);
and U14590 (N_14590,N_10773,N_10647);
nor U14591 (N_14591,N_9913,N_9071);
or U14592 (N_14592,N_9657,N_9975);
and U14593 (N_14593,N_9559,N_10673);
and U14594 (N_14594,N_10516,N_11347);
nor U14595 (N_14595,N_10321,N_10001);
nor U14596 (N_14596,N_9357,N_10784);
nor U14597 (N_14597,N_11502,N_11054);
and U14598 (N_14598,N_10543,N_11862);
nor U14599 (N_14599,N_10360,N_11842);
nor U14600 (N_14600,N_9084,N_9410);
and U14601 (N_14601,N_9149,N_10886);
or U14602 (N_14602,N_10478,N_9566);
nor U14603 (N_14603,N_10011,N_9531);
or U14604 (N_14604,N_9465,N_9609);
or U14605 (N_14605,N_11011,N_9980);
and U14606 (N_14606,N_11909,N_9457);
nand U14607 (N_14607,N_9420,N_10263);
nand U14608 (N_14608,N_11763,N_11758);
xnor U14609 (N_14609,N_11753,N_10055);
nor U14610 (N_14610,N_10354,N_9979);
nor U14611 (N_14611,N_11671,N_10223);
and U14612 (N_14612,N_10649,N_9182);
nor U14613 (N_14613,N_9782,N_10302);
and U14614 (N_14614,N_9059,N_9036);
nor U14615 (N_14615,N_10184,N_9758);
or U14616 (N_14616,N_9530,N_9414);
or U14617 (N_14617,N_11980,N_11548);
or U14618 (N_14618,N_11500,N_10281);
nor U14619 (N_14619,N_11183,N_10038);
and U14620 (N_14620,N_10366,N_9425);
nor U14621 (N_14621,N_9379,N_10460);
and U14622 (N_14622,N_9432,N_9318);
nor U14623 (N_14623,N_10617,N_11499);
or U14624 (N_14624,N_10738,N_9998);
nor U14625 (N_14625,N_9301,N_9948);
or U14626 (N_14626,N_10503,N_10569);
nand U14627 (N_14627,N_9552,N_11437);
nand U14628 (N_14628,N_9958,N_11032);
and U14629 (N_14629,N_10309,N_9907);
nor U14630 (N_14630,N_11061,N_11075);
or U14631 (N_14631,N_10843,N_11971);
nand U14632 (N_14632,N_10269,N_10174);
nand U14633 (N_14633,N_11592,N_10414);
and U14634 (N_14634,N_10617,N_10137);
nor U14635 (N_14635,N_9979,N_10389);
or U14636 (N_14636,N_10559,N_11702);
nand U14637 (N_14637,N_11212,N_9062);
nand U14638 (N_14638,N_10108,N_10506);
nor U14639 (N_14639,N_10044,N_10610);
nor U14640 (N_14640,N_11327,N_10272);
or U14641 (N_14641,N_11089,N_11300);
nand U14642 (N_14642,N_9753,N_10192);
nor U14643 (N_14643,N_9527,N_11061);
nand U14644 (N_14644,N_9198,N_11018);
nand U14645 (N_14645,N_11904,N_10036);
nand U14646 (N_14646,N_9053,N_10702);
nand U14647 (N_14647,N_9076,N_9617);
xor U14648 (N_14648,N_11943,N_11682);
or U14649 (N_14649,N_9094,N_11543);
and U14650 (N_14650,N_11394,N_11865);
nand U14651 (N_14651,N_10958,N_11259);
and U14652 (N_14652,N_9419,N_11502);
nor U14653 (N_14653,N_10576,N_10747);
or U14654 (N_14654,N_11695,N_10058);
nand U14655 (N_14655,N_11507,N_9199);
and U14656 (N_14656,N_9869,N_11995);
or U14657 (N_14657,N_11852,N_9677);
nor U14658 (N_14658,N_9119,N_9502);
nor U14659 (N_14659,N_11322,N_10954);
nor U14660 (N_14660,N_9445,N_11622);
nor U14661 (N_14661,N_11170,N_9965);
and U14662 (N_14662,N_10023,N_9338);
or U14663 (N_14663,N_10915,N_9038);
nand U14664 (N_14664,N_10649,N_10019);
nor U14665 (N_14665,N_9922,N_11290);
nand U14666 (N_14666,N_11110,N_10039);
or U14667 (N_14667,N_9315,N_10544);
or U14668 (N_14668,N_9551,N_9100);
or U14669 (N_14669,N_9148,N_10818);
nor U14670 (N_14670,N_10298,N_11663);
and U14671 (N_14671,N_11964,N_10745);
nand U14672 (N_14672,N_11167,N_9178);
or U14673 (N_14673,N_10834,N_11337);
and U14674 (N_14674,N_9811,N_9681);
xor U14675 (N_14675,N_9073,N_10674);
or U14676 (N_14676,N_9672,N_11412);
or U14677 (N_14677,N_11450,N_9503);
nor U14678 (N_14678,N_10599,N_10004);
nor U14679 (N_14679,N_11406,N_10716);
or U14680 (N_14680,N_10602,N_10527);
or U14681 (N_14681,N_11754,N_9327);
xnor U14682 (N_14682,N_9107,N_10206);
nand U14683 (N_14683,N_11532,N_10389);
nand U14684 (N_14684,N_11979,N_10633);
or U14685 (N_14685,N_11765,N_9734);
nor U14686 (N_14686,N_11755,N_11676);
nor U14687 (N_14687,N_9431,N_11313);
nand U14688 (N_14688,N_11433,N_10911);
and U14689 (N_14689,N_9059,N_10754);
nand U14690 (N_14690,N_9482,N_9928);
nor U14691 (N_14691,N_11041,N_9854);
nand U14692 (N_14692,N_10881,N_11577);
and U14693 (N_14693,N_9464,N_11940);
or U14694 (N_14694,N_11158,N_11406);
nor U14695 (N_14695,N_9727,N_11850);
or U14696 (N_14696,N_10308,N_9629);
nand U14697 (N_14697,N_10303,N_11764);
and U14698 (N_14698,N_9610,N_11073);
nor U14699 (N_14699,N_11434,N_10654);
nor U14700 (N_14700,N_10223,N_9973);
and U14701 (N_14701,N_9618,N_11107);
nor U14702 (N_14702,N_11046,N_9264);
nor U14703 (N_14703,N_9117,N_9507);
nor U14704 (N_14704,N_10947,N_10864);
or U14705 (N_14705,N_11050,N_10727);
xnor U14706 (N_14706,N_11411,N_11078);
nor U14707 (N_14707,N_10788,N_9993);
nor U14708 (N_14708,N_9124,N_9333);
or U14709 (N_14709,N_11332,N_11985);
or U14710 (N_14710,N_10960,N_11304);
or U14711 (N_14711,N_10505,N_11321);
or U14712 (N_14712,N_9266,N_10016);
or U14713 (N_14713,N_10410,N_11630);
nand U14714 (N_14714,N_9910,N_10016);
or U14715 (N_14715,N_11461,N_9733);
nor U14716 (N_14716,N_10200,N_10622);
or U14717 (N_14717,N_9289,N_11281);
or U14718 (N_14718,N_9861,N_11187);
and U14719 (N_14719,N_11286,N_11969);
nand U14720 (N_14720,N_11725,N_10739);
or U14721 (N_14721,N_10212,N_11192);
and U14722 (N_14722,N_11056,N_10938);
nor U14723 (N_14723,N_11265,N_9055);
xnor U14724 (N_14724,N_9594,N_10688);
nand U14725 (N_14725,N_9164,N_10534);
and U14726 (N_14726,N_10163,N_11460);
nand U14727 (N_14727,N_9804,N_10560);
or U14728 (N_14728,N_9667,N_10157);
or U14729 (N_14729,N_9919,N_11799);
nand U14730 (N_14730,N_10024,N_11696);
and U14731 (N_14731,N_9089,N_9152);
nor U14732 (N_14732,N_10645,N_11385);
and U14733 (N_14733,N_11835,N_10050);
or U14734 (N_14734,N_10858,N_11440);
and U14735 (N_14735,N_10911,N_10796);
or U14736 (N_14736,N_9045,N_10884);
nor U14737 (N_14737,N_10894,N_10149);
nor U14738 (N_14738,N_9383,N_9764);
or U14739 (N_14739,N_9691,N_9703);
or U14740 (N_14740,N_10740,N_9838);
nand U14741 (N_14741,N_10414,N_11350);
nand U14742 (N_14742,N_9311,N_9694);
nor U14743 (N_14743,N_9428,N_9292);
or U14744 (N_14744,N_9554,N_10311);
nor U14745 (N_14745,N_10524,N_9472);
nor U14746 (N_14746,N_9012,N_10419);
or U14747 (N_14747,N_9533,N_9201);
or U14748 (N_14748,N_10024,N_11144);
nand U14749 (N_14749,N_10616,N_9561);
or U14750 (N_14750,N_11738,N_11844);
nor U14751 (N_14751,N_9784,N_10710);
nor U14752 (N_14752,N_10402,N_10476);
and U14753 (N_14753,N_11140,N_11956);
nor U14754 (N_14754,N_9656,N_10686);
nand U14755 (N_14755,N_11025,N_10793);
nand U14756 (N_14756,N_10884,N_10569);
nor U14757 (N_14757,N_10345,N_9989);
or U14758 (N_14758,N_11704,N_11927);
and U14759 (N_14759,N_10910,N_10216);
xor U14760 (N_14760,N_10504,N_9564);
nand U14761 (N_14761,N_11322,N_10250);
or U14762 (N_14762,N_9310,N_9169);
and U14763 (N_14763,N_9441,N_9849);
nand U14764 (N_14764,N_10072,N_10782);
nor U14765 (N_14765,N_9311,N_10587);
or U14766 (N_14766,N_10695,N_11503);
xor U14767 (N_14767,N_9832,N_11145);
nand U14768 (N_14768,N_11626,N_11243);
nand U14769 (N_14769,N_9201,N_11281);
and U14770 (N_14770,N_9367,N_11173);
or U14771 (N_14771,N_11674,N_11103);
and U14772 (N_14772,N_9826,N_11027);
nand U14773 (N_14773,N_11824,N_10771);
nor U14774 (N_14774,N_10350,N_10950);
nor U14775 (N_14775,N_11747,N_9357);
nor U14776 (N_14776,N_10308,N_11601);
and U14777 (N_14777,N_10378,N_9534);
nor U14778 (N_14778,N_11258,N_11761);
and U14779 (N_14779,N_11410,N_10222);
nor U14780 (N_14780,N_10494,N_10776);
and U14781 (N_14781,N_9831,N_9585);
and U14782 (N_14782,N_9933,N_11852);
and U14783 (N_14783,N_9534,N_11793);
and U14784 (N_14784,N_10397,N_11626);
and U14785 (N_14785,N_11644,N_11720);
nand U14786 (N_14786,N_11527,N_11709);
and U14787 (N_14787,N_11788,N_11048);
nor U14788 (N_14788,N_10034,N_10407);
or U14789 (N_14789,N_11307,N_9264);
or U14790 (N_14790,N_11054,N_11907);
or U14791 (N_14791,N_10897,N_10808);
and U14792 (N_14792,N_11517,N_11146);
and U14793 (N_14793,N_9400,N_11183);
or U14794 (N_14794,N_9077,N_9125);
nand U14795 (N_14795,N_11460,N_9827);
nor U14796 (N_14796,N_10381,N_9634);
or U14797 (N_14797,N_11079,N_9685);
and U14798 (N_14798,N_10006,N_10110);
or U14799 (N_14799,N_10957,N_10038);
nor U14800 (N_14800,N_10409,N_10361);
nand U14801 (N_14801,N_10462,N_11145);
nand U14802 (N_14802,N_11686,N_9520);
and U14803 (N_14803,N_10010,N_9664);
or U14804 (N_14804,N_10094,N_11027);
and U14805 (N_14805,N_10000,N_9595);
or U14806 (N_14806,N_10927,N_10322);
nand U14807 (N_14807,N_10451,N_10537);
nand U14808 (N_14808,N_9190,N_9045);
nor U14809 (N_14809,N_10848,N_10647);
nand U14810 (N_14810,N_11541,N_10502);
nor U14811 (N_14811,N_11638,N_9156);
xnor U14812 (N_14812,N_11223,N_10573);
nand U14813 (N_14813,N_10842,N_11670);
nor U14814 (N_14814,N_11328,N_10312);
xnor U14815 (N_14815,N_10257,N_9811);
or U14816 (N_14816,N_11584,N_9323);
xnor U14817 (N_14817,N_11373,N_11528);
nand U14818 (N_14818,N_9411,N_10707);
nand U14819 (N_14819,N_9507,N_11937);
or U14820 (N_14820,N_11307,N_11332);
nand U14821 (N_14821,N_9147,N_11931);
or U14822 (N_14822,N_10022,N_11153);
nor U14823 (N_14823,N_11467,N_11548);
and U14824 (N_14824,N_10857,N_9980);
or U14825 (N_14825,N_9055,N_11150);
nor U14826 (N_14826,N_11960,N_10486);
nand U14827 (N_14827,N_11302,N_10696);
nand U14828 (N_14828,N_10163,N_9632);
nor U14829 (N_14829,N_10614,N_10578);
nand U14830 (N_14830,N_10265,N_11032);
and U14831 (N_14831,N_10864,N_11634);
or U14832 (N_14832,N_10935,N_10882);
nor U14833 (N_14833,N_9511,N_10739);
or U14834 (N_14834,N_10419,N_9224);
nor U14835 (N_14835,N_10175,N_11546);
or U14836 (N_14836,N_9381,N_11288);
or U14837 (N_14837,N_10082,N_9399);
or U14838 (N_14838,N_9559,N_11087);
or U14839 (N_14839,N_9410,N_11304);
and U14840 (N_14840,N_10222,N_10211);
or U14841 (N_14841,N_10668,N_11902);
nor U14842 (N_14842,N_11677,N_11150);
nor U14843 (N_14843,N_11581,N_11937);
nor U14844 (N_14844,N_10379,N_11457);
nand U14845 (N_14845,N_11656,N_11205);
or U14846 (N_14846,N_10677,N_11577);
nand U14847 (N_14847,N_11067,N_9048);
or U14848 (N_14848,N_9297,N_10816);
and U14849 (N_14849,N_10316,N_9339);
nand U14850 (N_14850,N_11669,N_9816);
or U14851 (N_14851,N_11256,N_10360);
and U14852 (N_14852,N_10128,N_10518);
nand U14853 (N_14853,N_11058,N_11402);
nand U14854 (N_14854,N_11922,N_10834);
nand U14855 (N_14855,N_11943,N_9342);
nor U14856 (N_14856,N_11285,N_10757);
nand U14857 (N_14857,N_11268,N_11361);
nand U14858 (N_14858,N_11372,N_9201);
nor U14859 (N_14859,N_10992,N_9537);
nor U14860 (N_14860,N_9679,N_10765);
or U14861 (N_14861,N_9530,N_9033);
nor U14862 (N_14862,N_11866,N_9017);
nor U14863 (N_14863,N_9590,N_11920);
nor U14864 (N_14864,N_11987,N_11448);
nor U14865 (N_14865,N_9378,N_10199);
nand U14866 (N_14866,N_10395,N_11449);
nor U14867 (N_14867,N_10031,N_10042);
nor U14868 (N_14868,N_11890,N_9076);
nor U14869 (N_14869,N_9624,N_9973);
or U14870 (N_14870,N_11102,N_9982);
and U14871 (N_14871,N_9427,N_9456);
and U14872 (N_14872,N_9206,N_10932);
and U14873 (N_14873,N_9138,N_10294);
or U14874 (N_14874,N_9754,N_10112);
nor U14875 (N_14875,N_9686,N_9002);
nor U14876 (N_14876,N_9680,N_11964);
and U14877 (N_14877,N_9143,N_9815);
or U14878 (N_14878,N_10061,N_9170);
nand U14879 (N_14879,N_10147,N_11783);
or U14880 (N_14880,N_11484,N_11810);
nor U14881 (N_14881,N_10388,N_10841);
nand U14882 (N_14882,N_9245,N_10781);
and U14883 (N_14883,N_10079,N_10919);
nor U14884 (N_14884,N_11481,N_9802);
and U14885 (N_14885,N_10638,N_9006);
or U14886 (N_14886,N_9590,N_11853);
nand U14887 (N_14887,N_9421,N_9275);
or U14888 (N_14888,N_11069,N_11218);
nor U14889 (N_14889,N_11593,N_9865);
nor U14890 (N_14890,N_10439,N_10253);
or U14891 (N_14891,N_10760,N_11630);
nand U14892 (N_14892,N_11652,N_11902);
and U14893 (N_14893,N_10136,N_10507);
and U14894 (N_14894,N_11289,N_10531);
nand U14895 (N_14895,N_9111,N_9916);
nand U14896 (N_14896,N_9870,N_11128);
and U14897 (N_14897,N_11847,N_11170);
or U14898 (N_14898,N_11833,N_9593);
nand U14899 (N_14899,N_11745,N_11720);
or U14900 (N_14900,N_10925,N_9884);
or U14901 (N_14901,N_9603,N_10402);
or U14902 (N_14902,N_9431,N_10714);
or U14903 (N_14903,N_9451,N_10705);
nand U14904 (N_14904,N_9655,N_9919);
or U14905 (N_14905,N_9492,N_9816);
nand U14906 (N_14906,N_10620,N_10140);
and U14907 (N_14907,N_9310,N_10886);
nand U14908 (N_14908,N_9210,N_9890);
nand U14909 (N_14909,N_10470,N_10808);
nor U14910 (N_14910,N_9011,N_9666);
nand U14911 (N_14911,N_9412,N_10607);
nor U14912 (N_14912,N_11841,N_10499);
and U14913 (N_14913,N_9564,N_9870);
or U14914 (N_14914,N_9202,N_10848);
nand U14915 (N_14915,N_10115,N_10800);
or U14916 (N_14916,N_9246,N_11934);
xor U14917 (N_14917,N_9655,N_10201);
nand U14918 (N_14918,N_11872,N_9128);
or U14919 (N_14919,N_11314,N_9532);
nor U14920 (N_14920,N_11876,N_9401);
or U14921 (N_14921,N_11244,N_11255);
nand U14922 (N_14922,N_11539,N_11522);
nand U14923 (N_14923,N_10875,N_10194);
and U14924 (N_14924,N_11776,N_10009);
nor U14925 (N_14925,N_9311,N_9394);
and U14926 (N_14926,N_11595,N_9052);
nand U14927 (N_14927,N_9563,N_9488);
or U14928 (N_14928,N_9109,N_11011);
and U14929 (N_14929,N_10561,N_10160);
or U14930 (N_14930,N_9698,N_9614);
and U14931 (N_14931,N_11616,N_11001);
nor U14932 (N_14932,N_10106,N_10174);
and U14933 (N_14933,N_11523,N_9078);
nand U14934 (N_14934,N_10195,N_9435);
or U14935 (N_14935,N_9564,N_10326);
nor U14936 (N_14936,N_11089,N_9159);
or U14937 (N_14937,N_11246,N_11671);
nand U14938 (N_14938,N_11860,N_11118);
or U14939 (N_14939,N_10915,N_10885);
nor U14940 (N_14940,N_11645,N_10097);
nand U14941 (N_14941,N_10398,N_9403);
nand U14942 (N_14942,N_11243,N_10643);
nand U14943 (N_14943,N_11727,N_10616);
nor U14944 (N_14944,N_10604,N_11020);
nand U14945 (N_14945,N_10856,N_11576);
and U14946 (N_14946,N_11063,N_10927);
or U14947 (N_14947,N_9201,N_11191);
or U14948 (N_14948,N_11187,N_10064);
or U14949 (N_14949,N_10454,N_10142);
and U14950 (N_14950,N_11121,N_11872);
nand U14951 (N_14951,N_9347,N_11333);
and U14952 (N_14952,N_10534,N_11241);
nor U14953 (N_14953,N_11744,N_11653);
nand U14954 (N_14954,N_9201,N_10264);
or U14955 (N_14955,N_9372,N_11488);
nand U14956 (N_14956,N_11404,N_11534);
and U14957 (N_14957,N_10331,N_11659);
and U14958 (N_14958,N_11330,N_10546);
and U14959 (N_14959,N_11328,N_10844);
nor U14960 (N_14960,N_11012,N_9045);
or U14961 (N_14961,N_10966,N_10792);
and U14962 (N_14962,N_9333,N_9740);
or U14963 (N_14963,N_10625,N_10209);
and U14964 (N_14964,N_11464,N_9069);
nand U14965 (N_14965,N_11550,N_9239);
nand U14966 (N_14966,N_10057,N_11286);
nand U14967 (N_14967,N_9923,N_9288);
nor U14968 (N_14968,N_9533,N_11297);
nor U14969 (N_14969,N_9383,N_10712);
and U14970 (N_14970,N_9378,N_9941);
or U14971 (N_14971,N_10289,N_9667);
nand U14972 (N_14972,N_9508,N_10088);
and U14973 (N_14973,N_9966,N_11024);
nor U14974 (N_14974,N_9196,N_11315);
or U14975 (N_14975,N_11350,N_10885);
and U14976 (N_14976,N_11148,N_9610);
nor U14977 (N_14977,N_11603,N_9356);
nor U14978 (N_14978,N_11053,N_10894);
and U14979 (N_14979,N_10899,N_10770);
and U14980 (N_14980,N_10918,N_11166);
or U14981 (N_14981,N_10526,N_9626);
nor U14982 (N_14982,N_9982,N_9769);
xor U14983 (N_14983,N_10707,N_10489);
or U14984 (N_14984,N_11233,N_10866);
and U14985 (N_14985,N_9680,N_9420);
nor U14986 (N_14986,N_9869,N_11564);
nand U14987 (N_14987,N_9266,N_9926);
nor U14988 (N_14988,N_10852,N_11166);
nor U14989 (N_14989,N_9495,N_11846);
nand U14990 (N_14990,N_11532,N_9474);
or U14991 (N_14991,N_11454,N_9330);
or U14992 (N_14992,N_11024,N_11459);
or U14993 (N_14993,N_11429,N_10723);
nor U14994 (N_14994,N_9827,N_11212);
nand U14995 (N_14995,N_11847,N_10961);
or U14996 (N_14996,N_11520,N_10069);
xor U14997 (N_14997,N_11203,N_9904);
or U14998 (N_14998,N_10397,N_9881);
and U14999 (N_14999,N_9535,N_9035);
and UO_0 (O_0,N_13660,N_12526);
and UO_1 (O_1,N_13295,N_14005);
nor UO_2 (O_2,N_14194,N_12497);
nand UO_3 (O_3,N_13484,N_12429);
and UO_4 (O_4,N_13069,N_13753);
or UO_5 (O_5,N_14956,N_14546);
nand UO_6 (O_6,N_12600,N_12758);
and UO_7 (O_7,N_14171,N_13692);
and UO_8 (O_8,N_12752,N_12495);
nor UO_9 (O_9,N_12264,N_12473);
and UO_10 (O_10,N_13280,N_12990);
nand UO_11 (O_11,N_13306,N_12289);
or UO_12 (O_12,N_14053,N_14148);
nand UO_13 (O_13,N_14300,N_12901);
nand UO_14 (O_14,N_13812,N_14353);
nand UO_15 (O_15,N_13234,N_13841);
nand UO_16 (O_16,N_14963,N_13767);
nand UO_17 (O_17,N_12207,N_12824);
or UO_18 (O_18,N_14891,N_14478);
nand UO_19 (O_19,N_12970,N_14422);
and UO_20 (O_20,N_14816,N_14346);
and UO_21 (O_21,N_12946,N_12193);
or UO_22 (O_22,N_12565,N_13070);
or UO_23 (O_23,N_14312,N_13560);
nor UO_24 (O_24,N_14611,N_12195);
or UO_25 (O_25,N_12118,N_13723);
and UO_26 (O_26,N_13887,N_12548);
nor UO_27 (O_27,N_12988,N_12062);
nor UO_28 (O_28,N_14810,N_13419);
nor UO_29 (O_29,N_13770,N_12575);
and UO_30 (O_30,N_13957,N_12808);
nor UO_31 (O_31,N_13495,N_12408);
nor UO_32 (O_32,N_12254,N_13130);
nor UO_33 (O_33,N_12219,N_14225);
and UO_34 (O_34,N_14626,N_13607);
or UO_35 (O_35,N_14561,N_13864);
nor UO_36 (O_36,N_13141,N_14117);
or UO_37 (O_37,N_13305,N_12609);
nor UO_38 (O_38,N_13489,N_14511);
nand UO_39 (O_39,N_12623,N_14771);
nand UO_40 (O_40,N_13014,N_13639);
and UO_41 (O_41,N_12120,N_13885);
or UO_42 (O_42,N_13217,N_14720);
nor UO_43 (O_43,N_12542,N_13325);
or UO_44 (O_44,N_14282,N_13226);
or UO_45 (O_45,N_14766,N_14387);
nand UO_46 (O_46,N_14994,N_14877);
and UO_47 (O_47,N_13566,N_12535);
or UO_48 (O_48,N_14083,N_13974);
nand UO_49 (O_49,N_14157,N_13010);
or UO_50 (O_50,N_12248,N_12260);
or UO_51 (O_51,N_13463,N_12133);
nand UO_52 (O_52,N_13046,N_12371);
nand UO_53 (O_53,N_12330,N_12423);
and UO_54 (O_54,N_13834,N_12868);
and UO_55 (O_55,N_14285,N_13034);
and UO_56 (O_56,N_13703,N_14125);
nand UO_57 (O_57,N_13230,N_13430);
and UO_58 (O_58,N_14883,N_12262);
nor UO_59 (O_59,N_13371,N_13162);
or UO_60 (O_60,N_14698,N_13365);
nand UO_61 (O_61,N_13921,N_14999);
or UO_62 (O_62,N_12259,N_12279);
nand UO_63 (O_63,N_14678,N_13129);
nor UO_64 (O_64,N_14719,N_12387);
or UO_65 (O_65,N_12492,N_14376);
nor UO_66 (O_66,N_14703,N_13643);
or UO_67 (O_67,N_12555,N_13867);
nand UO_68 (O_68,N_12945,N_13188);
nand UO_69 (O_69,N_12521,N_12991);
nand UO_70 (O_70,N_14863,N_13412);
nand UO_71 (O_71,N_13232,N_13790);
nor UO_72 (O_72,N_13003,N_14978);
and UO_73 (O_73,N_13299,N_14428);
and UO_74 (O_74,N_14363,N_14645);
or UO_75 (O_75,N_12577,N_12759);
or UO_76 (O_76,N_14872,N_12063);
nor UO_77 (O_77,N_13916,N_13826);
or UO_78 (O_78,N_13737,N_12782);
and UO_79 (O_79,N_14648,N_13939);
nand UO_80 (O_80,N_12208,N_12415);
xnor UO_81 (O_81,N_12608,N_13460);
nor UO_82 (O_82,N_13238,N_14458);
nor UO_83 (O_83,N_13761,N_12618);
nand UO_84 (O_84,N_12559,N_13290);
nand UO_85 (O_85,N_12541,N_13282);
nand UO_86 (O_86,N_14651,N_13661);
nand UO_87 (O_87,N_14588,N_12652);
nand UO_88 (O_88,N_12926,N_14178);
and UO_89 (O_89,N_12728,N_13652);
nor UO_90 (O_90,N_13634,N_12144);
nand UO_91 (O_91,N_12220,N_14276);
and UO_92 (O_92,N_14841,N_13387);
nand UO_93 (O_93,N_13145,N_12392);
or UO_94 (O_94,N_13592,N_13549);
and UO_95 (O_95,N_12523,N_12885);
nor UO_96 (O_96,N_13699,N_12880);
or UO_97 (O_97,N_13385,N_14525);
and UO_98 (O_98,N_14093,N_12238);
nor UO_99 (O_99,N_14094,N_14708);
xor UO_100 (O_100,N_14682,N_14560);
nand UO_101 (O_101,N_13468,N_14340);
and UO_102 (O_102,N_14038,N_14201);
xnor UO_103 (O_103,N_14949,N_13138);
nor UO_104 (O_104,N_12490,N_12025);
or UO_105 (O_105,N_13391,N_12230);
nand UO_106 (O_106,N_14523,N_14076);
nor UO_107 (O_107,N_14239,N_14031);
nand UO_108 (O_108,N_14254,N_12723);
or UO_109 (O_109,N_13808,N_13646);
and UO_110 (O_110,N_12302,N_14538);
and UO_111 (O_111,N_13722,N_13236);
or UO_112 (O_112,N_13392,N_14928);
and UO_113 (O_113,N_12560,N_13688);
or UO_114 (O_114,N_14008,N_14074);
nor UO_115 (O_115,N_13399,N_13594);
nand UO_116 (O_116,N_14494,N_14914);
and UO_117 (O_117,N_12750,N_13576);
nor UO_118 (O_118,N_12757,N_12378);
nand UO_119 (O_119,N_14469,N_14836);
nor UO_120 (O_120,N_13390,N_13860);
nand UO_121 (O_121,N_13383,N_14144);
or UO_122 (O_122,N_14137,N_12682);
xnor UO_123 (O_123,N_13076,N_14025);
nand UO_124 (O_124,N_13814,N_14681);
or UO_125 (O_125,N_14334,N_13479);
nand UO_126 (O_126,N_14327,N_12200);
xnor UO_127 (O_127,N_14654,N_12727);
or UO_128 (O_128,N_12799,N_14447);
nand UO_129 (O_129,N_12903,N_12742);
nor UO_130 (O_130,N_14871,N_12068);
and UO_131 (O_131,N_14461,N_12593);
nor UO_132 (O_132,N_14542,N_12566);
nand UO_133 (O_133,N_14236,N_12232);
or UO_134 (O_134,N_14661,N_13871);
and UO_135 (O_135,N_13769,N_13529);
xor UO_136 (O_136,N_14266,N_13298);
and UO_137 (O_137,N_14187,N_12852);
or UO_138 (O_138,N_13410,N_12810);
nand UO_139 (O_139,N_14901,N_12530);
nor UO_140 (O_140,N_13423,N_14910);
nor UO_141 (O_141,N_12563,N_13323);
nand UO_142 (O_142,N_13984,N_14037);
and UO_143 (O_143,N_13552,N_14641);
or UO_144 (O_144,N_14233,N_12453);
and UO_145 (O_145,N_14255,N_13047);
nand UO_146 (O_146,N_13296,N_14826);
nor UO_147 (O_147,N_14058,N_13170);
or UO_148 (O_148,N_14180,N_13820);
nand UO_149 (O_149,N_14457,N_13959);
and UO_150 (O_150,N_14289,N_12338);
or UO_151 (O_151,N_14106,N_14183);
nand UO_152 (O_152,N_13114,N_12962);
nand UO_153 (O_153,N_14134,N_12909);
or UO_154 (O_154,N_12224,N_12849);
or UO_155 (O_155,N_12659,N_14691);
or UO_156 (O_156,N_13096,N_13177);
nand UO_157 (O_157,N_13839,N_14534);
or UO_158 (O_158,N_14436,N_13263);
nand UO_159 (O_159,N_12143,N_12165);
nand UO_160 (O_160,N_13568,N_12536);
nand UO_161 (O_161,N_13376,N_14398);
nor UO_162 (O_162,N_14294,N_12212);
nor UO_163 (O_163,N_12789,N_12813);
or UO_164 (O_164,N_13780,N_14393);
or UO_165 (O_165,N_14743,N_14551);
xnor UO_166 (O_166,N_13085,N_12518);
nor UO_167 (O_167,N_14834,N_12983);
or UO_168 (O_168,N_14092,N_12053);
and UO_169 (O_169,N_12633,N_14499);
or UO_170 (O_170,N_13478,N_13264);
or UO_171 (O_171,N_14895,N_12491);
and UO_172 (O_172,N_14045,N_14797);
and UO_173 (O_173,N_14563,N_12639);
and UO_174 (O_174,N_12681,N_14403);
nand UO_175 (O_175,N_12456,N_12009);
and UO_176 (O_176,N_13697,N_13173);
or UO_177 (O_177,N_14659,N_14330);
or UO_178 (O_178,N_14596,N_14578);
nand UO_179 (O_179,N_12930,N_13992);
nor UO_180 (O_180,N_14411,N_14988);
and UO_181 (O_181,N_13740,N_13797);
and UO_182 (O_182,N_13905,N_14251);
nand UO_183 (O_183,N_12817,N_12936);
nor UO_184 (O_184,N_13098,N_12596);
or UO_185 (O_185,N_12240,N_13935);
and UO_186 (O_186,N_13513,N_14192);
and UO_187 (O_187,N_14380,N_13159);
and UO_188 (O_188,N_13459,N_13933);
nor UO_189 (O_189,N_14317,N_12046);
and UO_190 (O_190,N_12890,N_13176);
nor UO_191 (O_191,N_13150,N_14166);
and UO_192 (O_192,N_14685,N_13061);
or UO_193 (O_193,N_13635,N_14077);
and UO_194 (O_194,N_12142,N_14302);
and UO_195 (O_195,N_14498,N_13791);
nor UO_196 (O_196,N_13906,N_13185);
and UO_197 (O_197,N_12434,N_13914);
and UO_198 (O_198,N_13406,N_14684);
or UO_199 (O_199,N_14989,N_13804);
or UO_200 (O_200,N_14822,N_13457);
nand UO_201 (O_201,N_12999,N_12617);
nor UO_202 (O_202,N_13848,N_14026);
or UO_203 (O_203,N_12549,N_13413);
nor UO_204 (O_204,N_12987,N_12251);
nor UO_205 (O_205,N_13408,N_14196);
xnor UO_206 (O_206,N_14765,N_12614);
nor UO_207 (O_207,N_12801,N_13626);
nand UO_208 (O_208,N_12672,N_14540);
or UO_209 (O_209,N_13755,N_14814);
or UO_210 (O_210,N_13875,N_12329);
nand UO_211 (O_211,N_13800,N_14524);
or UO_212 (O_212,N_14844,N_12018);
nor UO_213 (O_213,N_13564,N_14604);
and UO_214 (O_214,N_12222,N_12601);
and UO_215 (O_215,N_13710,N_12496);
nand UO_216 (O_216,N_12398,N_14042);
or UO_217 (O_217,N_12942,N_14227);
nand UO_218 (O_218,N_14492,N_14853);
nor UO_219 (O_219,N_12964,N_13899);
and UO_220 (O_220,N_14761,N_14627);
or UO_221 (O_221,N_12627,N_14435);
nor UO_222 (O_222,N_13094,N_14549);
nor UO_223 (O_223,N_12380,N_14991);
and UO_224 (O_224,N_13053,N_14177);
and UO_225 (O_225,N_14869,N_14198);
nand UO_226 (O_226,N_13971,N_13718);
or UO_227 (O_227,N_12404,N_14679);
nor UO_228 (O_228,N_12564,N_13680);
nor UO_229 (O_229,N_13343,N_14262);
nand UO_230 (O_230,N_12997,N_14906);
nand UO_231 (O_231,N_13544,N_13977);
or UO_232 (O_232,N_14516,N_12960);
nor UO_233 (O_233,N_13813,N_13895);
nand UO_234 (O_234,N_13996,N_14636);
or UO_235 (O_235,N_12873,N_14060);
and UO_236 (O_236,N_14655,N_13008);
or UO_237 (O_237,N_12865,N_13907);
nor UO_238 (O_238,N_14874,N_14305);
and UO_239 (O_239,N_12592,N_13553);
or UO_240 (O_240,N_13980,N_14013);
nor UO_241 (O_241,N_14557,N_13714);
or UO_242 (O_242,N_13494,N_13036);
nor UO_243 (O_243,N_14114,N_14326);
and UO_244 (O_244,N_12707,N_13190);
nand UO_245 (O_245,N_12694,N_12961);
and UO_246 (O_246,N_14120,N_12335);
or UO_247 (O_247,N_13949,N_12011);
or UO_248 (O_248,N_14406,N_13677);
and UO_249 (O_249,N_13026,N_14948);
or UO_250 (O_250,N_12129,N_13208);
nand UO_251 (O_251,N_12275,N_13458);
nand UO_252 (O_252,N_14905,N_14760);
or UO_253 (O_253,N_13222,N_14472);
xnor UO_254 (O_254,N_13614,N_13080);
and UO_255 (O_255,N_14209,N_13777);
xor UO_256 (O_256,N_13128,N_14342);
nand UO_257 (O_257,N_14056,N_13912);
nor UO_258 (O_258,N_13218,N_14974);
nor UO_259 (O_259,N_14858,N_12414);
and UO_260 (O_260,N_14344,N_13055);
or UO_261 (O_261,N_13951,N_12000);
nand UO_262 (O_262,N_12459,N_13449);
or UO_263 (O_263,N_13429,N_13726);
and UO_264 (O_264,N_13893,N_12569);
or UO_265 (O_265,N_13774,N_14307);
nand UO_266 (O_266,N_13338,N_13588);
and UO_267 (O_267,N_14271,N_14744);
nor UO_268 (O_268,N_13171,N_12911);
nor UO_269 (O_269,N_14287,N_13013);
nor UO_270 (O_270,N_13843,N_13806);
nand UO_271 (O_271,N_13934,N_12151);
or UO_272 (O_272,N_12074,N_12699);
and UO_273 (O_273,N_12236,N_14202);
xor UO_274 (O_274,N_13133,N_12493);
nand UO_275 (O_275,N_12696,N_12692);
or UO_276 (O_276,N_12583,N_12020);
nor UO_277 (O_277,N_14371,N_13354);
and UO_278 (O_278,N_12695,N_14532);
nor UO_279 (O_279,N_12171,N_12393);
nor UO_280 (O_280,N_14559,N_13397);
and UO_281 (O_281,N_12673,N_14799);
nand UO_282 (O_282,N_14405,N_13438);
or UO_283 (O_283,N_14800,N_14543);
nor UO_284 (O_284,N_12540,N_14264);
xor UO_285 (O_285,N_14351,N_13653);
or UO_286 (O_286,N_12933,N_12572);
nand UO_287 (O_287,N_13702,N_12571);
and UO_288 (O_288,N_13088,N_12920);
and UO_289 (O_289,N_12858,N_14426);
nand UO_290 (O_290,N_14146,N_12202);
nand UO_291 (O_291,N_14859,N_12927);
or UO_292 (O_292,N_13411,N_12993);
nor UO_293 (O_293,N_14935,N_13771);
and UO_294 (O_294,N_12267,N_12738);
and UO_295 (O_295,N_13486,N_12221);
nor UO_296 (O_296,N_13727,N_13369);
and UO_297 (O_297,N_14709,N_14163);
or UO_298 (O_298,N_12114,N_14851);
nor UO_299 (O_299,N_13382,N_13361);
nand UO_300 (O_300,N_13712,N_14213);
and UO_301 (O_301,N_14860,N_12288);
nor UO_302 (O_302,N_14848,N_12625);
nor UO_303 (O_303,N_12745,N_12800);
and UO_304 (O_304,N_12538,N_12095);
nand UO_305 (O_305,N_14133,N_14795);
or UO_306 (O_306,N_12377,N_13203);
or UO_307 (O_307,N_13874,N_14211);
and UO_308 (O_308,N_12029,N_14983);
and UO_309 (O_309,N_14637,N_12857);
nand UO_310 (O_310,N_12989,N_14712);
nand UO_311 (O_311,N_14984,N_14442);
nor UO_312 (O_312,N_12741,N_13291);
nor UO_313 (O_313,N_13572,N_12923);
and UO_314 (O_314,N_13346,N_14110);
or UO_315 (O_315,N_12359,N_13969);
or UO_316 (O_316,N_13545,N_12823);
and UO_317 (O_317,N_13273,N_12110);
or UO_318 (O_318,N_13084,N_13816);
and UO_319 (O_319,N_13968,N_13890);
nor UO_320 (O_320,N_14181,N_12109);
and UO_321 (O_321,N_13310,N_13243);
or UO_322 (O_322,N_12273,N_13829);
nand UO_323 (O_323,N_13157,N_14047);
or UO_324 (O_324,N_12635,N_13204);
and UO_325 (O_325,N_12159,N_12767);
and UO_326 (O_326,N_13415,N_14129);
nor UO_327 (O_327,N_12904,N_12894);
or UO_328 (O_328,N_13444,N_13628);
nor UO_329 (O_329,N_13311,N_13002);
or UO_330 (O_330,N_13464,N_12995);
nor UO_331 (O_331,N_12096,N_13798);
or UO_332 (O_332,N_12299,N_13043);
nor UO_333 (O_333,N_12594,N_14812);
nand UO_334 (O_334,N_12950,N_13897);
nand UO_335 (O_335,N_12021,N_12528);
or UO_336 (O_336,N_13695,N_14382);
nor UO_337 (O_337,N_12051,N_13929);
nor UO_338 (O_338,N_14268,N_12715);
nor UO_339 (O_339,N_13372,N_13858);
or UO_340 (O_340,N_12486,N_12186);
or UO_341 (O_341,N_14040,N_14752);
and UO_342 (O_342,N_14899,N_12401);
nand UO_343 (O_343,N_13876,N_14855);
and UO_344 (O_344,N_14642,N_13551);
or UO_345 (O_345,N_12442,N_12086);
and UO_346 (O_346,N_12014,N_12336);
and UO_347 (O_347,N_13825,N_14575);
or UO_348 (O_348,N_13083,N_12550);
and UO_349 (O_349,N_14950,N_14758);
nor UO_350 (O_350,N_12725,N_13453);
and UO_351 (O_351,N_12313,N_12947);
nand UO_352 (O_352,N_12140,N_14606);
or UO_353 (O_353,N_14616,N_12737);
or UO_354 (O_354,N_12937,N_12113);
xnor UO_355 (O_355,N_14238,N_14452);
or UO_356 (O_356,N_13579,N_12155);
nand UO_357 (O_357,N_12718,N_13878);
or UO_358 (O_358,N_14904,N_13904);
and UO_359 (O_359,N_12843,N_12515);
xor UO_360 (O_360,N_13888,N_14833);
nand UO_361 (O_361,N_13152,N_14222);
or UO_362 (O_362,N_14728,N_14441);
and UO_363 (O_363,N_14212,N_14937);
and UO_364 (O_364,N_13042,N_13577);
nand UO_365 (O_365,N_14861,N_12866);
nor UO_366 (O_366,N_12355,N_12644);
nand UO_367 (O_367,N_14624,N_13331);
nor UO_368 (O_368,N_14842,N_13743);
nand UO_369 (O_369,N_14257,N_12658);
nor UO_370 (O_370,N_12877,N_12134);
nand UO_371 (O_371,N_12056,N_12726);
nand UO_372 (O_372,N_12705,N_12048);
nand UO_373 (O_373,N_13117,N_13180);
or UO_374 (O_374,N_14017,N_14725);
nand UO_375 (O_375,N_14359,N_12024);
nor UO_376 (O_376,N_13001,N_13401);
nand UO_377 (O_377,N_14296,N_14065);
or UO_378 (O_378,N_13927,N_14818);
nand UO_379 (O_379,N_13642,N_13210);
nor UO_380 (O_380,N_13105,N_14383);
and UO_381 (O_381,N_12765,N_14701);
nand UO_382 (O_382,N_13242,N_14581);
nor UO_383 (O_383,N_14666,N_13450);
and UO_384 (O_384,N_14357,N_12498);
and UO_385 (O_385,N_12116,N_14558);
and UO_386 (O_386,N_12520,N_12588);
or UO_387 (O_387,N_12931,N_12245);
and UO_388 (O_388,N_13960,N_14135);
nor UO_389 (O_389,N_12331,N_12769);
or UO_390 (O_390,N_12512,N_12590);
nor UO_391 (O_391,N_12478,N_12557);
nor UO_392 (O_392,N_13742,N_12882);
nand UO_393 (O_393,N_14769,N_13099);
and UO_394 (O_394,N_13955,N_13616);
nor UO_395 (O_395,N_13670,N_12318);
nor UO_396 (O_396,N_13507,N_12973);
or UO_397 (O_397,N_13694,N_12869);
xnor UO_398 (O_398,N_12332,N_12848);
nand UO_399 (O_399,N_12756,N_12735);
and UO_400 (O_400,N_13474,N_14787);
nand UO_401 (O_401,N_14235,N_14061);
or UO_402 (O_402,N_14495,N_12788);
or UO_403 (O_403,N_13973,N_13198);
and UO_404 (O_404,N_13095,N_14656);
or UO_405 (O_405,N_14052,N_13448);
nand UO_406 (O_406,N_12284,N_12959);
nor UO_407 (O_407,N_13562,N_13075);
nor UO_408 (O_408,N_14004,N_13205);
xnor UO_409 (O_409,N_13821,N_13368);
or UO_410 (O_410,N_13582,N_13400);
nor UO_411 (O_411,N_13414,N_14857);
or UO_412 (O_412,N_12704,N_12485);
or UO_413 (O_413,N_12345,N_14805);
or UO_414 (O_414,N_12762,N_14884);
or UO_415 (O_415,N_14786,N_12624);
nor UO_416 (O_416,N_13490,N_12851);
and UO_417 (O_417,N_14951,N_13522);
nand UO_418 (O_418,N_12832,N_12712);
nand UO_419 (O_419,N_14622,N_13669);
and UO_420 (O_420,N_12465,N_12666);
or UO_421 (O_421,N_14780,N_12397);
nand UO_422 (O_422,N_12806,N_13528);
and UO_423 (O_423,N_13689,N_12509);
nand UO_424 (O_424,N_14808,N_14085);
or UO_425 (O_425,N_14729,N_13881);
or UO_426 (O_426,N_14530,N_14754);
nor UO_427 (O_427,N_13667,N_13751);
nand UO_428 (O_428,N_13941,N_12416);
nor UO_429 (O_429,N_14349,N_13297);
nand UO_430 (O_430,N_14308,N_13279);
and UO_431 (O_431,N_12561,N_14484);
nand UO_432 (O_432,N_13758,N_13764);
or UO_433 (O_433,N_14158,N_14205);
nand UO_434 (O_434,N_14281,N_13165);
and UO_435 (O_435,N_14594,N_12483);
nor UO_436 (O_436,N_13902,N_12087);
nor UO_437 (O_437,N_13735,N_12304);
or UO_438 (O_438,N_13765,N_12527);
nand UO_439 (O_439,N_13097,N_14152);
or UO_440 (O_440,N_14550,N_13163);
or UO_441 (O_441,N_13597,N_13747);
or UO_442 (O_442,N_12778,N_14782);
and UO_443 (O_443,N_13750,N_14621);
or UO_444 (O_444,N_12427,N_13212);
and UO_445 (O_445,N_13420,N_12435);
nor UO_446 (O_446,N_13533,N_12437);
or UO_447 (O_447,N_14136,N_12383);
and UO_448 (O_448,N_12733,N_14942);
nand UO_449 (O_449,N_12117,N_14714);
or UO_450 (O_450,N_13025,N_12676);
or UO_451 (O_451,N_12754,N_12833);
nand UO_452 (O_452,N_14773,N_12237);
nand UO_453 (O_453,N_14630,N_14612);
nor UO_454 (O_454,N_12686,N_14062);
and UO_455 (O_455,N_12821,N_14223);
nand UO_456 (O_456,N_14587,N_14726);
or UO_457 (O_457,N_12119,N_13213);
and UO_458 (O_458,N_13684,N_12785);
nor UO_459 (O_459,N_12104,N_14759);
or UO_460 (O_460,N_13776,N_13144);
and UO_461 (O_461,N_14700,N_13051);
or UO_462 (O_462,N_13989,N_12949);
and UO_463 (O_463,N_12261,N_14938);
or UO_464 (O_464,N_12286,N_14420);
nand UO_465 (O_465,N_12123,N_14595);
nor UO_466 (O_466,N_13455,N_12385);
nand UO_467 (O_467,N_13550,N_12711);
and UO_468 (O_468,N_12255,N_13987);
or UO_469 (O_469,N_14030,N_13235);
nand UO_470 (O_470,N_13557,N_12090);
or UO_471 (O_471,N_13831,N_13779);
or UO_472 (O_472,N_12215,N_12085);
nor UO_473 (O_473,N_14794,N_14921);
and UO_474 (O_474,N_12534,N_14444);
nand UO_475 (O_475,N_12154,N_14835);
or UO_476 (O_476,N_12276,N_13155);
nor UO_477 (O_477,N_13883,N_12182);
nor UO_478 (O_478,N_13106,N_13501);
or UO_479 (O_479,N_12668,N_14482);
xor UO_480 (O_480,N_14735,N_13828);
nor UO_481 (O_481,N_13865,N_12337);
and UO_482 (O_482,N_12481,N_12402);
nor UO_483 (O_483,N_12524,N_13174);
nand UO_484 (O_484,N_13854,N_12305);
nor UO_485 (O_485,N_12729,N_14510);
and UO_486 (O_486,N_13351,N_12316);
or UO_487 (O_487,N_12910,N_12266);
or UO_488 (O_488,N_14897,N_12131);
nor UO_489 (O_489,N_14274,N_12854);
nand UO_490 (O_490,N_14241,N_13108);
or UO_491 (O_491,N_14035,N_13972);
nand UO_492 (O_492,N_14480,N_12010);
nand UO_493 (O_493,N_14509,N_13074);
nand UO_494 (O_494,N_14699,N_13530);
and UO_495 (O_495,N_14090,N_13915);
or UO_496 (O_496,N_13793,N_14896);
and UO_497 (O_497,N_13100,N_14506);
and UO_498 (O_498,N_14041,N_13134);
or UO_499 (O_499,N_14502,N_13123);
and UO_500 (O_500,N_13250,N_14690);
and UO_501 (O_501,N_13313,N_13649);
xnor UO_502 (O_502,N_14710,N_12158);
nand UO_503 (O_503,N_14977,N_14926);
nand UO_504 (O_504,N_13148,N_13062);
nor UO_505 (O_505,N_12688,N_13169);
or UO_506 (O_506,N_14845,N_14089);
nor UO_507 (O_507,N_12399,N_12653);
or UO_508 (O_508,N_13598,N_14936);
or UO_509 (O_509,N_14221,N_12791);
nand UO_510 (O_510,N_12683,N_12184);
nor UO_511 (O_511,N_14454,N_13621);
or UO_512 (O_512,N_12640,N_14068);
nand UO_513 (O_513,N_13645,N_12282);
or UO_514 (O_514,N_12457,N_13064);
nor UO_515 (O_515,N_13345,N_12145);
or UO_516 (O_516,N_12407,N_13307);
nand UO_517 (O_517,N_14903,N_13956);
or UO_518 (O_518,N_14341,N_12736);
and UO_519 (O_519,N_12722,N_12657);
nand UO_520 (O_520,N_12678,N_14547);
nor UO_521 (O_521,N_14500,N_14731);
and UO_522 (O_522,N_14039,N_12700);
nand UO_523 (O_523,N_14629,N_14643);
and UO_524 (O_524,N_12709,N_14096);
and UO_525 (O_525,N_12343,N_12774);
and UO_526 (O_526,N_12773,N_14356);
and UO_527 (O_527,N_12844,N_14464);
or UO_528 (O_528,N_14693,N_14172);
nor UO_529 (O_529,N_12629,N_13832);
and UO_530 (O_530,N_13254,N_13830);
and UO_531 (O_531,N_13518,N_12400);
and UO_532 (O_532,N_13581,N_14190);
nor UO_533 (O_533,N_13452,N_14807);
nor UO_534 (O_534,N_12646,N_12443);
and UO_535 (O_535,N_12779,N_13020);
or UO_536 (O_536,N_14483,N_12441);
nand UO_537 (O_537,N_14944,N_14751);
or UO_538 (O_538,N_14788,N_14811);
nand UO_539 (O_539,N_13216,N_13007);
nand UO_540 (O_540,N_12470,N_14508);
and UO_541 (O_541,N_13186,N_13471);
or UO_542 (O_542,N_14430,N_14695);
nand UO_543 (O_543,N_14980,N_13470);
or UO_544 (O_544,N_13436,N_13600);
or UO_545 (O_545,N_13112,N_14781);
or UO_546 (O_546,N_12772,N_14741);
and UO_547 (O_547,N_14465,N_14367);
nor UO_548 (O_548,N_13880,N_14019);
or UO_549 (O_549,N_12418,N_14003);
and UO_550 (O_550,N_13292,N_12980);
or UO_551 (O_551,N_14217,N_12231);
xnor UO_552 (O_552,N_13836,N_13179);
nand UO_553 (O_553,N_12645,N_13067);
xor UO_554 (O_554,N_13342,N_13251);
nor UO_555 (O_555,N_13000,N_13196);
nand UO_556 (O_556,N_14783,N_12553);
and UO_557 (O_557,N_14882,N_12032);
nand UO_558 (O_558,N_13807,N_13332);
or UO_559 (O_559,N_13066,N_13624);
nor UO_560 (O_560,N_14736,N_13659);
and UO_561 (O_561,N_14733,N_13195);
or UO_562 (O_562,N_13574,N_12023);
and UO_563 (O_563,N_14043,N_14939);
or UO_564 (O_564,N_12827,N_12748);
nor UO_565 (O_565,N_14467,N_13153);
and UO_566 (O_566,N_14071,N_12107);
and UO_567 (O_567,N_13432,N_14625);
nor UO_568 (O_568,N_13672,N_12693);
and UO_569 (O_569,N_14310,N_12507);
or UO_570 (O_570,N_14128,N_14108);
nor UO_571 (O_571,N_12522,N_13673);
nor UO_572 (O_572,N_14918,N_13244);
or UO_573 (O_573,N_14653,N_14311);
and UO_574 (O_574,N_12697,N_12420);
and UO_575 (O_575,N_14996,N_12615);
nand UO_576 (O_576,N_13149,N_13734);
xor UO_577 (O_577,N_13168,N_13241);
and UO_578 (O_578,N_13589,N_13884);
nand UO_579 (O_579,N_12544,N_12599);
nand UO_580 (O_580,N_13898,N_13850);
xor UO_581 (O_581,N_12296,N_12812);
or UO_582 (O_582,N_12619,N_14070);
nand UO_583 (O_583,N_12075,N_13328);
or UO_584 (O_584,N_13644,N_14474);
or UO_585 (O_585,N_13602,N_14569);
nand UO_586 (O_586,N_13559,N_13360);
nand UO_587 (O_587,N_13431,N_14941);
or UO_588 (O_588,N_14954,N_13433);
nor UO_589 (O_589,N_14421,N_14909);
nor UO_590 (O_590,N_13192,N_13315);
nor UO_591 (O_591,N_13610,N_14174);
or UO_592 (O_592,N_14732,N_13340);
and UO_593 (O_593,N_13838,N_12570);
or UO_594 (O_594,N_12034,N_12022);
and UO_595 (O_595,N_13037,N_13322);
and UO_596 (O_596,N_12390,N_13258);
or UO_597 (O_597,N_12822,N_14020);
nand UO_598 (O_598,N_14079,N_13056);
xnor UO_599 (O_599,N_14772,N_14553);
and UO_600 (O_600,N_12325,N_14001);
xor UO_601 (O_601,N_14730,N_13139);
or UO_602 (O_602,N_14111,N_13327);
or UO_603 (O_603,N_12862,N_13286);
or UO_604 (O_604,N_14409,N_14328);
nand UO_605 (O_605,N_14429,N_13146);
nand UO_606 (O_606,N_12992,N_14981);
xor UO_607 (O_607,N_14846,N_14424);
nand UO_608 (O_608,N_12341,N_12976);
nand UO_609 (O_609,N_13005,N_13394);
and UO_610 (O_610,N_13531,N_14431);
or UO_611 (O_611,N_13498,N_14246);
or UO_612 (O_612,N_12417,N_13543);
and UO_613 (O_613,N_14867,N_14652);
or UO_614 (O_614,N_13435,N_12846);
or UO_615 (O_615,N_12787,N_13833);
nand UO_616 (O_616,N_13508,N_12472);
nor UO_617 (O_617,N_14862,N_12545);
or UO_618 (O_618,N_13675,N_14838);
nand UO_619 (O_619,N_12743,N_14915);
and UO_620 (O_620,N_13454,N_12170);
and UO_621 (O_621,N_13795,N_13674);
or UO_622 (O_622,N_13082,N_12060);
nor UO_623 (O_623,N_14088,N_13405);
and UO_624 (O_624,N_13917,N_12939);
xor UO_625 (O_625,N_12744,N_14667);
nor UO_626 (O_626,N_12576,N_13161);
nor UO_627 (O_627,N_13294,N_12891);
nand UO_628 (O_628,N_12612,N_12631);
and UO_629 (O_629,N_14961,N_14348);
nor UO_630 (O_630,N_14737,N_13257);
and UO_631 (O_631,N_13439,N_14048);
nand UO_632 (O_632,N_13909,N_13632);
nor UO_633 (O_633,N_12647,N_13647);
nor UO_634 (O_634,N_13891,N_14024);
nand UO_635 (O_635,N_12396,N_14556);
nand UO_636 (O_636,N_14286,N_14138);
and UO_637 (O_637,N_13462,N_13936);
or UO_638 (O_638,N_12139,N_14375);
or UO_639 (O_639,N_12246,N_12746);
or UO_640 (O_640,N_14159,N_14658);
or UO_641 (O_641,N_13932,N_14162);
and UO_642 (O_642,N_14615,N_12146);
and UO_643 (O_643,N_13259,N_14063);
nor UO_644 (O_644,N_14668,N_13983);
nor UO_645 (O_645,N_12298,N_13931);
xor UO_646 (O_646,N_12256,N_12574);
or UO_647 (O_647,N_13719,N_14527);
nand UO_648 (O_648,N_12130,N_12469);
and UO_649 (O_649,N_12320,N_14477);
nor UO_650 (O_650,N_13503,N_14952);
nor UO_651 (O_651,N_12189,N_14628);
nor UO_652 (O_652,N_14601,N_14116);
and UO_653 (O_653,N_14945,N_13546);
and UO_654 (O_654,N_13260,N_13473);
nor UO_655 (O_655,N_12966,N_12050);
nor UO_656 (O_656,N_13116,N_12616);
nor UO_657 (O_657,N_14756,N_13536);
nor UO_658 (O_658,N_12606,N_14253);
nor UO_659 (O_659,N_12088,N_12176);
or UO_660 (O_660,N_12586,N_14554);
and UO_661 (O_661,N_13788,N_13679);
nor UO_662 (O_662,N_12838,N_13785);
nor UO_663 (O_663,N_12350,N_13604);
nor UO_664 (O_664,N_12227,N_12102);
nor UO_665 (O_665,N_12019,N_13613);
or UO_666 (O_666,N_12780,N_14505);
or UO_667 (O_667,N_12094,N_13154);
nor UO_668 (O_668,N_13089,N_13223);
nor UO_669 (O_669,N_14418,N_13525);
nand UO_670 (O_670,N_14433,N_14967);
nand UO_671 (O_671,N_14908,N_13640);
nand UO_672 (O_672,N_14107,N_12853);
nor UO_673 (O_673,N_14173,N_12306);
nor UO_674 (O_674,N_13285,N_12975);
or UO_675 (O_675,N_14318,N_14747);
or UO_676 (O_676,N_13749,N_13443);
nand UO_677 (O_677,N_12409,N_14248);
and UO_678 (O_678,N_13424,N_13252);
and UO_679 (O_679,N_12349,N_13946);
and UO_680 (O_680,N_12106,N_13754);
nor UO_681 (O_681,N_12043,N_14825);
nor UO_682 (O_682,N_12346,N_13827);
or UO_683 (O_683,N_12985,N_14131);
nor UO_684 (O_684,N_13009,N_13229);
nor UO_685 (O_685,N_12353,N_13608);
nand UO_686 (O_686,N_13300,N_13233);
nand UO_687 (O_687,N_12795,N_14432);
or UO_688 (O_688,N_14126,N_13961);
or UO_689 (O_689,N_13320,N_14191);
and UO_690 (O_690,N_12460,N_13118);
nand UO_691 (O_691,N_13447,N_14400);
nor UO_692 (O_692,N_13476,N_13851);
and UO_693 (O_693,N_12803,N_12505);
nor UO_694 (O_694,N_12183,N_14293);
nand UO_695 (O_695,N_12468,N_14054);
and UO_696 (O_696,N_12932,N_13206);
nor UO_697 (O_697,N_14168,N_13512);
nor UO_698 (O_698,N_14301,N_13500);
nor UO_699 (O_699,N_14219,N_12038);
nand UO_700 (O_700,N_13107,N_12137);
or UO_701 (O_701,N_14321,N_13491);
nor UO_702 (O_702,N_14369,N_14423);
nand UO_703 (O_703,N_14985,N_13011);
or UO_704 (O_704,N_14593,N_14571);
nor UO_705 (O_705,N_12938,N_12511);
nor UO_706 (O_706,N_12448,N_12953);
and UO_707 (O_707,N_12175,N_13965);
and UO_708 (O_708,N_12781,N_13261);
nor UO_709 (O_709,N_14032,N_14746);
or UO_710 (O_710,N_14689,N_14109);
nor UO_711 (O_711,N_14288,N_13981);
and UO_712 (O_712,N_13434,N_13802);
or UO_713 (O_713,N_14946,N_12876);
nand UO_714 (O_714,N_13416,N_13757);
nor UO_715 (O_715,N_13334,N_13181);
nor UO_716 (O_716,N_12214,N_12079);
or UO_717 (O_717,N_14396,N_12066);
nor UO_718 (O_718,N_12912,N_13587);
xor UO_719 (O_719,N_14459,N_13054);
and UO_720 (O_720,N_13132,N_13333);
nand UO_721 (O_721,N_12818,N_12105);
and UO_722 (O_722,N_14774,N_13569);
nor UO_723 (O_723,N_13789,N_13440);
xnor UO_724 (O_724,N_13759,N_14840);
nand UO_725 (O_725,N_14716,N_13184);
nand UO_726 (O_726,N_12792,N_14366);
and UO_727 (O_727,N_13337,N_12589);
nand UO_728 (O_728,N_13277,N_14609);
and UO_729 (O_729,N_13472,N_12467);
nand UO_730 (O_730,N_12917,N_14462);
nor UO_731 (O_731,N_12041,N_13606);
nand UO_732 (O_732,N_12831,N_13541);
nand UO_733 (O_733,N_12798,N_14493);
nor UO_734 (O_734,N_12297,N_12340);
and UO_735 (O_735,N_12840,N_14099);
or UO_736 (O_736,N_13738,N_13104);
nor UO_737 (O_737,N_14237,N_13926);
nor UO_738 (O_738,N_14879,N_12097);
and UO_739 (O_739,N_12516,N_12986);
nor UO_740 (O_740,N_12258,N_13685);
and UO_741 (O_741,N_14095,N_14907);
nor UO_742 (O_742,N_14603,N_12285);
nor UO_743 (O_743,N_14160,N_14446);
nand UO_744 (O_744,N_14304,N_13193);
nor UO_745 (O_745,N_14749,N_14320);
nor UO_746 (O_746,N_12956,N_13289);
and UO_747 (O_747,N_12091,N_14034);
nor UO_748 (O_748,N_13409,N_13609);
nand UO_749 (O_749,N_13304,N_13772);
or UO_750 (O_750,N_14990,N_12480);
nand UO_751 (O_751,N_12948,N_14303);
and UO_752 (O_752,N_14279,N_12552);
and UO_753 (O_753,N_14381,N_12764);
or UO_754 (O_754,N_13445,N_13136);
or UO_755 (O_755,N_12077,N_12166);
nand UO_756 (O_756,N_14269,N_12706);
and UO_757 (O_757,N_13923,N_13058);
nand UO_758 (O_758,N_13496,N_13822);
xor UO_759 (O_759,N_13732,N_12761);
and UO_760 (O_760,N_12027,N_12093);
nor UO_761 (O_761,N_13975,N_13676);
nor UO_762 (O_762,N_14837,N_13030);
nor UO_763 (O_763,N_12445,N_12364);
nand UO_764 (O_764,N_12136,N_14971);
or UO_765 (O_765,N_13514,N_14727);
nand UO_766 (O_766,N_14149,N_14112);
nor UO_767 (O_767,N_14583,N_12280);
or UO_768 (O_768,N_13156,N_12185);
or UO_769 (O_769,N_14982,N_14784);
nor UO_770 (O_770,N_14960,N_12368);
and UO_771 (O_771,N_14920,N_12887);
nor UO_772 (O_772,N_13121,N_12972);
or UO_773 (O_773,N_14831,N_14200);
nor UO_774 (O_774,N_13596,N_12598);
and UO_775 (O_775,N_13246,N_13783);
nand UO_776 (O_776,N_12430,N_14649);
nor UO_777 (O_777,N_14325,N_14998);
nand UO_778 (O_778,N_12169,N_14664);
nand UO_779 (O_779,N_14434,N_13985);
or UO_780 (O_780,N_14401,N_14992);
or UO_781 (O_781,N_12687,N_12875);
nand UO_782 (O_782,N_12287,N_13255);
nor UO_783 (O_783,N_14927,N_12979);
or UO_784 (O_784,N_14687,N_13301);
or UO_785 (O_785,N_13359,N_14449);
nor UO_786 (O_786,N_14101,N_14890);
or UO_787 (O_787,N_13668,N_14893);
and UO_788 (O_788,N_14723,N_13175);
xor UO_789 (O_789,N_14372,N_12874);
nand UO_790 (O_790,N_13319,N_14450);
nor UO_791 (O_791,N_12517,N_12126);
nand UO_792 (O_792,N_14460,N_12180);
or UO_793 (O_793,N_14574,N_14513);
nor UO_794 (O_794,N_13172,N_14384);
nand UO_795 (O_795,N_12819,N_14798);
and UO_796 (O_796,N_13815,N_12755);
nor UO_797 (O_797,N_13696,N_12651);
or UO_798 (O_798,N_12654,N_14979);
nor UO_799 (O_799,N_13272,N_14082);
nor UO_800 (O_800,N_13868,N_13077);
nand UO_801 (O_801,N_12229,N_14620);
nand UO_802 (O_802,N_13502,N_12026);
and UO_803 (O_803,N_12150,N_12573);
nor UO_804 (O_804,N_12749,N_14337);
nand UO_805 (O_805,N_12584,N_14002);
xor UO_806 (O_806,N_13681,N_13655);
nand UO_807 (O_807,N_12211,N_12253);
or UO_808 (O_808,N_13625,N_12499);
nand UO_809 (O_809,N_13705,N_12902);
and UO_810 (O_810,N_12815,N_12943);
and UO_811 (O_811,N_13823,N_13943);
nor UO_812 (O_812,N_12361,N_12978);
and UO_813 (O_813,N_13824,N_14394);
nand UO_814 (O_814,N_12076,N_12474);
nor UO_815 (O_815,N_13396,N_12602);
and UO_816 (O_816,N_13706,N_13584);
nor UO_817 (O_817,N_13752,N_14564);
or UO_818 (O_818,N_12015,N_13071);
nand UO_819 (O_819,N_13402,N_12698);
and UO_820 (O_820,N_12164,N_12049);
nor UO_821 (O_821,N_12081,N_14802);
nor UO_822 (O_822,N_12637,N_14817);
and UO_823 (O_823,N_13844,N_12213);
and UO_824 (O_824,N_14806,N_14154);
or UO_825 (O_825,N_12928,N_13485);
and UO_826 (O_826,N_12500,N_13182);
nor UO_827 (O_827,N_12872,N_13877);
or UO_828 (O_828,N_13335,N_12710);
nand UO_829 (O_829,N_14456,N_14419);
nor UO_830 (O_830,N_14657,N_12322);
xnor UO_831 (O_831,N_13027,N_12111);
nor UO_832 (O_832,N_12309,N_12099);
nand UO_833 (O_833,N_13633,N_12513);
and UO_834 (O_834,N_13641,N_12905);
nor UO_835 (O_835,N_14322,N_13330);
or UO_836 (O_836,N_12089,N_14000);
nand UO_837 (O_837,N_14352,N_14290);
nand UO_838 (O_838,N_13849,N_12065);
nand UO_839 (O_839,N_13995,N_12228);
or UO_840 (O_840,N_14228,N_14696);
and UO_841 (O_841,N_14329,N_12190);
or UO_842 (O_842,N_13511,N_14122);
nand UO_843 (O_843,N_13567,N_12008);
and UO_844 (O_844,N_12242,N_12719);
nand UO_845 (O_845,N_12845,N_12363);
or UO_846 (O_846,N_14912,N_13591);
or UO_847 (O_847,N_13925,N_12039);
or UO_848 (O_848,N_14229,N_14215);
or UO_849 (O_849,N_12157,N_14098);
nor UO_850 (O_850,N_13237,N_14663);
or UO_851 (O_851,N_12370,N_13922);
or UO_852 (O_852,N_14790,N_12971);
or UO_853 (O_853,N_13704,N_13663);
nor UO_854 (O_854,N_13889,N_12381);
xor UO_855 (O_855,N_14165,N_14930);
nand UO_856 (O_856,N_12895,N_12451);
and UO_857 (O_857,N_12580,N_13388);
or UO_858 (O_858,N_13142,N_13856);
or UO_859 (O_859,N_12354,N_13274);
nand UO_860 (O_860,N_14069,N_12770);
nand UO_861 (O_861,N_12045,N_12042);
nand UO_862 (O_862,N_13651,N_13215);
nand UO_863 (O_863,N_12103,N_13016);
and UO_864 (O_864,N_13720,N_12847);
and UO_865 (O_865,N_12249,N_14280);
nor UO_866 (O_866,N_13221,N_13638);
or UO_867 (O_867,N_12082,N_14335);
nand UO_868 (O_868,N_12127,N_13220);
nand UO_869 (O_869,N_13928,N_14244);
xor UO_870 (O_870,N_13381,N_14440);
or UO_871 (O_871,N_13708,N_13857);
nand UO_872 (O_872,N_13847,N_13748);
nor UO_873 (O_873,N_12784,N_13724);
nand UO_874 (O_874,N_12582,N_14355);
and UO_875 (O_875,N_12913,N_13837);
or UO_876 (O_876,N_12389,N_14203);
nand UO_877 (O_877,N_14821,N_14993);
or UO_878 (O_878,N_12546,N_12047);
and UO_879 (O_879,N_13021,N_12475);
nand UO_880 (O_880,N_13326,N_14924);
nor UO_881 (O_881,N_13869,N_12587);
and UO_882 (O_882,N_12897,N_14123);
or UO_883 (O_883,N_13189,N_14526);
nand UO_884 (O_884,N_13004,N_13963);
nor UO_885 (O_885,N_13690,N_13842);
or UO_886 (O_886,N_13539,N_14084);
nand UO_887 (O_887,N_14226,N_12452);
or UO_888 (O_888,N_14868,N_13324);
nor UO_889 (O_889,N_12428,N_14164);
or UO_890 (O_890,N_13137,N_12073);
xor UO_891 (O_891,N_12793,N_14210);
or UO_892 (O_892,N_14161,N_13362);
nand UO_893 (O_893,N_14973,N_14608);
and UO_894 (O_894,N_12811,N_14103);
nand UO_895 (O_895,N_14379,N_13442);
nand UO_896 (O_896,N_14273,N_12422);
and UO_897 (O_897,N_14175,N_12641);
or UO_898 (O_898,N_13475,N_13768);
and UO_899 (O_899,N_12036,N_12977);
and UO_900 (O_900,N_13357,N_14986);
or UO_901 (O_901,N_13919,N_13060);
nand UO_902 (O_902,N_14828,N_12181);
and UO_903 (O_903,N_13716,N_12324);
nor UO_904 (O_904,N_14156,N_12356);
and UO_905 (O_905,N_12055,N_12918);
and UO_906 (O_906,N_12662,N_12607);
or UO_907 (O_907,N_14408,N_12403);
or UO_908 (O_908,N_12567,N_13492);
nand UO_909 (O_909,N_14377,N_13386);
and UO_910 (O_910,N_14179,N_13620);
nor UO_911 (O_911,N_14917,N_13059);
nor UO_912 (O_912,N_12444,N_14873);
and UO_913 (O_913,N_13262,N_14057);
nand UO_914 (O_914,N_13465,N_14911);
and UO_915 (O_915,N_14292,N_12395);
nand UO_916 (O_916,N_14544,N_13038);
and UO_917 (O_917,N_13451,N_12790);
nand UO_918 (O_918,N_12716,N_14567);
and UO_919 (O_919,N_12916,N_14036);
and UO_920 (O_920,N_14476,N_12369);
and UO_921 (O_921,N_13739,N_14665);
or UO_922 (O_922,N_13356,N_13160);
and UO_923 (O_923,N_14866,N_14854);
nand UO_924 (O_924,N_13583,N_14957);
or UO_925 (O_925,N_14364,N_12649);
nand UO_926 (O_926,N_14819,N_12900);
and UO_927 (O_927,N_13762,N_13835);
nor UO_928 (O_928,N_13556,N_12940);
nor UO_929 (O_929,N_12239,N_12643);
nor UO_930 (O_930,N_14739,N_12632);
and UO_931 (O_931,N_14585,N_12017);
nand UO_932 (O_932,N_14323,N_13794);
xor UO_933 (O_933,N_14295,N_14339);
or UO_934 (O_934,N_14113,N_12783);
nor UO_935 (O_935,N_13686,N_12804);
or UO_936 (O_936,N_14829,N_13840);
or UO_937 (O_937,N_12163,N_14755);
or UO_938 (O_938,N_12796,N_13997);
nand UO_939 (O_939,N_13792,N_13124);
or UO_940 (O_940,N_12198,N_13023);
nand UO_941 (O_941,N_12829,N_14243);
or UO_942 (O_942,N_14529,N_13523);
nand UO_943 (O_943,N_12172,N_12272);
or UO_944 (O_944,N_13425,N_13519);
and UO_945 (O_945,N_13612,N_14704);
nand UO_946 (O_946,N_13773,N_13178);
nor UO_947 (O_947,N_13086,N_12837);
nand UO_948 (O_948,N_13866,N_12610);
or UO_949 (O_949,N_13187,N_12438);
nor UO_950 (O_950,N_14591,N_12747);
nand UO_951 (O_951,N_13380,N_13103);
or UO_952 (O_952,N_13120,N_14218);
nand UO_953 (O_953,N_12951,N_14439);
nor UO_954 (O_954,N_14011,N_14750);
nand UO_955 (O_955,N_12671,N_13317);
or UO_956 (O_956,N_13622,N_12455);
xnor UO_957 (O_957,N_12974,N_14496);
nand UO_958 (O_958,N_14539,N_12342);
xor UO_959 (O_959,N_13270,N_13461);
nor UO_960 (O_960,N_12775,N_13801);
nor UO_961 (O_961,N_13441,N_14267);
nand UO_962 (O_962,N_12464,N_12225);
and UO_963 (O_963,N_12859,N_12310);
and UO_964 (O_964,N_13637,N_13942);
nor UO_965 (O_965,N_13937,N_13873);
and UO_966 (O_966,N_12122,N_12001);
or UO_967 (O_967,N_13571,N_13982);
nand UO_968 (O_968,N_13268,N_13227);
or UO_969 (O_969,N_13713,N_14471);
nand UO_970 (O_970,N_14278,N_12112);
and UO_971 (O_971,N_14105,N_14966);
or UO_972 (O_972,N_14614,N_13344);
or UO_973 (O_973,N_13760,N_14360);
nand UO_974 (O_974,N_12376,N_14490);
nor UO_975 (O_975,N_12630,N_12375);
or UO_976 (O_976,N_14324,N_13805);
nor UO_977 (O_977,N_13366,N_14185);
or UO_978 (O_978,N_13456,N_14602);
or UO_979 (O_979,N_12433,N_14410);
nand UO_980 (O_980,N_14789,N_12234);
nor UO_981 (O_981,N_12454,N_13363);
and UO_982 (O_982,N_12458,N_13355);
and UO_983 (O_983,N_12915,N_12954);
nor UO_984 (O_984,N_12935,N_14521);
nand UO_985 (O_985,N_13962,N_13908);
and UO_986 (O_986,N_14900,N_12691);
or UO_987 (O_987,N_14204,N_13721);
or UO_988 (O_988,N_13745,N_13563);
and UO_989 (O_989,N_14470,N_13428);
nand UO_990 (O_990,N_14331,N_13418);
and UO_991 (O_991,N_14206,N_14014);
nand UO_992 (O_992,N_13018,N_13143);
nor UO_993 (O_993,N_14865,N_13988);
or UO_994 (O_994,N_14925,N_14548);
or UO_995 (O_995,N_14415,N_12620);
nand UO_996 (O_996,N_12479,N_13707);
and UO_997 (O_997,N_12360,N_12879);
nand UO_998 (O_998,N_12730,N_13818);
nand UO_999 (O_999,N_12825,N_14385);
nand UO_1000 (O_1000,N_12463,N_12334);
and UO_1001 (O_1001,N_14195,N_14150);
nor UO_1002 (O_1002,N_12826,N_12344);
and UO_1003 (O_1003,N_13158,N_13126);
and UO_1004 (O_1004,N_12621,N_14613);
or UO_1005 (O_1005,N_12432,N_14391);
and UO_1006 (O_1006,N_13846,N_13903);
nand UO_1007 (O_1007,N_14970,N_14734);
xnor UO_1008 (O_1008,N_13778,N_12058);
or UO_1009 (O_1009,N_13421,N_13781);
nand UO_1010 (O_1010,N_14717,N_13817);
or UO_1011 (O_1011,N_13682,N_12303);
nand UO_1012 (O_1012,N_12921,N_12425);
nand UO_1013 (O_1013,N_14055,N_14306);
nor UO_1014 (O_1014,N_12934,N_14338);
or UO_1015 (O_1015,N_13281,N_14940);
nor UO_1016 (O_1016,N_12503,N_14027);
or UO_1017 (O_1017,N_14404,N_12476);
or UO_1018 (O_1018,N_12391,N_12177);
and UO_1019 (O_1019,N_14445,N_14370);
nand UO_1020 (O_1020,N_12188,N_14572);
nand UO_1021 (O_1021,N_14597,N_12178);
nor UO_1022 (O_1022,N_13350,N_14706);
nor UO_1023 (O_1023,N_14451,N_14016);
xor UO_1024 (O_1024,N_14672,N_13349);
or UO_1025 (O_1025,N_13611,N_14208);
or UO_1026 (O_1026,N_14886,N_14792);
xor UO_1027 (O_1027,N_14503,N_14680);
or UO_1028 (O_1028,N_14425,N_13666);
nand UO_1029 (O_1029,N_12367,N_13239);
nand UO_1030 (O_1030,N_13367,N_13687);
nand UO_1031 (O_1031,N_13404,N_14958);
and UO_1032 (O_1032,N_14975,N_12850);
nand UO_1033 (O_1033,N_14875,N_13329);
nor UO_1034 (O_1034,N_12674,N_12003);
or UO_1035 (O_1035,N_13309,N_14976);
nor UO_1036 (O_1036,N_14674,N_12578);
nand UO_1037 (O_1037,N_14313,N_14475);
nor UO_1038 (O_1038,N_13678,N_14207);
nor UO_1039 (O_1039,N_13224,N_12786);
or UO_1040 (O_1040,N_14186,N_13945);
nand UO_1041 (O_1041,N_13480,N_14932);
nor UO_1042 (O_1042,N_14856,N_14374);
or UO_1043 (O_1043,N_13650,N_12373);
or UO_1044 (O_1044,N_13595,N_14823);
nand UO_1045 (O_1045,N_12197,N_13863);
xor UO_1046 (O_1046,N_12016,N_14193);
nand UO_1047 (O_1047,N_14453,N_14284);
and UO_1048 (O_1048,N_14007,N_12410);
and UO_1049 (O_1049,N_14722,N_13125);
nor UO_1050 (O_1050,N_12690,N_12078);
and UO_1051 (O_1051,N_14489,N_12969);
and UO_1052 (O_1052,N_13052,N_13316);
nand UO_1053 (O_1053,N_12753,N_13211);
nand UO_1054 (O_1054,N_12210,N_13481);
nand UO_1055 (O_1055,N_14809,N_13976);
nor UO_1056 (O_1056,N_14463,N_12372);
or UO_1057 (O_1057,N_14676,N_14968);
nor UO_1058 (O_1058,N_14582,N_13092);
or UO_1059 (O_1059,N_14427,N_13782);
nand UO_1060 (O_1060,N_13079,N_13746);
nand UO_1061 (O_1061,N_12591,N_12167);
or UO_1062 (O_1062,N_12362,N_14299);
nor UO_1063 (O_1063,N_13561,N_12828);
nor UO_1064 (O_1064,N_14881,N_13271);
and UO_1065 (O_1065,N_14552,N_12884);
nor UO_1066 (O_1066,N_14785,N_14176);
and UO_1067 (O_1067,N_14533,N_14518);
nor UO_1068 (O_1068,N_13231,N_12867);
nand UO_1069 (O_1069,N_14740,N_12080);
nor UO_1070 (O_1070,N_12092,N_13072);
nand UO_1071 (O_1071,N_14151,N_14006);
or UO_1072 (O_1072,N_12300,N_12160);
or UO_1073 (O_1073,N_13736,N_13393);
xnor UO_1074 (O_1074,N_13796,N_12740);
or UO_1075 (O_1075,N_12883,N_12820);
nand UO_1076 (O_1076,N_13341,N_14566);
and UO_1077 (O_1077,N_13766,N_13999);
or UO_1078 (O_1078,N_14801,N_12358);
nor UO_1079 (O_1079,N_14080,N_12717);
and UO_1080 (O_1080,N_14314,N_12263);
xnor UO_1081 (O_1081,N_14618,N_12461);
nand UO_1082 (O_1082,N_13284,N_12797);
and UO_1083 (O_1083,N_12366,N_14688);
or UO_1084 (O_1084,N_12634,N_14350);
nand UO_1085 (O_1085,N_14770,N_13427);
nor UO_1086 (O_1086,N_14072,N_14934);
and UO_1087 (O_1087,N_14605,N_14610);
and UO_1088 (O_1088,N_12864,N_14832);
nor UO_1089 (O_1089,N_13656,N_14466);
and UO_1090 (O_1090,N_14724,N_14898);
and UO_1091 (O_1091,N_14358,N_12192);
nand UO_1092 (O_1092,N_14104,N_13283);
and UO_1093 (O_1093,N_14876,N_14519);
nor UO_1094 (O_1094,N_14824,N_13524);
nand UO_1095 (O_1095,N_13930,N_12059);
or UO_1096 (O_1096,N_14389,N_13446);
nor UO_1097 (O_1097,N_13347,N_12626);
or UO_1098 (O_1098,N_12543,N_14075);
or UO_1099 (O_1099,N_14715,N_14216);
nand UO_1100 (O_1100,N_13532,N_12252);
or UO_1101 (O_1101,N_13352,N_12834);
and UO_1102 (O_1102,N_13775,N_14029);
or UO_1103 (O_1103,N_13336,N_14143);
nor UO_1104 (O_1104,N_12484,N_14839);
nand UO_1105 (O_1105,N_13570,N_14501);
or UO_1106 (O_1106,N_13312,N_12487);
or UO_1107 (O_1107,N_13379,N_12244);
and UO_1108 (O_1108,N_12514,N_13012);
xor UO_1109 (O_1109,N_14711,N_12650);
and UO_1110 (O_1110,N_12998,N_14536);
nor UO_1111 (O_1111,N_14010,N_13665);
and UO_1112 (O_1112,N_13247,N_12771);
or UO_1113 (O_1113,N_12243,N_14188);
xnor UO_1114 (O_1114,N_14913,N_13044);
nand UO_1115 (O_1115,N_12308,N_13093);
nor UO_1116 (O_1116,N_12379,N_12199);
nor UO_1117 (O_1117,N_14965,N_12595);
or UO_1118 (O_1118,N_13872,N_12605);
nand UO_1119 (O_1119,N_12914,N_12121);
and UO_1120 (O_1120,N_13671,N_12033);
and UO_1121 (O_1121,N_14033,N_13029);
nand UO_1122 (O_1122,N_12763,N_13482);
or UO_1123 (O_1123,N_12406,N_13537);
and UO_1124 (O_1124,N_14580,N_12777);
or UO_1125 (O_1125,N_12611,N_12713);
nand UO_1126 (O_1126,N_14779,N_12290);
and UO_1127 (O_1127,N_13520,N_14231);
nand UO_1128 (O_1128,N_13353,N_12899);
and UO_1129 (O_1129,N_12319,N_14437);
or UO_1130 (O_1130,N_14064,N_13542);
nand UO_1131 (O_1131,N_13910,N_12525);
nand UO_1132 (O_1132,N_13348,N_13717);
nor UO_1133 (O_1133,N_14820,N_14028);
nor UO_1134 (O_1134,N_12501,N_14397);
or UO_1135 (O_1135,N_12384,N_12863);
or UO_1136 (O_1136,N_14669,N_14230);
or UO_1137 (O_1137,N_12462,N_14916);
nand UO_1138 (O_1138,N_12768,N_14275);
nor UO_1139 (O_1139,N_14768,N_13201);
nand UO_1140 (O_1140,N_13048,N_12529);
nand UO_1141 (O_1141,N_14619,N_13787);
xor UO_1142 (O_1142,N_14748,N_12957);
nand UO_1143 (O_1143,N_14738,N_13786);
nand UO_1144 (O_1144,N_13437,N_12250);
and UO_1145 (O_1145,N_12664,N_14660);
nand UO_1146 (O_1146,N_12604,N_12162);
xor UO_1147 (O_1147,N_13375,N_14297);
nor UO_1148 (O_1148,N_14638,N_13228);
or UO_1149 (O_1149,N_14767,N_13979);
or UO_1150 (O_1150,N_14395,N_14443);
or UO_1151 (O_1151,N_14885,N_13115);
and UO_1152 (O_1152,N_13374,N_14345);
nand UO_1153 (O_1153,N_13245,N_13377);
nand UO_1154 (O_1154,N_12357,N_12871);
xor UO_1155 (O_1155,N_12070,N_12886);
and UO_1156 (O_1156,N_14537,N_14015);
or UO_1157 (O_1157,N_13535,N_14634);
and UO_1158 (O_1158,N_14713,N_13166);
nand UO_1159 (O_1159,N_14617,N_12670);
nand UO_1160 (O_1160,N_14887,N_14147);
or UO_1161 (O_1161,N_12531,N_13573);
nand UO_1162 (O_1162,N_13119,N_12628);
and UO_1163 (O_1163,N_12194,N_12321);
nor UO_1164 (O_1164,N_12878,N_12861);
and UO_1165 (O_1165,N_14309,N_12504);
nand UO_1166 (O_1166,N_14894,N_13040);
nor UO_1167 (O_1167,N_14507,N_13050);
nor UO_1168 (O_1168,N_12724,N_13041);
and UO_1169 (O_1169,N_14778,N_14517);
or UO_1170 (O_1170,N_13398,N_12283);
nand UO_1171 (O_1171,N_13015,N_12677);
nand UO_1172 (O_1172,N_14646,N_12955);
or UO_1173 (O_1173,N_13886,N_14199);
nand UO_1174 (O_1174,N_13057,N_13384);
and UO_1175 (O_1175,N_14413,N_12149);
nand UO_1176 (O_1176,N_12125,N_14448);
nor UO_1177 (O_1177,N_13318,N_12348);
or UO_1178 (O_1178,N_13920,N_12204);
nor UO_1179 (O_1179,N_12168,N_12562);
nand UO_1180 (O_1180,N_12187,N_12597);
nand UO_1181 (O_1181,N_13944,N_14265);
nor UO_1182 (O_1182,N_14675,N_12613);
nor UO_1183 (O_1183,N_13534,N_12135);
and UO_1184 (O_1184,N_14969,N_13662);
nand UO_1185 (O_1185,N_13516,N_12585);
nand UO_1186 (O_1186,N_12052,N_13127);
nor UO_1187 (O_1187,N_13855,N_12265);
xor UO_1188 (O_1188,N_13164,N_13615);
and UO_1189 (O_1189,N_12064,N_14130);
nand UO_1190 (O_1190,N_13028,N_13882);
and UO_1191 (O_1191,N_14520,N_14012);
nand UO_1192 (O_1192,N_14570,N_12994);
and UO_1193 (O_1193,N_13784,N_13488);
and UO_1194 (O_1194,N_12101,N_13467);
nor UO_1195 (O_1195,N_13870,N_13683);
nor UO_1196 (O_1196,N_14486,N_12533);
or UO_1197 (O_1197,N_14473,N_13700);
and UO_1198 (O_1198,N_14962,N_14579);
and UO_1199 (O_1199,N_14091,N_14753);
nor UO_1200 (O_1200,N_13122,N_12731);
nand UO_1201 (O_1201,N_14721,N_13590);
and UO_1202 (O_1202,N_14140,N_13256);
and UO_1203 (O_1203,N_12537,N_14880);
or UO_1204 (O_1204,N_12963,N_12147);
nand UO_1205 (O_1205,N_14515,N_14577);
xnor UO_1206 (O_1206,N_14141,N_12274);
or UO_1207 (O_1207,N_13950,N_14568);
and UO_1208 (O_1208,N_13269,N_14488);
and UO_1209 (O_1209,N_12209,N_12449);
or UO_1210 (O_1210,N_14623,N_12394);
nand UO_1211 (O_1211,N_12223,N_12907);
nor UO_1212 (O_1212,N_13627,N_13741);
xor UO_1213 (O_1213,N_13952,N_14870);
or UO_1214 (O_1214,N_14124,N_12138);
or UO_1215 (O_1215,N_12084,N_12339);
and UO_1216 (O_1216,N_12814,N_13321);
nor UO_1217 (O_1217,N_12148,N_14142);
nor UO_1218 (O_1218,N_12839,N_14632);
xnor UO_1219 (O_1219,N_14504,N_12860);
nand UO_1220 (O_1220,N_13151,N_14258);
nand UO_1221 (O_1221,N_13131,N_14263);
nand UO_1222 (O_1222,N_13691,N_12807);
and UO_1223 (O_1223,N_13924,N_13555);
and UO_1224 (O_1224,N_13859,N_14849);
nor UO_1225 (O_1225,N_12294,N_14050);
or UO_1226 (O_1226,N_13648,N_14416);
nor UO_1227 (O_1227,N_12268,N_13954);
or UO_1228 (O_1228,N_13978,N_14023);
or UO_1229 (O_1229,N_13900,N_12809);
or UO_1230 (O_1230,N_12446,N_14247);
nand UO_1231 (O_1231,N_13913,N_12307);
nand UO_1232 (O_1232,N_13517,N_13711);
nand UO_1233 (O_1233,N_13417,N_14100);
nor UO_1234 (O_1234,N_13407,N_14497);
nor UO_1235 (O_1235,N_12067,N_13019);
and UO_1236 (O_1236,N_14545,N_13664);
nor UO_1237 (O_1237,N_13811,N_13035);
or UO_1238 (O_1238,N_12217,N_12889);
and UO_1239 (O_1239,N_12898,N_14485);
nor UO_1240 (O_1240,N_13207,N_14333);
and UO_1241 (O_1241,N_13601,N_12896);
or UO_1242 (O_1242,N_14022,N_13032);
or UO_1243 (O_1243,N_13214,N_14673);
nand UO_1244 (O_1244,N_14888,N_13102);
and UO_1245 (O_1245,N_12739,N_14336);
or UO_1246 (O_1246,N_13861,N_13725);
nand UO_1247 (O_1247,N_12794,N_14153);
or UO_1248 (O_1248,N_13308,N_14512);
nand UO_1249 (O_1249,N_12323,N_13045);
nand UO_1250 (O_1250,N_12892,N_12069);
nor UO_1251 (O_1251,N_14972,N_14049);
nand UO_1252 (O_1252,N_12656,N_14277);
or UO_1253 (O_1253,N_14378,N_13266);
nand UO_1254 (O_1254,N_13558,N_14414);
xor UO_1255 (O_1255,N_13194,N_12241);
and UO_1256 (O_1256,N_12421,N_13763);
nand UO_1257 (O_1257,N_14214,N_12734);
nor UO_1258 (O_1258,N_13623,N_12281);
nor UO_1259 (O_1259,N_12642,N_14804);
or UO_1260 (O_1260,N_14169,N_13636);
or UO_1261 (O_1261,N_14639,N_13599);
and UO_1262 (O_1262,N_12315,N_12012);
nand UO_1263 (O_1263,N_12841,N_12386);
or UO_1264 (O_1264,N_14298,N_13364);
nor UO_1265 (O_1265,N_12547,N_13819);
and UO_1266 (O_1266,N_13469,N_12132);
or UO_1267 (O_1267,N_14943,N_14562);
nand UO_1268 (O_1268,N_13966,N_14252);
xor UO_1269 (O_1269,N_13693,N_14964);
and UO_1270 (O_1270,N_13395,N_14481);
and UO_1271 (O_1271,N_14115,N_12269);
and UO_1272 (O_1272,N_12579,N_14541);
nand UO_1273 (O_1273,N_14933,N_12179);
and UO_1274 (O_1274,N_14852,N_14635);
and UO_1275 (O_1275,N_12440,N_14671);
xor UO_1276 (O_1276,N_14182,N_14044);
nand UO_1277 (O_1277,N_12426,N_14078);
nor UO_1278 (O_1278,N_14796,N_14923);
and UO_1279 (O_1279,N_13483,N_12554);
nand UO_1280 (O_1280,N_13521,N_12277);
nand UO_1281 (O_1281,N_12028,N_13756);
nor UO_1282 (O_1282,N_12996,N_12660);
and UO_1283 (O_1283,N_13197,N_13403);
or UO_1284 (O_1284,N_13618,N_12013);
and UO_1285 (O_1285,N_14647,N_14491);
nand UO_1286 (O_1286,N_13022,N_13111);
nand UO_1287 (O_1287,N_13526,N_13275);
nor UO_1288 (O_1288,N_12291,N_13810);
or UO_1289 (O_1289,N_12701,N_12708);
nor UO_1290 (O_1290,N_13631,N_12292);
or UO_1291 (O_1291,N_13894,N_13033);
nand UO_1292 (O_1292,N_13658,N_12141);
nor UO_1293 (O_1293,N_12314,N_14407);
and UO_1294 (O_1294,N_13515,N_14847);
or UO_1295 (O_1295,N_12235,N_12388);
nand UO_1296 (O_1296,N_12098,N_12191);
or UO_1297 (O_1297,N_14059,N_14803);
nor UO_1298 (O_1298,N_14683,N_13733);
nor UO_1299 (O_1299,N_13219,N_12689);
and UO_1300 (O_1300,N_12278,N_13110);
xor UO_1301 (O_1301,N_12888,N_14763);
nor UO_1302 (O_1302,N_13265,N_14386);
and UO_1303 (O_1303,N_13911,N_13701);
and UO_1304 (O_1304,N_12412,N_13603);
and UO_1305 (O_1305,N_14388,N_12489);
and UO_1306 (O_1306,N_14878,N_12732);
xnor UO_1307 (O_1307,N_12035,N_13970);
and UO_1308 (O_1308,N_12044,N_14590);
and UO_1309 (O_1309,N_12466,N_14291);
nand UO_1310 (O_1310,N_14677,N_14127);
nand UO_1311 (O_1311,N_14343,N_12551);
and UO_1312 (O_1312,N_14272,N_14365);
and UO_1313 (O_1313,N_12295,N_12870);
nand UO_1314 (O_1314,N_13809,N_12655);
nor UO_1315 (O_1315,N_14097,N_12450);
and UO_1316 (O_1316,N_14354,N_12665);
nor UO_1317 (O_1317,N_13287,N_12327);
nand UO_1318 (O_1318,N_14850,N_13426);
nor UO_1319 (O_1319,N_12351,N_12216);
and UO_1320 (O_1320,N_13967,N_13586);
nand UO_1321 (O_1321,N_13709,N_14261);
and UO_1322 (O_1322,N_13091,N_13578);
nor UO_1323 (O_1323,N_14694,N_12233);
nor UO_1324 (O_1324,N_13862,N_14592);
nor UO_1325 (O_1325,N_12667,N_12836);
nor UO_1326 (O_1326,N_12072,N_14929);
and UO_1327 (O_1327,N_12982,N_12856);
nand UO_1328 (O_1328,N_14073,N_13901);
nor UO_1329 (O_1329,N_14889,N_14362);
or UO_1330 (O_1330,N_12031,N_13078);
and UO_1331 (O_1331,N_13031,N_14232);
nand UO_1332 (O_1332,N_13991,N_12002);
nor UO_1333 (O_1333,N_13466,N_13990);
nor UO_1334 (O_1334,N_14775,N_14522);
nand UO_1335 (O_1335,N_13575,N_14412);
xnor UO_1336 (O_1336,N_12328,N_14046);
nor UO_1337 (O_1337,N_14955,N_14633);
and UO_1338 (O_1338,N_12124,N_12247);
nand UO_1339 (O_1339,N_14644,N_14947);
or UO_1340 (O_1340,N_12347,N_13505);
and UO_1341 (O_1341,N_14102,N_14598);
or UO_1342 (O_1342,N_13728,N_12941);
nor UO_1343 (O_1343,N_12471,N_12965);
nand UO_1344 (O_1344,N_14368,N_14995);
or UO_1345 (O_1345,N_14250,N_14757);
nor UO_1346 (O_1346,N_13715,N_12502);
nand UO_1347 (O_1347,N_12004,N_12802);
nand UO_1348 (O_1348,N_12333,N_13302);
nand UO_1349 (O_1349,N_12005,N_13147);
nand UO_1350 (O_1350,N_12556,N_14260);
or UO_1351 (O_1351,N_13339,N_13049);
and UO_1352 (O_1352,N_12161,N_13509);
nand UO_1353 (O_1353,N_14189,N_14487);
or UO_1354 (O_1354,N_14931,N_14234);
or UO_1355 (O_1355,N_12685,N_14224);
nor UO_1356 (O_1356,N_13249,N_12855);
and UO_1357 (O_1357,N_12684,N_13948);
and UO_1358 (O_1358,N_13081,N_13140);
nor UO_1359 (O_1359,N_14347,N_12061);
and UO_1360 (O_1360,N_13248,N_14662);
or UO_1361 (O_1361,N_12083,N_13744);
and UO_1362 (O_1362,N_13964,N_14514);
and UO_1363 (O_1363,N_14531,N_12203);
or UO_1364 (O_1364,N_14631,N_13109);
nand UO_1365 (O_1365,N_12622,N_12680);
nand UO_1366 (O_1366,N_12981,N_13373);
nor UO_1367 (O_1367,N_14742,N_14705);
or UO_1368 (O_1368,N_13370,N_14777);
or UO_1369 (O_1369,N_12816,N_12636);
nor UO_1370 (O_1370,N_13947,N_12766);
nand UO_1371 (O_1371,N_14535,N_14316);
and UO_1372 (O_1372,N_12405,N_13065);
nor UO_1373 (O_1373,N_13389,N_12128);
nor UO_1374 (O_1374,N_12174,N_12952);
and UO_1375 (O_1375,N_14132,N_13565);
nand UO_1376 (O_1376,N_14402,N_14139);
or UO_1377 (O_1377,N_13958,N_12218);
nor UO_1378 (O_1378,N_14121,N_14256);
nand UO_1379 (O_1379,N_12201,N_13090);
or UO_1380 (O_1380,N_12805,N_12893);
or UO_1381 (O_1381,N_12413,N_14184);
nand UO_1382 (O_1382,N_12720,N_14399);
or UO_1383 (O_1383,N_13892,N_14319);
nand UO_1384 (O_1384,N_14242,N_12906);
or UO_1385 (O_1385,N_13068,N_14718);
nor UO_1386 (O_1386,N_13087,N_13017);
and UO_1387 (O_1387,N_13199,N_14959);
or UO_1388 (O_1388,N_12924,N_12007);
and UO_1389 (O_1389,N_12057,N_14119);
nand UO_1390 (O_1390,N_13986,N_12054);
or UO_1391 (O_1391,N_12271,N_14702);
or UO_1392 (O_1392,N_14145,N_13113);
and UO_1393 (O_1393,N_12153,N_14892);
or UO_1394 (O_1394,N_12703,N_12881);
nor UO_1395 (O_1395,N_13303,N_14555);
and UO_1396 (O_1396,N_13799,N_14815);
and UO_1397 (O_1397,N_13422,N_14997);
nor UO_1398 (O_1398,N_12424,N_14283);
and UO_1399 (O_1399,N_14864,N_14793);
and UO_1400 (O_1400,N_12352,N_14827);
nand UO_1401 (O_1401,N_13314,N_13619);
nor UO_1402 (O_1402,N_14118,N_12071);
and UO_1403 (O_1403,N_12714,N_13073);
nor UO_1404 (O_1404,N_12830,N_14417);
and UO_1405 (O_1405,N_12568,N_14565);
nand UO_1406 (O_1406,N_12751,N_14220);
nor UO_1407 (O_1407,N_14670,N_13278);
nor UO_1408 (O_1408,N_14170,N_13998);
and UO_1409 (O_1409,N_13605,N_12152);
or UO_1410 (O_1410,N_14902,N_13135);
and UO_1411 (O_1411,N_13698,N_14455);
nand UO_1412 (O_1412,N_12374,N_14599);
and UO_1413 (O_1413,N_13585,N_12638);
nor UO_1414 (O_1414,N_12984,N_14813);
nand UO_1415 (O_1415,N_14528,N_14830);
and UO_1416 (O_1416,N_12257,N_13378);
nor UO_1417 (O_1417,N_14987,N_13293);
and UO_1418 (O_1418,N_13209,N_13063);
nand UO_1419 (O_1419,N_14791,N_14707);
nor UO_1420 (O_1420,N_13896,N_14332);
nor UO_1421 (O_1421,N_12156,N_12040);
nand UO_1422 (O_1422,N_12326,N_14009);
nand UO_1423 (O_1423,N_14776,N_13547);
or UO_1424 (O_1424,N_12506,N_12382);
nor UO_1425 (O_1425,N_13938,N_12365);
nor UO_1426 (O_1426,N_12447,N_12494);
and UO_1427 (O_1427,N_14762,N_12419);
or UO_1428 (O_1428,N_14584,N_12508);
or UO_1429 (O_1429,N_13548,N_12115);
nor UO_1430 (O_1430,N_12663,N_12603);
nor UO_1431 (O_1431,N_13267,N_12488);
xnor UO_1432 (O_1432,N_12581,N_14373);
nor UO_1433 (O_1433,N_13731,N_12037);
nor UO_1434 (O_1434,N_12226,N_14081);
or UO_1435 (O_1435,N_14479,N_14167);
nor UO_1436 (O_1436,N_14692,N_12312);
or UO_1437 (O_1437,N_12760,N_14315);
or UO_1438 (O_1438,N_13358,N_12100);
or UO_1439 (O_1439,N_14640,N_14922);
nor UO_1440 (O_1440,N_12648,N_12835);
and UO_1441 (O_1441,N_12702,N_12196);
or UO_1442 (O_1442,N_12919,N_12929);
nor UO_1443 (O_1443,N_14686,N_12311);
and UO_1444 (O_1444,N_12431,N_14697);
nand UO_1445 (O_1445,N_13183,N_13006);
and UO_1446 (O_1446,N_13580,N_12776);
or UO_1447 (O_1447,N_12925,N_13994);
and UO_1448 (O_1448,N_14259,N_12661);
or UO_1449 (O_1449,N_13101,N_13253);
and UO_1450 (O_1450,N_14087,N_14468);
and UO_1451 (O_1451,N_13510,N_12944);
or UO_1452 (O_1452,N_14589,N_14392);
or UO_1453 (O_1453,N_14066,N_13729);
nor UO_1454 (O_1454,N_13024,N_12173);
nor UO_1455 (O_1455,N_13654,N_13493);
nor UO_1456 (O_1456,N_14438,N_12477);
or UO_1457 (O_1457,N_12922,N_14607);
or UO_1458 (O_1458,N_12205,N_13845);
nand UO_1459 (O_1459,N_13487,N_14764);
and UO_1460 (O_1460,N_12439,N_14843);
or UO_1461 (O_1461,N_13477,N_14240);
nor UO_1462 (O_1462,N_13202,N_12510);
or UO_1463 (O_1463,N_14650,N_14745);
nor UO_1464 (O_1464,N_14600,N_13167);
nand UO_1465 (O_1465,N_13497,N_13288);
xor UO_1466 (O_1466,N_12558,N_14018);
nor UO_1467 (O_1467,N_13852,N_12317);
or UO_1468 (O_1468,N_12721,N_13630);
nor UO_1469 (O_1469,N_13803,N_13730);
nand UO_1470 (O_1470,N_12301,N_13506);
nor UO_1471 (O_1471,N_13538,N_13240);
or UO_1472 (O_1472,N_12436,N_14919);
and UO_1473 (O_1473,N_12675,N_14361);
nor UO_1474 (O_1474,N_12108,N_13504);
or UO_1475 (O_1475,N_13879,N_13657);
and UO_1476 (O_1476,N_14953,N_13853);
or UO_1477 (O_1477,N_14051,N_14573);
or UO_1478 (O_1478,N_12030,N_14245);
or UO_1479 (O_1479,N_13039,N_13225);
nand UO_1480 (O_1480,N_12482,N_12532);
nand UO_1481 (O_1481,N_13200,N_14197);
or UO_1482 (O_1482,N_12293,N_13918);
and UO_1483 (O_1483,N_14576,N_12006);
or UO_1484 (O_1484,N_14586,N_14086);
and UO_1485 (O_1485,N_14390,N_12679);
or UO_1486 (O_1486,N_12967,N_12539);
nor UO_1487 (O_1487,N_12270,N_12842);
nand UO_1488 (O_1488,N_12908,N_13940);
and UO_1489 (O_1489,N_13499,N_13527);
nor UO_1490 (O_1490,N_12669,N_12206);
nand UO_1491 (O_1491,N_14067,N_12968);
nor UO_1492 (O_1492,N_12411,N_13629);
and UO_1493 (O_1493,N_13953,N_13593);
nor UO_1494 (O_1494,N_14021,N_13993);
nand UO_1495 (O_1495,N_13554,N_13276);
nand UO_1496 (O_1496,N_13540,N_12519);
nand UO_1497 (O_1497,N_14270,N_12958);
nand UO_1498 (O_1498,N_13617,N_13191);
nor UO_1499 (O_1499,N_14155,N_14249);
and UO_1500 (O_1500,N_14488,N_13686);
and UO_1501 (O_1501,N_13111,N_13642);
xor UO_1502 (O_1502,N_12660,N_12874);
or UO_1503 (O_1503,N_13334,N_14071);
and UO_1504 (O_1504,N_14878,N_12974);
and UO_1505 (O_1505,N_12357,N_12009);
or UO_1506 (O_1506,N_13161,N_12491);
nand UO_1507 (O_1507,N_13650,N_13856);
nand UO_1508 (O_1508,N_12144,N_13664);
and UO_1509 (O_1509,N_14757,N_13969);
nor UO_1510 (O_1510,N_13863,N_12956);
nand UO_1511 (O_1511,N_14856,N_12793);
nor UO_1512 (O_1512,N_12631,N_13272);
nand UO_1513 (O_1513,N_14751,N_14285);
or UO_1514 (O_1514,N_13956,N_14809);
and UO_1515 (O_1515,N_12293,N_12479);
and UO_1516 (O_1516,N_13163,N_14605);
nor UO_1517 (O_1517,N_14644,N_12771);
nor UO_1518 (O_1518,N_12441,N_12330);
nor UO_1519 (O_1519,N_13739,N_14090);
and UO_1520 (O_1520,N_14423,N_14573);
or UO_1521 (O_1521,N_13558,N_13643);
nand UO_1522 (O_1522,N_12716,N_14523);
nand UO_1523 (O_1523,N_14343,N_13938);
nand UO_1524 (O_1524,N_13820,N_14823);
or UO_1525 (O_1525,N_12083,N_13602);
or UO_1526 (O_1526,N_13209,N_14275);
and UO_1527 (O_1527,N_13969,N_12198);
nor UO_1528 (O_1528,N_14284,N_14079);
nand UO_1529 (O_1529,N_12302,N_14035);
nand UO_1530 (O_1530,N_12218,N_14162);
nor UO_1531 (O_1531,N_13513,N_13408);
or UO_1532 (O_1532,N_13293,N_14102);
nand UO_1533 (O_1533,N_13134,N_14854);
or UO_1534 (O_1534,N_14413,N_12115);
nor UO_1535 (O_1535,N_12700,N_12913);
nor UO_1536 (O_1536,N_13034,N_13428);
or UO_1537 (O_1537,N_13695,N_14283);
nand UO_1538 (O_1538,N_13658,N_14399);
and UO_1539 (O_1539,N_13807,N_13776);
or UO_1540 (O_1540,N_14935,N_12903);
nor UO_1541 (O_1541,N_13540,N_14872);
or UO_1542 (O_1542,N_13263,N_14931);
nor UO_1543 (O_1543,N_14429,N_13275);
or UO_1544 (O_1544,N_13671,N_13299);
and UO_1545 (O_1545,N_13073,N_13932);
nor UO_1546 (O_1546,N_13892,N_14613);
nand UO_1547 (O_1547,N_12160,N_12669);
nand UO_1548 (O_1548,N_12580,N_12863);
nand UO_1549 (O_1549,N_13446,N_12113);
nand UO_1550 (O_1550,N_14320,N_12759);
nor UO_1551 (O_1551,N_13529,N_14825);
and UO_1552 (O_1552,N_14375,N_12498);
nor UO_1553 (O_1553,N_14842,N_14785);
or UO_1554 (O_1554,N_12754,N_13596);
nand UO_1555 (O_1555,N_13255,N_13311);
or UO_1556 (O_1556,N_12703,N_12450);
and UO_1557 (O_1557,N_13278,N_12831);
or UO_1558 (O_1558,N_14700,N_13292);
or UO_1559 (O_1559,N_14328,N_13043);
nor UO_1560 (O_1560,N_12573,N_12521);
and UO_1561 (O_1561,N_12581,N_14023);
nand UO_1562 (O_1562,N_12983,N_13613);
or UO_1563 (O_1563,N_14863,N_12613);
or UO_1564 (O_1564,N_12985,N_13734);
and UO_1565 (O_1565,N_13271,N_14992);
xor UO_1566 (O_1566,N_14979,N_13929);
nor UO_1567 (O_1567,N_13891,N_13901);
or UO_1568 (O_1568,N_14389,N_12191);
and UO_1569 (O_1569,N_13746,N_14358);
nand UO_1570 (O_1570,N_13700,N_13645);
nor UO_1571 (O_1571,N_14567,N_14558);
xnor UO_1572 (O_1572,N_14039,N_13670);
and UO_1573 (O_1573,N_12283,N_14680);
nand UO_1574 (O_1574,N_12573,N_13052);
or UO_1575 (O_1575,N_13042,N_14984);
and UO_1576 (O_1576,N_12668,N_13941);
or UO_1577 (O_1577,N_14099,N_12462);
or UO_1578 (O_1578,N_13699,N_13158);
and UO_1579 (O_1579,N_14361,N_13738);
nand UO_1580 (O_1580,N_12331,N_13892);
or UO_1581 (O_1581,N_13188,N_14115);
xor UO_1582 (O_1582,N_12626,N_14561);
nor UO_1583 (O_1583,N_13208,N_12867);
nand UO_1584 (O_1584,N_12402,N_13173);
nor UO_1585 (O_1585,N_12018,N_12494);
or UO_1586 (O_1586,N_12432,N_13765);
or UO_1587 (O_1587,N_13220,N_12861);
nor UO_1588 (O_1588,N_12240,N_12159);
or UO_1589 (O_1589,N_12617,N_13188);
and UO_1590 (O_1590,N_12737,N_13592);
nand UO_1591 (O_1591,N_13364,N_12937);
nor UO_1592 (O_1592,N_12540,N_12544);
or UO_1593 (O_1593,N_12515,N_13582);
and UO_1594 (O_1594,N_14767,N_13846);
nand UO_1595 (O_1595,N_12895,N_14066);
and UO_1596 (O_1596,N_12843,N_12317);
and UO_1597 (O_1597,N_13698,N_13661);
xor UO_1598 (O_1598,N_13173,N_13955);
nand UO_1599 (O_1599,N_13854,N_12035);
or UO_1600 (O_1600,N_14620,N_12969);
nand UO_1601 (O_1601,N_14641,N_12409);
or UO_1602 (O_1602,N_13386,N_14074);
and UO_1603 (O_1603,N_12625,N_13559);
and UO_1604 (O_1604,N_13164,N_14509);
or UO_1605 (O_1605,N_12868,N_13174);
or UO_1606 (O_1606,N_13606,N_14405);
and UO_1607 (O_1607,N_14296,N_14785);
nand UO_1608 (O_1608,N_14708,N_12520);
nand UO_1609 (O_1609,N_12749,N_14096);
nor UO_1610 (O_1610,N_12352,N_12811);
or UO_1611 (O_1611,N_12186,N_13916);
or UO_1612 (O_1612,N_13162,N_13948);
and UO_1613 (O_1613,N_14884,N_12826);
or UO_1614 (O_1614,N_12755,N_13182);
or UO_1615 (O_1615,N_13619,N_12930);
nand UO_1616 (O_1616,N_12240,N_14691);
nand UO_1617 (O_1617,N_13027,N_12921);
nor UO_1618 (O_1618,N_14623,N_14528);
nor UO_1619 (O_1619,N_14182,N_13562);
and UO_1620 (O_1620,N_14252,N_14275);
and UO_1621 (O_1621,N_14383,N_14148);
nand UO_1622 (O_1622,N_13699,N_14563);
or UO_1623 (O_1623,N_12687,N_14831);
nand UO_1624 (O_1624,N_13736,N_13696);
nor UO_1625 (O_1625,N_14539,N_14872);
nor UO_1626 (O_1626,N_14697,N_12868);
nand UO_1627 (O_1627,N_14962,N_14178);
nand UO_1628 (O_1628,N_13542,N_13176);
and UO_1629 (O_1629,N_12936,N_14807);
or UO_1630 (O_1630,N_14620,N_12745);
nor UO_1631 (O_1631,N_12831,N_13824);
or UO_1632 (O_1632,N_14108,N_14751);
and UO_1633 (O_1633,N_13037,N_14708);
nor UO_1634 (O_1634,N_14613,N_13544);
or UO_1635 (O_1635,N_12023,N_14992);
and UO_1636 (O_1636,N_13597,N_14922);
nand UO_1637 (O_1637,N_14193,N_12009);
nand UO_1638 (O_1638,N_13501,N_12292);
and UO_1639 (O_1639,N_13206,N_12287);
or UO_1640 (O_1640,N_14485,N_14802);
nor UO_1641 (O_1641,N_14771,N_13682);
nand UO_1642 (O_1642,N_13389,N_12569);
or UO_1643 (O_1643,N_13634,N_13620);
nor UO_1644 (O_1644,N_14656,N_14311);
and UO_1645 (O_1645,N_14254,N_12372);
and UO_1646 (O_1646,N_12258,N_14200);
nor UO_1647 (O_1647,N_12972,N_13451);
and UO_1648 (O_1648,N_14312,N_14243);
or UO_1649 (O_1649,N_14438,N_13340);
nand UO_1650 (O_1650,N_12551,N_14647);
and UO_1651 (O_1651,N_13616,N_13857);
nor UO_1652 (O_1652,N_14211,N_12112);
nor UO_1653 (O_1653,N_13162,N_13074);
and UO_1654 (O_1654,N_14680,N_14027);
or UO_1655 (O_1655,N_13130,N_14968);
and UO_1656 (O_1656,N_12996,N_14183);
and UO_1657 (O_1657,N_14667,N_12607);
nor UO_1658 (O_1658,N_13590,N_12936);
or UO_1659 (O_1659,N_14043,N_12356);
or UO_1660 (O_1660,N_14105,N_13753);
nor UO_1661 (O_1661,N_14903,N_14339);
or UO_1662 (O_1662,N_13698,N_14924);
nand UO_1663 (O_1663,N_14574,N_12338);
nor UO_1664 (O_1664,N_13442,N_13841);
nand UO_1665 (O_1665,N_14384,N_12384);
and UO_1666 (O_1666,N_12814,N_13772);
nor UO_1667 (O_1667,N_14952,N_12264);
xnor UO_1668 (O_1668,N_13430,N_14130);
nand UO_1669 (O_1669,N_12898,N_14490);
nand UO_1670 (O_1670,N_12236,N_14513);
and UO_1671 (O_1671,N_12732,N_14699);
or UO_1672 (O_1672,N_12708,N_13927);
and UO_1673 (O_1673,N_14597,N_13160);
and UO_1674 (O_1674,N_14717,N_12593);
or UO_1675 (O_1675,N_14816,N_14199);
nand UO_1676 (O_1676,N_12217,N_14293);
or UO_1677 (O_1677,N_14167,N_12124);
nand UO_1678 (O_1678,N_14961,N_12589);
and UO_1679 (O_1679,N_12071,N_14103);
nand UO_1680 (O_1680,N_12487,N_12704);
or UO_1681 (O_1681,N_13662,N_12673);
and UO_1682 (O_1682,N_14727,N_13306);
or UO_1683 (O_1683,N_12727,N_13473);
xnor UO_1684 (O_1684,N_14389,N_14317);
or UO_1685 (O_1685,N_13259,N_14502);
nand UO_1686 (O_1686,N_13953,N_14309);
or UO_1687 (O_1687,N_12052,N_12505);
and UO_1688 (O_1688,N_12184,N_14277);
nand UO_1689 (O_1689,N_13009,N_13715);
or UO_1690 (O_1690,N_12617,N_13660);
nand UO_1691 (O_1691,N_13457,N_12358);
or UO_1692 (O_1692,N_13966,N_14758);
and UO_1693 (O_1693,N_14229,N_14438);
nand UO_1694 (O_1694,N_12095,N_13713);
or UO_1695 (O_1695,N_13215,N_12004);
nand UO_1696 (O_1696,N_13798,N_14225);
or UO_1697 (O_1697,N_13844,N_13172);
nor UO_1698 (O_1698,N_12768,N_14859);
nor UO_1699 (O_1699,N_13571,N_14962);
nand UO_1700 (O_1700,N_14388,N_12691);
and UO_1701 (O_1701,N_12141,N_14098);
nand UO_1702 (O_1702,N_14938,N_13141);
and UO_1703 (O_1703,N_12459,N_14139);
and UO_1704 (O_1704,N_13383,N_13694);
nand UO_1705 (O_1705,N_13506,N_14209);
nor UO_1706 (O_1706,N_12343,N_12828);
nand UO_1707 (O_1707,N_14066,N_14567);
or UO_1708 (O_1708,N_13876,N_14532);
or UO_1709 (O_1709,N_12446,N_14918);
nor UO_1710 (O_1710,N_13646,N_14780);
or UO_1711 (O_1711,N_13546,N_12604);
nand UO_1712 (O_1712,N_14764,N_14506);
nand UO_1713 (O_1713,N_14770,N_13441);
and UO_1714 (O_1714,N_14082,N_12044);
and UO_1715 (O_1715,N_12518,N_12539);
and UO_1716 (O_1716,N_14410,N_14496);
or UO_1717 (O_1717,N_13585,N_14956);
nor UO_1718 (O_1718,N_13460,N_12682);
and UO_1719 (O_1719,N_14860,N_13104);
and UO_1720 (O_1720,N_13185,N_12611);
or UO_1721 (O_1721,N_13772,N_13483);
nand UO_1722 (O_1722,N_14133,N_14338);
nor UO_1723 (O_1723,N_12891,N_12886);
or UO_1724 (O_1724,N_12186,N_13215);
nand UO_1725 (O_1725,N_12002,N_14840);
and UO_1726 (O_1726,N_14182,N_12509);
and UO_1727 (O_1727,N_13110,N_14527);
and UO_1728 (O_1728,N_12018,N_14860);
and UO_1729 (O_1729,N_14605,N_14562);
nor UO_1730 (O_1730,N_14873,N_13609);
or UO_1731 (O_1731,N_13657,N_14265);
nand UO_1732 (O_1732,N_14328,N_13773);
and UO_1733 (O_1733,N_13332,N_13284);
nor UO_1734 (O_1734,N_13455,N_14437);
nor UO_1735 (O_1735,N_12212,N_13467);
or UO_1736 (O_1736,N_14980,N_12423);
and UO_1737 (O_1737,N_13361,N_13617);
nand UO_1738 (O_1738,N_12452,N_13864);
and UO_1739 (O_1739,N_13336,N_13644);
nand UO_1740 (O_1740,N_14241,N_13903);
nand UO_1741 (O_1741,N_12729,N_13753);
or UO_1742 (O_1742,N_14196,N_13584);
or UO_1743 (O_1743,N_13066,N_12637);
nand UO_1744 (O_1744,N_12380,N_13833);
nor UO_1745 (O_1745,N_13789,N_12002);
nand UO_1746 (O_1746,N_14677,N_14829);
or UO_1747 (O_1747,N_12205,N_13914);
or UO_1748 (O_1748,N_14122,N_13308);
and UO_1749 (O_1749,N_13866,N_14549);
nor UO_1750 (O_1750,N_13897,N_14145);
nand UO_1751 (O_1751,N_14133,N_14135);
or UO_1752 (O_1752,N_12856,N_12811);
or UO_1753 (O_1753,N_13776,N_14166);
and UO_1754 (O_1754,N_12590,N_12062);
and UO_1755 (O_1755,N_12564,N_13959);
and UO_1756 (O_1756,N_14600,N_12723);
nor UO_1757 (O_1757,N_12531,N_12941);
nand UO_1758 (O_1758,N_13704,N_12976);
nor UO_1759 (O_1759,N_14375,N_13226);
and UO_1760 (O_1760,N_14896,N_14174);
nor UO_1761 (O_1761,N_14125,N_13797);
and UO_1762 (O_1762,N_13679,N_14832);
nand UO_1763 (O_1763,N_12495,N_14659);
nor UO_1764 (O_1764,N_12502,N_12022);
and UO_1765 (O_1765,N_14675,N_13785);
and UO_1766 (O_1766,N_13450,N_14121);
nor UO_1767 (O_1767,N_13848,N_13180);
nor UO_1768 (O_1768,N_12906,N_13319);
and UO_1769 (O_1769,N_14041,N_14383);
or UO_1770 (O_1770,N_12040,N_14710);
or UO_1771 (O_1771,N_12524,N_13915);
nand UO_1772 (O_1772,N_14632,N_13675);
nand UO_1773 (O_1773,N_12980,N_12098);
nor UO_1774 (O_1774,N_14846,N_12856);
nor UO_1775 (O_1775,N_14453,N_13748);
nand UO_1776 (O_1776,N_13287,N_13137);
and UO_1777 (O_1777,N_12578,N_12119);
or UO_1778 (O_1778,N_12000,N_13919);
nor UO_1779 (O_1779,N_13550,N_12743);
or UO_1780 (O_1780,N_13968,N_13912);
nor UO_1781 (O_1781,N_14863,N_14137);
and UO_1782 (O_1782,N_12034,N_12757);
nand UO_1783 (O_1783,N_13356,N_13956);
or UO_1784 (O_1784,N_13511,N_14256);
and UO_1785 (O_1785,N_13302,N_13264);
or UO_1786 (O_1786,N_14368,N_14634);
or UO_1787 (O_1787,N_14995,N_12296);
and UO_1788 (O_1788,N_13706,N_14566);
nand UO_1789 (O_1789,N_12824,N_14431);
and UO_1790 (O_1790,N_13004,N_13695);
nor UO_1791 (O_1791,N_13701,N_12508);
or UO_1792 (O_1792,N_12773,N_13215);
and UO_1793 (O_1793,N_14338,N_14424);
nor UO_1794 (O_1794,N_13754,N_13532);
or UO_1795 (O_1795,N_12783,N_13015);
nand UO_1796 (O_1796,N_13753,N_14907);
nor UO_1797 (O_1797,N_12343,N_12200);
and UO_1798 (O_1798,N_13062,N_13825);
or UO_1799 (O_1799,N_12143,N_14512);
or UO_1800 (O_1800,N_12726,N_14790);
or UO_1801 (O_1801,N_13025,N_14448);
or UO_1802 (O_1802,N_12984,N_12588);
and UO_1803 (O_1803,N_12872,N_14058);
and UO_1804 (O_1804,N_12014,N_14703);
nand UO_1805 (O_1805,N_13403,N_12114);
nor UO_1806 (O_1806,N_13685,N_13206);
and UO_1807 (O_1807,N_12814,N_14923);
and UO_1808 (O_1808,N_12205,N_12484);
nor UO_1809 (O_1809,N_12451,N_13120);
nor UO_1810 (O_1810,N_12876,N_14177);
nor UO_1811 (O_1811,N_14024,N_12716);
nand UO_1812 (O_1812,N_13601,N_14702);
or UO_1813 (O_1813,N_13747,N_13571);
or UO_1814 (O_1814,N_14821,N_14290);
and UO_1815 (O_1815,N_14123,N_13912);
nor UO_1816 (O_1816,N_12053,N_12719);
nand UO_1817 (O_1817,N_13930,N_14313);
nand UO_1818 (O_1818,N_12710,N_13198);
nor UO_1819 (O_1819,N_14262,N_14258);
and UO_1820 (O_1820,N_14269,N_13030);
nand UO_1821 (O_1821,N_14672,N_14060);
and UO_1822 (O_1822,N_14944,N_12467);
nand UO_1823 (O_1823,N_13352,N_12250);
nor UO_1824 (O_1824,N_14520,N_13041);
nor UO_1825 (O_1825,N_14772,N_14489);
and UO_1826 (O_1826,N_12406,N_14658);
nor UO_1827 (O_1827,N_14472,N_12537);
nor UO_1828 (O_1828,N_13004,N_12010);
nor UO_1829 (O_1829,N_13219,N_13499);
or UO_1830 (O_1830,N_12697,N_13491);
nand UO_1831 (O_1831,N_14231,N_14828);
nor UO_1832 (O_1832,N_13749,N_13817);
nand UO_1833 (O_1833,N_14000,N_12250);
or UO_1834 (O_1834,N_12360,N_12959);
nand UO_1835 (O_1835,N_14045,N_13463);
or UO_1836 (O_1836,N_12777,N_12943);
nor UO_1837 (O_1837,N_13905,N_13018);
or UO_1838 (O_1838,N_14678,N_13514);
nor UO_1839 (O_1839,N_12987,N_13295);
nor UO_1840 (O_1840,N_12390,N_12362);
nor UO_1841 (O_1841,N_12685,N_13285);
or UO_1842 (O_1842,N_13221,N_14296);
nor UO_1843 (O_1843,N_12975,N_14743);
or UO_1844 (O_1844,N_14025,N_13865);
nor UO_1845 (O_1845,N_12805,N_12765);
and UO_1846 (O_1846,N_12688,N_12343);
or UO_1847 (O_1847,N_12570,N_14875);
and UO_1848 (O_1848,N_14942,N_12186);
xnor UO_1849 (O_1849,N_14076,N_14828);
and UO_1850 (O_1850,N_13710,N_13921);
nand UO_1851 (O_1851,N_13777,N_13803);
and UO_1852 (O_1852,N_12920,N_13149);
or UO_1853 (O_1853,N_12808,N_12984);
and UO_1854 (O_1854,N_12626,N_12939);
and UO_1855 (O_1855,N_13695,N_14108);
nor UO_1856 (O_1856,N_12033,N_12128);
nand UO_1857 (O_1857,N_12990,N_12167);
nand UO_1858 (O_1858,N_14585,N_13607);
and UO_1859 (O_1859,N_13128,N_12403);
nand UO_1860 (O_1860,N_12077,N_13256);
nor UO_1861 (O_1861,N_14770,N_12669);
nand UO_1862 (O_1862,N_14726,N_14075);
and UO_1863 (O_1863,N_14114,N_14151);
nor UO_1864 (O_1864,N_13534,N_13574);
nor UO_1865 (O_1865,N_12918,N_14749);
nor UO_1866 (O_1866,N_14010,N_13955);
nor UO_1867 (O_1867,N_14219,N_13171);
nor UO_1868 (O_1868,N_13591,N_14688);
and UO_1869 (O_1869,N_13464,N_13243);
nor UO_1870 (O_1870,N_13215,N_13375);
nand UO_1871 (O_1871,N_13839,N_13077);
or UO_1872 (O_1872,N_14532,N_13032);
or UO_1873 (O_1873,N_12741,N_13411);
and UO_1874 (O_1874,N_13209,N_13921);
nand UO_1875 (O_1875,N_14119,N_12083);
nor UO_1876 (O_1876,N_14212,N_14361);
and UO_1877 (O_1877,N_13444,N_12578);
nand UO_1878 (O_1878,N_14738,N_14377);
or UO_1879 (O_1879,N_13941,N_14203);
and UO_1880 (O_1880,N_13937,N_14508);
or UO_1881 (O_1881,N_14406,N_12561);
or UO_1882 (O_1882,N_13951,N_12234);
or UO_1883 (O_1883,N_13835,N_12269);
nor UO_1884 (O_1884,N_13803,N_12457);
or UO_1885 (O_1885,N_14805,N_12459);
nand UO_1886 (O_1886,N_14097,N_12571);
nor UO_1887 (O_1887,N_14233,N_12903);
nand UO_1888 (O_1888,N_14179,N_12353);
nand UO_1889 (O_1889,N_14281,N_13937);
nand UO_1890 (O_1890,N_13551,N_12499);
and UO_1891 (O_1891,N_12805,N_12250);
or UO_1892 (O_1892,N_14429,N_14345);
or UO_1893 (O_1893,N_14016,N_13259);
nor UO_1894 (O_1894,N_12391,N_14499);
nand UO_1895 (O_1895,N_13505,N_14477);
nor UO_1896 (O_1896,N_14860,N_12849);
and UO_1897 (O_1897,N_13560,N_14907);
or UO_1898 (O_1898,N_13206,N_13073);
or UO_1899 (O_1899,N_14562,N_12468);
and UO_1900 (O_1900,N_13665,N_12094);
and UO_1901 (O_1901,N_13691,N_12154);
nand UO_1902 (O_1902,N_14761,N_13550);
or UO_1903 (O_1903,N_12409,N_14496);
nand UO_1904 (O_1904,N_14897,N_13729);
nor UO_1905 (O_1905,N_13177,N_14482);
or UO_1906 (O_1906,N_13170,N_14393);
nor UO_1907 (O_1907,N_13815,N_12764);
nand UO_1908 (O_1908,N_13963,N_14433);
nand UO_1909 (O_1909,N_12090,N_13071);
and UO_1910 (O_1910,N_12103,N_14365);
or UO_1911 (O_1911,N_13941,N_14068);
and UO_1912 (O_1912,N_13979,N_14028);
nor UO_1913 (O_1913,N_13213,N_14899);
or UO_1914 (O_1914,N_14857,N_14345);
or UO_1915 (O_1915,N_14871,N_13180);
nand UO_1916 (O_1916,N_13196,N_12396);
and UO_1917 (O_1917,N_12700,N_13086);
nand UO_1918 (O_1918,N_14209,N_14733);
nor UO_1919 (O_1919,N_13812,N_14620);
nor UO_1920 (O_1920,N_13314,N_14082);
and UO_1921 (O_1921,N_13970,N_14014);
or UO_1922 (O_1922,N_12777,N_12704);
nor UO_1923 (O_1923,N_12341,N_12562);
and UO_1924 (O_1924,N_13434,N_14129);
and UO_1925 (O_1925,N_13483,N_14377);
and UO_1926 (O_1926,N_14017,N_13261);
and UO_1927 (O_1927,N_13671,N_12758);
and UO_1928 (O_1928,N_12520,N_14466);
or UO_1929 (O_1929,N_13695,N_12995);
and UO_1930 (O_1930,N_12297,N_14226);
or UO_1931 (O_1931,N_14669,N_14657);
or UO_1932 (O_1932,N_13495,N_14267);
and UO_1933 (O_1933,N_12853,N_13722);
nand UO_1934 (O_1934,N_12072,N_13377);
or UO_1935 (O_1935,N_14586,N_13115);
nand UO_1936 (O_1936,N_14546,N_14190);
and UO_1937 (O_1937,N_12908,N_14335);
nor UO_1938 (O_1938,N_12342,N_13842);
and UO_1939 (O_1939,N_13583,N_14433);
nand UO_1940 (O_1940,N_14282,N_12783);
nand UO_1941 (O_1941,N_12362,N_12270);
nand UO_1942 (O_1942,N_12816,N_12918);
and UO_1943 (O_1943,N_13945,N_12852);
nand UO_1944 (O_1944,N_14530,N_14575);
and UO_1945 (O_1945,N_14216,N_14528);
or UO_1946 (O_1946,N_14919,N_14111);
and UO_1947 (O_1947,N_12993,N_12794);
nand UO_1948 (O_1948,N_13935,N_12923);
nor UO_1949 (O_1949,N_13011,N_12915);
and UO_1950 (O_1950,N_14772,N_12155);
and UO_1951 (O_1951,N_12968,N_13102);
nor UO_1952 (O_1952,N_12716,N_14616);
or UO_1953 (O_1953,N_12353,N_13460);
and UO_1954 (O_1954,N_13860,N_14203);
nor UO_1955 (O_1955,N_13921,N_14960);
nand UO_1956 (O_1956,N_13349,N_13011);
nand UO_1957 (O_1957,N_13434,N_13662);
nor UO_1958 (O_1958,N_13254,N_14390);
nand UO_1959 (O_1959,N_14228,N_12224);
nand UO_1960 (O_1960,N_12387,N_12960);
nand UO_1961 (O_1961,N_14178,N_13415);
nor UO_1962 (O_1962,N_14221,N_12474);
or UO_1963 (O_1963,N_14824,N_14603);
nand UO_1964 (O_1964,N_13934,N_14634);
nand UO_1965 (O_1965,N_12579,N_14434);
or UO_1966 (O_1966,N_13826,N_12965);
and UO_1967 (O_1967,N_12735,N_13172);
or UO_1968 (O_1968,N_12971,N_13432);
and UO_1969 (O_1969,N_12095,N_12880);
nand UO_1970 (O_1970,N_12238,N_14071);
nand UO_1971 (O_1971,N_12510,N_12646);
nand UO_1972 (O_1972,N_12761,N_14075);
and UO_1973 (O_1973,N_14351,N_13062);
or UO_1974 (O_1974,N_12554,N_13074);
nand UO_1975 (O_1975,N_14161,N_13166);
or UO_1976 (O_1976,N_13435,N_13499);
nand UO_1977 (O_1977,N_14397,N_13863);
or UO_1978 (O_1978,N_13466,N_13426);
or UO_1979 (O_1979,N_12885,N_12140);
nand UO_1980 (O_1980,N_14286,N_12611);
and UO_1981 (O_1981,N_12317,N_14269);
or UO_1982 (O_1982,N_14240,N_14084);
and UO_1983 (O_1983,N_12112,N_12922);
and UO_1984 (O_1984,N_14198,N_12293);
nand UO_1985 (O_1985,N_14782,N_14321);
nor UO_1986 (O_1986,N_14028,N_12446);
nand UO_1987 (O_1987,N_14454,N_14876);
and UO_1988 (O_1988,N_14221,N_12194);
nor UO_1989 (O_1989,N_13423,N_13262);
or UO_1990 (O_1990,N_12722,N_12047);
nand UO_1991 (O_1991,N_12382,N_13902);
or UO_1992 (O_1992,N_14454,N_14119);
nor UO_1993 (O_1993,N_13095,N_12850);
nor UO_1994 (O_1994,N_12314,N_12014);
or UO_1995 (O_1995,N_13329,N_12298);
nand UO_1996 (O_1996,N_12692,N_14374);
or UO_1997 (O_1997,N_12047,N_13333);
nand UO_1998 (O_1998,N_13827,N_12764);
nor UO_1999 (O_1999,N_12411,N_13343);
endmodule